##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 01:18:08 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_single
  CLASS BLOCK ;
  SIZE 210.2200 BY 30.2600 ;
  FOREIGN S_term_single 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.632 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 29.5400 14.2200 30.2600 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21295 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.427 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.1708 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.7765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 29.5400 12.8400 30.2600 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.74 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.582 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 29.5400 11.4600 30.2600 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.92695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.1606 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.766 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 29.5400 10.5400 30.2600 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.738 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 29.5400 25.2600 30.2600 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1684 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6704 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.116 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 29.5400 23.8800 30.2600 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.356 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 29.5400 22.5000 30.2600 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.841 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.504 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 29.5400 21.1200 30.2600 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.836 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 29.5400 19.7400 30.2600 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.652 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 29.5400 18.3600 30.2600 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.938 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 29.5400 16.9800 30.2600 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.09735 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.291 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.8684 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.2645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.93 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 29.5400 15.6000 30.2600 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.49 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.818 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 29.5400 35.8400 30.2600 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.46455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 29.5400 34.4600 30.2600 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3324 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.184 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 29.5400 33.5400 30.2600 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.894 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 29.5400 32.1600 30.2600 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 29.5400 30.7800 30.2600 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.642 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.1325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.816 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.844 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 29.5400 29.4000 30.2600 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.154 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 29.5400 28.0200 30.2600 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.1128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.072 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 29.5400 26.6400 30.2600 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.202 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 29.5400 57.4600 30.2600 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3368 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.448 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 29.5400 56.5400 30.2600 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.2728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.333 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.547 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 29.5400 55.1600 30.2600 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.8168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.16 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 29.5400 53.7800 30.2600 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.6292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 63.0315 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.798 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 29.5400 52.4000 30.2600 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.358 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.322 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 29.5400 51.0200 30.2600 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9336 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.5905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 29.5400 49.6400 30.2600 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1852 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.952 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 29.5400 48.2600 30.2600 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.8384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 69.1145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.084 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 29.5400 46.8800 30.2600 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5264 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 29.5400 45.5000 30.2600 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 29.5400 44.1200 30.2600 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.296 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 29.5400 42.7400 30.2600 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.5428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.032 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 29.5400 41.3600 30.2600 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.552 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.642 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 29.5400 39.9800 30.2600 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.2116 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.9805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.846 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 29.5400 38.6000 30.2600 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.4056 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.9135 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5378 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 29.5400 37.2200 30.2600 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.984 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 29.5400 79.5400 30.2600 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.26695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.667 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.494 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 29.5400 78.1600 30.2600 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.723 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 29.5400 76.7800 30.2600 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.1572 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.7085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.284 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 29.5400 75.4000 30.2600 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.8136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 29.5400 74.0200 30.2600 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.414 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 29.5400 72.6400 30.2600 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.632 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 29.5400 71.2600 30.2600 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.522 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 29.5400 69.8800 30.2600 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.438 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 29.5400 68.5000 30.2600 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.988 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 29.5400 67.1200 30.2600 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 29.5400 65.7400 30.2600 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 29.5400 64.3600 30.2600 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.49 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.104 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 29.5400 62.9800 30.2600 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.466 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.094 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 29.5400 61.6000 30.2600 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.038 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 29.5400 60.2200 30.2600 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6265 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.9676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 29.5400 58.8400 30.2600 ;
    END
  END NN4BEG[0]
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2895 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.6388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.544 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 177.1400 29.5400 177.5200 30.2600 ;
    END
  END Co
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.62 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.67516 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.9277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 29.5400 84.6000 30.2600 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.97075 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.4057 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 29.5400 83.2200 30.2600 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.4739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.9214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 29.5400 81.8400 30.2600 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.808 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 32.2186 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 155.903 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 29.5400 80.4600 30.2600 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8348 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.0225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.772 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.0943 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 29.5400 106.2200 30.2600 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.584 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.367 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.3868 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 29.5400 104.8400 30.2600 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.5446 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 40.8714 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.333 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 29.5400 103.4600 30.2600 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 28.1632 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.84 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 29.5400 102.5400 30.2600 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.42 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.0676 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.664 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 29.5400 101.1600 30.2600 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2948 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3595 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 24.35 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.415 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 29.5400 99.7800 30.2600 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.082 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.8333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 29.5400 98.4000 30.2600 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.4173 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.8962 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 29.5400 97.0200 30.2600 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.392 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.7494 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.9811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 29.5400 95.6400 30.2600 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.844 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.3959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 29.5400 94.2600 30.2600 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 57.0984 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.409 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 29.5400 92.8800 30.2600 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.4739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.9214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 29.5400 91.5000 30.2600 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.39 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.6123 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 29.5400 90.1200 30.2600 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.25 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.055 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.5094 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 29.5400 88.7400 30.2600 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.95 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.3428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 29.5400 87.3600 30.2600 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.474 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.4752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.9277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 29.5400 85.9800 30.2600 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.48195 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.567 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.096 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.8664 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.8836 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 29.5400 127.8400 30.2600 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.14755 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.703 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.0915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.1038 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 29.5400 126.4600 30.2600 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.0896 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 52.1085 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.314 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 29.5400 125.5400 30.2600 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.8223 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.248 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 29.5400 124.1600 30.2600 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.40723 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.5881 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 29.5400 122.7800 30.2600 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42715 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.679 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.718 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.6072 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 119.588 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 29.5400 121.4000 30.2600 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.7305 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.7893 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 29.5400 120.0200 30.2600 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.17255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.203 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.78711 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.4874 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 29.5400 118.6400 30.2600 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.101 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 57.6142 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 310.013 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 29.5400 117.2600 30.2600 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.49 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.466 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.67138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.9088 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 29.5400 115.8800 30.2600 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.976 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.8186 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.9025 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 29.5400 114.5000 30.2600 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 42.9921 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.557 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 29.5400 113.1200 30.2600 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5129 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.3742 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 29.5400 111.7400 30.2600 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.19214 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.5126 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 29.5400 110.3600 30.2600 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.572 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.5821 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 102.72 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 29.5400 108.9800 30.2600 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.096 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.9192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.1478 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 29.5400 107.6000 30.2600 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.798 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3066 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.5094 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 29.5400 149.4600 30.2600 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.862 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.2325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.52296 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.7516 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 29.5400 148.5400 30.2600 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.474 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3431 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.2767 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 29.5400 147.1600 30.2600 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.27 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 16.8079 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 91.0283 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 29.5400 145.7800 30.2600 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.7708 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.7765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.62 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.67516 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.9277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 29.5400 144.4000 30.2600 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.0978 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.0409 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 29.5400 143.0200 30.2600 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.643 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 70.2959 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.214 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 29.5400 141.6400 30.2600 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.594 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.7607 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.613 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 29.5400 140.2600 30.2600 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19635 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.4828 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.81 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.2689 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 130.412 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 29.5400 138.8800 30.2600 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.86887 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.8962 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 29.5400 137.5000 30.2600 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6475 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.276 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.7318 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.7264 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 29.5400 136.1200 30.2600 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.05995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.438 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.8852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.4025 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 29.5400 134.7400 30.2600 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.27075 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.495 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.072 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.0575 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 29.5400 133.3600 30.2600 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.976 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.8774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 29.5400 131.9800 30.2600 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.27075 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.495 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.3657 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.0629 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 29.5400 130.6000 30.2600 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.128 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.1918 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 29.5400 129.2200 30.2600 ;
    END
  END SS4END[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2496 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.176 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.9024 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 74.4345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1708 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.195 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 57.1016 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 278.035 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.377 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.7086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 90.2467 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 474.157 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.96 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.7225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.038 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.31918 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.5723 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7548 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 63.4025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0123 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.6132 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 59.0393 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 315.516 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.7608 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 58.7265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.55317 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 71.7035 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 375.403 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.96905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.493 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.8512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 84.1785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4922 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.343 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.616 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.6321 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.34 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.889 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.0526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 58.1425 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 313.349 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5406 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.636 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.3544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.7444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 50.8456 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.698 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.4996 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 67.4205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.403 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.72799 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.1918 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.1612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.277 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 54.0909 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.723 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 49.3525 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 249.346 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.703 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.4478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.192 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 84.2456 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 439.629 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.217 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4756 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.3005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.3459 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2342 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.452 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 47.3645 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 232.374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 55.394 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.843 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.857 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.615 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 27.994 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.233 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.5588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 36.2494 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.05 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.729 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 64.6777 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 315.236 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.7298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.7724 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 36.9009 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 202.204 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.9588 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 111.642 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.0094 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7789 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.283 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 76.4085 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 377.657 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.758 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4399 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.0723 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5733 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.829 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 20.111 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 107.969 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.3968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 39.6381 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.855 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5211 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.4874 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7387 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.799 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6962 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.255 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2324 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.2296 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.34 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.173 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 28.6600 210.2200 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9612 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 26.6200 210.2200 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.267 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 24.9200 210.2200 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.3568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.04 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 22.8800 210.2200 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.672 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 21.1800 210.2200 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.562 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 19.1400 210.2200 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 17.4400 210.2200 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 15.7400 210.2200 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.6658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.688 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 13.7000 210.2200 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.5068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.84 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 12.0000 210.2200 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 10.3000 210.2200 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.8778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.152 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 8.2600 210.2200 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.2908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.688 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 6.5600 210.2200 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.002 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 4.5200 210.2200 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.888 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.9304 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 2.8200 210.2200 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.1928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.832 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 1.1200 210.2200 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.9268 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.5565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.9644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.888 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 27.6250 210.2200 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.081 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.754 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.6925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5374 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.944 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 25.9250 210.2200 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6596 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.776 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.5028 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.4365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.19 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 24.2250 210.2200 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.4062 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.9535 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1026 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.488 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 22.5250 210.2200 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.0368 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.0695 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.832 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 20.8250 210.2200 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.168 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 19.1250 210.2200 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.856 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.36 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.8154 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 58.9995 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 17.4250 210.2200 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.6848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.456 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 15.7250 210.2200 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6562 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.772 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.31 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 14.0250 210.2200 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.6448 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 88.0355 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 12.3250 210.2200 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.8728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 10.6250 210.2200 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8873 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 8.9250 210.2200 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3672 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.432 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.233 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4134 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.616 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 7.2250 210.2200 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.1504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.6745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 5.5250 210.2200 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.0956 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 75.4005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.43 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 3.8250 210.2200 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.4364 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 57.0675 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.463 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 2.1250 210.2200 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.0425 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.9969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 149.5400 0.0000 149.9200 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.537 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.4035 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.3145 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 144.0200 0.0000 144.4000 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.597 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.6664 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.2044 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 138.9600 0.0000 139.3400 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.367 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 32.6915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 159.072 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 133.4400 0.0000 133.8200 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7292 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.1038 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 128.3800 0.0000 128.7600 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.11 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.9292 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 133.714 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 123.3200 0.0000 123.7000 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.319 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.9053 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.1164 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 117.8000 0.0000 118.1800 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.893 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3041 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.978 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 112.2800 0.0000 112.6600 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.607 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 34.4865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 165.022 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 107.6800 0.0000 108.0600 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.929 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.2097 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.248 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 102.1600 0.0000 102.5400 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7947 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.8459 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 97.1000 0.0000 97.4800 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.467 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 28.7896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 133.664 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.5800 0.0000 91.9600 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.511 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.4676 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.211 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 86.0600 0.0000 86.4400 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.285 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 38.1324 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 204.409 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 81.4600 0.0000 81.8400 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.999 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.91289 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.1792 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 75.9400 0.0000 76.3200 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.319 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.6009 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 130.594 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 70.8800 0.0000 71.2600 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.799 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.4676 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.211 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 65.8200 0.0000 66.2000 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.119 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.528 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.77 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 60.3000 0.0000 60.6800 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.25 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.0802 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.978 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 55.2400 0.0000 55.6200 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6035 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.8648 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.1800 0.0000 50.5600 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.061 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.7224 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 199.2200 29.5400 199.6000 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.45 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 197.3800 29.5400 197.7600 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.449 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 195.0800 29.5400 195.4600 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.6098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.056 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 192.7800 29.5400 193.1600 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.749 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.4800 29.5400 190.8600 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.1800 29.5400 188.5600 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.391 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 185.8800 29.5400 186.2600 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.2344 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.328 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 184.0400 29.5400 184.4200 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 181.7400 29.5400 182.1200 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.149 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 179.4400 29.5400 179.8200 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0778 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.281 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.8400 29.5400 175.2200 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2262 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.787 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 172.5400 29.5400 172.9200 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.965 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 170.2400 29.5400 170.6200 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4378 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.963 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 168.4000 29.5400 168.7800 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.752 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 166.1000 29.5400 166.4800 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.839 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 163.8000 29.5400 164.1800 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.059 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.5000 29.5400 161.8800 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1416 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.246 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.2000 29.5400 159.5800 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.569 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 156.9000 29.5400 157.2800 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.768 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 155.0600 29.5400 155.4400 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 204.6600 6.0700 ;
        RECT 5.5600 23.0000 204.6600 25.0000 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 202.6600 15.0600 204.6600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 202.6600 9.6200 204.6600 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 202.6600 20.5000 204.6600 20.9800 ;
      LAYER met4 ;
        RECT 202.6600 4.0700 204.6600 25.0000 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 207.6600 3.0700 ;
        RECT 2.5600 26.0000 207.6600 28.0000 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 205.6600 6.9000 207.6600 7.3800 ;
        RECT 205.6600 12.3400 207.6600 12.8200 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 205.6600 17.7800 207.6600 18.2600 ;
      LAYER met4 ;
        RECT 205.6600 1.0700 207.6600 28.0000 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.6300 29.3700 210.2200 30.2600 ;
      RECT 148.7100 29.3700 148.9100 30.2600 ;
      RECT 147.3300 29.3700 147.9900 30.2600 ;
      RECT 145.9500 29.3700 146.6100 30.2600 ;
      RECT 144.5700 29.3700 145.2300 30.2600 ;
      RECT 143.1900 29.3700 143.8500 30.2600 ;
      RECT 141.8100 29.3700 142.4700 30.2600 ;
      RECT 140.4300 29.3700 141.0900 30.2600 ;
      RECT 139.0500 29.3700 139.7100 30.2600 ;
      RECT 137.6700 29.3700 138.3300 30.2600 ;
      RECT 136.2900 29.3700 136.9500 30.2600 ;
      RECT 134.9100 29.3700 135.5700 30.2600 ;
      RECT 133.5300 29.3700 134.1900 30.2600 ;
      RECT 132.1500 29.3700 132.8100 30.2600 ;
      RECT 130.7700 29.3700 131.4300 30.2600 ;
      RECT 129.3900 29.3700 130.0500 30.2600 ;
      RECT 128.0100 29.3700 128.6700 30.2600 ;
      RECT 126.6300 29.3700 127.2900 30.2600 ;
      RECT 125.7100 29.3700 125.9100 30.2600 ;
      RECT 124.3300 29.3700 124.9900 30.2600 ;
      RECT 122.9500 29.3700 123.6100 30.2600 ;
      RECT 121.5700 29.3700 122.2300 30.2600 ;
      RECT 120.1900 29.3700 120.8500 30.2600 ;
      RECT 118.8100 29.3700 119.4700 30.2600 ;
      RECT 117.4300 29.3700 118.0900 30.2600 ;
      RECT 116.0500 29.3700 116.7100 30.2600 ;
      RECT 114.6700 29.3700 115.3300 30.2600 ;
      RECT 113.2900 29.3700 113.9500 30.2600 ;
      RECT 111.9100 29.3700 112.5700 30.2600 ;
      RECT 110.5300 29.3700 111.1900 30.2600 ;
      RECT 109.1500 29.3700 109.8100 30.2600 ;
      RECT 107.7700 29.3700 108.4300 30.2600 ;
      RECT 106.3900 29.3700 107.0500 30.2600 ;
      RECT 105.0100 29.3700 105.6700 30.2600 ;
      RECT 103.6300 29.3700 104.2900 30.2600 ;
      RECT 102.7100 29.3700 102.9100 30.2600 ;
      RECT 101.3300 29.3700 101.9900 30.2600 ;
      RECT 99.9500 29.3700 100.6100 30.2600 ;
      RECT 98.5700 29.3700 99.2300 30.2600 ;
      RECT 97.1900 29.3700 97.8500 30.2600 ;
      RECT 95.8100 29.3700 96.4700 30.2600 ;
      RECT 94.4300 29.3700 95.0900 30.2600 ;
      RECT 93.0500 29.3700 93.7100 30.2600 ;
      RECT 91.6700 29.3700 92.3300 30.2600 ;
      RECT 90.2900 29.3700 90.9500 30.2600 ;
      RECT 88.9100 29.3700 89.5700 30.2600 ;
      RECT 87.5300 29.3700 88.1900 30.2600 ;
      RECT 86.1500 29.3700 86.8100 30.2600 ;
      RECT 84.7700 29.3700 85.4300 30.2600 ;
      RECT 83.3900 29.3700 84.0500 30.2600 ;
      RECT 82.0100 29.3700 82.6700 30.2600 ;
      RECT 80.6300 29.3700 81.2900 30.2600 ;
      RECT 79.7100 29.3700 79.9100 30.2600 ;
      RECT 78.3300 29.3700 78.9900 30.2600 ;
      RECT 76.9500 29.3700 77.6100 30.2600 ;
      RECT 75.5700 29.3700 76.2300 30.2600 ;
      RECT 74.1900 29.3700 74.8500 30.2600 ;
      RECT 72.8100 29.3700 73.4700 30.2600 ;
      RECT 71.4300 29.3700 72.0900 30.2600 ;
      RECT 70.0500 29.3700 70.7100 30.2600 ;
      RECT 68.6700 29.3700 69.3300 30.2600 ;
      RECT 67.2900 29.3700 67.9500 30.2600 ;
      RECT 65.9100 29.3700 66.5700 30.2600 ;
      RECT 64.5300 29.3700 65.1900 30.2600 ;
      RECT 63.1500 29.3700 63.8100 30.2600 ;
      RECT 61.7700 29.3700 62.4300 30.2600 ;
      RECT 60.3900 29.3700 61.0500 30.2600 ;
      RECT 59.0100 29.3700 59.6700 30.2600 ;
      RECT 57.6300 29.3700 58.2900 30.2600 ;
      RECT 56.7100 29.3700 56.9100 30.2600 ;
      RECT 55.3300 29.3700 55.9900 30.2600 ;
      RECT 53.9500 29.3700 54.6100 30.2600 ;
      RECT 52.5700 29.3700 53.2300 30.2600 ;
      RECT 51.1900 29.3700 51.8500 30.2600 ;
      RECT 49.8100 29.3700 50.4700 30.2600 ;
      RECT 48.4300 29.3700 49.0900 30.2600 ;
      RECT 47.0500 29.3700 47.7100 30.2600 ;
      RECT 45.6700 29.3700 46.3300 30.2600 ;
      RECT 44.2900 29.3700 44.9500 30.2600 ;
      RECT 42.9100 29.3700 43.5700 30.2600 ;
      RECT 41.5300 29.3700 42.1900 30.2600 ;
      RECT 40.1500 29.3700 40.8100 30.2600 ;
      RECT 38.7700 29.3700 39.4300 30.2600 ;
      RECT 37.3900 29.3700 38.0500 30.2600 ;
      RECT 36.0100 29.3700 36.6700 30.2600 ;
      RECT 34.6300 29.3700 35.2900 30.2600 ;
      RECT 33.7100 29.3700 33.9100 30.2600 ;
      RECT 32.3300 29.3700 32.9900 30.2600 ;
      RECT 30.9500 29.3700 31.6100 30.2600 ;
      RECT 29.5700 29.3700 30.2300 30.2600 ;
      RECT 28.1900 29.3700 28.8500 30.2600 ;
      RECT 26.8100 29.3700 27.4700 30.2600 ;
      RECT 25.4300 29.3700 26.0900 30.2600 ;
      RECT 24.0500 29.3700 24.7100 30.2600 ;
      RECT 22.6700 29.3700 23.3300 30.2600 ;
      RECT 21.2900 29.3700 21.9500 30.2600 ;
      RECT 19.9100 29.3700 20.5700 30.2600 ;
      RECT 18.5300 29.3700 19.1900 30.2600 ;
      RECT 17.1500 29.3700 17.8100 30.2600 ;
      RECT 15.7700 29.3700 16.4300 30.2600 ;
      RECT 14.3900 29.3700 15.0500 30.2600 ;
      RECT 13.0100 29.3700 13.6700 30.2600 ;
      RECT 11.6300 29.3700 12.2900 30.2600 ;
      RECT 10.7100 29.3700 10.9100 30.2600 ;
      RECT 0.0000 29.3700 9.9900 30.2600 ;
      RECT 0.0000 28.9850 210.2200 29.3700 ;
      RECT 0.5000 28.4750 210.2200 28.9850 ;
      RECT 0.0000 27.9650 210.2200 28.4750 ;
      RECT 0.0000 27.4550 209.7200 27.9650 ;
      RECT 0.0000 26.9450 210.2200 27.4550 ;
      RECT 0.5000 26.4350 210.2200 26.9450 ;
      RECT 0.0000 26.2650 210.2200 26.4350 ;
      RECT 0.0000 25.7550 209.7200 26.2650 ;
      RECT 0.0000 25.2450 210.2200 25.7550 ;
      RECT 0.5000 24.7350 210.2200 25.2450 ;
      RECT 0.0000 24.5650 210.2200 24.7350 ;
      RECT 0.0000 24.0550 209.7200 24.5650 ;
      RECT 0.0000 23.2050 210.2200 24.0550 ;
      RECT 0.5000 22.8650 210.2200 23.2050 ;
      RECT 0.5000 22.6950 209.7200 22.8650 ;
      RECT 0.0000 22.3550 209.7200 22.6950 ;
      RECT 0.0000 21.5050 210.2200 22.3550 ;
      RECT 0.5000 21.1650 210.2200 21.5050 ;
      RECT 0.5000 20.9950 209.7200 21.1650 ;
      RECT 0.0000 20.6550 209.7200 20.9950 ;
      RECT 0.0000 19.4650 210.2200 20.6550 ;
      RECT 0.5000 18.9550 209.7200 19.4650 ;
      RECT 0.0000 17.7650 210.2200 18.9550 ;
      RECT 0.5000 17.2550 209.7200 17.7650 ;
      RECT 0.0000 16.0650 210.2200 17.2550 ;
      RECT 0.5000 15.5550 209.7200 16.0650 ;
      RECT 0.0000 14.3650 210.2200 15.5550 ;
      RECT 0.0000 14.0250 209.7200 14.3650 ;
      RECT 0.5000 13.8550 209.7200 14.0250 ;
      RECT 0.5000 13.5150 210.2200 13.8550 ;
      RECT 0.0000 12.6650 210.2200 13.5150 ;
      RECT 0.0000 12.3250 209.7200 12.6650 ;
      RECT 0.5000 12.1550 209.7200 12.3250 ;
      RECT 0.5000 11.8150 210.2200 12.1550 ;
      RECT 0.0000 10.9650 210.2200 11.8150 ;
      RECT 0.0000 10.6250 209.7200 10.9650 ;
      RECT 0.5000 10.4550 209.7200 10.6250 ;
      RECT 0.5000 10.1150 210.2200 10.4550 ;
      RECT 0.0000 9.2650 210.2200 10.1150 ;
      RECT 0.0000 8.7550 209.7200 9.2650 ;
      RECT 0.0000 8.5850 210.2200 8.7550 ;
      RECT 0.5000 8.0750 210.2200 8.5850 ;
      RECT 0.0000 7.5650 210.2200 8.0750 ;
      RECT 0.0000 7.0550 209.7200 7.5650 ;
      RECT 0.0000 6.8850 210.2200 7.0550 ;
      RECT 0.5000 6.3750 210.2200 6.8850 ;
      RECT 0.0000 5.8650 210.2200 6.3750 ;
      RECT 0.0000 5.3550 209.7200 5.8650 ;
      RECT 0.0000 4.8450 210.2200 5.3550 ;
      RECT 0.5000 4.3350 210.2200 4.8450 ;
      RECT 0.0000 4.1650 210.2200 4.3350 ;
      RECT 0.0000 3.6550 209.7200 4.1650 ;
      RECT 0.0000 3.1450 210.2200 3.6550 ;
      RECT 0.5000 2.6350 210.2200 3.1450 ;
      RECT 0.0000 2.4650 210.2200 2.6350 ;
      RECT 0.0000 1.9550 209.7200 2.4650 ;
      RECT 0.0000 1.4450 210.2200 1.9550 ;
      RECT 0.5000 0.9350 210.2200 1.4450 ;
      RECT 0.0000 0.0000 210.2200 0.9350 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 210.2200 30.2600 ;
    LAYER met2 ;
      RECT 199.7400 29.4000 210.2200 30.2600 ;
      RECT 197.9000 29.4000 199.0800 30.2600 ;
      RECT 195.6000 29.4000 197.2400 30.2600 ;
      RECT 193.3000 29.4000 194.9400 30.2600 ;
      RECT 191.0000 29.4000 192.6400 30.2600 ;
      RECT 188.7000 29.4000 190.3400 30.2600 ;
      RECT 186.4000 29.4000 188.0400 30.2600 ;
      RECT 184.5600 29.4000 185.7400 30.2600 ;
      RECT 182.2600 29.4000 183.9000 30.2600 ;
      RECT 179.9600 29.4000 181.6000 30.2600 ;
      RECT 177.6600 29.4000 179.3000 30.2600 ;
      RECT 175.3600 29.4000 177.0000 30.2600 ;
      RECT 173.0600 29.4000 174.7000 30.2600 ;
      RECT 170.7600 29.4000 172.4000 30.2600 ;
      RECT 168.9200 29.4000 170.1000 30.2600 ;
      RECT 166.6200 29.4000 168.2600 30.2600 ;
      RECT 164.3200 29.4000 165.9600 30.2600 ;
      RECT 162.0200 29.4000 163.6600 30.2600 ;
      RECT 159.7200 29.4000 161.3600 30.2600 ;
      RECT 157.4200 29.4000 159.0600 30.2600 ;
      RECT 155.5800 29.4000 156.7600 30.2600 ;
      RECT 0.0000 29.4000 154.9200 30.2600 ;
      RECT 0.0000 28.9400 210.2200 29.4000 ;
      RECT 0.0000 28.5200 209.5950 28.9400 ;
      RECT 0.0000 27.9200 210.2200 28.5200 ;
      RECT 0.6250 27.5000 210.2200 27.9200 ;
      RECT 0.0000 26.9000 210.2200 27.5000 ;
      RECT 0.0000 26.4800 209.5950 26.9000 ;
      RECT 0.0000 26.2200 210.2200 26.4800 ;
      RECT 0.6250 25.8000 210.2200 26.2200 ;
      RECT 0.0000 25.2000 210.2200 25.8000 ;
      RECT 0.0000 24.7800 209.5950 25.2000 ;
      RECT 0.0000 24.5200 210.2200 24.7800 ;
      RECT 0.6250 24.1000 210.2200 24.5200 ;
      RECT 0.0000 23.1600 210.2200 24.1000 ;
      RECT 0.0000 22.8200 209.5950 23.1600 ;
      RECT 0.6250 22.7400 209.5950 22.8200 ;
      RECT 0.6250 22.4000 210.2200 22.7400 ;
      RECT 0.0000 21.4600 210.2200 22.4000 ;
      RECT 0.0000 21.1200 209.5950 21.4600 ;
      RECT 0.6250 21.0400 209.5950 21.1200 ;
      RECT 0.6250 20.7000 210.2200 21.0400 ;
      RECT 0.0000 19.4200 210.2200 20.7000 ;
      RECT 0.6250 19.0000 209.5950 19.4200 ;
      RECT 0.0000 17.7200 210.2200 19.0000 ;
      RECT 0.6250 17.3000 209.5950 17.7200 ;
      RECT 0.0000 16.0200 210.2200 17.3000 ;
      RECT 0.6250 15.6000 209.5950 16.0200 ;
      RECT 0.0000 14.3200 210.2200 15.6000 ;
      RECT 0.6250 13.9800 210.2200 14.3200 ;
      RECT 0.6250 13.9000 209.5950 13.9800 ;
      RECT 0.0000 13.5600 209.5950 13.9000 ;
      RECT 0.0000 12.6200 210.2200 13.5600 ;
      RECT 0.6250 12.2800 210.2200 12.6200 ;
      RECT 0.6250 12.2000 209.5950 12.2800 ;
      RECT 0.0000 11.8600 209.5950 12.2000 ;
      RECT 0.0000 10.9200 210.2200 11.8600 ;
      RECT 0.6250 10.5800 210.2200 10.9200 ;
      RECT 0.6250 10.5000 209.5950 10.5800 ;
      RECT 0.0000 10.1600 209.5950 10.5000 ;
      RECT 0.0000 9.2200 210.2200 10.1600 ;
      RECT 0.6250 8.8000 210.2200 9.2200 ;
      RECT 0.0000 8.5400 210.2200 8.8000 ;
      RECT 0.0000 8.1200 209.5950 8.5400 ;
      RECT 0.0000 7.5200 210.2200 8.1200 ;
      RECT 0.6250 7.1000 210.2200 7.5200 ;
      RECT 0.0000 6.8400 210.2200 7.1000 ;
      RECT 0.0000 6.4200 209.5950 6.8400 ;
      RECT 0.0000 5.8200 210.2200 6.4200 ;
      RECT 0.6250 5.4000 210.2200 5.8200 ;
      RECT 0.0000 4.8000 210.2200 5.4000 ;
      RECT 0.0000 4.3800 209.5950 4.8000 ;
      RECT 0.0000 4.1200 210.2200 4.3800 ;
      RECT 0.6250 3.7000 210.2200 4.1200 ;
      RECT 0.0000 3.1000 210.2200 3.7000 ;
      RECT 0.0000 2.6800 209.5950 3.1000 ;
      RECT 0.0000 2.4200 210.2200 2.6800 ;
      RECT 0.6250 2.0000 210.2200 2.4200 ;
      RECT 0.0000 1.4000 210.2200 2.0000 ;
      RECT 0.0000 0.9800 209.5950 1.4000 ;
      RECT 0.0000 0.8600 210.2200 0.9800 ;
      RECT 150.0600 0.0000 210.2200 0.8600 ;
      RECT 144.5400 0.0000 149.4000 0.8600 ;
      RECT 139.4800 0.0000 143.8800 0.8600 ;
      RECT 133.9600 0.0000 138.8200 0.8600 ;
      RECT 128.9000 0.0000 133.3000 0.8600 ;
      RECT 123.8400 0.0000 128.2400 0.8600 ;
      RECT 118.3200 0.0000 123.1800 0.8600 ;
      RECT 112.8000 0.0000 117.6600 0.8600 ;
      RECT 108.2000 0.0000 112.1400 0.8600 ;
      RECT 102.6800 0.0000 107.5400 0.8600 ;
      RECT 97.6200 0.0000 102.0200 0.8600 ;
      RECT 92.1000 0.0000 96.9600 0.8600 ;
      RECT 86.5800 0.0000 91.4400 0.8600 ;
      RECT 81.9800 0.0000 85.9200 0.8600 ;
      RECT 76.4600 0.0000 81.3200 0.8600 ;
      RECT 71.4000 0.0000 75.8000 0.8600 ;
      RECT 66.3400 0.0000 70.7400 0.8600 ;
      RECT 60.8200 0.0000 65.6800 0.8600 ;
      RECT 55.7600 0.0000 60.1600 0.8600 ;
      RECT 50.7000 0.0000 55.1000 0.8600 ;
      RECT 0.0000 0.0000 50.0400 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 210.2200 30.2600 ;
      RECT 207.9600 25.7000 210.2200 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 210.2200 25.7000 ;
      RECT 204.9600 22.7000 210.2200 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 210.2200 22.7000 ;
      RECT 204.9600 20.2000 210.2200 21.2800 ;
      RECT 7.8600 20.2000 202.3600 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 210.2200 20.2000 ;
      RECT 207.9600 17.4800 210.2200 18.5600 ;
      RECT 4.8600 17.4800 205.3600 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 210.2200 17.4800 ;
      RECT 204.9600 14.7600 210.2200 15.8400 ;
      RECT 7.8600 14.7600 202.3600 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 210.2200 14.7600 ;
      RECT 207.9600 12.0400 210.2200 13.1200 ;
      RECT 4.8600 12.0400 205.3600 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 210.2200 12.0400 ;
      RECT 204.9600 9.3200 210.2200 10.4000 ;
      RECT 7.8600 9.3200 202.3600 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 210.2200 9.3200 ;
      RECT 207.9600 6.6000 210.2200 7.6800 ;
      RECT 4.8600 6.6000 205.3600 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 210.2200 6.6000 ;
      RECT 204.9600 3.7700 210.2200 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 210.2200 3.7700 ;
      RECT 207.9600 0.7700 210.2200 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 210.2200 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 210.2200 30.2600 ;
      RECT 4.8600 25.3000 205.3600 28.3000 ;
      RECT 204.9600 3.7700 205.3600 25.3000 ;
      RECT 7.8600 3.7700 202.3600 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 207.9600 0.7700 210.2200 28.3000 ;
      RECT 4.8600 0.7700 205.3600 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 210.2200 0.7700 ;
  END
END S_term_single

END LIBRARY
