magic
tech sky130A
magscale 1 2
timestamp 1762063561
<< obsli1 >>
rect 1104 2159 21988 22865
<< obsm1 >>
rect 1104 2128 21988 22896
<< metal2 >>
rect 5170 24475 5226 25275
rect 5814 24475 5870 25275
rect 7102 24475 7158 25275
rect 7746 24475 7802 25275
rect 9034 24475 9090 25275
rect 9678 24475 9734 25275
rect 10966 24475 11022 25275
rect 11610 24475 11666 25275
rect 12254 24475 12310 25275
rect 12898 24475 12954 25275
rect 13542 24475 13598 25275
rect 14186 24475 14242 25275
rect 14830 24475 14886 25275
rect 16118 24475 16174 25275
rect 16762 24475 16818 25275
rect 17406 24475 17462 25275
rect 18050 24475 18106 25275
rect 19338 24475 19394 25275
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
<< obsm2 >>
rect 1122 24419 5114 24562
rect 5282 24419 5758 24562
rect 5926 24419 7046 24562
rect 7214 24419 7690 24562
rect 7858 24419 8978 24562
rect 9146 24419 9622 24562
rect 9790 24419 10910 24562
rect 11078 24419 11554 24562
rect 11722 24419 12198 24562
rect 12366 24419 12842 24562
rect 13010 24419 13486 24562
rect 13654 24419 14130 24562
rect 14298 24419 14774 24562
rect 14942 24419 16062 24562
rect 16230 24419 16706 24562
rect 16874 24419 17350 24562
rect 17518 24419 17994 24562
rect 18162 24419 19282 24562
rect 19450 24419 21692 24562
rect 1122 856 21692 24419
rect 1122 734 3182 856
rect 3350 734 3826 856
rect 3994 734 4470 856
rect 4638 734 5114 856
rect 5282 734 5758 856
rect 5926 734 6402 856
rect 6570 734 7046 856
rect 7214 734 7690 856
rect 7858 734 8334 856
rect 8502 734 8978 856
rect 9146 734 9622 856
rect 9790 734 10266 856
rect 10434 734 10910 856
rect 11078 734 11554 856
rect 11722 734 12198 856
rect 12366 734 12842 856
rect 13010 734 13486 856
rect 13654 734 14130 856
rect 14298 734 14774 856
rect 14942 734 15418 856
rect 15586 734 16062 856
rect 16230 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17994 856
rect 18162 734 18638 856
rect 18806 734 21692 856
<< metal3 >>
rect 0 21768 800 21888
rect 22331 21768 23131 21888
rect 0 21088 800 21208
rect 22331 21088 23131 21208
rect 0 20408 800 20528
rect 22331 20408 23131 20528
rect 0 19728 800 19848
rect 22331 19728 23131 19848
rect 0 19048 800 19168
rect 22331 19048 23131 19168
rect 0 18368 800 18488
rect 22331 18368 23131 18488
rect 0 17688 800 17808
rect 22331 17688 23131 17808
rect 0 17008 800 17128
rect 22331 17008 23131 17128
rect 0 16328 800 16448
rect 22331 16328 23131 16448
rect 0 15648 800 15768
rect 22331 15648 23131 15768
rect 0 14968 800 15088
rect 22331 14968 23131 15088
rect 0 14288 800 14408
rect 22331 14288 23131 14408
rect 0 13608 800 13728
rect 22331 13608 23131 13728
rect 0 12928 800 13048
rect 22331 12928 23131 13048
rect 0 12248 800 12368
rect 22331 12248 23131 12368
rect 0 11568 800 11688
rect 22331 11568 23131 11688
rect 0 10888 800 11008
rect 22331 10888 23131 11008
rect 0 10208 800 10328
rect 22331 10208 23131 10328
rect 0 9528 800 9648
rect 22331 9528 23131 9648
rect 0 8848 800 8968
rect 22331 8848 23131 8968
rect 0 8168 800 8288
rect 22331 8168 23131 8288
rect 0 7488 800 7608
rect 22331 7488 23131 7608
rect 0 6808 800 6928
rect 22331 6808 23131 6928
rect 0 6128 800 6248
rect 22331 6128 23131 6248
rect 0 5448 800 5568
rect 22331 5448 23131 5568
rect 0 4768 800 4888
rect 22331 4768 23131 4888
rect 0 4088 800 4208
rect 22331 4088 23131 4208
rect 0 3408 800 3528
rect 22331 3408 23131 3528
rect 0 2728 800 2848
rect 0 2048 800 2168
rect 0 1368 800 1488
rect 0 688 800 808
<< obsm3 >>
rect 800 21968 22331 22881
rect 880 21688 22251 21968
rect 800 21288 22331 21688
rect 880 21008 22251 21288
rect 800 20608 22331 21008
rect 880 20328 22251 20608
rect 800 19928 22331 20328
rect 880 19648 22251 19928
rect 800 19248 22331 19648
rect 880 18968 22251 19248
rect 800 18568 22331 18968
rect 880 18288 22251 18568
rect 800 17888 22331 18288
rect 880 17608 22251 17888
rect 800 17208 22331 17608
rect 880 16928 22251 17208
rect 800 16528 22331 16928
rect 880 16248 22251 16528
rect 800 15848 22331 16248
rect 880 15568 22251 15848
rect 800 15168 22331 15568
rect 880 14888 22251 15168
rect 800 14488 22331 14888
rect 880 14208 22251 14488
rect 800 13808 22331 14208
rect 880 13528 22251 13808
rect 800 13128 22331 13528
rect 880 12848 22251 13128
rect 800 12448 22331 12848
rect 880 12168 22251 12448
rect 800 11768 22331 12168
rect 880 11488 22251 11768
rect 800 11088 22331 11488
rect 880 10808 22251 11088
rect 800 10408 22331 10808
rect 880 10128 22251 10408
rect 800 9728 22331 10128
rect 880 9448 22251 9728
rect 800 9048 22331 9448
rect 880 8768 22251 9048
rect 800 8368 22331 8768
rect 880 8088 22251 8368
rect 800 7688 22331 8088
rect 880 7408 22251 7688
rect 800 7008 22331 7408
rect 880 6728 22251 7008
rect 800 6328 22331 6728
rect 880 6048 22251 6328
rect 800 5648 22331 6048
rect 880 5368 22251 5648
rect 800 4968 22331 5368
rect 880 4688 22251 4968
rect 800 4288 22331 4688
rect 880 4008 22251 4288
rect 800 3608 22331 4008
rect 880 3328 22251 3608
rect 800 2928 22331 3328
rect 880 2648 22331 2928
rect 800 2248 22331 2648
rect 880 1968 22331 2248
rect 800 1568 22331 1968
rect 880 1288 22331 1568
rect 800 888 22331 1288
rect 880 718 22331 888
<< metal4 >>
rect 3554 2128 3874 22896
rect 4214 2128 4534 22896
rect 8775 2128 9095 22896
rect 9435 2128 9755 22896
rect 13996 2128 14316 22896
rect 14656 2128 14976 22896
rect 19217 2128 19537 22896
rect 19877 2128 20197 22896
<< obsm4 >>
rect 3003 6427 3474 21181
rect 3954 6427 4134 21181
rect 4614 6427 8695 21181
rect 9175 6427 9355 21181
rect 9835 6427 13916 21181
rect 14396 6427 14576 21181
rect 15056 6427 17789 21181
<< metal5 >>
rect 1056 20764 22036 21084
rect 1056 20104 22036 20424
rect 1056 15596 22036 15916
rect 1056 14936 22036 15256
rect 1056 10428 22036 10748
rect 1056 9768 22036 10088
rect 1056 5260 22036 5580
rect 1056 4600 22036 4920
<< labels >>
rlabel metal3 s 0 19728 800 19848 6 spi_cs_n
port 1 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 spi_miso
port 2 nsew signal output
rlabel metal2 s 16762 24475 16818 25275 6 spi_mosi
port 3 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 spi_sck
port 4 nsew signal input
rlabel metal4 s 3554 2128 3874 22896 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 8775 2128 9095 22896 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 13996 2128 14316 22896 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 19217 2128 19537 22896 6 vccd1
port 5 nsew power bidirectional
rlabel metal5 s 1056 4600 22036 4920 6 vccd1
port 5 nsew power bidirectional
rlabel metal5 s 1056 9768 22036 10088 6 vccd1
port 5 nsew power bidirectional
rlabel metal5 s 1056 14936 22036 15256 6 vccd1
port 5 nsew power bidirectional
rlabel metal5 s 1056 20104 22036 20424 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 4214 2128 4534 22896 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 9435 2128 9755 22896 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 14656 2128 14976 22896 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 19877 2128 20197 22896 6 vssd1
port 6 nsew ground bidirectional
rlabel metal5 s 1056 5260 22036 5580 6 vssd1
port 6 nsew ground bidirectional
rlabel metal5 s 1056 10428 22036 10748 6 vssd1
port 6 nsew ground bidirectional
rlabel metal5 s 1056 15596 22036 15916 6 vssd1
port 6 nsew ground bidirectional
rlabel metal5 s 1056 20764 22036 21084 6 vssd1
port 6 nsew ground bidirectional
rlabel metal2 s 17406 24475 17462 25275 6 wbs_adr_o[0]
port 7 nsew signal output
rlabel metal2 s 12254 24475 12310 25275 6 wbs_adr_o[10]
port 8 nsew signal output
rlabel metal2 s 9034 24475 9090 25275 6 wbs_adr_o[11]
port 9 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 wbs_adr_o[12]
port 10 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 wbs_adr_o[13]
port 11 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 wbs_adr_o[14]
port 12 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 wbs_adr_o[15]
port 13 nsew signal output
rlabel metal2 s 19338 24475 19394 25275 6 wbs_adr_o[16]
port 14 nsew signal output
rlabel metal3 s 22331 19048 23131 19168 6 wbs_adr_o[17]
port 15 nsew signal output
rlabel metal3 s 22331 20408 23131 20528 6 wbs_adr_o[18]
port 16 nsew signal output
rlabel metal3 s 22331 21088 23131 21208 6 wbs_adr_o[19]
port 17 nsew signal output
rlabel metal3 s 22331 16328 23131 16448 6 wbs_adr_o[1]
port 18 nsew signal output
rlabel metal2 s 18050 24475 18106 25275 6 wbs_adr_o[20]
port 19 nsew signal output
rlabel metal3 s 22331 19728 23131 19848 6 wbs_adr_o[21]
port 20 nsew signal output
rlabel metal3 s 22331 18368 23131 18488 6 wbs_adr_o[22]
port 21 nsew signal output
rlabel metal3 s 22331 17008 23131 17128 6 wbs_adr_o[23]
port 22 nsew signal output
rlabel metal2 s 16118 24475 16174 25275 6 wbs_adr_o[24]
port 23 nsew signal output
rlabel metal3 s 22331 17688 23131 17808 6 wbs_adr_o[25]
port 24 nsew signal output
rlabel metal2 s 12898 24475 12954 25275 6 wbs_adr_o[26]
port 25 nsew signal output
rlabel metal2 s 10966 24475 11022 25275 6 wbs_adr_o[27]
port 26 nsew signal output
rlabel metal2 s 5814 24475 5870 25275 6 wbs_adr_o[28]
port 27 nsew signal output
rlabel metal2 s 5170 24475 5226 25275 6 wbs_adr_o[29]
port 28 nsew signal output
rlabel metal2 s 14830 24475 14886 25275 6 wbs_adr_o[2]
port 29 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 wbs_adr_o[30]
port 30 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 wbs_adr_o[31]
port 31 nsew signal output
rlabel metal2 s 9678 24475 9734 25275 6 wbs_adr_o[3]
port 32 nsew signal output
rlabel metal2 s 7102 24475 7158 25275 6 wbs_adr_o[4]
port 33 nsew signal output
rlabel metal2 s 7746 24475 7802 25275 6 wbs_adr_o[5]
port 34 nsew signal output
rlabel metal2 s 11610 24475 11666 25275 6 wbs_adr_o[6]
port 35 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 wbs_adr_o[7]
port 36 nsew signal output
rlabel metal2 s 14186 24475 14242 25275 6 wbs_adr_o[8]
port 37 nsew signal output
rlabel metal2 s 13542 24475 13598 25275 6 wbs_adr_o[9]
port 38 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 wbs_cyc_o
port 39 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[0]
port 40 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_dat_i[10]
port 41 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[11]
port 42 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 wbs_dat_i[12]
port 43 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wbs_dat_i[13]
port 44 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wbs_dat_i[14]
port 45 nsew signal input
rlabel metal3 s 0 688 800 808 6 wbs_dat_i[15]
port 46 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 wbs_dat_i[16]
port 47 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_i[17]
port 48 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[18]
port 49 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[19]
port 50 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 wbs_dat_i[1]
port 51 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 wbs_dat_i[20]
port 52 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_dat_i[21]
port 53 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 wbs_dat_i[22]
port 54 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 wbs_dat_i[23]
port 55 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 wbs_dat_i[24]
port 56 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[25]
port 57 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[26]
port 58 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[27]
port 59 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_i[28]
port 60 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wbs_dat_i[29]
port 61 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[2]
port 62 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wbs_dat_i[30]
port 63 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wbs_dat_i[31]
port 64 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[3]
port 65 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wbs_dat_i[4]
port 66 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_dat_i[5]
port 67 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wbs_dat_i[6]
port 68 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 wbs_dat_i[7]
port 69 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wbs_dat_i[8]
port 70 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[9]
port 71 nsew signal input
rlabel metal3 s 22331 4088 23131 4208 6 wbs_dat_o[0]
port 72 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[10]
port 73 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[11]
port 74 nsew signal output
rlabel metal3 s 22331 10888 23131 11008 6 wbs_dat_o[12]
port 75 nsew signal output
rlabel metal3 s 22331 10208 23131 10328 6 wbs_dat_o[13]
port 76 nsew signal output
rlabel metal3 s 22331 11568 23131 11688 6 wbs_dat_o[14]
port 77 nsew signal output
rlabel metal3 s 22331 9528 23131 9648 6 wbs_dat_o[15]
port 78 nsew signal output
rlabel metal3 s 22331 12928 23131 13048 6 wbs_dat_o[16]
port 79 nsew signal output
rlabel metal3 s 22331 12248 23131 12368 6 wbs_dat_o[17]
port 80 nsew signal output
rlabel metal3 s 22331 13608 23131 13728 6 wbs_dat_o[18]
port 81 nsew signal output
rlabel metal3 s 22331 14288 23131 14408 6 wbs_dat_o[19]
port 82 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[1]
port 83 nsew signal output
rlabel metal3 s 22331 15648 23131 15768 6 wbs_dat_o[20]
port 84 nsew signal output
rlabel metal3 s 22331 14968 23131 15088 6 wbs_dat_o[21]
port 85 nsew signal output
rlabel metal3 s 22331 6808 23131 6928 6 wbs_dat_o[22]
port 86 nsew signal output
rlabel metal3 s 22331 8168 23131 8288 6 wbs_dat_o[23]
port 87 nsew signal output
rlabel metal3 s 22331 7488 23131 7608 6 wbs_dat_o[24]
port 88 nsew signal output
rlabel metal3 s 22331 5448 23131 5568 6 wbs_dat_o[25]
port 89 nsew signal output
rlabel metal3 s 22331 3408 23131 3528 6 wbs_dat_o[26]
port 90 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[27]
port 91 nsew signal output
rlabel metal3 s 22331 8848 23131 8968 6 wbs_dat_o[28]
port 92 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[29]
port 93 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[2]
port 94 nsew signal output
rlabel metal3 s 22331 4768 23131 4888 6 wbs_dat_o[30]
port 95 nsew signal output
rlabel metal3 s 22331 6128 23131 6248 6 wbs_dat_o[31]
port 96 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[3]
port 97 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[4]
port 98 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[5]
port 99 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[6]
port 100 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[7]
port 101 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_o[8]
port 102 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[9]
port 103 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 wbs_stb_o
port 104 nsew signal output
rlabel metal3 s 22331 21768 23131 21888 6 wbs_we_o
port 105 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 23131 25275
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1926560
string GDS_FILE /openlane/designs/spi_to_wbs/runs/RUN_2025.11.02_06.05.16/results/signoff/spi_to_wbs.magic.gds
string GDS_START 326696
<< end >>

