##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 01:26:46 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_DSP
  CLASS BLOCK ;
  SIZE 210.2200 BY 30.2600 ;
  FOREIGN S_term_DSP 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.692 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 29.5400 14.2200 30.2600 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 29.5400 12.8400 30.2600 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4654 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 29.5400 11.4600 30.2600 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.484 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 29.5400 10.5400 30.2600 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.466 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 29.5400 25.2600 30.2600 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.566 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 29.5400 23.8800 30.2600 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 29.5400 22.5000 30.2600 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.519 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.9784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.296 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 29.5400 21.1200 30.2600 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.9318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.44 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 29.5400 19.7400 30.2600 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.3556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.504 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 29.5400 18.3600 30.2600 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2972 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.304 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 29.5400 16.9800 30.2600 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 29.5400 15.6000 30.2600 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 29.5400 35.8400 30.2600 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.39 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 29.5400 34.4600 30.2600 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.3472 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 46.6585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 29.5400 33.5400 30.2600 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.2872 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 66.3215 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 29.5400 32.1600 30.2600 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8768 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.102 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 29.5400 30.7800 30.2600 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.1164 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.5045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.286 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 29.5400 29.4000 30.2600 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.226 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 29.5400 28.0200 30.2600 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 29.5400 26.6400 30.2600 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.6116 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.9805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 29.5400 57.4600 30.2600 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.19 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 29.5400 56.5400 30.2600 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.584 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.8425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.476 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 29.5400 55.1600 30.2600 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.286 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 29.5400 53.7800 30.2600 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.02 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 29.5400 52.4000 30.2600 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5094 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 29.5400 51.0200 30.2600 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.1437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 29.5400 49.6400 30.2600 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.071 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.862 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.2325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.038 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 29.5400 48.2600 30.2600 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.274 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 29.5400 46.8800 30.2600 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.6216 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.0305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 29.5400 45.5000 30.2600 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.507 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 29.5400 44.1200 30.2600 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.723 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 29.5400 42.7400 30.2600 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.312 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 29.5400 41.3600 30.2600 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.9872 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 64.8585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.74 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.582 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 29.5400 39.9800 30.2600 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.572 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 29.5400 38.6000 30.2600 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.714 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.818 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 29.5400 37.2200 30.2600 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.44755 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.703 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.377 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.048 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 29.5400 79.5400 30.2600 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18875 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.575 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3677 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 29.5400 78.1600 30.2600 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.63495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.747 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.9456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 29.5400 76.7800 30.2600 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.548 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 29.5400 75.4000 30.2600 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 29.5400 74.0200 30.2600 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.277 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 29.5400 72.6400 30.2600 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 29.5400 71.2600 30.2600 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.024 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 29.5400 69.8800 30.2600 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.592 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 29.5400 68.5000 30.2600 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 29.5400 67.1200 30.2600 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.616 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 29.5400 65.7400 30.2600 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.048 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 29.5400 64.3600 30.2600 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 29.5400 62.9800 30.2600 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 29.5400 61.6000 30.2600 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9844 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.686 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 29.5400 60.2200 30.2600 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.228 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 29.5400 58.8400 30.2600 ;
    END
  END NN4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.342 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8362 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.7327 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 29.5400 84.6000 30.2600 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 33.3393 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.833 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 29.5400 83.2200 30.2600 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.6865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.5692 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 29.5400 81.8400 30.2600 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.978 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.16572 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.0629 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 29.5400 80.4600 30.2600 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.762 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.0035 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.9937 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 29.5400 106.2200 30.2600 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7469 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.2862 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 29.5400 104.8400 30.2600 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.316 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.173 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 29.5400 103.4600 30.2600 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.9088 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 29.5400 102.5400 30.2600 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.064 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2055 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.572 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.0412 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 95.0157 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 29.5400 101.1600 30.2600 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5469 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.2862 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 29.5400 99.7800 30.2600 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.75 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.326 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1506 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.0786 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 29.5400 98.4000 30.2600 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6815 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2198 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.9088 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 29.5400 97.0200 30.2600 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.4097 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.1855 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 29.5400 95.6400 30.2600 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6877 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.9906 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 29.5400 94.2600 30.2600 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.094 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.1947 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.9497 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 29.5400 92.8800 30.2600 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.8774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 29.5400 91.5000 30.2600 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.42762 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 23.4038 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 130.145 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 29.5400 90.1200 30.2600 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.02987 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.2862 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 29.5400 88.7400 30.2600 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.95 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7481 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.2924 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 29.5400 87.3600 30.2600 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.0739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.437 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 29.5400 85.9800 30.2600 ;
    END
  END S2END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2328 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.9506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 66.4884 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 351.453 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 29.5400 149.4600 30.2600 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.80835 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.951 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.1845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.50283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.4906 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 29.5400 148.5400 30.2600 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75055 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.883 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4903 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.978 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 29.5400 147.1600 30.2600 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.10786 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.5157 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 29.5400 145.7800 30.2600 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.74 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.582 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0349 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.7264 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 29.5400 144.4000 30.2600 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.8444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 98.4494 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 527.34 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 29.5400 143.0200 30.2600 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.549 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 76.872 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.541 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 29.5400 141.6400 30.2600 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8335 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.49403 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.022 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 29.5400 140.2600 30.2600 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 46.5368 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 228.236 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 29.5400 138.8800 30.2600 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.798 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.0311 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.965 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 29.5400 137.5000 30.2600 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.63495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.747 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.46761 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.8899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 29.5400 136.1200 30.2600 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 41.4481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 224.462 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 29.5400 134.7400 30.2600 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.3628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 49.1752 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 255.296 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 29.5400 133.3600 30.2600 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7406 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.2547 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 29.5400 131.9800 30.2600 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6953 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.0283 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 29.5400 130.6000 30.2600 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.67138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.9088 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 29.5400 129.2200 30.2600 ;
    END
  END SS4END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.12075 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 92.8355 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 490.761 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 29.5400 127.8400 30.2600 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7259 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1974 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 56.1569 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 301.371 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 29.5400 126.4600 30.2600 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.844 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.3959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 29.5400 125.5400 30.2600 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.032 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.58333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.4686 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 29.5400 124.1600 30.2600 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.7318 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 116.984 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 29.5400 122.7800 30.2600 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.19214 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.5126 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 29.5400 121.4000 30.2600 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.7959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 29.5400 120.0200 30.2600 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.52275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.615 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.342 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8362 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.7327 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 29.5400 118.6400 30.2600 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.4022 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.5629 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 29.5400 117.2600 30.2600 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2572 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1715 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9393 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.2233 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 29.5400 115.8800 30.2600 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5488 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.952 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.9843 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 29.5400 114.5000 30.2600 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.284 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.8777 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.2547 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 29.5400 113.1200 30.2600 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.224 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.5116 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 113.11 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 29.5400 111.7400 30.2600 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.2365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5116 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.7296 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 29.5400 110.3600 30.2600 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1964 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8675 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.224 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.1858 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 111.481 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 29.5400 108.9800 30.2600 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.62484 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.261 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 29.5400 107.6000 30.2600 ;
    END
  END S4END[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8126 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.956 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.8212 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 74.0285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.486 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.9214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0498 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.588 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.5442 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.684 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 60.8525 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 300.811 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.49 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.43 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.284 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.8491 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.6164 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.9675 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 37.2079 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.73 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.633 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.0875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0653 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.8008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 92.1915 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 480.849 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 56.467 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 296.189 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1998 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.588 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 18.3156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.5005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7217 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.7453 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.622 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 28.706 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 148.585 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.1848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.177 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 19.4657 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 104.267 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.9848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.658 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.1352 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.708 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 79.8009 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 393.814 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.4188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 54.7726 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.415 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6562 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.772 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.7372 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.6085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 55.345 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 284.824 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.2556 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.2005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.844 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 64.8135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 314.714 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.262 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.7204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.9969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9336 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.5905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 33.9267 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 162.16 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.335 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 55.4129 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 296.421 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.105 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 29.2645 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.509 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 43.5198 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.289 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.734 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7406 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.5755 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1946 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.629 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 28.6915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.588 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8995 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 40.6506 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 193.616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4244 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 75.9186 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.918 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.448 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.1242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.4937 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 29.1877 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 148.302 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 16.9978 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 90.9277 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.627 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 35.9475 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 183.113 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.0332 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 81.1035 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 439.862 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.685 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 26.467 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 141.358 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 93.9487 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 487.195 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.9575 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.9182 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.9848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 74.1418 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 384.296 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 28.6600 210.2200 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.499 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.4108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.328 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 26.6200 210.2200 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.99 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 24.9200 210.2200 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6962 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.255 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 22.8800 210.2200 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.682 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.496 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 21.1800 210.2200 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 19.1400 210.2200 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.465 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 17.4400 210.2200 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.641 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 15.7400 210.2200 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.0118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 13.7000 210.2200 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3305 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 12.0000 210.2200 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4115 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 10.3000 210.2200 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.228 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 8.2600 210.2200 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.257 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 6.5600 210.2200 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.326 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 4.5200 210.2200 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4904 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.36 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 2.8200 210.2200 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.168 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 1.1200 210.2200 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.34 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.6084 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.9645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 27.6250 210.2200 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.081 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.2488 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.1665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.504 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 25.9250 210.2200 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.6896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.3705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 24.2250 210.2200 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.76925 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.905 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 18.0748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 90.2965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.724 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 22.5250 210.2200 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.1876 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.8605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.2518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 20.8250 210.2200 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.545 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 19.1250 210.2200 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2172 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.432 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.264 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 17.4250 210.2200 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.6392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.122 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 15.7250 210.2200 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.098 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3755 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.062 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 14.0250 210.2200 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.4488 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.692 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 12.3250 210.2200 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1046 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.476 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.1064 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.3435 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9708 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.264 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 10.6250 210.2200 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 11.9732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 59.829 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 8.9250 210.2200 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.838 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2484 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.736 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 7.2250 210.2200 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8397 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 5.5250 210.2200 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.2384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 76.1145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 3.8250 210.2200 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.3744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.18 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 209.8900 2.1250 210.2200 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0602 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.119 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.489 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.9969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 149.5400 0.0000 149.9200 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.503 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.37 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.1079 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.676 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 144.0200 0.0000 144.4000 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0898 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.01 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.4214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 138.9600 0.0000 139.3400 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2186 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.948 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.9214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 133.4400 0.0000 133.8200 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1166 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.438 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.1544 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.2987 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 128.3800 0.0000 128.7600 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0674 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.155 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.168 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.4676 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.5723 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 123.3200 0.0000 123.7000 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.75 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7116 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.0849 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 117.8000 0.0000 118.1800 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.709 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.437 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.833 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.811 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.7381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 112.7400 0.0000 113.1200 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.485 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.317 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 33.2223 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 158.638 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 107.6800 0.0000 108.0600 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6138 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.961 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.2802 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.1478 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 102.1600 0.0000 102.5400 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5494 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.942 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.777 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.9528 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 97.1000 0.0000 97.4800 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0522 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.116 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.0211 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.2421 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 91.5800 0.0000 91.9600 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4206 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.995 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.082 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.8425 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.764 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 86.5200 0.0000 86.9000 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6138 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.961 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5022 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.151 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 81.4600 0.0000 81.8400 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.964 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.88145 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.9591 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 75.9400 0.0000 76.3200 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.709 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.437 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6814 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.544 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 70.8800 0.0000 71.2600 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6824 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.304 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 83.194 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.384 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 65.8200 0.0000 66.2000 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.571 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.71 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.6311 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 95.6824 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 60.3000 0.0000 60.6800 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.817 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.866 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.048 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3506 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.7453 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 55.2400 0.0000 55.6200 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5494 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.668 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.4462 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 102.626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 50.1800 0.0000 50.5600 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.237 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 199.6800 29.5400 200.0600 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.203 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 196.9200 29.5400 197.3000 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.6200 29.5400 195.0000 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.7158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.288 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 192.3200 29.5400 192.7000 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 190.0200 29.5400 190.4000 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.965 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 187.7200 29.5400 188.1000 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.663 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 185.4200 29.5400 185.8000 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.1200 29.5400 183.5000 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.011 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.8200 29.5400 181.2000 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.6342 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 178.5200 29.5400 178.9000 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.509 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 175.7600 29.5400 176.1400 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.473 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 173.4600 29.5400 173.8400 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.245 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 171.1600 29.5400 171.5400 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.617 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 168.8600 29.5400 169.2400 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.311 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.9424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.104 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 166.5600 29.5400 166.9400 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.8328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.912 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 164.2600 29.5400 164.6400 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.869 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.9600 29.5400 162.3400 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.2628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.872 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 159.6600 29.5400 160.0400 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.122 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.3600 29.5400 157.7400 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.58 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.0600 29.5400 155.4400 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 204.6600 6.0700 ;
        RECT 5.5600 23.0000 204.6600 25.0000 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 202.6600 15.0600 204.6600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 202.6600 9.6200 204.6600 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 202.6600 20.5000 204.6600 20.9800 ;
      LAYER met4 ;
        RECT 202.6600 4.0700 204.6600 25.0000 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 207.6600 3.0700 ;
        RECT 2.5600 26.0000 207.6600 28.0000 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 205.6600 6.9000 207.6600 7.3800 ;
        RECT 205.6600 12.3400 207.6600 12.8200 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 205.6600 17.7800 207.6600 18.2600 ;
      LAYER met4 ;
        RECT 205.6600 1.0700 207.6600 28.0000 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.6300 29.3700 210.2200 30.2600 ;
      RECT 148.7100 29.3700 148.9100 30.2600 ;
      RECT 147.3300 29.3700 147.9900 30.2600 ;
      RECT 145.9500 29.3700 146.6100 30.2600 ;
      RECT 144.5700 29.3700 145.2300 30.2600 ;
      RECT 143.1900 29.3700 143.8500 30.2600 ;
      RECT 141.8100 29.3700 142.4700 30.2600 ;
      RECT 140.4300 29.3700 141.0900 30.2600 ;
      RECT 139.0500 29.3700 139.7100 30.2600 ;
      RECT 137.6700 29.3700 138.3300 30.2600 ;
      RECT 136.2900 29.3700 136.9500 30.2600 ;
      RECT 134.9100 29.3700 135.5700 30.2600 ;
      RECT 133.5300 29.3700 134.1900 30.2600 ;
      RECT 132.1500 29.3700 132.8100 30.2600 ;
      RECT 130.7700 29.3700 131.4300 30.2600 ;
      RECT 129.3900 29.3700 130.0500 30.2600 ;
      RECT 128.0100 29.3700 128.6700 30.2600 ;
      RECT 126.6300 29.3700 127.2900 30.2600 ;
      RECT 125.7100 29.3700 125.9100 30.2600 ;
      RECT 124.3300 29.3700 124.9900 30.2600 ;
      RECT 122.9500 29.3700 123.6100 30.2600 ;
      RECT 121.5700 29.3700 122.2300 30.2600 ;
      RECT 120.1900 29.3700 120.8500 30.2600 ;
      RECT 118.8100 29.3700 119.4700 30.2600 ;
      RECT 117.4300 29.3700 118.0900 30.2600 ;
      RECT 116.0500 29.3700 116.7100 30.2600 ;
      RECT 114.6700 29.3700 115.3300 30.2600 ;
      RECT 113.2900 29.3700 113.9500 30.2600 ;
      RECT 111.9100 29.3700 112.5700 30.2600 ;
      RECT 110.5300 29.3700 111.1900 30.2600 ;
      RECT 109.1500 29.3700 109.8100 30.2600 ;
      RECT 107.7700 29.3700 108.4300 30.2600 ;
      RECT 106.3900 29.3700 107.0500 30.2600 ;
      RECT 105.0100 29.3700 105.6700 30.2600 ;
      RECT 103.6300 29.3700 104.2900 30.2600 ;
      RECT 102.7100 29.3700 102.9100 30.2600 ;
      RECT 101.3300 29.3700 101.9900 30.2600 ;
      RECT 99.9500 29.3700 100.6100 30.2600 ;
      RECT 98.5700 29.3700 99.2300 30.2600 ;
      RECT 97.1900 29.3700 97.8500 30.2600 ;
      RECT 95.8100 29.3700 96.4700 30.2600 ;
      RECT 94.4300 29.3700 95.0900 30.2600 ;
      RECT 93.0500 29.3700 93.7100 30.2600 ;
      RECT 91.6700 29.3700 92.3300 30.2600 ;
      RECT 90.2900 29.3700 90.9500 30.2600 ;
      RECT 88.9100 29.3700 89.5700 30.2600 ;
      RECT 87.5300 29.3700 88.1900 30.2600 ;
      RECT 86.1500 29.3700 86.8100 30.2600 ;
      RECT 84.7700 29.3700 85.4300 30.2600 ;
      RECT 83.3900 29.3700 84.0500 30.2600 ;
      RECT 82.0100 29.3700 82.6700 30.2600 ;
      RECT 80.6300 29.3700 81.2900 30.2600 ;
      RECT 79.7100 29.3700 79.9100 30.2600 ;
      RECT 78.3300 29.3700 78.9900 30.2600 ;
      RECT 76.9500 29.3700 77.6100 30.2600 ;
      RECT 75.5700 29.3700 76.2300 30.2600 ;
      RECT 74.1900 29.3700 74.8500 30.2600 ;
      RECT 72.8100 29.3700 73.4700 30.2600 ;
      RECT 71.4300 29.3700 72.0900 30.2600 ;
      RECT 70.0500 29.3700 70.7100 30.2600 ;
      RECT 68.6700 29.3700 69.3300 30.2600 ;
      RECT 67.2900 29.3700 67.9500 30.2600 ;
      RECT 65.9100 29.3700 66.5700 30.2600 ;
      RECT 64.5300 29.3700 65.1900 30.2600 ;
      RECT 63.1500 29.3700 63.8100 30.2600 ;
      RECT 61.7700 29.3700 62.4300 30.2600 ;
      RECT 60.3900 29.3700 61.0500 30.2600 ;
      RECT 59.0100 29.3700 59.6700 30.2600 ;
      RECT 57.6300 29.3700 58.2900 30.2600 ;
      RECT 56.7100 29.3700 56.9100 30.2600 ;
      RECT 55.3300 29.3700 55.9900 30.2600 ;
      RECT 53.9500 29.3700 54.6100 30.2600 ;
      RECT 52.5700 29.3700 53.2300 30.2600 ;
      RECT 51.1900 29.3700 51.8500 30.2600 ;
      RECT 49.8100 29.3700 50.4700 30.2600 ;
      RECT 48.4300 29.3700 49.0900 30.2600 ;
      RECT 47.0500 29.3700 47.7100 30.2600 ;
      RECT 45.6700 29.3700 46.3300 30.2600 ;
      RECT 44.2900 29.3700 44.9500 30.2600 ;
      RECT 42.9100 29.3700 43.5700 30.2600 ;
      RECT 41.5300 29.3700 42.1900 30.2600 ;
      RECT 40.1500 29.3700 40.8100 30.2600 ;
      RECT 38.7700 29.3700 39.4300 30.2600 ;
      RECT 37.3900 29.3700 38.0500 30.2600 ;
      RECT 36.0100 29.3700 36.6700 30.2600 ;
      RECT 34.6300 29.3700 35.2900 30.2600 ;
      RECT 33.7100 29.3700 33.9100 30.2600 ;
      RECT 32.3300 29.3700 32.9900 30.2600 ;
      RECT 30.9500 29.3700 31.6100 30.2600 ;
      RECT 29.5700 29.3700 30.2300 30.2600 ;
      RECT 28.1900 29.3700 28.8500 30.2600 ;
      RECT 26.8100 29.3700 27.4700 30.2600 ;
      RECT 25.4300 29.3700 26.0900 30.2600 ;
      RECT 24.0500 29.3700 24.7100 30.2600 ;
      RECT 22.6700 29.3700 23.3300 30.2600 ;
      RECT 21.2900 29.3700 21.9500 30.2600 ;
      RECT 19.9100 29.3700 20.5700 30.2600 ;
      RECT 18.5300 29.3700 19.1900 30.2600 ;
      RECT 17.1500 29.3700 17.8100 30.2600 ;
      RECT 15.7700 29.3700 16.4300 30.2600 ;
      RECT 14.3900 29.3700 15.0500 30.2600 ;
      RECT 13.0100 29.3700 13.6700 30.2600 ;
      RECT 11.6300 29.3700 12.2900 30.2600 ;
      RECT 10.7100 29.3700 10.9100 30.2600 ;
      RECT 0.0000 29.3700 9.9900 30.2600 ;
      RECT 0.0000 28.9850 210.2200 29.3700 ;
      RECT 0.5000 28.4750 210.2200 28.9850 ;
      RECT 0.0000 27.9650 210.2200 28.4750 ;
      RECT 0.0000 27.4550 209.7200 27.9650 ;
      RECT 0.0000 26.9450 210.2200 27.4550 ;
      RECT 0.5000 26.4350 210.2200 26.9450 ;
      RECT 0.0000 26.2650 210.2200 26.4350 ;
      RECT 0.0000 25.7550 209.7200 26.2650 ;
      RECT 0.0000 25.2450 210.2200 25.7550 ;
      RECT 0.5000 24.7350 210.2200 25.2450 ;
      RECT 0.0000 24.5650 210.2200 24.7350 ;
      RECT 0.0000 24.0550 209.7200 24.5650 ;
      RECT 0.0000 23.2050 210.2200 24.0550 ;
      RECT 0.5000 22.8650 210.2200 23.2050 ;
      RECT 0.5000 22.6950 209.7200 22.8650 ;
      RECT 0.0000 22.3550 209.7200 22.6950 ;
      RECT 0.0000 21.5050 210.2200 22.3550 ;
      RECT 0.5000 21.1650 210.2200 21.5050 ;
      RECT 0.5000 20.9950 209.7200 21.1650 ;
      RECT 0.0000 20.6550 209.7200 20.9950 ;
      RECT 0.0000 19.4650 210.2200 20.6550 ;
      RECT 0.5000 18.9550 209.7200 19.4650 ;
      RECT 0.0000 17.7650 210.2200 18.9550 ;
      RECT 0.5000 17.2550 209.7200 17.7650 ;
      RECT 0.0000 16.0650 210.2200 17.2550 ;
      RECT 0.5000 15.5550 209.7200 16.0650 ;
      RECT 0.0000 14.3650 210.2200 15.5550 ;
      RECT 0.0000 14.0250 209.7200 14.3650 ;
      RECT 0.5000 13.8550 209.7200 14.0250 ;
      RECT 0.5000 13.5150 210.2200 13.8550 ;
      RECT 0.0000 12.6650 210.2200 13.5150 ;
      RECT 0.0000 12.3250 209.7200 12.6650 ;
      RECT 0.5000 12.1550 209.7200 12.3250 ;
      RECT 0.5000 11.8150 210.2200 12.1550 ;
      RECT 0.0000 10.9650 210.2200 11.8150 ;
      RECT 0.0000 10.6250 209.7200 10.9650 ;
      RECT 0.5000 10.4550 209.7200 10.6250 ;
      RECT 0.5000 10.1150 210.2200 10.4550 ;
      RECT 0.0000 9.2650 210.2200 10.1150 ;
      RECT 0.0000 8.7550 209.7200 9.2650 ;
      RECT 0.0000 8.5850 210.2200 8.7550 ;
      RECT 0.5000 8.0750 210.2200 8.5850 ;
      RECT 0.0000 7.5650 210.2200 8.0750 ;
      RECT 0.0000 7.0550 209.7200 7.5650 ;
      RECT 0.0000 6.8850 210.2200 7.0550 ;
      RECT 0.5000 6.3750 210.2200 6.8850 ;
      RECT 0.0000 5.8650 210.2200 6.3750 ;
      RECT 0.0000 5.3550 209.7200 5.8650 ;
      RECT 0.0000 4.8450 210.2200 5.3550 ;
      RECT 0.5000 4.3350 210.2200 4.8450 ;
      RECT 0.0000 4.1650 210.2200 4.3350 ;
      RECT 0.0000 3.6550 209.7200 4.1650 ;
      RECT 0.0000 3.1450 210.2200 3.6550 ;
      RECT 0.5000 2.6350 210.2200 3.1450 ;
      RECT 0.0000 2.4650 210.2200 2.6350 ;
      RECT 0.0000 1.9550 209.7200 2.4650 ;
      RECT 0.0000 1.4450 210.2200 1.9550 ;
      RECT 0.5000 0.9350 210.2200 1.4450 ;
      RECT 0.0000 0.0000 210.2200 0.9350 ;
    LAYER met1 ;
      RECT 0.0000 0.8600 210.2200 30.2600 ;
      RECT 150.0600 0.0000 210.2200 0.8600 ;
      RECT 144.5400 0.0000 149.4000 0.8600 ;
      RECT 139.4800 0.0000 143.8800 0.8600 ;
      RECT 133.9600 0.0000 138.8200 0.8600 ;
      RECT 128.9000 0.0000 133.3000 0.8600 ;
      RECT 123.8400 0.0000 128.2400 0.8600 ;
      RECT 118.3200 0.0000 123.1800 0.8600 ;
      RECT 113.2600 0.0000 117.6600 0.8600 ;
      RECT 108.2000 0.0000 112.6000 0.8600 ;
      RECT 102.6800 0.0000 107.5400 0.8600 ;
      RECT 97.6200 0.0000 102.0200 0.8600 ;
      RECT 92.1000 0.0000 96.9600 0.8600 ;
      RECT 87.0400 0.0000 91.4400 0.8600 ;
      RECT 81.9800 0.0000 86.3800 0.8600 ;
      RECT 76.4600 0.0000 81.3200 0.8600 ;
      RECT 71.4000 0.0000 75.8000 0.8600 ;
      RECT 66.3400 0.0000 70.7400 0.8600 ;
      RECT 60.8200 0.0000 65.6800 0.8600 ;
      RECT 55.7600 0.0000 60.1600 0.8600 ;
      RECT 50.7000 0.0000 55.1000 0.8600 ;
      RECT 0.0000 0.0000 50.0400 0.8600 ;
    LAYER met2 ;
      RECT 200.2000 29.4000 210.2200 30.2600 ;
      RECT 197.4400 29.4000 199.5400 30.2600 ;
      RECT 195.1400 29.4000 196.7800 30.2600 ;
      RECT 192.8400 29.4000 194.4800 30.2600 ;
      RECT 190.5400 29.4000 192.1800 30.2600 ;
      RECT 188.2400 29.4000 189.8800 30.2600 ;
      RECT 185.9400 29.4000 187.5800 30.2600 ;
      RECT 183.6400 29.4000 185.2800 30.2600 ;
      RECT 181.3400 29.4000 182.9800 30.2600 ;
      RECT 179.0400 29.4000 180.6800 30.2600 ;
      RECT 176.2800 29.4000 178.3800 30.2600 ;
      RECT 173.9800 29.4000 175.6200 30.2600 ;
      RECT 171.6800 29.4000 173.3200 30.2600 ;
      RECT 169.3800 29.4000 171.0200 30.2600 ;
      RECT 167.0800 29.4000 168.7200 30.2600 ;
      RECT 164.7800 29.4000 166.4200 30.2600 ;
      RECT 162.4800 29.4000 164.1200 30.2600 ;
      RECT 160.1800 29.4000 161.8200 30.2600 ;
      RECT 157.8800 29.4000 159.5200 30.2600 ;
      RECT 155.5800 29.4000 157.2200 30.2600 ;
      RECT 0.0000 29.4000 154.9200 30.2600 ;
      RECT 0.0000 28.9400 210.2200 29.4000 ;
      RECT 0.0000 28.5200 209.5950 28.9400 ;
      RECT 0.0000 27.9200 210.2200 28.5200 ;
      RECT 0.6250 27.5000 210.2200 27.9200 ;
      RECT 0.0000 26.9000 210.2200 27.5000 ;
      RECT 0.0000 26.4800 209.5950 26.9000 ;
      RECT 0.0000 26.2200 210.2200 26.4800 ;
      RECT 0.6250 25.8000 210.2200 26.2200 ;
      RECT 0.0000 25.2000 210.2200 25.8000 ;
      RECT 0.0000 24.7800 209.5950 25.2000 ;
      RECT 0.0000 24.5200 210.2200 24.7800 ;
      RECT 0.6250 24.1000 210.2200 24.5200 ;
      RECT 0.0000 23.1600 210.2200 24.1000 ;
      RECT 0.0000 22.8200 209.5950 23.1600 ;
      RECT 0.6250 22.7400 209.5950 22.8200 ;
      RECT 0.6250 22.4000 210.2200 22.7400 ;
      RECT 0.0000 21.4600 210.2200 22.4000 ;
      RECT 0.0000 21.1200 209.5950 21.4600 ;
      RECT 0.6250 21.0400 209.5950 21.1200 ;
      RECT 0.6250 20.7000 210.2200 21.0400 ;
      RECT 0.0000 19.4200 210.2200 20.7000 ;
      RECT 0.6250 19.0000 209.5950 19.4200 ;
      RECT 0.0000 17.7200 210.2200 19.0000 ;
      RECT 0.6250 17.3000 209.5950 17.7200 ;
      RECT 0.0000 16.0200 210.2200 17.3000 ;
      RECT 0.6250 15.6000 209.5950 16.0200 ;
      RECT 0.0000 14.3200 210.2200 15.6000 ;
      RECT 0.6250 13.9800 210.2200 14.3200 ;
      RECT 0.6250 13.9000 209.5950 13.9800 ;
      RECT 0.0000 13.5600 209.5950 13.9000 ;
      RECT 0.0000 12.6200 210.2200 13.5600 ;
      RECT 0.6250 12.2800 210.2200 12.6200 ;
      RECT 0.6250 12.2000 209.5950 12.2800 ;
      RECT 0.0000 11.8600 209.5950 12.2000 ;
      RECT 0.0000 10.9200 210.2200 11.8600 ;
      RECT 0.6250 10.5800 210.2200 10.9200 ;
      RECT 0.6250 10.5000 209.5950 10.5800 ;
      RECT 0.0000 10.1600 209.5950 10.5000 ;
      RECT 0.0000 9.2200 210.2200 10.1600 ;
      RECT 0.6250 8.8000 210.2200 9.2200 ;
      RECT 0.0000 8.5400 210.2200 8.8000 ;
      RECT 0.0000 8.1200 209.5950 8.5400 ;
      RECT 0.0000 7.5200 210.2200 8.1200 ;
      RECT 0.6250 7.1000 210.2200 7.5200 ;
      RECT 0.0000 6.8400 210.2200 7.1000 ;
      RECT 0.0000 6.4200 209.5950 6.8400 ;
      RECT 0.0000 5.8200 210.2200 6.4200 ;
      RECT 0.6250 5.4000 210.2200 5.8200 ;
      RECT 0.0000 4.8000 210.2200 5.4000 ;
      RECT 0.0000 4.3800 209.5950 4.8000 ;
      RECT 0.0000 4.1200 210.2200 4.3800 ;
      RECT 0.6250 3.7000 210.2200 4.1200 ;
      RECT 0.0000 3.1000 210.2200 3.7000 ;
      RECT 0.0000 2.6800 209.5950 3.1000 ;
      RECT 0.0000 2.4200 210.2200 2.6800 ;
      RECT 0.6250 2.0000 210.2200 2.4200 ;
      RECT 0.0000 1.4000 210.2200 2.0000 ;
      RECT 0.0000 0.9800 209.5950 1.4000 ;
      RECT 0.0000 0.0000 210.2200 0.9800 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 210.2200 30.2600 ;
      RECT 207.9600 25.7000 210.2200 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 210.2200 25.7000 ;
      RECT 204.9600 22.7000 210.2200 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 210.2200 22.7000 ;
      RECT 204.9600 20.2000 210.2200 21.2800 ;
      RECT 7.8600 20.2000 202.3600 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 210.2200 20.2000 ;
      RECT 207.9600 17.4800 210.2200 18.5600 ;
      RECT 4.8600 17.4800 205.3600 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 210.2200 17.4800 ;
      RECT 204.9600 14.7600 210.2200 15.8400 ;
      RECT 7.8600 14.7600 202.3600 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 210.2200 14.7600 ;
      RECT 207.9600 12.0400 210.2200 13.1200 ;
      RECT 4.8600 12.0400 205.3600 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 210.2200 12.0400 ;
      RECT 204.9600 9.3200 210.2200 10.4000 ;
      RECT 7.8600 9.3200 202.3600 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 210.2200 9.3200 ;
      RECT 207.9600 6.6000 210.2200 7.6800 ;
      RECT 4.8600 6.6000 205.3600 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 210.2200 6.6000 ;
      RECT 204.9600 3.7700 210.2200 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 210.2200 3.7700 ;
      RECT 207.9600 0.7700 210.2200 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 210.2200 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 210.2200 30.2600 ;
      RECT 4.8600 25.3000 205.3600 28.3000 ;
      RECT 204.9600 3.7700 205.3600 25.3000 ;
      RECT 7.8600 3.7700 202.3600 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 207.9600 0.7700 210.2200 28.3000 ;
      RECT 4.8600 0.7700 205.3600 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 210.2200 0.7700 ;
  END
END S_term_DSP

END LIBRARY
