##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 00:21:33 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO W_IO
  CLASS BLOCK ;
  SIZE 69.9200 BY 219.6400 ;
  FOREIGN W_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 0.7368 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.647 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 84.6400 69.9200 85.0200 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2742 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2665 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 83.2800 69.9200 83.6600 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.409 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.937 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.4098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.656 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 81.5800 69.9200 81.9600 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.784 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 80.2200 69.9200 80.6000 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.152 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 96.5400 69.9200 96.9200 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.6 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 94.8400 69.9200 95.2200 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0702 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.243 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 93.4800 69.9200 93.8600 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.311 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.447 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8119 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.8 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 92.1200 69.9200 92.5000 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.6604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.184 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 90.4200 69.9200 90.8000 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5994 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.889 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.4318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.44 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 89.0600 69.9200 89.4400 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6775 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 87.7000 69.9200 88.0800 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5146 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.698 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 86.0000 69.9200 86.3800 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3754 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.769 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.286 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 108.4400 69.9200 108.8200 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.481 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.5608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.128 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 107.7600 69.9200 108.1400 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.4874 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3325 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 105.3800 69.9200 105.7600 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.992 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 103.3400 69.9200 103.7200 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.3428 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6095 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 102.3200 69.9200 102.7000 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8294 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.039 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.0568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.44 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 101.3000 69.9200 101.6800 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6022 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.903 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.1845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.352 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 100.6200 69.9200 101.0000 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.5095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 97.9000 69.9200 98.2800 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.5466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5915 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 131.9000 69.9200 132.2800 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5994 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.889 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 129.8600 69.9200 130.2400 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5686 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.56 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 128.8400 69.9200 129.2200 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.418 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.88 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 127.4800 69.9200 127.8600 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.5586 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.756 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 125.7800 69.9200 126.1600 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.4688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.304 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 124.4200 69.9200 124.8000 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8938 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.968 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 123.0600 69.9200 123.4400 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8126 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.955 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 121.3600 69.9200 121.7400 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1514 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.649 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8988 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.376 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 120.0000 69.9200 120.3800 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0366 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.08 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 118.6400 69.9200 119.0200 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7881 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.0568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.166 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 116.9400 69.9200 117.3200 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.726 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 115.5800 69.9200 115.9600 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.311 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.447 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.7408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.088 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 114.2200 69.9200 114.6000 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1822 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.803 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 112.5200 69.9200 112.9000 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.794 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8655 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 111.1600 69.9200 111.5400 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0534 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.3498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.336 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 109.8000 69.9200 110.1800 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.481 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.568 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 149.5800 69.9200 149.9600 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.311 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.447 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.6 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 147.8800 69.9200 148.2600 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.358 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 146.5200 69.9200 146.9000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.633 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.057 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.3528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.352 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 145.1600 69.9200 145.5400 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.4538 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1645 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 143.4600 69.9200 143.8400 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9378 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.581 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.416 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 142.1000 69.9200 142.4800 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.25 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 140.7400 69.9200 141.1200 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.087 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.327 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.9408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.488 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 139.0400 69.9200 139.4200 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0842 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.419 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 137.3400 69.9200 137.7200 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6974 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.379 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.7788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.624 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 136.3200 69.9200 136.7000 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8294 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.039 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 133.9400 69.9200 134.3200 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7562 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.636 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 133.2600 69.9200 133.6400 ;
    END
  END E6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0404 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.094 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.3951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.8045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.2436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 38.2834 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 202.411 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.348374 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 13.9200 69.9200 14.3000 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9654 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.719 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.4348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.712 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 88.6079 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 423.742 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 12.5600 69.9200 12.9400 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4226 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.4755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.817 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.1138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 44.879 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.874 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.267073 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 11.2000 69.9200 11.5800 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.832 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 113.327 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 547.849 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.646541 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 9.8400 69.9200 10.2200 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.423 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.007 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.3284 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.056 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 25.8200 69.9200 26.2000 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.755 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.667 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.9895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 24.4600 69.9200 24.8400 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.145 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.617 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.9725 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.456 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 22.7600 69.9200 23.1400 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.468 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.936 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.8116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.936 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 21.4000 69.9200 21.7800 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9504 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.5611 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.536 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 20.0400 69.9200 20.4200 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3074 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.429 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.1376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.99 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 18.3400 69.9200 18.7200 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2462 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.123 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.9275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4085 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.448 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 16.9800 69.9200 17.3600 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.199 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.887 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.936 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.9898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.416 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 15.6200 69.9200 16.0000 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.955 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.667 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7596 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 37.7200 69.9200 38.1000 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1786 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.2045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.0965 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.784 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 36.0200 69.9200 36.4000 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.515 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4433 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.7015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.0277 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.28 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 34.6600 69.9200 35.0400 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0154 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.969 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.9949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9327 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.44 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 33.3000 69.9200 33.6800 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.853 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.157 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9468 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.1776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.318 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 31.6000 69.9200 31.9800 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3714 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.749 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.344 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 30.2400 69.9200 30.6200 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0802 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.293 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.9575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.1417 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.888 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 28.8800 69.9200 29.2600 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9818 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.801 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7524 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.7405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.24 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 27.1800 69.9200 27.5600 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8602 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.193 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.4419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 61.5200 69.9200 61.9000 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2158 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.971 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.7628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.872 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 59.8200 69.9200 60.2000 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2402 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.093 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8654 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.36 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 58.4600 69.9200 58.8400 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.06 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.9828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.712 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 57.7800 69.9200 58.1600 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9378 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.581 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.6388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.544 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 54.7200 69.9200 55.1000 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.5472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.274 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 53.7000 69.9200 54.0800 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8566 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.175 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.4194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.648 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 52.3400 69.9200 52.7200 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.164 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.675 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.784 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 50.9800 69.9200 51.3600 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8258 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.021 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.6164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.512 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 49.2800 69.9200 49.6600 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.1256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.944 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 47.9200 69.9200 48.3000 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8598 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.191 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.0678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.832 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 46.9000 69.9200 47.2800 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5378 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.581 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.9128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.672 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 46.2200 69.9200 46.6000 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8598 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.191 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.264 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 43.5000 69.9200 43.8800 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.501 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.397 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5724 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.457 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 42.1400 69.9200 42.5200 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.9288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.424 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 40.7800 69.9200 41.1600 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3786 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.8218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.52 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 39.0800 69.9200 39.4600 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2802 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.293 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7355 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.192 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 78.8600 69.9200 79.2400 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4996 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.353 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.5593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 77.5000 69.9200 77.8800 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.885 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.8048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.096 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 75.8000 69.9200 76.1800 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5718 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.751 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.5998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.336 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 74.4400 69.9200 74.8200 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.711 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.447 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.134 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.016 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 73.0800 69.9200 73.4600 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3786 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.1649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.6535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 71.3800 69.9200 71.7600 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4806 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.7926 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.168 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 70.0200 69.9200 70.4000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0534 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.408 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 68.6600 69.9200 69.0400 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1412 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2783 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.224 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 67.6400 69.9200 68.0200 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0646 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.178 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.1105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9504 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.2948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.376 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 65.6000 69.9200 65.9800 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7114 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.449 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.451 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.0728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.192 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 64.2400 69.9200 64.6200 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.989 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.9607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.6325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.608 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.2000 62.5400 69.9200 62.9200 ;
    END
  END W6END[0]
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.706 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.3699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.6785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 100.2800 0.7200 100.6600 ;
    END
  END A_I_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1514 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.649 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.9755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 98.2400 0.7200 98.6200 ;
    END
  END A_T_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6523 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.8485 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 56.4775 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.651 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 95.8600 0.7200 96.2400 ;
    END
  END A_O_top
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.0636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 289.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 12.264 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 64.7362 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 45.5800 0.0000 45.9600 0.7200 ;
    END
  END UserCLK
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.219 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 84.3000 0.7200 84.6800 ;
    END
  END B_I_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.4083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.8705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.376 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 81.9200 0.7200 82.3000 ;
    END
  END B_T_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.515 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.4474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met3  ;
    ANTENNAMAXAREACAR 46.0353 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.455 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.602111 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 48.5965 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.876 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.602111 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 79.8800 0.7200 80.2600 ;
    END
  END B_O_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.6004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8975 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 102.6600 0.7200 103.0400 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.389 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8405 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 105.0400 0.7200 105.4200 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5182 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.483 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.2441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.0495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.1468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.92 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 107.4200 0.7200 107.8000 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.765 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.717 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.8733 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.0775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.1448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.576 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 109.8000 0.7200 110.1800 ;
    END
  END A_config_C_bit3
  PIN B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.3554 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6725 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 86.6800 0.7200 87.0600 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6638 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.211 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.336 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 89.0600 0.7200 89.4400 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.4538 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.1645 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 91.1000 0.7200 91.4800 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.572 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.094 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 93.4800 0.7200 93.8600 ;
    END
  END B_config_C_bit3
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 20.2647 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.3594 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 209.3100 0.7200 209.6900 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 11.0217 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 52.6436 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 207.4800 0.7200 207.8600 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 29.0061 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.651 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 205.6500 0.7200 206.0300 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 23.515 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 118.046 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352288 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 203.8200 0.7200 204.2000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 18.5576 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.4015 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352288 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 201.9900 0.7200 202.3700 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 9.44345 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.9234 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352288 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 200.1600 0.7200 200.5400 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.3468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 29.9392 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.289 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.381305 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 198.3300 0.7200 198.7100 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.5578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 44.0257 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 228.715 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.60386 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 196.5000 0.7200 196.8800 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.8258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 32.6288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.244 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 195.2800 0.7200 195.6600 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.0588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 43.4403 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.512 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 193.4500 0.7200 193.8300 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.8518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 51.9375 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.968 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.60386 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 191.6200 0.7200 192.0000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9996 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.6298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 36.8501 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.764 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 189.7900 0.7200 190.1700 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.6078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 38.5184 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 197.834 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 187.9600 0.7200 188.3400 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9406 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.1728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 35.3038 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 177.19 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 186.1300 0.7200 186.5100 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 24.4437 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 121.229 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 184.3000 0.7200 184.6800 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 20.8526 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.672 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 182.4700 0.7200 182.8500 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8168 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.4992 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 181.2500 0.7200 181.6300 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 21.8518 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 105.551 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 179.4200 0.7200 179.8000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 14.2673 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.1218 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 177.5900 0.7200 177.9700 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 8.42098 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 38.4039 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.356071 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 175.7600 0.7200 176.1400 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 11.0821 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.1116 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.356071 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 173.9300 0.7200 174.3100 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 8.48085 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.9435 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.356071 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 172.1000 0.7200 172.4800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.4168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 23.29 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.146 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 170.2700 0.7200 170.6500 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.8288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 42.2198 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 212.372 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.859215 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 168.4400 0.7200 168.8200 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 14.8141 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 70.233 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 167.2200 0.7200 167.6000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 28.6749 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 138.861 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 165.3900 0.7200 165.7700 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.6538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 39.3876 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.726 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 163.5600 0.7200 163.9400 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.0646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 47.4504 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 242.648 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 161.7300 0.7200 162.1100 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 22.2867 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 108.985 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 159.9000 0.7200 160.2800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.6538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 33.6488 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 172.15 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 158.0700 0.7200 158.4500 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 19.4317 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.81 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 156.2400 0.7200 156.6200 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 15.9225 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 81.2247 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.356071 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 155.0200 0.7200 155.4000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.9204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 209.3100 69.9200 209.6900 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.7464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 207.4800 69.9200 207.8600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 205.6500 69.9200 206.0300 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 203.8200 69.9200 204.2000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.8096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.592 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 201.9900 69.9200 202.3700 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.0036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.96 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 200.1600 69.9200 200.5400 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.6798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.096 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 198.3300 69.9200 198.7100 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.1348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.856 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 196.5000 69.9200 196.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.185 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.5968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.32 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 195.2800 69.9200 195.6600 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7806 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.8668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 193.4500 69.9200 193.8300 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.688 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 191.6200 69.9200 192.0000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.4398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.816 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 189.7900 69.9200 190.1700 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6086 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.3788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.824 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 187.9600 69.9200 188.3400 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.5488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.064 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 186.1300 69.9200 186.5100 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 184.3000 69.9200 184.6800 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 182.4700 69.9200 182.8500 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.7684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.76 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 181.2500 69.9200 181.6300 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.1314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.696 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 179.4200 69.9200 179.8000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 177.5900 69.9200 177.9700 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.3064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 175.7600 69.9200 176.1400 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.88 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 173.9300 69.9200 174.3100 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 172.1000 69.9200 172.4800 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.6726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.528 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 170.8800 69.9200 171.2600 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 169.6600 69.9200 170.0400 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.5778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 115.552 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 168.4400 69.9200 168.8200 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.1918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 167.2200 69.9200 167.6000 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.4968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.12 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 166.0000 69.9200 166.3800 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.888 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 162.9500 69.9200 163.3300 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.616 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 159.9000 69.9200 160.2800 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9106 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.2078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 158.0700 69.9200 158.4500 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 156.2400 69.9200 156.6200 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.944 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.2000 155.0200 69.9200 155.4000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.98397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.5253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 59.3800 0.0000 59.7600 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.80835 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.951 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6796 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.23892 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.89091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 56.6200 0.0000 57.0000 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4845 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.8668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 67.8327 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 359.162 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 53.8600 0.0000 54.2400 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.02236 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.71717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 51.1000 0.0000 51.4800 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.39569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.5838 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 48.3400 0.0000 48.7200 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.1104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.478 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 8.52579 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 41.398 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 42.8200 0.0000 43.2000 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.8538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.7758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.065 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 40.0600 0.0000 40.4400 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.9 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 144.382 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 42.1473 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 208.646 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 37.3000 0.0000 37.6800 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.5037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.3528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.6121 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 329.662 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 34.5400 0.0000 34.9200 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.40013 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 5.60606 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 0.0000 32.1600 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.7204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.528 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 10.6941 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 52.2397 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 29.4800 0.0000 29.8600 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.78343 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.5226 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 26.7200 0.0000 27.1000 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.2936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.19205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.56566 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 23.9600 0.0000 24.3400 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 27.122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.492 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 39.0502 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 193.857 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 21.2000 0.0000 21.5800 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.8196 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.024 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 6.96936 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 32.9199 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 18.4400 0.0000 18.8200 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.964 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.5534 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.3724 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 15.6800 0.0000 16.0600 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3616 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 26.3799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5815 LAYER met2  ;
    ANTENNAMAXAREACAR 34.2113 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 165.71 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.49577 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.2056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.704 LAYER met3  ;
    ANTENNAGATEAREA 3.0585 LAYER met3  ;
    ANTENNAMAXAREACAR 35.9133 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.094 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 12.9200 0.0000 13.3000 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.5844 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 140.287 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8995 LAYER met2  ;
    ANTENNAMAXAREACAR 34.1515 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 164.864 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.661471 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.944 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 38.0924 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 186.237 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.669182 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 0.0000 10.5400 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 24.0363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.311 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met2  ;
    ANTENNAMAXAREACAR 22.2111 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.459 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.477858 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.1796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.232 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 24.3934 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.883 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 7.4000 0.0000 7.7800 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 24.3707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2175 LAYER met2  ;
    ANTENNAMAXAREACAR 30.3021 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 140.872 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.631153 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.5963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.44 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 33.4427 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 157.881 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.642228 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 5.1000 0.0000 5.4800 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.6596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.224 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 59.3800 218.9200 59.7600 219.6400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.2088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 218.9200 56.5400 219.6400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 218.9200 53.7800 219.6400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.5051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.7448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.776 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 218.9200 51.0200 219.6400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.86615 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.019 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.7019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.3385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.0198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.576 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 218.9200 48.2600 219.6400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 44.6600 218.9200 45.0400 219.6400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 41.9000 218.9200 42.2800 219.6400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.1400 218.9200 39.5200 219.6400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.3800 218.9200 36.7600 219.6400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.2207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.0348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.6200 218.9200 34.0000 219.6400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 218.9200 30.7800 219.6400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.5399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.2178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 193.632 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 218.9200 28.0200 219.6400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.1745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.1958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 218.9200 25.2600 219.6400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9412 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.248 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 218.9200 22.5000 219.6400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.176 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 218.9200 19.7400 219.6400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.7861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.1328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.512 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.1400 218.9200 16.5200 219.6400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.052 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 13.3800 218.9200 13.7600 219.6400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.1858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.6200 218.9200 11.0000 219.6400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2124 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.988 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 7.8600 218.9200 8.2400 219.6400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.5047 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.535 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.8316 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.121 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 5.1000 218.9200 5.4800 219.6400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 3.3900 5.3300 66.5300 6.3300 ;
        RECT 3.3900 212.6300 66.5300 213.6300 ;
        RECT 3.3900 12.3400 4.3900 12.8200 ;
        RECT 3.3900 23.2200 4.3900 23.7000 ;
        RECT 3.3900 17.7800 4.3900 18.2600 ;
        RECT 3.3900 39.5400 4.3900 40.0200 ;
        RECT 3.3900 34.1000 4.3900 34.5800 ;
        RECT 3.3900 28.6600 4.3900 29.1400 ;
        RECT 3.3900 50.4200 4.3900 50.9000 ;
        RECT 3.3900 44.9800 4.3900 45.4600 ;
        RECT 3.3900 66.7400 4.3900 67.2200 ;
        RECT 3.3900 61.3000 4.3900 61.7800 ;
        RECT 3.3900 55.8600 4.3900 56.3400 ;
        RECT 3.3900 77.6200 4.3900 78.1000 ;
        RECT 3.3900 72.1800 4.3900 72.6600 ;
        RECT 3.3900 93.9400 4.3900 94.4200 ;
        RECT 3.3900 88.5000 4.3900 88.9800 ;
        RECT 3.3900 83.0600 4.3900 83.5400 ;
        RECT 3.3900 104.8200 4.3900 105.3000 ;
        RECT 3.3900 99.3800 4.3900 99.8600 ;
        RECT 65.5300 12.3400 66.5300 12.8200 ;
        RECT 65.5300 23.2200 66.5300 23.7000 ;
        RECT 65.5300 17.7800 66.5300 18.2600 ;
        RECT 65.5300 39.5400 66.5300 40.0200 ;
        RECT 65.5300 34.1000 66.5300 34.5800 ;
        RECT 65.5300 28.6600 66.5300 29.1400 ;
        RECT 65.5300 50.4200 66.5300 50.9000 ;
        RECT 65.5300 44.9800 66.5300 45.4600 ;
        RECT 65.5300 66.7400 66.5300 67.2200 ;
        RECT 65.5300 61.3000 66.5300 61.7800 ;
        RECT 65.5300 55.8600 66.5300 56.3400 ;
        RECT 65.5300 77.6200 66.5300 78.1000 ;
        RECT 65.5300 72.1800 66.5300 72.6600 ;
        RECT 65.5300 93.9400 66.5300 94.4200 ;
        RECT 65.5300 88.5000 66.5300 88.9800 ;
        RECT 65.5300 83.0600 66.5300 83.5400 ;
        RECT 65.5300 104.8200 66.5300 105.3000 ;
        RECT 65.5300 99.3800 66.5300 99.8600 ;
        RECT 3.3900 164.6600 4.3900 165.1400 ;
        RECT 3.3900 121.1400 4.3900 121.6200 ;
        RECT 3.3900 115.7000 4.3900 116.1800 ;
        RECT 3.3900 110.2600 4.3900 110.7400 ;
        RECT 3.3900 132.0200 4.3900 132.5000 ;
        RECT 3.3900 126.5800 4.3900 127.0600 ;
        RECT 3.3900 148.3400 4.3900 148.8200 ;
        RECT 3.3900 142.9000 4.3900 143.3800 ;
        RECT 3.3900 137.4600 4.3900 137.9400 ;
        RECT 3.3900 159.2200 4.3900 159.7000 ;
        RECT 3.3900 153.7800 4.3900 154.2600 ;
        RECT 3.3900 191.8600 4.3900 192.3400 ;
        RECT 3.3900 175.5400 4.3900 176.0200 ;
        RECT 3.3900 170.1000 4.3900 170.5800 ;
        RECT 3.3900 186.4200 4.3900 186.9000 ;
        RECT 3.3900 180.9800 4.3900 181.4600 ;
        RECT 3.3900 202.7400 4.3900 203.2200 ;
        RECT 3.3900 197.3000 4.3900 197.7800 ;
        RECT 3.3900 208.1800 4.3900 208.6600 ;
        RECT 65.5300 164.6600 66.5300 165.1400 ;
        RECT 65.5300 121.1400 66.5300 121.6200 ;
        RECT 65.5300 115.7000 66.5300 116.1800 ;
        RECT 65.5300 110.2600 66.5300 110.7400 ;
        RECT 65.5300 132.0200 66.5300 132.5000 ;
        RECT 65.5300 126.5800 66.5300 127.0600 ;
        RECT 65.5300 148.3400 66.5300 148.8200 ;
        RECT 65.5300 142.9000 66.5300 143.3800 ;
        RECT 65.5300 137.4600 66.5300 137.9400 ;
        RECT 65.5300 159.2200 66.5300 159.7000 ;
        RECT 65.5300 153.7800 66.5300 154.2600 ;
        RECT 65.5300 191.8600 66.5300 192.3400 ;
        RECT 65.5300 175.5400 66.5300 176.0200 ;
        RECT 65.5300 170.1000 66.5300 170.5800 ;
        RECT 65.5300 186.4200 66.5300 186.9000 ;
        RECT 65.5300 180.9800 66.5300 181.4600 ;
        RECT 65.5300 202.7400 66.5300 203.2200 ;
        RECT 65.5300 197.3000 66.5300 197.7800 ;
        RECT 65.5300 208.1800 66.5300 208.6600 ;
      LAYER met4 ;
        RECT 3.3900 5.3300 4.3900 213.6300 ;
        RECT 65.5300 5.3300 66.5300 213.6300 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 1.5900 3.5300 68.3300 4.5300 ;
        RECT 1.5900 214.4300 68.3300 215.4300 ;
        RECT 1.5900 9.6200 2.5900 10.1000 ;
        RECT 1.5900 25.9400 2.5900 26.4200 ;
        RECT 1.5900 20.5000 2.5900 20.9800 ;
        RECT 1.5900 15.0600 2.5900 15.5400 ;
        RECT 1.5900 36.8200 2.5900 37.3000 ;
        RECT 1.5900 31.3800 2.5900 31.8600 ;
        RECT 1.5900 53.1400 2.5900 53.6200 ;
        RECT 1.5900 47.7000 2.5900 48.1800 ;
        RECT 1.5900 42.2600 2.5900 42.7400 ;
        RECT 1.5900 64.0200 2.5900 64.5000 ;
        RECT 1.5900 58.5800 2.5900 59.0600 ;
        RECT 1.5900 80.3400 2.5900 80.8200 ;
        RECT 1.5900 74.9000 2.5900 75.3800 ;
        RECT 1.5900 69.4600 2.5900 69.9400 ;
        RECT 1.5900 91.2200 2.5900 91.7000 ;
        RECT 1.5900 85.7800 2.5900 86.2600 ;
        RECT 1.5900 107.5400 2.5900 108.0200 ;
        RECT 1.5900 102.1000 2.5900 102.5800 ;
        RECT 1.5900 96.6600 2.5900 97.1400 ;
        RECT 67.3300 9.6200 68.3300 10.1000 ;
        RECT 67.3300 25.9400 68.3300 26.4200 ;
        RECT 67.3300 20.5000 68.3300 20.9800 ;
        RECT 67.3300 15.0600 68.3300 15.5400 ;
        RECT 67.3300 36.8200 68.3300 37.3000 ;
        RECT 67.3300 31.3800 68.3300 31.8600 ;
        RECT 67.3300 53.1400 68.3300 53.6200 ;
        RECT 67.3300 47.7000 68.3300 48.1800 ;
        RECT 67.3300 42.2600 68.3300 42.7400 ;
        RECT 67.3300 64.0200 68.3300 64.5000 ;
        RECT 67.3300 58.5800 68.3300 59.0600 ;
        RECT 67.3300 80.3400 68.3300 80.8200 ;
        RECT 67.3300 74.9000 68.3300 75.3800 ;
        RECT 67.3300 69.4600 68.3300 69.9400 ;
        RECT 67.3300 91.2200 68.3300 91.7000 ;
        RECT 67.3300 85.7800 68.3300 86.2600 ;
        RECT 67.3300 107.5400 68.3300 108.0200 ;
        RECT 67.3300 102.1000 68.3300 102.5800 ;
        RECT 67.3300 96.6600 68.3300 97.1400 ;
        RECT 1.5900 118.4200 2.5900 118.9000 ;
        RECT 1.5900 112.9800 2.5900 113.4600 ;
        RECT 1.5900 134.7400 2.5900 135.2200 ;
        RECT 1.5900 129.3000 2.5900 129.7800 ;
        RECT 1.5900 123.8600 2.5900 124.3400 ;
        RECT 1.5900 145.6200 2.5900 146.1000 ;
        RECT 1.5900 140.1800 2.5900 140.6600 ;
        RECT 1.5900 161.9400 2.5900 162.4200 ;
        RECT 1.5900 156.5000 2.5900 156.9800 ;
        RECT 1.5900 151.0600 2.5900 151.5400 ;
        RECT 1.5900 178.2600 2.5900 178.7400 ;
        RECT 1.5900 172.8200 2.5900 173.3000 ;
        RECT 1.5900 167.3800 2.5900 167.8600 ;
        RECT 1.5900 189.1400 2.5900 189.6200 ;
        RECT 1.5900 183.7000 2.5900 184.1800 ;
        RECT 1.5900 205.4600 2.5900 205.9400 ;
        RECT 1.5900 200.0200 2.5900 200.5000 ;
        RECT 1.5900 194.5800 2.5900 195.0600 ;
        RECT 67.3300 118.4200 68.3300 118.9000 ;
        RECT 67.3300 112.9800 68.3300 113.4600 ;
        RECT 67.3300 134.7400 68.3300 135.2200 ;
        RECT 67.3300 129.3000 68.3300 129.7800 ;
        RECT 67.3300 123.8600 68.3300 124.3400 ;
        RECT 67.3300 145.6200 68.3300 146.1000 ;
        RECT 67.3300 140.1800 68.3300 140.6600 ;
        RECT 67.3300 161.9400 68.3300 162.4200 ;
        RECT 67.3300 156.5000 68.3300 156.9800 ;
        RECT 67.3300 151.0600 68.3300 151.5400 ;
        RECT 67.3300 178.2600 68.3300 178.7400 ;
        RECT 67.3300 172.8200 68.3300 173.3000 ;
        RECT 67.3300 167.3800 68.3300 167.8600 ;
        RECT 67.3300 189.1400 68.3300 189.6200 ;
        RECT 67.3300 183.7000 68.3300 184.1800 ;
        RECT 67.3300 205.4600 68.3300 205.9400 ;
        RECT 67.3300 200.0200 68.3300 200.5000 ;
        RECT 67.3300 194.5800 68.3300 195.0600 ;
      LAYER met4 ;
        RECT 1.5900 3.5300 2.5900 215.4300 ;
        RECT 67.3300 3.5300 68.3300 215.4300 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 59.9300 218.7500 69.9200 219.6400 ;
      RECT 56.7100 218.7500 59.2100 219.6400 ;
      RECT 53.9500 218.7500 55.9900 219.6400 ;
      RECT 51.1900 218.7500 53.2300 219.6400 ;
      RECT 48.4300 218.7500 50.4700 219.6400 ;
      RECT 45.2100 218.7500 47.7100 219.6400 ;
      RECT 42.4500 218.7500 44.4900 219.6400 ;
      RECT 39.6900 218.7500 41.7300 219.6400 ;
      RECT 36.9300 218.7500 38.9700 219.6400 ;
      RECT 34.1700 218.7500 36.2100 219.6400 ;
      RECT 30.9500 218.7500 33.4500 219.6400 ;
      RECT 28.1900 218.7500 30.2300 219.6400 ;
      RECT 25.4300 218.7500 27.4700 219.6400 ;
      RECT 22.6700 218.7500 24.7100 219.6400 ;
      RECT 19.9100 218.7500 21.9500 219.6400 ;
      RECT 16.6900 218.7500 19.1900 219.6400 ;
      RECT 13.9300 218.7500 15.9700 219.6400 ;
      RECT 11.1700 218.7500 13.2100 219.6400 ;
      RECT 8.4100 218.7500 10.4500 219.6400 ;
      RECT 5.6500 218.7500 7.6900 219.6400 ;
      RECT 0.0000 218.7500 4.9300 219.6400 ;
      RECT 0.0000 0.8900 69.9200 218.7500 ;
      RECT 59.9300 0.0000 69.9200 0.8900 ;
      RECT 57.1700 0.0000 59.2100 0.8900 ;
      RECT 54.4100 0.0000 56.4500 0.8900 ;
      RECT 51.6500 0.0000 53.6900 0.8900 ;
      RECT 48.8900 0.0000 50.9300 0.8900 ;
      RECT 46.1300 0.0000 48.1700 0.8900 ;
      RECT 43.3700 0.0000 45.4100 0.8900 ;
      RECT 40.6100 0.0000 42.6500 0.8900 ;
      RECT 37.8500 0.0000 39.8900 0.8900 ;
      RECT 35.0900 0.0000 37.1300 0.8900 ;
      RECT 32.3300 0.0000 34.3700 0.8900 ;
      RECT 30.0300 0.0000 31.6100 0.8900 ;
      RECT 27.2700 0.0000 29.3100 0.8900 ;
      RECT 24.5100 0.0000 26.5500 0.8900 ;
      RECT 21.7500 0.0000 23.7900 0.8900 ;
      RECT 18.9900 0.0000 21.0300 0.8900 ;
      RECT 16.2300 0.0000 18.2700 0.8900 ;
      RECT 13.4700 0.0000 15.5100 0.8900 ;
      RECT 10.7100 0.0000 12.7500 0.8900 ;
      RECT 7.9500 0.0000 9.9900 0.8900 ;
      RECT 5.6500 0.0000 7.2300 0.8900 ;
      RECT 0.0000 0.0000 4.9300 0.8900 ;
    LAYER met1 ;
      RECT 0.0000 150.1000 69.9200 219.6400 ;
      RECT 0.0000 149.4400 69.0600 150.1000 ;
      RECT 0.0000 148.4000 69.9200 149.4400 ;
      RECT 0.0000 147.7400 69.0600 148.4000 ;
      RECT 0.0000 147.0400 69.9200 147.7400 ;
      RECT 0.0000 146.3800 69.0600 147.0400 ;
      RECT 0.0000 145.6800 69.9200 146.3800 ;
      RECT 0.0000 145.0200 69.0600 145.6800 ;
      RECT 0.0000 143.9800 69.9200 145.0200 ;
      RECT 0.0000 143.3200 69.0600 143.9800 ;
      RECT 0.0000 142.6200 69.9200 143.3200 ;
      RECT 0.0000 141.9600 69.0600 142.6200 ;
      RECT 0.0000 141.2600 69.9200 141.9600 ;
      RECT 0.0000 140.6000 69.0600 141.2600 ;
      RECT 0.0000 139.5600 69.9200 140.6000 ;
      RECT 0.0000 138.9000 69.0600 139.5600 ;
      RECT 0.0000 137.8600 69.9200 138.9000 ;
      RECT 0.0000 137.2000 69.0600 137.8600 ;
      RECT 0.0000 136.8400 69.9200 137.2000 ;
      RECT 0.0000 136.1800 69.0600 136.8400 ;
      RECT 0.0000 134.4600 69.9200 136.1800 ;
      RECT 0.0000 133.8000 69.0600 134.4600 ;
      RECT 0.0000 133.7800 69.9200 133.8000 ;
      RECT 0.0000 133.1200 69.0600 133.7800 ;
      RECT 0.0000 132.4200 69.9200 133.1200 ;
      RECT 0.0000 131.7600 69.0600 132.4200 ;
      RECT 0.0000 130.3800 69.9200 131.7600 ;
      RECT 0.0000 129.7200 69.0600 130.3800 ;
      RECT 0.0000 129.3600 69.9200 129.7200 ;
      RECT 0.0000 128.7000 69.0600 129.3600 ;
      RECT 0.0000 128.0000 69.9200 128.7000 ;
      RECT 0.0000 127.3400 69.0600 128.0000 ;
      RECT 0.0000 126.3000 69.9200 127.3400 ;
      RECT 0.0000 125.6400 69.0600 126.3000 ;
      RECT 0.0000 124.9400 69.9200 125.6400 ;
      RECT 0.0000 124.2800 69.0600 124.9400 ;
      RECT 0.0000 123.5800 69.9200 124.2800 ;
      RECT 0.0000 122.9200 69.0600 123.5800 ;
      RECT 0.0000 121.8800 69.9200 122.9200 ;
      RECT 0.0000 121.2200 69.0600 121.8800 ;
      RECT 0.0000 120.5200 69.9200 121.2200 ;
      RECT 0.0000 119.8600 69.0600 120.5200 ;
      RECT 0.0000 119.1600 69.9200 119.8600 ;
      RECT 0.0000 118.5000 69.0600 119.1600 ;
      RECT 0.0000 117.4600 69.9200 118.5000 ;
      RECT 0.0000 116.8000 69.0600 117.4600 ;
      RECT 0.0000 116.1000 69.9200 116.8000 ;
      RECT 0.0000 115.4400 69.0600 116.1000 ;
      RECT 0.0000 114.7400 69.9200 115.4400 ;
      RECT 0.0000 114.0800 69.0600 114.7400 ;
      RECT 0.0000 113.0400 69.9200 114.0800 ;
      RECT 0.0000 112.3800 69.0600 113.0400 ;
      RECT 0.0000 111.6800 69.9200 112.3800 ;
      RECT 0.0000 111.0200 69.0600 111.6800 ;
      RECT 0.0000 110.3200 69.9200 111.0200 ;
      RECT 0.8600 109.6600 69.0600 110.3200 ;
      RECT 0.0000 108.9600 69.9200 109.6600 ;
      RECT 0.0000 108.3000 69.0600 108.9600 ;
      RECT 0.0000 108.2800 69.9200 108.3000 ;
      RECT 0.0000 107.9400 69.0600 108.2800 ;
      RECT 0.8600 107.6200 69.0600 107.9400 ;
      RECT 0.8600 107.2800 69.9200 107.6200 ;
      RECT 0.0000 105.9000 69.9200 107.2800 ;
      RECT 0.0000 105.5600 69.0600 105.9000 ;
      RECT 0.8600 105.2400 69.0600 105.5600 ;
      RECT 0.8600 104.9000 69.9200 105.2400 ;
      RECT 0.0000 103.8600 69.9200 104.9000 ;
      RECT 0.0000 103.2000 69.0600 103.8600 ;
      RECT 0.0000 103.1800 69.9200 103.2000 ;
      RECT 0.8600 102.8400 69.9200 103.1800 ;
      RECT 0.8600 102.5200 69.0600 102.8400 ;
      RECT 0.0000 102.1800 69.0600 102.5200 ;
      RECT 0.0000 101.8200 69.9200 102.1800 ;
      RECT 0.0000 101.1600 69.0600 101.8200 ;
      RECT 0.0000 101.1400 69.9200 101.1600 ;
      RECT 0.0000 100.8000 69.0600 101.1400 ;
      RECT 0.8600 100.4800 69.0600 100.8000 ;
      RECT 0.8600 100.1400 69.9200 100.4800 ;
      RECT 0.0000 98.7600 69.9200 100.1400 ;
      RECT 0.8600 98.4200 69.9200 98.7600 ;
      RECT 0.8600 98.1000 69.0600 98.4200 ;
      RECT 0.0000 97.7600 69.0600 98.1000 ;
      RECT 0.0000 97.0600 69.9200 97.7600 ;
      RECT 0.0000 96.4000 69.0600 97.0600 ;
      RECT 0.0000 96.3800 69.9200 96.4000 ;
      RECT 0.8600 95.7200 69.9200 96.3800 ;
      RECT 0.0000 95.3600 69.9200 95.7200 ;
      RECT 0.0000 94.7000 69.0600 95.3600 ;
      RECT 0.0000 94.0000 69.9200 94.7000 ;
      RECT 0.8600 93.3400 69.0600 94.0000 ;
      RECT 0.0000 92.6400 69.9200 93.3400 ;
      RECT 0.0000 91.9800 69.0600 92.6400 ;
      RECT 0.0000 91.6200 69.9200 91.9800 ;
      RECT 0.8600 90.9600 69.9200 91.6200 ;
      RECT 0.0000 90.9400 69.9200 90.9600 ;
      RECT 0.0000 90.2800 69.0600 90.9400 ;
      RECT 0.0000 89.5800 69.9200 90.2800 ;
      RECT 0.8600 88.9200 69.0600 89.5800 ;
      RECT 0.0000 88.2200 69.9200 88.9200 ;
      RECT 0.0000 87.5600 69.0600 88.2200 ;
      RECT 0.0000 87.2000 69.9200 87.5600 ;
      RECT 0.8600 86.5400 69.9200 87.2000 ;
      RECT 0.0000 86.5200 69.9200 86.5400 ;
      RECT 0.0000 85.8600 69.0600 86.5200 ;
      RECT 0.0000 85.1600 69.9200 85.8600 ;
      RECT 0.0000 84.8200 69.0600 85.1600 ;
      RECT 0.8600 84.5000 69.0600 84.8200 ;
      RECT 0.8600 84.1600 69.9200 84.5000 ;
      RECT 0.0000 83.8000 69.9200 84.1600 ;
      RECT 0.0000 83.1400 69.0600 83.8000 ;
      RECT 0.0000 82.4400 69.9200 83.1400 ;
      RECT 0.8600 82.1000 69.9200 82.4400 ;
      RECT 0.8600 81.7800 69.0600 82.1000 ;
      RECT 0.0000 81.4400 69.0600 81.7800 ;
      RECT 0.0000 80.7400 69.9200 81.4400 ;
      RECT 0.0000 80.4000 69.0600 80.7400 ;
      RECT 0.8600 80.0800 69.0600 80.4000 ;
      RECT 0.8600 79.7400 69.9200 80.0800 ;
      RECT 0.0000 79.3800 69.9200 79.7400 ;
      RECT 0.0000 78.7200 69.0600 79.3800 ;
      RECT 0.0000 78.0200 69.9200 78.7200 ;
      RECT 0.0000 77.3600 69.0600 78.0200 ;
      RECT 0.0000 76.3200 69.9200 77.3600 ;
      RECT 0.0000 75.6600 69.0600 76.3200 ;
      RECT 0.0000 74.9600 69.9200 75.6600 ;
      RECT 0.0000 74.3000 69.0600 74.9600 ;
      RECT 0.0000 73.6000 69.9200 74.3000 ;
      RECT 0.0000 72.9400 69.0600 73.6000 ;
      RECT 0.0000 71.9000 69.9200 72.9400 ;
      RECT 0.0000 71.2400 69.0600 71.9000 ;
      RECT 0.0000 70.5400 69.9200 71.2400 ;
      RECT 0.0000 69.8800 69.0600 70.5400 ;
      RECT 0.0000 69.1800 69.9200 69.8800 ;
      RECT 0.0000 68.5200 69.0600 69.1800 ;
      RECT 0.0000 68.1600 69.9200 68.5200 ;
      RECT 0.0000 67.5000 69.0600 68.1600 ;
      RECT 0.0000 66.1200 69.9200 67.5000 ;
      RECT 0.0000 65.4600 69.0600 66.1200 ;
      RECT 0.0000 64.7600 69.9200 65.4600 ;
      RECT 0.0000 64.1000 69.0600 64.7600 ;
      RECT 0.0000 63.0600 69.9200 64.1000 ;
      RECT 0.0000 62.4000 69.0600 63.0600 ;
      RECT 0.0000 62.0400 69.9200 62.4000 ;
      RECT 0.0000 61.3800 69.0600 62.0400 ;
      RECT 0.0000 60.3400 69.9200 61.3800 ;
      RECT 0.0000 59.6800 69.0600 60.3400 ;
      RECT 0.0000 58.9800 69.9200 59.6800 ;
      RECT 0.0000 58.3200 69.0600 58.9800 ;
      RECT 0.0000 58.3000 69.9200 58.3200 ;
      RECT 0.0000 57.6400 69.0600 58.3000 ;
      RECT 0.0000 55.2400 69.9200 57.6400 ;
      RECT 0.0000 54.5800 69.0600 55.2400 ;
      RECT 0.0000 54.2200 69.9200 54.5800 ;
      RECT 0.0000 53.5600 69.0600 54.2200 ;
      RECT 0.0000 52.8600 69.9200 53.5600 ;
      RECT 0.0000 52.2000 69.0600 52.8600 ;
      RECT 0.0000 51.5000 69.9200 52.2000 ;
      RECT 0.0000 50.8400 69.0600 51.5000 ;
      RECT 0.0000 49.8000 69.9200 50.8400 ;
      RECT 0.0000 49.1400 69.0600 49.8000 ;
      RECT 0.0000 48.4400 69.9200 49.1400 ;
      RECT 0.0000 47.7800 69.0600 48.4400 ;
      RECT 0.0000 47.4200 69.9200 47.7800 ;
      RECT 0.0000 46.7600 69.0600 47.4200 ;
      RECT 0.0000 46.7400 69.9200 46.7600 ;
      RECT 0.0000 46.0800 69.0600 46.7400 ;
      RECT 0.0000 44.0200 69.9200 46.0800 ;
      RECT 0.0000 43.3600 69.0600 44.0200 ;
      RECT 0.0000 42.6600 69.9200 43.3600 ;
      RECT 0.0000 42.0000 69.0600 42.6600 ;
      RECT 0.0000 41.3000 69.9200 42.0000 ;
      RECT 0.0000 40.6400 69.0600 41.3000 ;
      RECT 0.0000 39.6000 69.9200 40.6400 ;
      RECT 0.0000 38.9400 69.0600 39.6000 ;
      RECT 0.0000 38.2400 69.9200 38.9400 ;
      RECT 0.0000 37.5800 69.0600 38.2400 ;
      RECT 0.0000 36.5400 69.9200 37.5800 ;
      RECT 0.0000 35.8800 69.0600 36.5400 ;
      RECT 0.0000 35.1800 69.9200 35.8800 ;
      RECT 0.0000 34.5200 69.0600 35.1800 ;
      RECT 0.0000 33.8200 69.9200 34.5200 ;
      RECT 0.0000 33.1600 69.0600 33.8200 ;
      RECT 0.0000 32.1200 69.9200 33.1600 ;
      RECT 0.0000 31.4600 69.0600 32.1200 ;
      RECT 0.0000 30.7600 69.9200 31.4600 ;
      RECT 0.0000 30.1000 69.0600 30.7600 ;
      RECT 0.0000 29.4000 69.9200 30.1000 ;
      RECT 0.0000 28.7400 69.0600 29.4000 ;
      RECT 0.0000 27.7000 69.9200 28.7400 ;
      RECT 0.0000 27.0400 69.0600 27.7000 ;
      RECT 0.0000 26.3400 69.9200 27.0400 ;
      RECT 0.0000 25.6800 69.0600 26.3400 ;
      RECT 0.0000 24.9800 69.9200 25.6800 ;
      RECT 0.0000 24.3200 69.0600 24.9800 ;
      RECT 0.0000 23.2800 69.9200 24.3200 ;
      RECT 0.0000 22.6200 69.0600 23.2800 ;
      RECT 0.0000 21.9200 69.9200 22.6200 ;
      RECT 0.0000 21.2600 69.0600 21.9200 ;
      RECT 0.0000 20.5600 69.9200 21.2600 ;
      RECT 0.0000 19.9000 69.0600 20.5600 ;
      RECT 0.0000 18.8600 69.9200 19.9000 ;
      RECT 0.0000 18.2000 69.0600 18.8600 ;
      RECT 0.0000 17.5000 69.9200 18.2000 ;
      RECT 0.0000 16.8400 69.0600 17.5000 ;
      RECT 0.0000 16.1400 69.9200 16.8400 ;
      RECT 0.0000 15.4800 69.0600 16.1400 ;
      RECT 0.0000 14.4400 69.9200 15.4800 ;
      RECT 0.0000 13.7800 69.0600 14.4400 ;
      RECT 0.0000 13.0800 69.9200 13.7800 ;
      RECT 0.0000 12.4200 69.0600 13.0800 ;
      RECT 0.0000 11.7200 69.9200 12.4200 ;
      RECT 0.0000 11.0600 69.0600 11.7200 ;
      RECT 0.0000 10.3600 69.9200 11.0600 ;
      RECT 0.0000 9.7000 69.0600 10.3600 ;
      RECT 0.0000 0.0000 69.9200 9.7000 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 69.9200 219.6400 ;
    LAYER met3 ;
      RECT 0.0000 215.7300 69.9200 219.6400 ;
      RECT 68.6300 214.1300 69.9200 215.7300 ;
      RECT 0.0000 214.1300 1.2900 215.7300 ;
      RECT 0.0000 213.9300 69.9200 214.1300 ;
      RECT 66.8300 212.3300 69.9200 213.9300 ;
      RECT 0.0000 212.3300 3.0900 213.9300 ;
      RECT 0.0000 209.9900 69.9200 212.3300 ;
      RECT 1.0200 209.0100 68.9000 209.9900 ;
      RECT 0.0000 208.9600 69.9200 209.0100 ;
      RECT 66.8300 208.1600 69.9200 208.9600 ;
      RECT 0.0000 208.1600 3.0900 208.9600 ;
      RECT 66.8300 207.8800 68.9000 208.1600 ;
      RECT 4.6900 207.8800 65.2300 208.9600 ;
      RECT 1.0200 207.8800 3.0900 208.1600 ;
      RECT 1.0200 207.1800 68.9000 207.8800 ;
      RECT 0.0000 206.3300 69.9200 207.1800 ;
      RECT 1.0200 206.2400 68.9000 206.3300 ;
      RECT 68.6300 205.3500 68.9000 206.2400 ;
      RECT 1.0200 205.3500 1.2900 206.2400 ;
      RECT 68.6300 205.1600 69.9200 205.3500 ;
      RECT 2.8900 205.1600 67.0300 206.2400 ;
      RECT 0.0000 205.1600 1.2900 205.3500 ;
      RECT 0.0000 204.5000 69.9200 205.1600 ;
      RECT 1.0200 203.5200 68.9000 204.5000 ;
      RECT 66.8300 202.6700 69.9200 203.5200 ;
      RECT 0.0000 202.6700 3.0900 203.5200 ;
      RECT 66.8300 202.4400 68.9000 202.6700 ;
      RECT 4.6900 202.4400 65.2300 203.5200 ;
      RECT 1.0200 202.4400 3.0900 202.6700 ;
      RECT 1.0200 201.6900 68.9000 202.4400 ;
      RECT 0.0000 200.8400 69.9200 201.6900 ;
      RECT 1.0200 200.8000 68.9000 200.8400 ;
      RECT 68.6300 199.8600 68.9000 200.8000 ;
      RECT 1.0200 199.8600 1.2900 200.8000 ;
      RECT 68.6300 199.7200 69.9200 199.8600 ;
      RECT 2.8900 199.7200 67.0300 200.8000 ;
      RECT 0.0000 199.7200 1.2900 199.8600 ;
      RECT 0.0000 199.0100 69.9200 199.7200 ;
      RECT 1.0200 198.0800 68.9000 199.0100 ;
      RECT 66.8300 198.0300 68.9000 198.0800 ;
      RECT 1.0200 198.0300 3.0900 198.0800 ;
      RECT 66.8300 197.1800 69.9200 198.0300 ;
      RECT 0.0000 197.1800 3.0900 198.0300 ;
      RECT 66.8300 197.0000 68.9000 197.1800 ;
      RECT 4.6900 197.0000 65.2300 198.0800 ;
      RECT 1.0200 197.0000 3.0900 197.1800 ;
      RECT 1.0200 196.2000 68.9000 197.0000 ;
      RECT 0.0000 195.9600 69.9200 196.2000 ;
      RECT 1.0200 195.3600 68.9000 195.9600 ;
      RECT 68.6300 194.9800 68.9000 195.3600 ;
      RECT 1.0200 194.9800 1.2900 195.3600 ;
      RECT 68.6300 194.2800 69.9200 194.9800 ;
      RECT 2.8900 194.2800 67.0300 195.3600 ;
      RECT 0.0000 194.2800 1.2900 194.9800 ;
      RECT 0.0000 194.1300 69.9200 194.2800 ;
      RECT 1.0200 193.1500 68.9000 194.1300 ;
      RECT 0.0000 192.6400 69.9200 193.1500 ;
      RECT 66.8300 192.3000 69.9200 192.6400 ;
      RECT 0.0000 192.3000 3.0900 192.6400 ;
      RECT 66.8300 191.5600 68.9000 192.3000 ;
      RECT 4.6900 191.5600 65.2300 192.6400 ;
      RECT 1.0200 191.5600 3.0900 192.3000 ;
      RECT 1.0200 191.3200 68.9000 191.5600 ;
      RECT 0.0000 190.4700 69.9200 191.3200 ;
      RECT 1.0200 189.9200 68.9000 190.4700 ;
      RECT 68.6300 189.4900 68.9000 189.9200 ;
      RECT 1.0200 189.4900 1.2900 189.9200 ;
      RECT 68.6300 188.8400 69.9200 189.4900 ;
      RECT 2.8900 188.8400 67.0300 189.9200 ;
      RECT 0.0000 188.8400 1.2900 189.4900 ;
      RECT 0.0000 188.6400 69.9200 188.8400 ;
      RECT 1.0200 187.6600 68.9000 188.6400 ;
      RECT 0.0000 187.2000 69.9200 187.6600 ;
      RECT 66.8300 186.8100 69.9200 187.2000 ;
      RECT 0.0000 186.8100 3.0900 187.2000 ;
      RECT 66.8300 186.1200 68.9000 186.8100 ;
      RECT 4.6900 186.1200 65.2300 187.2000 ;
      RECT 1.0200 186.1200 3.0900 186.8100 ;
      RECT 1.0200 185.8300 68.9000 186.1200 ;
      RECT 0.0000 184.9800 69.9200 185.8300 ;
      RECT 1.0200 184.4800 68.9000 184.9800 ;
      RECT 68.6300 184.0000 68.9000 184.4800 ;
      RECT 1.0200 184.0000 1.2900 184.4800 ;
      RECT 68.6300 183.4000 69.9200 184.0000 ;
      RECT 2.8900 183.4000 67.0300 184.4800 ;
      RECT 0.0000 183.4000 1.2900 184.0000 ;
      RECT 0.0000 183.1500 69.9200 183.4000 ;
      RECT 1.0200 182.1700 68.9000 183.1500 ;
      RECT 0.0000 181.9300 69.9200 182.1700 ;
      RECT 1.0200 181.7600 68.9000 181.9300 ;
      RECT 66.8300 180.9500 68.9000 181.7600 ;
      RECT 1.0200 180.9500 3.0900 181.7600 ;
      RECT 66.8300 180.6800 69.9200 180.9500 ;
      RECT 4.6900 180.6800 65.2300 181.7600 ;
      RECT 0.0000 180.6800 3.0900 180.9500 ;
      RECT 0.0000 180.1000 69.9200 180.6800 ;
      RECT 1.0200 179.1200 68.9000 180.1000 ;
      RECT 0.0000 179.0400 69.9200 179.1200 ;
      RECT 68.6300 178.2700 69.9200 179.0400 ;
      RECT 0.0000 178.2700 1.2900 179.0400 ;
      RECT 68.6300 177.9600 68.9000 178.2700 ;
      RECT 2.8900 177.9600 67.0300 179.0400 ;
      RECT 1.0200 177.9600 1.2900 178.2700 ;
      RECT 1.0200 177.2900 68.9000 177.9600 ;
      RECT 0.0000 176.4400 69.9200 177.2900 ;
      RECT 1.0200 176.3200 68.9000 176.4400 ;
      RECT 66.8300 175.4600 68.9000 176.3200 ;
      RECT 1.0200 175.4600 3.0900 176.3200 ;
      RECT 66.8300 175.2400 69.9200 175.4600 ;
      RECT 4.6900 175.2400 65.2300 176.3200 ;
      RECT 0.0000 175.2400 3.0900 175.4600 ;
      RECT 0.0000 174.6100 69.9200 175.2400 ;
      RECT 1.0200 173.6300 68.9000 174.6100 ;
      RECT 0.0000 173.6000 69.9200 173.6300 ;
      RECT 68.6300 172.7800 69.9200 173.6000 ;
      RECT 0.0000 172.7800 1.2900 173.6000 ;
      RECT 68.6300 172.5200 68.9000 172.7800 ;
      RECT 2.8900 172.5200 67.0300 173.6000 ;
      RECT 1.0200 172.5200 1.2900 172.7800 ;
      RECT 1.0200 171.8000 68.9000 172.5200 ;
      RECT 0.0000 171.5600 69.9200 171.8000 ;
      RECT 0.0000 170.9500 68.9000 171.5600 ;
      RECT 1.0200 170.8800 68.9000 170.9500 ;
      RECT 66.8300 170.5800 68.9000 170.8800 ;
      RECT 66.8300 170.3400 69.9200 170.5800 ;
      RECT 1.0200 169.9700 3.0900 170.8800 ;
      RECT 66.8300 169.8000 68.9000 170.3400 ;
      RECT 4.6900 169.8000 65.2300 170.8800 ;
      RECT 0.0000 169.8000 3.0900 169.9700 ;
      RECT 0.0000 169.3600 68.9000 169.8000 ;
      RECT 0.0000 169.1200 69.9200 169.3600 ;
      RECT 1.0200 168.1600 68.9000 169.1200 ;
      RECT 68.6300 168.1400 68.9000 168.1600 ;
      RECT 1.0200 168.1400 1.2900 168.1600 ;
      RECT 68.6300 167.9000 69.9200 168.1400 ;
      RECT 0.0000 167.9000 1.2900 168.1400 ;
      RECT 68.6300 167.0800 68.9000 167.9000 ;
      RECT 2.8900 167.0800 67.0300 168.1600 ;
      RECT 1.0200 167.0800 1.2900 167.9000 ;
      RECT 1.0200 166.9200 68.9000 167.0800 ;
      RECT 0.0000 166.6800 69.9200 166.9200 ;
      RECT 0.0000 166.0700 68.9000 166.6800 ;
      RECT 1.0200 165.7000 68.9000 166.0700 ;
      RECT 1.0200 165.4400 69.9200 165.7000 ;
      RECT 1.0200 165.0900 3.0900 165.4400 ;
      RECT 66.8300 164.3600 69.9200 165.4400 ;
      RECT 4.6900 164.3600 65.2300 165.4400 ;
      RECT 0.0000 164.3600 3.0900 165.0900 ;
      RECT 0.0000 164.2400 69.9200 164.3600 ;
      RECT 1.0200 163.6300 69.9200 164.2400 ;
      RECT 1.0200 163.2600 68.9000 163.6300 ;
      RECT 0.0000 162.7200 68.9000 163.2600 ;
      RECT 68.6300 162.6500 68.9000 162.7200 ;
      RECT 0.0000 162.4100 1.2900 162.7200 ;
      RECT 68.6300 161.6400 69.9200 162.6500 ;
      RECT 2.8900 161.6400 67.0300 162.7200 ;
      RECT 1.0200 161.6400 1.2900 162.4100 ;
      RECT 1.0200 161.4300 69.9200 161.6400 ;
      RECT 0.0000 160.5800 69.9200 161.4300 ;
      RECT 1.0200 160.0000 68.9000 160.5800 ;
      RECT 66.8300 159.6000 68.9000 160.0000 ;
      RECT 1.0200 159.6000 3.0900 160.0000 ;
      RECT 66.8300 158.9200 69.9200 159.6000 ;
      RECT 4.6900 158.9200 65.2300 160.0000 ;
      RECT 0.0000 158.9200 3.0900 159.6000 ;
      RECT 0.0000 158.7500 69.9200 158.9200 ;
      RECT 1.0200 157.7700 68.9000 158.7500 ;
      RECT 0.0000 157.2800 69.9200 157.7700 ;
      RECT 68.6300 156.9200 69.9200 157.2800 ;
      RECT 0.0000 156.9200 1.2900 157.2800 ;
      RECT 68.6300 156.2000 68.9000 156.9200 ;
      RECT 2.8900 156.2000 67.0300 157.2800 ;
      RECT 1.0200 156.2000 1.2900 156.9200 ;
      RECT 1.0200 155.9400 68.9000 156.2000 ;
      RECT 0.0000 155.7000 69.9200 155.9400 ;
      RECT 1.0200 154.7200 68.9000 155.7000 ;
      RECT 0.0000 154.5600 69.9200 154.7200 ;
      RECT 66.8300 153.4800 69.9200 154.5600 ;
      RECT 4.6900 153.4800 65.2300 154.5600 ;
      RECT 0.0000 153.4800 3.0900 154.5600 ;
      RECT 0.0000 151.8400 69.9200 153.4800 ;
      RECT 68.6300 150.7600 69.9200 151.8400 ;
      RECT 2.8900 150.7600 67.0300 151.8400 ;
      RECT 0.0000 150.7600 1.2900 151.8400 ;
      RECT 0.0000 149.1200 69.9200 150.7600 ;
      RECT 66.8300 148.0400 69.9200 149.1200 ;
      RECT 4.6900 148.0400 65.2300 149.1200 ;
      RECT 0.0000 148.0400 3.0900 149.1200 ;
      RECT 0.0000 146.4000 69.9200 148.0400 ;
      RECT 68.6300 145.3200 69.9200 146.4000 ;
      RECT 2.8900 145.3200 67.0300 146.4000 ;
      RECT 0.0000 145.3200 1.2900 146.4000 ;
      RECT 0.0000 143.6800 69.9200 145.3200 ;
      RECT 66.8300 142.6000 69.9200 143.6800 ;
      RECT 4.6900 142.6000 65.2300 143.6800 ;
      RECT 0.0000 142.6000 3.0900 143.6800 ;
      RECT 0.0000 140.9600 69.9200 142.6000 ;
      RECT 68.6300 139.8800 69.9200 140.9600 ;
      RECT 2.8900 139.8800 67.0300 140.9600 ;
      RECT 0.0000 139.8800 1.2900 140.9600 ;
      RECT 0.0000 138.2400 69.9200 139.8800 ;
      RECT 66.8300 137.1600 69.9200 138.2400 ;
      RECT 4.6900 137.1600 65.2300 138.2400 ;
      RECT 0.0000 137.1600 3.0900 138.2400 ;
      RECT 0.0000 135.5200 69.9200 137.1600 ;
      RECT 68.6300 134.4400 69.9200 135.5200 ;
      RECT 2.8900 134.4400 67.0300 135.5200 ;
      RECT 0.0000 134.4400 1.2900 135.5200 ;
      RECT 0.0000 132.8000 69.9200 134.4400 ;
      RECT 66.8300 131.7200 69.9200 132.8000 ;
      RECT 4.6900 131.7200 65.2300 132.8000 ;
      RECT 0.0000 131.7200 3.0900 132.8000 ;
      RECT 0.0000 130.0800 69.9200 131.7200 ;
      RECT 68.6300 129.0000 69.9200 130.0800 ;
      RECT 2.8900 129.0000 67.0300 130.0800 ;
      RECT 0.0000 129.0000 1.2900 130.0800 ;
      RECT 0.0000 127.3600 69.9200 129.0000 ;
      RECT 66.8300 126.2800 69.9200 127.3600 ;
      RECT 4.6900 126.2800 65.2300 127.3600 ;
      RECT 0.0000 126.2800 3.0900 127.3600 ;
      RECT 0.0000 124.6400 69.9200 126.2800 ;
      RECT 68.6300 123.5600 69.9200 124.6400 ;
      RECT 2.8900 123.5600 67.0300 124.6400 ;
      RECT 0.0000 123.5600 1.2900 124.6400 ;
      RECT 0.0000 121.9200 69.9200 123.5600 ;
      RECT 66.8300 120.8400 69.9200 121.9200 ;
      RECT 4.6900 120.8400 65.2300 121.9200 ;
      RECT 0.0000 120.8400 3.0900 121.9200 ;
      RECT 0.0000 119.2000 69.9200 120.8400 ;
      RECT 68.6300 118.1200 69.9200 119.2000 ;
      RECT 2.8900 118.1200 67.0300 119.2000 ;
      RECT 0.0000 118.1200 1.2900 119.2000 ;
      RECT 0.0000 116.4800 69.9200 118.1200 ;
      RECT 66.8300 115.4000 69.9200 116.4800 ;
      RECT 4.6900 115.4000 65.2300 116.4800 ;
      RECT 0.0000 115.4000 3.0900 116.4800 ;
      RECT 0.0000 113.7600 69.9200 115.4000 ;
      RECT 68.6300 112.6800 69.9200 113.7600 ;
      RECT 2.8900 112.6800 67.0300 113.7600 ;
      RECT 0.0000 112.6800 1.2900 113.7600 ;
      RECT 0.0000 111.0400 69.9200 112.6800 ;
      RECT 66.8300 109.9600 69.9200 111.0400 ;
      RECT 4.6900 109.9600 65.2300 111.0400 ;
      RECT 0.0000 109.9600 3.0900 111.0400 ;
      RECT 0.0000 108.3200 69.9200 109.9600 ;
      RECT 68.6300 107.2400 69.9200 108.3200 ;
      RECT 2.8900 107.2400 67.0300 108.3200 ;
      RECT 0.0000 107.2400 1.2900 108.3200 ;
      RECT 0.0000 105.6000 69.9200 107.2400 ;
      RECT 66.8300 104.5200 69.9200 105.6000 ;
      RECT 4.6900 104.5200 65.2300 105.6000 ;
      RECT 0.0000 104.5200 3.0900 105.6000 ;
      RECT 0.0000 102.8800 69.9200 104.5200 ;
      RECT 68.6300 101.8000 69.9200 102.8800 ;
      RECT 2.8900 101.8000 67.0300 102.8800 ;
      RECT 0.0000 101.8000 1.2900 102.8800 ;
      RECT 0.0000 100.1600 69.9200 101.8000 ;
      RECT 66.8300 99.0800 69.9200 100.1600 ;
      RECT 4.6900 99.0800 65.2300 100.1600 ;
      RECT 0.0000 99.0800 3.0900 100.1600 ;
      RECT 0.0000 97.4400 69.9200 99.0800 ;
      RECT 68.6300 96.3600 69.9200 97.4400 ;
      RECT 2.8900 96.3600 67.0300 97.4400 ;
      RECT 0.0000 96.3600 1.2900 97.4400 ;
      RECT 0.0000 94.7200 69.9200 96.3600 ;
      RECT 66.8300 93.6400 69.9200 94.7200 ;
      RECT 4.6900 93.6400 65.2300 94.7200 ;
      RECT 0.0000 93.6400 3.0900 94.7200 ;
      RECT 0.0000 92.0000 69.9200 93.6400 ;
      RECT 68.6300 90.9200 69.9200 92.0000 ;
      RECT 2.8900 90.9200 67.0300 92.0000 ;
      RECT 0.0000 90.9200 1.2900 92.0000 ;
      RECT 0.0000 89.2800 69.9200 90.9200 ;
      RECT 66.8300 88.2000 69.9200 89.2800 ;
      RECT 4.6900 88.2000 65.2300 89.2800 ;
      RECT 0.0000 88.2000 3.0900 89.2800 ;
      RECT 0.0000 86.5600 69.9200 88.2000 ;
      RECT 68.6300 85.4800 69.9200 86.5600 ;
      RECT 2.8900 85.4800 67.0300 86.5600 ;
      RECT 0.0000 85.4800 1.2900 86.5600 ;
      RECT 0.0000 83.8400 69.9200 85.4800 ;
      RECT 66.8300 82.7600 69.9200 83.8400 ;
      RECT 4.6900 82.7600 65.2300 83.8400 ;
      RECT 0.0000 82.7600 3.0900 83.8400 ;
      RECT 0.0000 81.1200 69.9200 82.7600 ;
      RECT 68.6300 80.0400 69.9200 81.1200 ;
      RECT 2.8900 80.0400 67.0300 81.1200 ;
      RECT 0.0000 80.0400 1.2900 81.1200 ;
      RECT 0.0000 78.4000 69.9200 80.0400 ;
      RECT 66.8300 77.3200 69.9200 78.4000 ;
      RECT 4.6900 77.3200 65.2300 78.4000 ;
      RECT 0.0000 77.3200 3.0900 78.4000 ;
      RECT 0.0000 75.6800 69.9200 77.3200 ;
      RECT 68.6300 74.6000 69.9200 75.6800 ;
      RECT 2.8900 74.6000 67.0300 75.6800 ;
      RECT 0.0000 74.6000 1.2900 75.6800 ;
      RECT 0.0000 72.9600 69.9200 74.6000 ;
      RECT 66.8300 71.8800 69.9200 72.9600 ;
      RECT 4.6900 71.8800 65.2300 72.9600 ;
      RECT 0.0000 71.8800 3.0900 72.9600 ;
      RECT 0.0000 70.2400 69.9200 71.8800 ;
      RECT 68.6300 69.1600 69.9200 70.2400 ;
      RECT 2.8900 69.1600 67.0300 70.2400 ;
      RECT 0.0000 69.1600 1.2900 70.2400 ;
      RECT 0.0000 67.5200 69.9200 69.1600 ;
      RECT 66.8300 66.4400 69.9200 67.5200 ;
      RECT 4.6900 66.4400 65.2300 67.5200 ;
      RECT 0.0000 66.4400 3.0900 67.5200 ;
      RECT 0.0000 64.8000 69.9200 66.4400 ;
      RECT 68.6300 63.7200 69.9200 64.8000 ;
      RECT 2.8900 63.7200 67.0300 64.8000 ;
      RECT 0.0000 63.7200 1.2900 64.8000 ;
      RECT 0.0000 62.0800 69.9200 63.7200 ;
      RECT 66.8300 61.0000 69.9200 62.0800 ;
      RECT 4.6900 61.0000 65.2300 62.0800 ;
      RECT 0.0000 61.0000 3.0900 62.0800 ;
      RECT 0.0000 59.3600 69.9200 61.0000 ;
      RECT 68.6300 58.2800 69.9200 59.3600 ;
      RECT 2.8900 58.2800 67.0300 59.3600 ;
      RECT 0.0000 58.2800 1.2900 59.3600 ;
      RECT 0.0000 56.6400 69.9200 58.2800 ;
      RECT 66.8300 55.5600 69.9200 56.6400 ;
      RECT 4.6900 55.5600 65.2300 56.6400 ;
      RECT 0.0000 55.5600 3.0900 56.6400 ;
      RECT 0.0000 53.9200 69.9200 55.5600 ;
      RECT 68.6300 52.8400 69.9200 53.9200 ;
      RECT 2.8900 52.8400 67.0300 53.9200 ;
      RECT 0.0000 52.8400 1.2900 53.9200 ;
      RECT 0.0000 51.2000 69.9200 52.8400 ;
      RECT 66.8300 50.1200 69.9200 51.2000 ;
      RECT 4.6900 50.1200 65.2300 51.2000 ;
      RECT 0.0000 50.1200 3.0900 51.2000 ;
      RECT 0.0000 48.4800 69.9200 50.1200 ;
      RECT 68.6300 47.4000 69.9200 48.4800 ;
      RECT 2.8900 47.4000 67.0300 48.4800 ;
      RECT 0.0000 47.4000 1.2900 48.4800 ;
      RECT 0.0000 45.7600 69.9200 47.4000 ;
      RECT 66.8300 44.6800 69.9200 45.7600 ;
      RECT 4.6900 44.6800 65.2300 45.7600 ;
      RECT 0.0000 44.6800 3.0900 45.7600 ;
      RECT 0.0000 43.0400 69.9200 44.6800 ;
      RECT 68.6300 41.9600 69.9200 43.0400 ;
      RECT 2.8900 41.9600 67.0300 43.0400 ;
      RECT 0.0000 41.9600 1.2900 43.0400 ;
      RECT 0.0000 40.3200 69.9200 41.9600 ;
      RECT 66.8300 39.2400 69.9200 40.3200 ;
      RECT 4.6900 39.2400 65.2300 40.3200 ;
      RECT 0.0000 39.2400 3.0900 40.3200 ;
      RECT 0.0000 37.6000 69.9200 39.2400 ;
      RECT 68.6300 36.5200 69.9200 37.6000 ;
      RECT 2.8900 36.5200 67.0300 37.6000 ;
      RECT 0.0000 36.5200 1.2900 37.6000 ;
      RECT 0.0000 34.8800 69.9200 36.5200 ;
      RECT 66.8300 33.8000 69.9200 34.8800 ;
      RECT 4.6900 33.8000 65.2300 34.8800 ;
      RECT 0.0000 33.8000 3.0900 34.8800 ;
      RECT 0.0000 32.1600 69.9200 33.8000 ;
      RECT 68.6300 31.0800 69.9200 32.1600 ;
      RECT 2.8900 31.0800 67.0300 32.1600 ;
      RECT 0.0000 31.0800 1.2900 32.1600 ;
      RECT 0.0000 29.4400 69.9200 31.0800 ;
      RECT 66.8300 28.3600 69.9200 29.4400 ;
      RECT 4.6900 28.3600 65.2300 29.4400 ;
      RECT 0.0000 28.3600 3.0900 29.4400 ;
      RECT 0.0000 26.7200 69.9200 28.3600 ;
      RECT 68.6300 25.6400 69.9200 26.7200 ;
      RECT 2.8900 25.6400 67.0300 26.7200 ;
      RECT 0.0000 25.6400 1.2900 26.7200 ;
      RECT 0.0000 24.0000 69.9200 25.6400 ;
      RECT 66.8300 22.9200 69.9200 24.0000 ;
      RECT 4.6900 22.9200 65.2300 24.0000 ;
      RECT 0.0000 22.9200 3.0900 24.0000 ;
      RECT 0.0000 21.2800 69.9200 22.9200 ;
      RECT 68.6300 20.2000 69.9200 21.2800 ;
      RECT 2.8900 20.2000 67.0300 21.2800 ;
      RECT 0.0000 20.2000 1.2900 21.2800 ;
      RECT 0.0000 18.5600 69.9200 20.2000 ;
      RECT 66.8300 17.4800 69.9200 18.5600 ;
      RECT 4.6900 17.4800 65.2300 18.5600 ;
      RECT 0.0000 17.4800 3.0900 18.5600 ;
      RECT 0.0000 15.8400 69.9200 17.4800 ;
      RECT 68.6300 14.7600 69.9200 15.8400 ;
      RECT 2.8900 14.7600 67.0300 15.8400 ;
      RECT 0.0000 14.7600 1.2900 15.8400 ;
      RECT 0.0000 13.1200 69.9200 14.7600 ;
      RECT 66.8300 12.0400 69.9200 13.1200 ;
      RECT 4.6900 12.0400 65.2300 13.1200 ;
      RECT 0.0000 12.0400 3.0900 13.1200 ;
      RECT 0.0000 10.4000 69.9200 12.0400 ;
      RECT 68.6300 9.3200 69.9200 10.4000 ;
      RECT 2.8900 9.3200 67.0300 10.4000 ;
      RECT 0.0000 9.3200 1.2900 10.4000 ;
      RECT 0.0000 6.6300 69.9200 9.3200 ;
      RECT 66.8300 5.0300 69.9200 6.6300 ;
      RECT 0.0000 5.0300 3.0900 6.6300 ;
      RECT 0.0000 4.8300 69.9200 5.0300 ;
      RECT 68.6300 3.2300 69.9200 4.8300 ;
      RECT 0.0000 3.2300 1.2900 4.8300 ;
      RECT 0.0000 0.0000 69.9200 3.2300 ;
    LAYER met4 ;
      RECT 0.0000 215.7300 69.9200 219.6400 ;
      RECT 2.8900 213.9300 67.0300 215.7300 ;
      RECT 66.8300 5.0300 67.0300 213.9300 ;
      RECT 4.6900 5.0300 65.2300 213.9300 ;
      RECT 2.8900 5.0300 3.0900 213.9300 ;
      RECT 68.6300 3.2300 69.9200 215.7300 ;
      RECT 2.8900 3.2300 67.0300 5.0300 ;
      RECT 0.0000 3.2300 1.2900 215.7300 ;
      RECT 0.0000 0.0000 69.9200 3.2300 ;
  END
END W_IO

END LIBRARY
