* NGSPICE file created from spi_to_wbs.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

.subckt spi_to_wbs spi_cs_n spi_miso spi_mosi spi_sck vccd1 vssd1 wbs_adr_o[0] wbs_adr_o[10]
+ wbs_adr_o[11] wbs_adr_o[12] wbs_adr_o[13] wbs_adr_o[14] wbs_adr_o[15] wbs_adr_o[16]
+ wbs_adr_o[17] wbs_adr_o[18] wbs_adr_o[19] wbs_adr_o[1] wbs_adr_o[20] wbs_adr_o[21]
+ wbs_adr_o[22] wbs_adr_o[23] wbs_adr_o[24] wbs_adr_o[25] wbs_adr_o[26] wbs_adr_o[27]
+ wbs_adr_o[28] wbs_adr_o[29] wbs_adr_o[2] wbs_adr_o[30] wbs_adr_o[31] wbs_adr_o[3]
+ wbs_adr_o[4] wbs_adr_o[5] wbs_adr_o[6] wbs_adr_o[7] wbs_adr_o[8] wbs_adr_o[9] wbs_cyc_o
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_o wbs_we_o
XTAP_TAPCELL_ROW_32_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0985_ clknet_4_1_0_spi_sck _0040_ vssd1 vssd1 vccd1 vccd1 data_out\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ _0390_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_11_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0968_ clknet_4_3_0_spi_sck _0023_ vssd1 vssd1 vccd1 vccd1 shift_out\[3\] sky130_fd_sc_hd__dfxtp_2
X_0899_ wbs_dat_o[30] data_in\[30\] _0443_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__mux2_2
X_0753_ addr\[30\] addr\[14\] _0216_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Left_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0822_ _0412_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__buf_1
X_0684_ _0335_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__buf_1
X_1098_ clknet_4_14_0_spi_sck _0153_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0736_ _0368_ wbs_adr_o[8] _0356_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0805_ _0403_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__buf_1
X_1021_ clknet_4_15_0_spi_sck _0076_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[0] sky130_fd_sc_hd__dfxtp_2
X_0667_ _0326_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__buf_1
XFILLER_0_24_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0598_ _0252_ _0253_ _0286_ _0287_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__or4_2
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0521_ addr\[30\] _0223_ _0227_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__mux2_2
X_1004_ clknet_4_4_0_spi_sck _0059_ vssd1 vssd1 vccd1 vccd1 addr\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0719_ _0357_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__buf_1
XFILLER_0_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0504_ state\[2\] state\[1\] state\[0\] state\[3\] vssd1 vssd1 vccd1 vccd1 _0215_
+ sky130_fd_sc_hd__and4bb_2
XTAP_TAPCELL_ROW_23_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0984_ clknet_4_2_0_spi_sck _0039_ vssd1 vssd1 vccd1 vccd1 data_out\[19\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_37_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0898_ _0451_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__buf_1
X_0967_ clknet_4_2_0_spi_sck _0022_ vssd1 vssd1 vccd1 vccd1 shift_out\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0752_ _0379_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0821_ _0236_ data_in\[10\] _0409_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1097_ clknet_4_11_0_spi_sck _0152_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__dfxtp_2
X_0683_ _0242_ data_in\[5\] _0329_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__mux2_2
XFILLER_0_10_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0735_ addr\[24\] addr\[8\] _0348_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__mux2_2
X_0666_ addr\[13\] _0242_ _0320_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__mux2_2
X_0804_ addr\[2\] _0236_ _0400_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__mux2_2
X_1020_ clknet_4_14_0_spi_sck _0075_ vssd1 vssd1 vccd1 vccd1 addr\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0597_ data_out\[23\] _0194_ _0247_ wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__a22o_2
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1003_ clknet_4_4_0_spi_sck _0058_ vssd1 vssd1 vccd1 vccd1 addr\[14\] sky130_fd_sc_hd__dfxtp_2
X_0520_ _0226_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0718_ _0355_ wbs_adr_o[2] _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__mux2_2
X_0649_ wbs_dat_i[30] data_out\[30\] _0291_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0503_ bit_count\[1\] bit_count\[0\] bit_count\[2\] vssd1 vssd1 vccd1 vccd1 _0214_
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_14_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ clknet_4_2_0_spi_sck _0038_ vssd1 vssd1 vccd1 vccd1 data_out\[18\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_3_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0897_ wbs_dat_o[29] data_in\[29\] _0443_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0966_ clknet_4_2_0_spi_sck _0021_ vssd1 vssd1 vccd1 vccd1 shift_out\[1\] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_1_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0751_ _0378_ wbs_adr_o[13] _0350_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1096_ clknet_4_9_0_spi_sck _0151_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__dfxtp_2
X_0682_ _0334_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0820_ _0411_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__buf_1
X_0949_ _0474_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__buf_1
X_0665_ _0325_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__buf_1
XFILLER_0_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0803_ _0402_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__buf_1
X_0734_ _0367_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__buf_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1079_ clknet_4_15_0_spi_sck _0134_ vssd1 vssd1 vccd1 vccd1 wbs_we_o sky130_fd_sc_hd__dfxtp_2
XFILLER_0_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0596_ data_out\[31\] _0198_ _0249_ data_out\[15\] vssd1 vssd1 vccd1 vccd1 _0286_
+ sky130_fd_sc_hd__a22o_2
Xhold10 addr\[20\] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__dlygate4sd3_1
X_0717_ _0350_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__clkbuf_4
X_1002_ clknet_4_5_0_spi_sck _0057_ vssd1 vssd1 vccd1 vccd1 addr\[13\] sky130_fd_sc_hd__dfxtp_2
X_0648_ _0315_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__buf_1
X_0579_ data_out\[28\] _0198_ _0249_ data_out\[12\] vssd1 vssd1 vccd1 vccd1 _0272_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0502_ _0196_ _0202_ _0213_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0982_ clknet_4_0_0_spi_sck _0037_ vssd1 vssd1 vccd1 vccd1 data_out\[17\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_37_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0965_ clknet_4_10_0_spi_sck _0020_ vssd1 vssd1 vccd1 vccd1 data_in\[31\] sky130_fd_sc_hd__dfxtp_2
X_0896_ _0450_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__buf_1
XFILLER_0_37_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_5_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0750_ addr\[29\] addr\[13\] _0216_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1095_ clknet_4_11_0_spi_sck _0150_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_0_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0681_ _0240_ data_in\[4\] _0329_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__mux2_2
X_0948_ addr\[26\] shift_in\[1\] _0227_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__mux2_2
XFILLER_0_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0879_ _0441_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__buf_1
XFILLER_0_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0802_ addr\[1\] _0234_ _0400_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0664_ addr\[12\] _0240_ _0320_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__mux2_2
X_0733_ _0366_ wbs_adr_o[7] _0356_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1078_ clknet_4_1_0_spi_sck _0133_ _0003_ vssd1 vssd1 vccd1 vccd1 wbs_cyc_o sky130_fd_sc_hd__dfrtp_2
X_0595_ _0246_ _0250_ shift_out\[6\] vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__a21o_2
Xhold11 addr\[19\] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__dlygate4sd3_1
X_1001_ clknet_4_5_0_spi_sck _0056_ vssd1 vssd1 vccd1 vccd1 addr\[12\] sky130_fd_sc_hd__dfxtp_2
X_0716_ shift_in\[1\] addr\[2\] _0348_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0647_ wbs_dat_i[29] data_out\[29\] _0291_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0578_ data_out\[20\] _0194_ _0247_ wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__a22o_2
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0501_ _0202_ _0210_ _0196_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_17_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0981_ clknet_4_0_0_spi_sck _0036_ vssd1 vssd1 vccd1 vccd1 data_out\[16\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_37_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0895_ wbs_dat_o[28] data_in\[28\] _0443_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__mux2_2
X_0964_ clknet_4_10_0_spi_sck _0019_ vssd1 vssd1 vccd1 vccd1 data_in\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
X_0680_ _0333_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0947_ _0473_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__buf_1
X_0878_ wbs_dat_o[20] data_in\[20\] _0432_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__mux2_2
X_1094_ clknet_4_11_0_spi_sck _0149_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0663_ _0324_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__buf_1
X_0801_ _0401_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__buf_1
X_0732_ shift_in\[6\] addr\[7\] _0348_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1077_ clknet_4_3_0_spi_sck _0132_ vssd1 vssd1 vccd1 vccd1 spi_miso sky130_fd_sc_hd__dfxtp_2
X_0594_ _0003_ _0280_ _0283_ _0284_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__a31o_2
Xhold12 addr\[23\] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dlygate4sd3_1
X_1000_ clknet_4_7_0_spi_sck _0055_ vssd1 vssd1 vccd1 vccd1 addr\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0715_ _0354_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1129_ clknet_4_9_0_spi_sck _0181_ vssd1 vssd1 vccd1 vccd1 command\[2\] sky130_fd_sc_hd__dfxtp_2
X_0646_ _0314_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__buf_1
X_0577_ _0246_ _0250_ shift_out\[3\] vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0500_ _0212_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0629_ wbs_dat_i[20] data_out\[20\] _0303_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_37_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0980_ clknet_4_0_0_spi_sck _0035_ vssd1 vssd1 vccd1 vccd1 data_out\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_24_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0894_ _0449_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__buf_1
X_0963_ clknet_4_10_0_spi_sck _0018_ vssd1 vssd1 vccd1 vccd1 data_in\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0946_ addr\[25\] shift_in\[0\] _0227_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__mux2_2
X_0877_ _0440_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__buf_1
XFILLER_0_19_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1093_ clknet_4_11_0_spi_sck _0148_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0662_ addr\[11\] _0238_ _0320_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__mux2_2
X_0800_ addr\[0\] _0231_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__mux2_2
X_0731_ _0365_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__buf_1
X_0593_ _0263_ shift_out\[6\] vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__and2_2
XFILLER_0_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold13 addr\[28\] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__dlygate4sd3_1
X_0929_ _0464_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__buf_1
X_1076_ clknet_4_11_0_spi_sck _0131_ vssd1 vssd1 vccd1 vccd1 data_in\[15\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_29_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1059_ clknet_4_6_0_spi_sck _0114_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[30] sky130_fd_sc_hd__dfxtp_2
X_0714_ _0353_ wbs_adr_o[1] _0351_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1128_ clknet_4_9_0_spi_sck _0180_ vssd1 vssd1 vccd1 vccd1 command\[1\] sky130_fd_sc_hd__dfxtp_2
X_0576_ _0257_ _0267_ _0268_ _0269_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__o31a_2
X_0645_ wbs_dat_i[28] data_out\[28\] _0291_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__mux2_2
X_0628_ _0305_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__buf_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0559_ data_out\[17\] _0194_ _0247_ wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_8_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0962_ clknet_4_9_0_spi_sck _0017_ vssd1 vssd1 vccd1 vccd1 data_in\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0893_ wbs_dat_o[27] data_in\[27\] _0443_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0945_ _0472_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__buf_1
X_0876_ wbs_dat_o[19] data_in\[19\] _0432_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1092_ clknet_4_9_0_spi_sck _0147_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0661_ _0323_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__buf_1
X_0730_ _0364_ wbs_adr_o[6] _0356_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__mux2_2
X_0592_ _0252_ _0253_ _0281_ _0282_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__or4_2
Xhold14 addr\[26\] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1075_ clknet_4_11_0_spi_sck _0130_ vssd1 vssd1 vccd1 vccd1 data_in\[14\] sky130_fd_sc_hd__dfxtp_2
X_0928_ command\[0\] _0231_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__mux2_2
X_0859_ wbs_dat_o[11] data_in\[11\] _0421_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1058_ clknet_4_7_0_spi_sck _0113_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[29] sky130_fd_sc_hd__dfxtp_2
X_0713_ shift_in\[0\] addr\[1\] _0348_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__mux2_2
X_1127_ clknet_4_9_0_spi_sck _0179_ vssd1 vssd1 vccd1 vccd1 command\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0644_ _0313_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__buf_1
X_0575_ _0003_ shift_out\[3\] vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0489_ _0203_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__buf_1
X_0558_ data_out\[25\] _0198_ _0249_ data_out\[9\] vssd1 vssd1 vccd1 vccd1 _0254_
+ sky130_fd_sc_hd__a22o_2
X_0627_ wbs_dat_i[19] data_out\[19\] _0303_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0961_ clknet_4_10_0_spi_sck _0016_ vssd1 vssd1 vccd1 vccd1 data_in\[27\] sky130_fd_sc_hd__dfxtp_2
X_0892_ _0448_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__buf_1
X_0944_ addr\[24\] _0231_ _0227_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__mux2_2
XFILLER_0_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1091_ clknet_4_8_0_spi_sck _0146_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_15_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0875_ _0439_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__buf_1
X_0660_ addr\[10\] _0236_ _0320_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__mux2_2
X_0591_ wbs_dat_i[6] _0247_ _0249_ data_out\[14\] vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a22o_2
XFILLER_0_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0789_ wbs_adr_o[23] _0394_ _0398_ net13 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__a22o_2
X_0927_ _0205_ _0318_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__nor2b_2
X_1074_ clknet_4_11_0_spi_sck _0129_ vssd1 vssd1 vccd1 vccd1 data_in\[13\] sky130_fd_sc_hd__dfxtp_2
X_0858_ _0430_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__buf_1
Xhold15 addr\[25\] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Left_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0712_ _0352_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__buf_1
X_1126_ clknet_4_4_0_spi_sck _0178_ _0010_ vssd1 vssd1 vccd1 vccd1 state\[3\] sky130_fd_sc_hd__dfrtp_2
X_0643_ wbs_dat_i[27] data_out\[27\] _0303_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__mux2_2
X_0574_ _0252_ _0253_ shift_out\[2\] vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__o21a_2
X_1057_ clknet_4_5_0_spi_sck _0112_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[28] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0488_ state\[3\] _0199_ _0202_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0557_ _0193_ net1 _0247_ _0248_ _0214_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__o41ai_4
X_0626_ _0304_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__buf_1
XFILLER_0_4_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1109_ clknet_4_10_0_spi_sck _0164_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_36_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0609_ _0295_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_20_Left_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0960_ clknet_4_10_0_spi_sck _0015_ vssd1 vssd1 vccd1 vccd1 data_in\[26\] sky130_fd_sc_hd__dfxtp_2
X_0891_ wbs_dat_o[26] data_in\[26\] _0443_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1090_ clknet_4_8_0_spi_sck _0145_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0874_ wbs_dat_o[18] data_in\[18\] _0432_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__mux2_2
X_0943_ _0471_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__buf_1
XFILLER_0_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_spi_sck spi_sck vssd1 vssd1 vccd1 vccd1 clknet_0_spi_sck sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_23_Left_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0926_ _0257_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__inv_2
X_0590_ data_out\[22\] _0193_ _0198_ data_out\[30\] vssd1 vssd1 vccd1 vccd1 _0281_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1073_ clknet_4_9_0_spi_sck _0128_ vssd1 vssd1 vccd1 vccd1 data_in\[12\] sky130_fd_sc_hd__dfxtp_2
X_0857_ wbs_dat_o[10] data_in\[10\] _0421_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold16 addr\[31\] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ wbs_adr_o[22] _0394_ _0398_ net5 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__a22o_2
XFILLER_0_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0711_ _0349_ wbs_adr_o[0] _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0642_ _0312_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__buf_1
X_0573_ _0265_ _0266_ _0246_ _0250_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__o211a_2
X_1056_ clknet_4_7_0_spi_sck _0111_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[27] sky130_fd_sc_hd__dfxtp_2
X_0909_ _0231_ _0234_ _0263_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__mux2_2
X_1125_ clknet_4_6_0_spi_sck _0177_ _0009_ vssd1 vssd1 vccd1 vccd1 state\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0487_ _0200_ _0201_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__nor2_2
X_1039_ clknet_4_14_0_spi_sck _0094_ vssd1 vssd1 vccd1 vccd1 data_in\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0556_ _0207_ _0208_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__or2_2
X_1108_ clknet_4_11_0_spi_sck _0163_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__dfxtp_2
X_0625_ wbs_dat_i[18] data_out\[18\] _0303_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0539_ shift_in\[3\] vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__buf_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0608_ wbs_dat_i[10] data_out\[10\] _0292_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__mux2_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0890_ _0447_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__buf_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0942_ command\[7\] _0229_ _0463_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__mux2_2
X_0873_ _0438_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__buf_1
XFILLER_0_2_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1141_ wbs_cyc_o vssd1 vssd1 vccd1 vccd1 wbs_stb_o sky130_fd_sc_hd__buf_2
X_1072_ clknet_4_8_0_spi_sck _0127_ vssd1 vssd1 vccd1 vccd1 data_in\[11\] sky130_fd_sc_hd__dfxtp_2
Xhold17 addr\[27\] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__dlygate4sd3_1
X_0787_ wbs_adr_o[21] _0394_ _0398_ net8 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__a22o_2
X_0925_ _0257_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0856_ _0429_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__buf_1
X_0710_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__clkbuf_4
X_0641_ wbs_dat_i[26] data_out\[26\] _0303_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__mux2_2
X_1055_ clknet_4_13_0_spi_sck _0110_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[26] sky130_fd_sc_hd__dfxtp_2
X_1124_ clknet_4_6_0_spi_sck _0176_ _0008_ vssd1 vssd1 vccd1 vccd1 state\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0908_ _0257_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__inv_2
X_0839_ _0420_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__buf_1
X_0572_ data_out\[27\] _0198_ _0249_ data_out\[11\] vssd1 vssd1 vccd1 vccd1 _0266_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0486_ state\[2\] _0195_ state\[3\] vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__o21a_2
X_0624_ _0291_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_4
X_0555_ _0246_ _0250_ shift_out\[0\] vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__a21o_2
X_1038_ clknet_4_11_0_spi_sck _0093_ vssd1 vssd1 vccd1 vccd1 data_in\[17\] sky130_fd_sc_hd__dfxtp_2
X_1107_ clknet_4_10_0_spi_sck _0162_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0607_ _0294_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__buf_1
X_0538_ _0239_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__buf_1
XFILLER_0_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0941_ _0470_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__buf_1
X_0872_ wbs_dat_o[17] data_in\[17\] _0432_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_0_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1140_ clknet_4_5_0_spi_sck _0192_ vssd1 vssd1 vccd1 vccd1 addr\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1071_ clknet_4_8_0_spi_sck _0126_ vssd1 vssd1 vccd1 vccd1 data_in\[10\] sky130_fd_sc_hd__dfxtp_2
X_0786_ wbs_adr_o[20] _0394_ _0398_ net11 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__a22o_2
X_0924_ _0257_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0855_ wbs_dat_o[9] data_in\[9\] _0421_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__mux2_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1054_ clknet_4_12_0_spi_sck _0109_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[25] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0907_ _0257_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__inv_2
X_1123_ clknet_4_3_0_spi_sck _0175_ _0007_ vssd1 vssd1 vccd1 vccd1 state\[0\] sky130_fd_sc_hd__dfrtp_2
X_0640_ _0311_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__buf_1
X_0571_ data_out\[19\] _0194_ _0247_ wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__a22o_2
X_0769_ data_in\[20\] _0240_ _0385_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__mux2_2
X_0838_ wbs_dat_o[1] data_in\[1\] _0397_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__mux2_2
X_0554_ _0194_ _0198_ _0247_ _0249_ _0214_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__o41a_2
X_0623_ _0302_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__buf_1
X_0485_ bit_count\[1\] bit_count\[0\] bit_count\[2\] vssd1 vssd1 vccd1 vccd1 _0200_
+ sky130_fd_sc_hd__nand3_2
X_1037_ clknet_4_12_0_spi_sck _0092_ vssd1 vssd1 vccd1 vccd1 data_in\[16\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1106_ clknet_4_10_0_spi_sck _0161_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_37_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_0_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0537_ _0238_ data_in\[27\] _0232_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__mux2_2
X_0606_ wbs_dat_i[9] data_out\[9\] _0292_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0940_ command\[6\] shift_in\[5\] _0463_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__mux2_2
X_0871_ _0437_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0785_ wbs_adr_o[19] _0394_ _0398_ net12 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__a22o_2
X_0923_ _0257_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1070_ clknet_4_8_0_spi_sck _0125_ vssd1 vssd1 vccd1 vccd1 data_in\[9\] sky130_fd_sc_hd__dfxtp_2
X_0854_ _0428_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__buf_1
X_1053_ clknet_4_15_0_spi_sck _0108_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[24] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_27_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1122_ clknet_4_6_0_spi_sck _0174_ vssd1 vssd1 vccd1 vccd1 shift_in\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0570_ _0003_ _0259_ _0262_ _0264_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__a31o_2
X_0699_ addr\[20\] _0240_ _0339_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__mux2_2
X_0906_ _0257_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__inv_2
X_0768_ _0389_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__buf_1
X_0837_ _0419_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__buf_1
XFILLER_0_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1036_ clknet_4_4_0_spi_sck _0091_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[15] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0484_ _0194_ _0198_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__or2_2
X_0553_ _0248_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_4
X_0622_ wbs_dat_i[17] data_out\[17\] _0292_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__mux2_2
X_1105_ clknet_4_10_0_spi_sck _0160_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_14_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ shift_in\[2\] vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0605_ _0293_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__buf_1
X_1019_ clknet_4_14_0_spi_sck _0074_ vssd1 vssd1 vccd1 vccd1 addr\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Left_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0519_ _0209_ _0225_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__and2_2
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0870_ wbs_dat_o[16] data_in\[16\] _0432_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_0_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0999_ clknet_4_13_0_spi_sck _0054_ vssd1 vssd1 vccd1 vccd1 addr\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0784_ wbs_adr_o[18] _0394_ _0398_ net10 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__a22o_2
X_0922_ _0462_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__buf_1
X_0853_ wbs_dat_o[8] data_in\[8\] _0421_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1052_ clknet_4_14_0_spi_sck _0107_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[23] sky130_fd_sc_hd__dfxtp_2
X_1121_ clknet_4_6_0_spi_sck _0173_ vssd1 vssd1 vccd1 vccd1 shift_in\[5\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_2_Left_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0698_ _0343_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__buf_1
X_0767_ data_in\[19\] _0238_ _0385_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__mux2_2
X_0836_ wbs_dat_o[0] data_in\[0\] _0397_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0905_ _0246_ _0225_ _0455_ net3 _0257_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__a32o_2
XFILLER_0_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1035_ clknet_4_5_0_spi_sck _0090_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[14] sky130_fd_sc_hd__dfxtp_2
X_0552_ state\[3\] _0196_ _0195_ state\[2\] vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__and4bb_2
X_0483_ net1 vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_4
X_0621_ _0301_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__buf_1
X_1104_ clknet_4_10_0_spi_sck _0159_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0819_ _0234_ data_in\[9\] _0409_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0604_ wbs_dat_i[8] data_out\[8\] _0292_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__mux2_2
Xclkbuf_4_8_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1018_ clknet_4_15_0_spi_sck _0073_ vssd1 vssd1 vccd1 vccd1 addr\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0535_ _0237_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__buf_1
X_0518_ _0224_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__buf_1
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0998_ clknet_4_12_0_spi_sck _0053_ vssd1 vssd1 vccd1 vccd1 addr\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0783_ wbs_adr_o[17] _0394_ _0398_ net6 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__a22o_2
X_0921_ _0223_ _0229_ spi_cs_n vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0852_ _0427_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__buf_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0697_ addr\[19\] _0238_ _0339_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__mux2_2
X_0835_ wbs_we_o _0394_ _0398_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__a21o_2
X_1120_ clknet_4_7_0_spi_sck _0172_ vssd1 vssd1 vccd1 vccd1 shift_in\[4\] sky130_fd_sc_hd__dfxtp_2
X_1051_ clknet_4_15_0_spi_sck _0106_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[22] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_28_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0766_ _0388_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__buf_1
X_0904_ wbs_dat_i[0] _0247_ _0249_ data_out\[8\] _0454_ vssd1 vssd1 vccd1 vccd1 _0455_
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_34_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1034_ clknet_4_5_0_spi_sck _0089_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[13] sky130_fd_sc_hd__dfxtp_2
X_0482_ state\[2\] _0195_ _0196_ state\[3\] vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__nor4b_1
XTAP_TAPCELL_ROW_17_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0551_ _0209_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_4
X_1103_ clknet_4_11_0_spi_sck _0158_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__dfxtp_2
X_0620_ wbs_dat_i[16] data_out\[16\] _0292_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__mux2_2
X_0749_ _0377_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0818_ _0410_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__buf_1
X_1017_ clknet_4_13_0_spi_sck _0072_ vssd1 vssd1 vccd1 vccd1 addr\[20\] sky130_fd_sc_hd__dfxtp_2
X_0603_ _0291_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0534_ _0236_ data_in\[26\] _0232_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__mux2_2
X_0517_ spi_cs_n bit_count\[2\] bit_count\[0\] bit_count\[1\] vssd1 vssd1 vccd1 vccd1
+ _0224_ sky130_fd_sc_hd__and4b_2
X_0997_ clknet_4_13_0_spi_sck _0052_ vssd1 vssd1 vccd1 vccd1 addr\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0920_ _0461_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__buf_1
X_0782_ wbs_adr_o[16] _0394_ _0398_ net7 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0851_ wbs_dat_o[7] data_in\[7\] _0421_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0696_ _0342_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__buf_1
X_1050_ clknet_4_15_0_spi_sck _0105_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[21] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0765_ data_in\[18\] _0236_ _0385_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0834_ _0418_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__buf_1
X_0903_ data_out\[16\] _0194_ _0198_ data_out\[24\] vssd1 vssd1 vccd1 vccd1 _0454_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0481_ state\[0\] vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__buf_1
X_0550_ _0207_ _0208_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__nor2_2
X_1102_ clknet_4_11_0_spi_sck _0157_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__dfxtp_2
X_0748_ _0376_ wbs_adr_o[12] _0350_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__mux2_2
X_1033_ clknet_4_5_0_spi_sck _0088_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[12] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0817_ _0231_ data_in\[8\] _0409_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__mux2_2
X_0679_ _0238_ data_in\[3\] _0329_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_8_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1016_ clknet_4_15_0_spi_sck _0071_ vssd1 vssd1 vccd1 vccd1 addr\[19\] sky130_fd_sc_hd__dfxtp_2
X_0533_ shift_in\[1\] vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0602_ _0290_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__buf_1
Xclkbuf_4_10_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
X_0516_ shift_in\[5\] vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_18_Left_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0996_ clknet_4_0_0_spi_sck _0051_ vssd1 vssd1 vccd1 vccd1 data_out\[31\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0781_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__buf_1
XFILLER_0_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0850_ _0426_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__buf_1
XFILLER_0_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0979_ clknet_4_1_0_spi_sck _0034_ vssd1 vssd1 vccd1 vccd1 data_out\[14\] sky130_fd_sc_hd__dfxtp_2
X_0902_ _0453_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__buf_1
X_0833_ shift_out\[7\] spi_miso _0263_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__mux2_2
X_0695_ addr\[18\] _0236_ _0339_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__mux2_2
X_0764_ _0387_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__buf_1
X_0480_ state\[1\] vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1032_ clknet_4_7_0_spi_sck _0087_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[11] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0747_ addr\[28\] addr\[12\] _0216_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1101_ clknet_4_14_0_spi_sck _0156_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__dfxtp_2
X_0816_ _0194_ _0225_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__nand2_2
X_0678_ _0332_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1015_ clknet_4_15_0_spi_sck _0070_ vssd1 vssd1 vccd1 vccd1 addr\[18\] sky130_fd_sc_hd__dfxtp_2
X_0601_ spi_cs_n _0200_ _0210_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__or3_2
X_0532_ _0235_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__buf_1
Xclkbuf_4_14_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0515_ _0214_ _0222_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_35_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0995_ clknet_4_1_0_spi_sck _0050_ vssd1 vssd1 vccd1 vccd1 data_out\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0780_ _0396_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__clkbuf_4
X_0978_ clknet_4_1_0_spi_sck _0033_ vssd1 vssd1 vccd1 vccd1 data_out\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0694_ _0341_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_22_Left_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0763_ data_in\[17\] _0234_ _0385_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__mux2_2
X_0832_ _0417_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__buf_1
X_0901_ wbs_dat_o[31] data_in\[31\] _0443_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__mux2_2
X_0746_ _0375_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__buf_1
X_1031_ clknet_4_7_0_spi_sck _0086_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[10] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_31_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0815_ _0408_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__buf_1
X_1100_ clknet_4_14_0_spi_sck _0155_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0677_ _0236_ data_in\[2\] _0329_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__mux2_2
X_0600_ _0003_ _0285_ _0288_ _0289_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__a31o_2
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0531_ _0234_ data_in\[25\] _0232_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__mux2_2
X_1014_ clknet_4_14_0_spi_sck _0069_ vssd1 vssd1 vccd1 vccd1 addr\[17\] sky130_fd_sc_hd__dfxtp_2
X_0729_ shift_in\[5\] addr\[6\] _0348_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_10_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0514_ bit_count\[1\] bit_count\[0\] bit_count\[2\] vssd1 vssd1 vccd1 vccd1 _0222_
+ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_4_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0994_ clknet_4_1_0_spi_sck _0049_ vssd1 vssd1 vccd1 vccd1 data_out\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0977_ clknet_4_1_0_spi_sck _0032_ vssd1 vssd1 vccd1 vccd1 data_out\[12\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0693_ addr\[17\] _0234_ _0339_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0762_ _0386_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__buf_1
X_0831_ _0229_ data_in\[15\] _0409_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__mux2_2
X_0900_ _0452_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_34_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ clknet_4_12_0_spi_sck _0085_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[9] sky130_fd_sc_hd__dfxtp_2
X_0814_ addr\[7\] _0229_ _0400_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__mux2_2
X_0745_ _0374_ wbs_adr_o[11] _0356_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0676_ _0331_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__buf_1
X_0530_ shift_in\[0\] vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_36_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1013_ clknet_4_15_0_spi_sck _0068_ vssd1 vssd1 vccd1 vccd1 addr\[16\] sky130_fd_sc_hd__dfxtp_2
X_0728_ _0363_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__buf_1
X_0659_ _0322_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__buf_1
XFILLER_0_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0513_ bit_count\[1\] bit_count\[0\] vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_4_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0993_ clknet_4_1_0_spi_sck _0048_ vssd1 vssd1 vccd1 vccd1 data_out\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0976_ clknet_4_2_0_spi_sck _0031_ vssd1 vssd1 vccd1 vccd1 data_out\[11\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_1_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0692_ _0340_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__buf_1
X_0761_ data_in\[16\] _0231_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__mux2_2
X_0830_ _0416_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_34_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0959_ clknet_4_10_0_spi_sck _0014_ vssd1 vssd1 vccd1 vccd1 data_in\[25\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0744_ addr\[27\] addr\[11\] _0216_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__mux2_2
X_0813_ _0407_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_22_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0675_ _0234_ data_in\[1\] _0329_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__mux2_2
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1089_ clknet_4_8_0_spi_sck _0144_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0727_ _0362_ wbs_adr_o[5] _0356_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1012_ clknet_4_8_0_spi_sck _0067_ vssd1 vssd1 vccd1 vccd1 data_in\[7\] sky130_fd_sc_hd__dfxtp_2
X_0658_ addr\[9\] _0234_ _0320_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__mux2_2
X_0589_ _0246_ _0250_ shift_out\[5\] vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_10_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0512_ bit_count\[0\] vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0992_ clknet_4_2_0_spi_sck _0047_ vssd1 vssd1 vccd1 vccd1 data_out\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ clknet_4_2_0_spi_sck _0030_ vssd1 vssd1 vccd1 vccd1 data_out\[10\] sky130_fd_sc_hd__dfxtp_2
X_0691_ addr\[16\] _0231_ _0339_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__mux2_2
X_0760_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__buf_1
XFILLER_0_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0958_ clknet_4_11_0_spi_sck _0013_ vssd1 vssd1 vccd1 vccd1 data_in\[24\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0889_ wbs_dat_o[25] data_in\[25\] _0443_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_25_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0743_ _0373_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__buf_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0812_ addr\[6\] _0223_ _0400_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_26_Left_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0674_ _0330_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__buf_1
XFILLER_0_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1088_ clknet_4_8_0_spi_sck _0143_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_36_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ clknet_4_8_0_spi_sck _0066_ vssd1 vssd1 vccd1 vccd1 data_in\[6\] sky130_fd_sc_hd__dfxtp_2
X_0657_ _0321_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__buf_1
X_0726_ shift_in\[4\] addr\[5\] _0348_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__mux2_2
X_0588_ _0003_ _0275_ _0278_ _0279_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a31o_2
X_0511_ _0214_ _0221_ wbs_cyc_o vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_4_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0709_ _0210_ _0217_ _0220_ _0200_ spi_cs_n vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__a2111o_2
XPHY_EDGE_ROW_13_Left_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0991_ clknet_4_2_0_spi_sck _0046_ vssd1 vssd1 vccd1 vccd1 data_out\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0974_ clknet_4_0_0_spi_sck _0029_ vssd1 vssd1 vccd1 vccd1 data_out\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0690_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__buf_1
XFILLER_0_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0957_ clknet_4_4_0_spi_sck _0012_ vssd1 vssd1 vccd1 vccd1 addr\[31\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0888_ _0446_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__buf_1
XFILLER_0_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_25_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0742_ _0372_ wbs_adr_o[10] _0356_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__mux2_2
X_0811_ _0406_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__buf_1
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0673_ _0231_ data_in\[0\] _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__mux2_2
X_1087_ clknet_4_8_0_spi_sck _0142_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_36_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ clknet_4_2_0_spi_sck _0065_ vssd1 vssd1 vccd1 vccd1 data_in\[5\] sky130_fd_sc_hd__dfxtp_2
X_0725_ _0361_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__buf_1
X_1139_ clknet_4_5_0_spi_sck _0191_ vssd1 vssd1 vccd1 vccd1 addr\[28\] sky130_fd_sc_hd__dfxtp_2
X_0656_ addr\[8\] _0231_ _0320_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__mux2_2
X_0587_ _0263_ shift_out\[5\] vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__and2_2
Xhold1 addr\[29\] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0510_ _0210_ _0217_ _0220_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0708_ spi_mosi addr\[0\] _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__mux2_2
X_0639_ wbs_dat_i[25] data_out\[25\] _0303_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__mux2_2
X_0990_ clknet_4_0_0_spi_sck _0045_ vssd1 vssd1 vccd1 vccd1 data_out\[25\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0973_ clknet_4_0_0_spi_sck _0028_ vssd1 vssd1 vccd1 vccd1 data_out\[8\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_28_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_7_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
X_0956_ clknet_4_5_0_spi_sck _0011_ vssd1 vssd1 vccd1 vccd1 addr\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0887_ wbs_dat_o[24] data_in\[24\] _0443_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__mux2_2
X_0741_ addr\[26\] addr\[10\] _0216_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__mux2_2
X_0810_ addr\[5\] _0242_ _0400_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_16_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0672_ _0225_ _0249_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0939_ _0469_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__buf_1
X_1086_ clknet_4_8_0_spi_sck _0141_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_7_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0724_ _0360_ wbs_adr_o[4] _0356_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__mux2_2
X_0655_ _0319_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0586_ _0252_ _0253_ _0276_ _0277_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__or4_2
X_1138_ clknet_4_7_0_spi_sck _0190_ vssd1 vssd1 vccd1 vccd1 addr\[27\] sky130_fd_sc_hd__dfxtp_2
X_1069_ clknet_4_9_0_spi_sck _0124_ vssd1 vssd1 vccd1 vccd1 data_in\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2 shift_out\[0\] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__dlygate4sd3_1
X_0707_ _0216_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__clkbuf_4
X_0638_ _0310_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__buf_1
X_0569_ _0263_ shift_out\[2\] vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__and2_2
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0972_ clknet_4_3_0_spi_sck _0027_ vssd1 vssd1 vccd1 vccd1 shift_out\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0955_ _0477_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__buf_1
XFILLER_0_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0886_ _0445_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__buf_1
X_0740_ _0371_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0671_ _0328_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__buf_1
X_0938_ command\[5\] _0242_ _0463_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__mux2_2
X_0869_ _0436_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1085_ clknet_4_2_0_spi_sck _0140_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0723_ shift_in\[3\] addr\[4\] _0348_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0654_ _0196_ _0318_ _0195_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__and3b_2
X_0585_ wbs_dat_i[5] _0247_ _0249_ data_out\[13\] vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__a22o_2
X_1137_ clknet_4_13_0_spi_sck _0189_ vssd1 vssd1 vccd1 vccd1 addr\[26\] sky130_fd_sc_hd__dfxtp_2
X_1068_ clknet_4_6_0_spi_sck _0123_ vssd1 vssd1 vccd1 vccd1 addr\[7\] sky130_fd_sc_hd__dfxtp_2
Xhold3 addr\[30\] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0706_ _0347_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__buf_1
X_0568_ spi_cs_n vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_4
X_0499_ _0195_ _0211_ _0202_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__mux2_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0637_ wbs_dat_i[24] data_out\[24\] _0303_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__mux2_2
XFILLER_0_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0971_ clknet_4_3_0_spi_sck _0026_ vssd1 vssd1 vccd1 vccd1 shift_out\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0954_ addr\[29\] shift_in\[4\] _0227_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_19_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0885_ wbs_dat_o[23] data_in\[23\] _0443_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_16_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0670_ addr\[15\] _0229_ _0320_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__mux2_2
X_1084_ clknet_4_3_0_spi_sck _0139_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_30_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0799_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_4
X_0937_ _0468_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__buf_1
X_0868_ wbs_dat_o[15] data_in\[15\] _0432_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_7_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0722_ _0359_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__buf_1
X_0653_ state\[3\] state\[2\] _0225_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nor3b_2
XPHY_EDGE_ROW_5_Left_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1136_ clknet_4_12_0_spi_sck _0188_ vssd1 vssd1 vccd1 vccd1 addr\[25\] sky130_fd_sc_hd__dfxtp_2
X_1067_ clknet_4_6_0_spi_sck _0122_ vssd1 vssd1 vccd1 vccd1 addr\[6\] sky130_fd_sc_hd__dfxtp_2
X_0584_ data_out\[21\] _0194_ _0198_ data_out\[29\] vssd1 vssd1 vccd1 vccd1 _0276_
+ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_31_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 addr\[22\] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__dlygate4sd3_1
X_0705_ addr\[23\] _0229_ _0339_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0498_ _0205_ _0206_ _0210_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a21bo_2
X_0567_ _0252_ _0253_ _0260_ _0261_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__or4_2
X_0636_ _0309_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__buf_1
X_1119_ clknet_4_7_0_spi_sck _0171_ vssd1 vssd1 vccd1 vccd1 shift_in\[3\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0619_ _0300_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_34_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0970_ clknet_4_3_0_spi_sck _0025_ vssd1 vssd1 vccd1 vccd1 shift_out\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0953_ _0476_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_19_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0884_ _0444_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__buf_1
Xclkbuf_4_13_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
X_1083_ clknet_4_2_0_spi_sck _0138_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_30_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0798_ _0195_ _0196_ _0318_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__and3b_2
X_0936_ command\[4\] _0240_ _0463_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__mux2_2
X_0867_ _0435_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_21_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1135_ clknet_4_13_0_spi_sck _0187_ vssd1 vssd1 vccd1 vccd1 addr\[24\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0721_ _0358_ wbs_adr_o[3] _0356_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__mux2_2
X_1066_ clknet_4_7_0_spi_sck _0121_ vssd1 vssd1 vccd1 vccd1 addr\[5\] sky130_fd_sc_hd__dfxtp_2
X_0919_ _0242_ _0223_ spi_cs_n vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0583_ _0246_ _0250_ shift_out\[4\] vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__a21o_2
X_0652_ _0317_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__buf_1
Xhold5 addr\[17\] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__dlygate4sd3_1
X_0704_ _0346_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__buf_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0566_ wbs_dat_i[2] _0247_ _0249_ data_out\[10\] vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__a22o_2
X_0635_ wbs_dat_i[23] data_out\[23\] _0303_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__mux2_2
X_1049_ clknet_4_13_0_spi_sck _0104_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[20] sky130_fd_sc_hd__dfxtp_2
X_1118_ clknet_4_7_0_spi_sck _0170_ vssd1 vssd1 vccd1 vccd1 shift_in\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0497_ _0207_ _0208_ _0209_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__or3b_2
X_0549_ spi_cs_n vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__inv_2
X_0618_ wbs_dat_i[15] data_out\[15\] _0292_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0952_ addr\[28\] shift_in\[3\] _0227_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_19_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0883_ wbs_dat_o[22] data_in\[22\] _0443_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0797_ wbs_adr_o[31] _0351_ _0397_ net17 vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__a22o_2
X_0866_ wbs_dat_o[14] data_in\[14\] _0432_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__mux2_2
X_0935_ _0467_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__buf_1
X_1082_ clknet_4_8_0_spi_sck _0137_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_21_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1065_ clknet_4_7_0_spi_sck _0120_ vssd1 vssd1 vccd1 vccd1 addr\[4\] sky130_fd_sc_hd__dfxtp_2
X_0720_ shift_in\[2\] addr\[3\] _0348_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__mux2_2
X_1134_ clknet_4_12_0_spi_sck _0186_ vssd1 vssd1 vccd1 vccd1 command\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0651_ wbs_dat_i[31] data_out\[31\] _0291_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__mux2_2
X_0582_ _0003_ _0270_ _0273_ _0274_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__a31o_2
X_0918_ _0460_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__buf_1
X_0849_ wbs_dat_o[6] data_in\[6\] _0421_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__mux2_2
Xhold6 addr\[16\] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__dlygate4sd3_1
X_0703_ addr\[22\] _0223_ _0339_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__mux2_2
X_1048_ clknet_4_15_0_spi_sck _0103_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[19] sky130_fd_sc_hd__dfxtp_2
X_1117_ clknet_4_13_0_spi_sck _0169_ vssd1 vssd1 vccd1 vccd1 shift_in\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0496_ state\[3\] state\[1\] state\[0\] state\[2\] vssd1 vssd1 vccd1 vccd1 _0209_
+ sky130_fd_sc_hd__nor4b_2
X_0634_ _0308_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__buf_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0565_ data_out\[18\] _0194_ _0198_ data_out\[26\] vssd1 vssd1 vccd1 vccd1 _0260_
+ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0479_ _0193_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_4
X_0617_ _0299_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__buf_1
X_0548_ _0245_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__buf_1
XFILLER_0_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0951_ _0475_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__buf_1
X_0882_ _0396_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0796_ wbs_adr_o[30] _0351_ _0397_ net4 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0934_ command\[3\] _0238_ _0463_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__mux2_2
X_0865_ _0434_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__buf_1
X_1081_ clknet_4_9_0_spi_sck _0136_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_21_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1064_ clknet_4_7_0_spi_sck _0119_ vssd1 vssd1 vccd1 vccd1 addr\[3\] sky130_fd_sc_hd__dfxtp_2
X_1133_ clknet_4_6_0_spi_sck _0185_ vssd1 vssd1 vccd1 vccd1 command\[6\] sky130_fd_sc_hd__dfxtp_2
X_0650_ _0316_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0581_ _0263_ shift_out\[4\] vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__and2_2
X_0917_ _0240_ _0242_ spi_cs_n vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__mux2_2
X_0779_ _0395_ _0232_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__nor2_2
X_0848_ _0425_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_9_Left_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7 addr\[21\] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__dlygate4sd3_1
X_1047_ clknet_4_15_0_spi_sck _0102_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[18] sky130_fd_sc_hd__dfxtp_2
X_0702_ _0345_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__buf_1
XFILLER_0_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1116_ clknet_4_12_0_spi_sck _0168_ vssd1 vssd1 vccd1 vccd1 shift_in\[0\] sky130_fd_sc_hd__dfxtp_2
X_0495_ command\[0\] command\[3\] command\[2\] command\[1\] vssd1 vssd1 vccd1 vccd1
+ _0208_ sky130_fd_sc_hd__or4b_2
X_0633_ wbs_dat_i[22] data_out\[22\] _0303_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0564_ _0246_ _0250_ shift_out\[1\] vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0616_ wbs_dat_i[14] data_out\[14\] _0292_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0478_ state\[3\] state\[2\] state\[1\] state\[0\] vssd1 vssd1 vccd1 vccd1 _0193_
+ sky130_fd_sc_hd__and4b_2
X_0547_ _0229_ data_in\[31\] _0232_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0950_ addr\[27\] shift_in\[2\] _0227_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__mux2_2
X_0881_ _0442_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__buf_1
XFILLER_0_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0795_ wbs_adr_o[29] _0351_ _0397_ net2 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0864_ wbs_dat_o[13] data_in\[13\] _0432_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__mux2_2
X_0933_ _0466_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__buf_1
X_1080_ clknet_4_9_0_spi_sck _0135_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_12_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0580_ _0252_ _0253_ _0271_ _0272_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_35_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0916_ _0459_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__buf_1
X_1063_ clknet_4_13_0_spi_sck _0118_ vssd1 vssd1 vccd1 vccd1 addr\[2\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_25_Left_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1132_ clknet_4_12_0_spi_sck _0184_ vssd1 vssd1 vccd1 vccd1 command\[5\] sky130_fd_sc_hd__dfxtp_2
X_0778_ command\[1\] _0218_ _0207_ _0219_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__or4_2
X_0847_ wbs_dat_o[5] data_in\[5\] _0421_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__mux2_2
Xhold8 addr\[24\] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__dlygate4sd3_1
X_0701_ addr\[21\] _0242_ _0339_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__mux2_2
XFILLER_0_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1046_ clknet_4_14_0_spi_sck _0101_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[17] sky130_fd_sc_hd__dfxtp_2
X_0494_ command\[5\] command\[4\] command\[7\] command\[6\] vssd1 vssd1 vccd1 vccd1
+ _0207_ sky130_fd_sc_hd__or4_2
X_1115_ clknet_4_4_0_spi_sck _0002_ _0006_ vssd1 vssd1 vccd1 vccd1 bit_count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_0632_ _0307_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__buf_1
X_0563_ _0003_ _0251_ _0256_ _0258_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__a31o_2
XFILLER_0_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1029_ clknet_4_13_0_spi_sck _0084_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[8] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0615_ _0298_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_12_Left_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0546_ _0244_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__buf_1
XFILLER_0_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0529_ _0233_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__buf_1
XFILLER_0_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0880_ wbs_dat_o[21] data_in\[21\] _0432_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__mux2_2
XFILLER_0_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ command\[2\] _0236_ _0463_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__mux2_2
X_0794_ wbs_adr_o[28] _0351_ _0397_ net14 vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__a22o_2
X_0863_ _0433_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0915_ _0238_ _0240_ _0263_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__mux2_2
X_0777_ _0351_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__buf_1
X_1062_ clknet_4_14_0_spi_sck _0117_ vssd1 vssd1 vccd1 vccd1 addr\[1\] sky130_fd_sc_hd__dfxtp_2
X_1131_ clknet_4_12_0_spi_sck _0183_ vssd1 vssd1 vccd1 vccd1 command\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_18_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0846_ _0424_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__buf_1
Xhold9 addr\[18\] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__dlygate4sd3_1
X_0700_ _0344_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__buf_1
XFILLER_0_31_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0493_ _0195_ _0196_ state\[3\] vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1114_ clknet_4_4_0_spi_sck _0001_ _0005_ vssd1 vssd1 vccd1 vccd1 bit_count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_0631_ wbs_dat_i[21] data_out\[21\] _0303_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__mux2_2
X_0562_ _0257_ shift_out\[1\] vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__and2_2
X_1045_ clknet_4_15_0_spi_sck _0100_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[16] sky130_fd_sc_hd__dfxtp_2
X_0829_ _0223_ data_in\[14\] _0409_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1028_ clknet_4_6_0_spi_sck _0083_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[7] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0614_ wbs_dat_i[13] data_out\[13\] _0292_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__mux2_2
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_2_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0545_ _0223_ data_in\[30\] _0232_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__mux2_2
XFILLER_0_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0528_ _0231_ data_in\[24\] _0232_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0793_ wbs_adr_o[27] _0351_ _0397_ net18 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a22o_2
X_0931_ _0465_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__buf_1
X_0862_ wbs_dat_o[12] data_in\[12\] _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_15_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1061_ clknet_4_13_0_spi_sck _0116_ vssd1 vssd1 vccd1 vccd1 addr\[0\] sky130_fd_sc_hd__dfxtp_2
X_0914_ _0458_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__buf_1
XFILLER_0_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1130_ clknet_4_3_0_spi_sck _0182_ vssd1 vssd1 vccd1 vccd1 command\[3\] sky130_fd_sc_hd__dfxtp_2
X_0845_ wbs_dat_o[4] data_in\[4\] _0421_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__mux2_2
X_0776_ _0393_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__buf_1
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0561_ spi_cs_n vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__buf_4
X_0492_ _0195_ _0196_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__or2_2
X_0630_ _0306_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__buf_1
X_1113_ clknet_4_4_0_spi_sck _0000_ _0004_ vssd1 vssd1 vccd1 vccd1 bit_count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_0759_ _0197_ _0225_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__and2_2
X_0828_ _0415_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__buf_1
X_1044_ clknet_4_11_0_spi_sck _0099_ vssd1 vssd1 vccd1 vccd1 data_in\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1027_ clknet_4_6_0_spi_sck _0082_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[6] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0613_ _0297_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__buf_1
X_0544_ _0243_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__buf_1
Xclkbuf_4_6_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0527_ _0216_ _0225_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__nand2_2
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0792_ wbs_adr_o[26] _0351_ _0397_ net15 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0930_ command\[1\] _0234_ _0463_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_15_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0861_ _0396_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1060_ clknet_4_4_0_spi_sck _0115_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[31] sky130_fd_sc_hd__dfxtp_2
X_0913_ _0236_ _0238_ _0263_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__mux2_2
X_0775_ data_in\[23\] _0229_ _0385_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__mux2_2
X_0844_ _0423_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__buf_1
XFILLER_0_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_29_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0758_ _0383_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__buf_1
X_0491_ state\[2\] _0204_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__xor2_2
X_0827_ _0242_ data_in\[13\] _0409_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__mux2_2
X_1043_ clknet_4_11_0_spi_sck _0098_ vssd1 vssd1 vccd1 vccd1 data_in\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0560_ _0252_ _0253_ _0254_ _0255_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__or4_2
X_1112_ clknet_4_0_0_spi_sck _0167_ vssd1 vssd1 vccd1 vccd1 shift_out\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0689_ _0195_ _0196_ _0318_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__and3_2
X_0612_ wbs_dat_i[12] data_out\[12\] _0292_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__mux2_2
X_0543_ _0242_ data_in\[29\] _0232_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__mux2_2
X_1026_ clknet_4_6_0_spi_sck _0081_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[5] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0526_ spi_mosi vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_16_Left_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1009_ clknet_4_3_0_spi_sck _0064_ vssd1 vssd1 vccd1 vccd1 data_in\[4\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_27_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0509_ command\[1\] _0218_ _0207_ _0219_ _0216_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__o41a_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0791_ wbs_adr_o[25] _0351_ _0397_ net16 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0860_ _0431_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__buf_1
X_0989_ clknet_4_0_0_spi_sck _0044_ vssd1 vssd1 vccd1 vccd1 data_out\[24\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0912_ _0457_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__buf_1
X_0774_ _0392_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__buf_1
X_0843_ wbs_dat_o[3] data_in\[3\] _0421_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1042_ clknet_4_14_0_spi_sck _0097_ vssd1 vssd1 vccd1 vccd1 data_in\[21\] sky130_fd_sc_hd__dfxtp_2
X_0490_ _0195_ _0196_ _0202_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__and3_2
Xmax_cap1 _0197_ vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
X_1111_ clknet_4_10_0_spi_sck _0166_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_30_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0757_ _0382_ wbs_adr_o[15] _0350_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__mux2_2
X_0826_ _0414_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__buf_1
XFILLER_0_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0688_ _0337_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__buf_1
XFILLER_0_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0542_ shift_in\[4\] vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0611_ _0296_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__buf_1
X_1025_ clknet_4_5_0_spi_sck _0080_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[4] sky130_fd_sc_hd__dfxtp_2
X_0809_ _0405_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0525_ _0230_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__buf_1
X_1008_ clknet_4_2_0_spi_sck _0063_ vssd1 vssd1 vccd1 vccd1 data_in\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0508_ command\[3\] command\[2\] vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__or2_2
X_0790_ wbs_adr_o[24] _0394_ _0398_ net9 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0988_ clknet_4_0_0_spi_sck _0043_ vssd1 vssd1 vccd1 vccd1 data_out\[23\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_20_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0911_ _0234_ _0236_ _0263_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__mux2_2
X_0773_ data_in\[22\] _0223_ _0385_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__mux2_2
X_0842_ _0422_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__buf_1
XFILLER_0_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1041_ clknet_4_12_0_spi_sck _0096_ vssd1 vssd1 vccd1 vccd1 data_in\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1110_ clknet_4_10_0_spi_sck _0165_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0756_ addr\[31\] addr\[15\] _0216_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0825_ _0240_ data_in\[12\] _0409_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0687_ _0229_ data_in\[7\] _0329_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_5_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0808_ addr\[4\] _0240_ _0400_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__mux2_2
X_1024_ clknet_4_7_0_spi_sck _0079_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[3] sky130_fd_sc_hd__dfxtp_2
X_0610_ wbs_dat_i[11] data_out\[11\] _0292_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__mux2_2
X_0541_ _0241_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__buf_1
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0739_ _0370_ wbs_adr_o[9] _0356_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__mux2_2
Xclkbuf_4_12_0_spi_sck clknet_0_spi_sck vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_spi_sck
+ sky130_fd_sc_hd__clkbuf_8
X_0524_ addr\[31\] _0229_ _0227_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__mux2_2
X_1007_ clknet_4_8_0_spi_sck _0062_ vssd1 vssd1 vccd1 vccd1 data_in\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0507_ command\[0\] vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0987_ clknet_4_1_0_spi_sck _0042_ vssd1 vssd1 vccd1 vccd1 data_out\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0910_ _0456_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__buf_1
X_0772_ _0391_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0841_ wbs_dat_o[2] data_in\[2\] _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1040_ clknet_4_14_0_spi_sck _0095_ vssd1 vssd1 vccd1 vccd1 data_in\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0755_ _0381_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__buf_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0824_ _0413_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__buf_1
XFILLER_0_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0686_ _0336_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__buf_1
XFILLER_0_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1023_ clknet_4_13_0_spi_sck _0078_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[2] sky130_fd_sc_hd__dfxtp_2
X_0540_ _0240_ data_in\[28\] _0232_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_5_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0807_ _0404_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__buf_1
X_0738_ addr\[25\] addr\[9\] _0348_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__mux2_2
X_0669_ _0327_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__buf_1
XFILLER_0_1_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0523_ shift_in\[6\] vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__buf_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1006_ clknet_4_9_0_spi_sck _0061_ vssd1 vssd1 vccd1 vccd1 data_in\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0506_ _0216_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0986_ clknet_4_1_0_spi_sck _0041_ vssd1 vssd1 vccd1 vccd1 data_out\[21\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_20_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0771_ data_in\[21\] _0242_ _0385_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__mux2_2
X_0840_ _0396_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0969_ clknet_4_3_0_spi_sck _0024_ vssd1 vssd1 vccd1 vccd1 shift_out\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0754_ _0380_ wbs_adr_o[14] _0350_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__mux2_2
X_0823_ _0238_ data_in\[11\] _0409_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__mux2_2
X_0685_ _0223_ data_in\[6\] _0329_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1099_ clknet_4_14_0_spi_sck _0154_ vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1022_ clknet_4_12_0_spi_sck _0077_ vssd1 vssd1 vccd1 vccd1 wbs_adr_o[1] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_5_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0737_ _0369_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__buf_1
X_0806_ addr\[3\] _0238_ _0400_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__mux2_2
X_0668_ addr\[14\] _0223_ _0320_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0599_ _0263_ shift_out\[7\] vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__and2_2
XFILLER_0_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0522_ _0228_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1005_ clknet_4_9_0_spi_sck _0060_ vssd1 vssd1 vccd1 vccd1 data_in\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0505_ _0215_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__buf_4
.ends

