##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 00:12:49 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LUT4AB
  CLASS BLOCK ;
  SIZE 210.2200 BY 219.6400 ;
  FOREIGN LUT4AB 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.5386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 218.9200 14.2200 219.6400 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 30.1638 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 150.745 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 218.9200 12.8400 219.6400 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.27075 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.495 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.3936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 96.8905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 218.9200 11.4600 219.6400 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.9658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.288 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 218.9200 10.5400 219.6400 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.4574 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.213 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 218.9200 25.2600 219.6400 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4872 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.2681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.1695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.0914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 218.9200 23.8800 219.6400 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.1216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 105.49 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 218.9200 22.5000 219.6400 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.9234 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 218.9200 21.1200 219.6400 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.4792 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.3185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.2126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.408 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 218.9200 19.7400 219.6400 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.686 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.3525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2744 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 218.9200 18.3600 219.6400 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.2835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.2465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.775 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6634 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.616 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 218.9200 16.9800 219.6400 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 229.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 218.9200 15.6000 219.6400 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.4712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.728 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 218.9200 35.8400 219.6400 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.6048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.696 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 218.9200 34.4600 219.6400 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.5192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 102.519 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.0906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.424 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 218.9200 33.5400 219.6400 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.4388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.958 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 218.9200 32.1600 219.6400 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.2698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.576 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 218.9200 30.7800 219.6400 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.636 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.1512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.638 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 218.9200 29.4000 219.6400 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.2932 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 218.9200 28.0200 219.6400 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.8644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 304.688 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 218.9200 26.6400 219.6400 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 218.9200 57.4600 219.6400 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.19 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 218.9200 56.5400 219.6400 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.2416 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 218.9200 55.1600 219.6400 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.40675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.2244 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 76.0445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.8178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 218.9200 53.7800 219.6400 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.8408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 218.9200 52.4000 219.6400 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.6 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 218.9200 51.0200 219.6400 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.8148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.816 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 218.9200 49.6400 219.6400 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.724 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.721 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 218.9200 48.2600 219.6400 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 218.9200 46.8800 219.6400 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.124 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 218.9200 45.5000 219.6400 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.8372 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.68 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 218.9200 44.1200 219.6400 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.105 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.3678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.432 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 218.9200 42.7400 219.6400 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.284 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 218.9200 41.3600 219.6400 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.3676 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.7605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.3386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.08 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 218.9200 39.9800 219.6400 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 218.9200 38.6000 219.6400 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.2066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.728 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 218.9200 37.2200 219.6400 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6124 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.944 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 218.9200 79.5400 219.6400 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.0594 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.728 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 218.9200 78.1600 219.6400 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.2912 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 218.9200 76.7800 219.6400 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.9426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.968 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 218.9200 75.4000 219.6400 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.69275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.815 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.416 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 218.9200 74.0200 219.6400 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 67.1825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.51 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 218.9200 72.6400 219.6400 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.9978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 218.9200 71.2600 219.6400 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7354 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 218.9200 69.8800 219.6400 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.32 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.5225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.318 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 218.9200 68.5000 219.6400 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.9496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.6705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 218.9200 67.1200 219.6400 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.844 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 218.9200 65.7400 219.6400 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.5788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 218.9200 64.3600 219.6400 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.0508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.408 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 218.9200 62.9800 219.6400 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.6968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.52 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 218.9200 61.6000 219.6400 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.0442 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.784 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 218.9200 60.2200 219.6400 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21295 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.427 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.9328 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.5865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 218.9200 58.8400 219.6400 ;
    END
  END NN4BEG[0]
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0209 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.067 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.6538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 177.1400 218.9200 177.5200 219.6400 ;
    END
  END Co
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.3144 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.4575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.337 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 0.0000 14.2200 0.7200 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.4976 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.2747 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 115.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.144 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 0.0000 12.8400 0.7200 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9412 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.2655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.1565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.2432 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.512 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 0.0000 11.4600 0.7200 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.9202 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.456 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 0.0000 10.5400 0.7200 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.63495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.747 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.3168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.5065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7488 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.4824 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.724 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.9892 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.3468 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 0.0000 25.2600 0.7200 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.6252 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.0485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.064 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.0552 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 0.0000 23.8800 0.7200 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7744 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.2113 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 128.475 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 0.0000 22.5000 0.7200 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.426 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.9504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 49.7024 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.563 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.284714 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 0.0000 21.1200 0.7200 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7488 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.2024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.442 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 15.8123 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.0579 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 0.0000 19.7400 0.7200 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.2616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.793 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 19.082 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.4808 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.243 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.096 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 32.8773 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 167.684 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 38.706 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.404 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 0.0000 18.3600 0.7200 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.3456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.6135 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.265 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.1274 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 12.8663 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 67.6633 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 0.0000 16.9800 0.7200 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.163 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.2035 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 29.7917 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 156.461 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 0.0000 15.6000 0.7200 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.0934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.576 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 0.0000 35.8400 0.7200 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.8791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.2245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.9886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.88 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 0.0000 34.4600 0.7200 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.2902 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.096 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 0.0000 33.5400 0.7200 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.6648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 103.246 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.7639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.9705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.672 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 0.0000 32.1600 0.7200 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.4418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.512 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 0.0000 30.7800 0.7200 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.096 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 0.0000 29.4000 0.7200 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.3999 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 0.0000 28.0200 0.7200 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.5977 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 0.0000 26.6400 0.7200 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1616 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.462 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.84242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.8175 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 0.0000 57.4600 0.7200 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.3678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.5762 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 402.178 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 0.0000 56.5400 0.7200 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.4534 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.1895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.13414 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.2761 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 0.0000 55.1600 0.7200 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.4025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.676 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2048 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.6296 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 0.0000 53.7800 0.7200 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.4646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7977 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 398.089 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 0.0000 52.4000 0.7200 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.4036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.2306 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 374.271 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 0.0000 51.0200 0.7200 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.8832 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 71.3537 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 380.854 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 0.0000 49.6400 0.7200 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.9716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.7435 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.864 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.13751 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.3838 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 0.0000 48.2600 0.7200 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.2848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.8392 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 417.706 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 0.0000 46.8800 0.7200 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.9264 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.5545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.82189 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.0189 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 0.0000 45.5000 0.7200 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.0329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.4918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.3156 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 383.108 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 0.0000 44.1200 0.7200 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.262 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.4864 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.7259 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 0.0000 42.7400 0.7200 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 0.0000 41.3600 0.7200 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.6695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.33 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.6174 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 0.0000 39.9800 0.7200 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.3054 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 0.0000 38.6000 0.7200 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.63795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.9808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.368 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 0.0000 37.2200 0.7200 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.2936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.2565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.4035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.7676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.7574 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 95.3892 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 0.0000 79.5400 0.7200 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.7208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 73.4895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.1128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.7032 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 400.535 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 0.0000 78.1600 0.7200 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75055 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.883 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.93 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.32465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.0761 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 0.0000 76.7800 0.7200 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48835 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.751 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.1464 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 70.6545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5343 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.6766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 49.1242 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 260.962 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 0.0000 75.4000 0.7200 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.69275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.815 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.8818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.6065 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.67 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 0.0000 74.0200 0.7200 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.9936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.8905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.244 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.2369 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.7401 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 0.0000 72.6400 0.7200 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.40675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.4903 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 125.296 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 0.0000 71.2600 0.7200 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3608 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.686 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.5185 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.198 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 0.0000 69.8800 0.7200 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.2538 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.1545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.602 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.76566 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.4337 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 0.0000 68.5000 0.7200 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.59832 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.6034 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 0.0000 67.1200 0.7200 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.659 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.2412 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 76.1285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.38 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.15556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.3832 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 0.0000 65.7400 0.7200 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.3134 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 73.7345 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 391.992 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 0.0000 64.3600 0.7200 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.6058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.368 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 0.0000 62.9800 0.7200 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0602 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.536 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 0.0000 61.6000 0.7200 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.9422 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 220.24 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 0.0000 60.2200 0.7200 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.1414 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 0.0000 58.8400 0.7200 ;
    END
  END NN4END[0]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.7244 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met4  ;
    ANTENNAMAXAREACAR 67.6433 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.958 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.800698 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 177.1400 0.0000 177.5200 0.7200 ;
    END
  END Ci
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5333 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.1696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 84.6400 210.2200 85.0200 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.2575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.184 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 83.2800 210.2200 83.6600 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 81.5800 210.2200 81.9600 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.139 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 80.2200 210.2200 80.6000 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.7956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.184 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 96.5400 210.2200 96.9200 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.7168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.96 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 94.8400 210.2200 95.2200 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 49.7898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 266.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 93.4800 210.2200 93.8600 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.4184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 92.1200 210.2200 92.5000 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 90.4200 210.2200 90.8000 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.1968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.2326 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 89.0600 210.2200 89.4400 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 87.7000 210.2200 88.0800 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 86.0000 210.2200 86.3800 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.639 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.6266 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.616 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 108.1000 210.2200 108.4800 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.2314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 106.7400 210.2200 107.1200 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 105.3800 210.2200 105.7600 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 267.984 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 103.6800 210.2200 104.0600 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.7658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.2876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.808 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 102.3200 210.2200 102.7000 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 100.9600 210.2200 101.3400 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 99.2600 210.2200 99.6400 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2873 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.1575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.7218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.32 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 97.9000 210.2200 98.2800 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.045 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 131.9000 210.2200 132.2800 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 42.6288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 227.824 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 130.2000 210.2200 130.5800 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.2288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 128.8400 210.2200 129.2200 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.52 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 127.4800 210.2200 127.8600 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 125.7800 210.2200 126.1600 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.9805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.6408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 124.4200 210.2200 124.8000 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.2826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 123.0600 210.2200 123.4400 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.933 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 121.3600 210.2200 121.7400 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.647 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.368 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 120.0000 210.2200 120.3800 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.5358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 118.6400 210.2200 119.0200 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.2522 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 116.9400 210.2200 117.3200 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 115.5800 210.2200 115.9600 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 114.2200 210.2200 114.6000 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 112.5200 210.2200 112.9000 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.025 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 111.1600 210.2200 111.5400 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 109.8000 210.2200 110.1800 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 149.5800 210.2200 149.9600 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.0094 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 147.8800 210.2200 148.2600 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.56 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 146.5200 210.2200 146.9000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 145.1600 210.2200 145.5400 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.191 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 143.4600 210.2200 143.8400 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.763 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 142.1000 210.2200 142.4800 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 140.7400 210.2200 141.1200 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 139.0400 210.2200 139.4200 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 137.6800 210.2200 138.0600 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.1525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 136.3200 210.2200 136.7000 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 134.6200 210.2200 135.0000 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 133.2600 210.2200 133.6400 ;
    END
  END E6BEG[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.8045 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 332.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.6400 0.7200 85.0200 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.6615 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.7856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.2800 0.7200 83.6600 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5817 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.643 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.2254 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.5800 0.7200 81.9600 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.2424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.2200 0.7200 80.6000 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.4214 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.7988 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 123.869 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.5400 0.7200 96.9200 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.7856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 43.469 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 225.115 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.8400 0.7200 95.2200 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 25.7482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.313 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.237576 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.4800 0.7200 93.8600 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0615 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.24229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.4047 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.96687 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 28.8976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 8.50505 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 43.7017 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.1200 0.7200 92.5000 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4467 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.8365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.17347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.9515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.992 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 16.386 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 83.3852 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.4200 0.7200 90.8000 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.41785 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.4842 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.497 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.784 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 24.9424 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 129.244 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 25.5954 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.36 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.0600 0.7200 89.4400 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.7017 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 371.82 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.7000 0.7200 88.0800 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6725 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.0808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.1916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 22.6995 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.422 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.0000 0.7200 86.3800 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4624 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.699 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.2223 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.1000 0.7200 108.4800 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1448 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.7400 0.7200 107.1200 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1448 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.544 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.3800 0.7200 105.7600 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.6800 0.7200 104.0600 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.5043 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3284 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.3200 0.7200 102.7000 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 215.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.332 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.6993 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.136 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 100.9600 0.7200 101.3400 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.541 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.0462 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.2600 0.7200 99.6400 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.0025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.9000 0.7200 98.2800 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.397 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.0216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 20.9881 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 108.284 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 131.9000 0.7200 132.2800 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.99731 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.701 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.2000 0.7200 130.5800 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.166 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2635 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.9293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.8400 0.7200 129.2200 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.07 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 23.8518 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.009 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.4800 0.7200 127.8600 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.25643 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.8512 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.7800 0.7200 126.1600 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.7763 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.4505 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.4200 0.7200 124.8000 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.68889 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.0135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.0600 0.7200 123.4400 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.217 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.6124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 60.9572 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 324.853 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.3600 0.7200 121.7400 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1625 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.5104 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 45.6726 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 242.624 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.0000 0.7200 120.3800 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.0155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5012 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 17.5029 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 94.1576 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.6400 0.7200 119.0200 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.1625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.3442 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 18.9916 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 102.302 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 116.9400 0.7200 117.3200 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 16.0408 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 85.4101 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.5800 0.7200 115.9600 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6874 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.2200 0.7200 114.6000 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.8516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.5200 0.7200 112.9000 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.5314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.1600 0.7200 111.5400 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.001 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.592 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.8000 0.7200 110.1800 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6865 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.9798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.94667 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 19.8949 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.5800 0.7200 149.9600 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.45 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.7536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 19.0873 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 100.734 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 147.8800 0.7200 148.2600 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.3945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.086 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 17.6628 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 94.8956 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.5200 0.7200 146.9000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.8768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 33.3639 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.466 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.1600 0.7200 145.5400 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.613 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.9331 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 134.963 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.4600 0.7200 143.8400 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.1342 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 53.0344 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.657 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.1000 0.7200 142.4800 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.3888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 232.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.8256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 15.2038 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 79.3306 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.7400 0.7200 141.1200 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.693 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.338 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.0400 0.7200 139.4200 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 22.0745 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.7 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.6800 0.7200 138.0600 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.306 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 42.3009 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 225.002 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.3200 0.7200 136.7000 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.699 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.2644 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.352 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.6200 0.7200 135.0000 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.1555 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.2600 0.7200 133.6400 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.4692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 260.384 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 0.0000 84.6000 0.7200 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.0472 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.8 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 0.0000 83.2200 0.7200 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.7684 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 320.176 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 0.0000 81.8400 0.7200 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.1892 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8315 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0693 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.14635 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.6922 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.24 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 0.0000 80.4600 0.7200 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.1478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 230.592 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 0.0000 106.2200 0.7200 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.6358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.528 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 0.0000 104.8400 0.7200 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.5338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 0.0000 103.4600 0.7200 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.77095 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.907 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.1888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.144 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 0.0000 102.5400 0.7200 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.1224 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 0.0000 101.1600 0.7200 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.5794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.168 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 0.0000 99.7800 0.7200 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.3444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 0.0000 98.4000 0.7200 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.998 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.3844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 0.0000 97.0200 0.7200 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 0.0000 95.6400 0.7200 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 0.0000 94.2600 0.7200 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.5592 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 0.0000 92.8800 0.7200 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.212 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.1658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.688 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 0.0000 91.5000 0.7200 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.3036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.282 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 0.0000 90.1200 0.7200 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.303 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.0374 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.944 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 0.0000 88.7400 0.7200 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2974 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.664 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 0.0000 87.3600 0.7200 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.978 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 0.0000 85.9800 0.7200 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2608 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.9028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.042 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 0.0000 127.8400 0.7200 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.1458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 0.0000 126.4600 0.7200 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.2718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 0.0000 125.5400 0.7200 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.9656 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.7135 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1601 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.9868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.4 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 0.0000 124.1600 0.7200 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.7794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 309.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 0.0000 122.7800 0.7200 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.354 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.6925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.9058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.968 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 0.0000 121.4000 0.7200 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.91 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.4725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.224 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 0.0000 120.0200 0.7200 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.016 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 0.0000 118.6400 0.7200 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.012 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.484 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 0.0000 117.2600 0.7200 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.2728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 0.0000 115.8800 0.7200 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.4849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.2686 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 0.0000 114.5000 0.7200 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.2728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 0.0000 113.1200 0.7200 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.69275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.815 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.9236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.5405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.98 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.782 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 0.0000 111.7400 0.7200 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.1064 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.4545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.77 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 0.0000 110.3600 0.7200 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.856 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.3458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 0.0000 108.9800 0.7200 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.6768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.08 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 0.0000 107.6000 0.7200 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8601 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.1882 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 0.0000 149.4600 0.7200 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.1842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 0.0000 148.5400 0.7200 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8483 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.1158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.088 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 0.0000 147.1600 0.7200 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.7007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.1808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 0.0000 145.7800 0.7200 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.60095 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.707 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.2996 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 46.4205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.2129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.2506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.944 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 0.0000 144.4000 0.7200 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.63495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.747 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.2216 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.0305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.752 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 0.0000 143.0200 0.7200 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.6752 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.168 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 0.0000 141.6400 0.7200 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.5748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 0.0000 140.2600 0.7200 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.339 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 0.0000 138.8800 0.7200 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 0.0000 137.5000 0.7200 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 0.0000 136.1200 0.7200 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.799 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 305.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 0.0000 134.7400 0.7200 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.6745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.2478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 0.0000 133.3600 0.7200 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 358.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 0.0000 131.9800 0.7200 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.8108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 348.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 0.0000 130.6000 0.7200 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.5334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 260.256 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 0.0000 129.2200 0.7200 ;
    END
  END SS4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.756 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.0343 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.0965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.1867 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 218.9200 84.6000 219.6400 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.0936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.44 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 218.9200 83.2200 219.6400 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.5942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.456 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.5012 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.744 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 218.9200 81.8400 219.6400 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.6669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 218.9200 80.4600 219.6400 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9962 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9035 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.8948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 84.0158 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 441.001 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 218.9200 106.2200 219.6400 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.8818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.226 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 402.341 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 218.9200 104.8400 219.6400 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.4719 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.2543 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 336.062 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 218.9200 103.4600 219.6400 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.1528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.3987 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 337.468 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 218.9200 102.5400 219.6400 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.5696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 217.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 58.0276 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 308.929 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 218.9200 101.1600 219.6400 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.6798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.9609 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 378.03 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 218.9200 99.7800 219.6400 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.89 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.4008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.4859 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 409.046 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 218.9200 98.4000 219.6400 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.0328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.899 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 380.442 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 218.9200 97.0200 219.6400 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.1304 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.2424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.708 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 218.9200 95.6400 219.6400 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.56 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 218.9200 94.2600 219.6400 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4008 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.296 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 218.9200 92.8800 219.6400 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.7064 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.512 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 218.9200 91.5000 219.6400 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9468 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.1997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.8185 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 218.9200 90.1200 219.6400 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.422 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.0225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.8235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 218.9200 88.7400 219.6400 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.42415 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.499 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6132 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9515 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.7032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.632 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 218.9200 87.3600 219.6400 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.176 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 218.9200 85.9800 219.6400 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.6724 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 8.39394 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.3724 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 218.9200 127.8400 219.6400 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.3336 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.5905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.48485 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.0296 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 218.9200 126.4600 219.6400 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.3828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.8681 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 413.7 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 218.9200 125.5400 219.6400 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.8345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.4908 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.3138 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 218.9200 124.1600 219.6400 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.3414 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 291.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.8206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.622 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 218.9200 122.7800 219.6400 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.193 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.2686 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.4117 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.74 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 218.9200 121.4000 219.6400 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.867 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.342 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.46256 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.2222 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 218.9200 120.0200 219.6400 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.3012 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 291.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.8288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 416.172 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 218.9200 118.6400 219.6400 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.5204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.9965 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 431.709 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 218.9200 117.2600 219.6400 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9336 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.5905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.6508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.6641 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.413 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 218.9200 115.8800 219.6400 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.40715 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.479 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.3468 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.6565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.162 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.56 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.4054 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 218.9200 114.5000 219.6400 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.58055 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.683 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.4488 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 72.1665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.628 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.96067 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.4088 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 218.9200 113.1200 219.6400 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9468 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.896 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.458 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 218.9200 111.7400 219.6400 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.80835 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.951 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.0635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.9865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.9536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.36 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 218.9200 110.3600 219.6400 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.3445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 218.9200 108.9800 219.6400 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.4676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 218.9200 107.6000 219.6400 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.681 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.9014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.9075 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 125.841 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 218.9200 149.4600 219.6400 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.5315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.9626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 15.8395 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.0721 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 218.9200 148.5400 219.6400 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2992 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.352 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1254 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.58485 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.3569 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 218.9200 147.1600 219.6400 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19635 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.2978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 79.0902 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.593 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 218.9200 145.7800 219.6400 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1375 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.0148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 251.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 65.8997 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.543 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 218.9200 144.4000 219.6400 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.4008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 46.6189 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 237.284 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 218.9200 143.0200 219.6400 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.03 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.9112 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 416.815 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 218.9200 141.6400 219.6400 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.9304 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.5745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8144 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.6774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 218.9200 140.2600 219.6400 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.5136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.4905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.01 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.25549 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.8828 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 218.9200 138.8800 219.6400 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.61755 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.903 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 76.2825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.84754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.8431 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 218.9200 137.5000 219.6400 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.8076 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 68.9605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.796 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.3569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.231 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 218.9200 136.1200 219.6400 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.75 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 88.676 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 31.3214 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 128.155 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 218.9200 134.7400 219.6400 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.6486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.4 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 218.9200 133.3600 219.6400 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.6334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.469 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 218.9200 131.9800 219.6400 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.9208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.099 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.4 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 218.9200 130.6000 219.6400 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.35 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 218.9200 129.2200 219.6400 ;
    END
  END SS4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.505 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.6786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 196.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 13.9200 0.7200 14.3000 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.368 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.5600 0.7200 12.9400 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.473 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.9812 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 11.2000 0.7200 11.5800 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.7206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.8400 0.7200 10.2200 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.1828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.8200 0.7200 26.2000 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.352 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.4600 0.7200 24.8400 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.013 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.839 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.7600 0.7200 23.1400 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.8688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.4000 0.7200 21.7800 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.0118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.0400 0.7200 20.4200 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.5928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.3400 0.7200 18.7200 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.9800 0.7200 17.3600 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5495 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.369 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.2188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.6200 0.7200 16.0000 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.7200 0.7200 38.1000 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.5608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.0200 0.7200 36.4000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.6588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.6600 0.7200 35.0400 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.3000 0.7200 33.6800 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.6000 0.7200 31.9800 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.2400 0.7200 30.6200 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.572 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 28.8800 0.7200 29.2600 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.1800 0.7200 27.5600 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.152 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.1800 0.7200 61.5600 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.584 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.8200 0.7200 60.2000 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.6448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.576 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.1200 0.7200 58.5000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.1968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.7600 0.7200 57.1400 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5878 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.713 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.4000 0.7200 55.7800 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.1308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.7000 0.7200 54.0800 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4221 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.2938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 220.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.3400 0.7200 52.7200 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.5914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 50.9800 0.7200 51.3600 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7692 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.2800 0.7200 49.6600 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 47.9200 0.7200 48.3000 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.7202 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.5600 0.7200 46.9400 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 149.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.8976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.8600 0.7200 45.2400 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.831 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.9858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.5000 0.7200 43.8800 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.643 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.9518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.88 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.1400 0.7200 42.5200 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.221 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.4400 0.7200 40.8200 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.921 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.184 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.0800 0.7200 39.4600 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.162 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.8600 0.7200 79.2400 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.7878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.672 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.5000 0.7200 77.8800 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.8000 0.7200 76.1800 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.031 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.4400 0.7200 74.8200 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.1384 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.0800 0.7200 73.4600 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.3800 0.7200 71.7600 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.0200 0.7200 70.4000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.5012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.388 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.6600 0.7200 69.0400 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.4407 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 66.9600 0.7200 67.3400 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.6665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.0614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.072 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.6000 0.7200 65.9800 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.328 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.2400 0.7200 64.6200 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.5400 0.7200 62.9200 ;
    END
  END W6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.871 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.1642 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 13.9200 210.2200 14.3000 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.4112 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.408 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 12.5600 210.2200 12.9400 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 67.8099 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 366.352 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 11.2000 210.2200 11.5800 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.5725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.5222 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 9.8400 210.2200 10.2200 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.095 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8672 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 15.9197 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 84.2081 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 25.8200 210.2200 26.2000 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.4798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 205.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 62.0412 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 325.972 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 24.4600 210.2200 24.8400 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.457 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.3005 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.48 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.3534 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.3279 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 22.7600 210.2200 23.1400 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 35.4121 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.863 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 21.4000 210.2200 21.7800 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.45 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.7234 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 28.103 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.228 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 20.0400 210.2200 20.4200 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.7818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.1922 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.492 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 18.3400 210.2200 18.7200 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.864 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.64377 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 29.0135 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 16.9800 210.2200 17.3600 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.731 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 31.2245 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 153.497 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 15.6200 210.2200 16.0000 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.881 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.6876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 37.7200 210.2200 38.1000 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.2248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.9024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 36.0200 210.2200 36.4000 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.3716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 34.6600 210.2200 35.0400 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.7485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.3176 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.9456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.504 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 33.3000 210.2200 33.6800 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.994 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.58 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 31.6000 210.2200 31.9800 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.0194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 230.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 30.2400 210.2200 30.6200 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.611 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.9094 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 28.8800 210.2200 29.2600 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.715 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.1918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 27.1800 210.2200 27.5600 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.4326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.463 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 38.8338 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.374 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 61.1800 210.2200 61.5600 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.64296 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.7838 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 59.8200 210.2200 60.2000 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.5308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3327 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 297.554 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 58.1200 210.2200 58.5000 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.65091 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.8236 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 56.7600 210.2200 57.1400 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.3968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 12.6447 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 64.365 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 55.4000 210.2200 55.7800 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.243 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 57.6823 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 304.498 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 53.7000 210.2200 54.0800 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.3082 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.315 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 25.0659 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.88 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 52.3400 210.2200 52.7200 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.829 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.44566 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.8471 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 50.9800 210.2200 51.3600 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.73899 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.264 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 49.2800 210.2200 49.6600 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2993 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.115 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.7158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 64.9496 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.774 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 47.9200 210.2200 48.3000 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.258 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4572 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.8976 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 46.5600 210.2200 46.9400 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.3528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 56.149 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 296.326 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 44.8600 210.2200 45.2400 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.5754 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 43.5000 210.2200 43.8800 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.183 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7596 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.7316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 42.1400 210.2200 42.5200 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.998 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 98.938 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 40.4400 210.2200 40.8200 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.6864 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 181.072 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 39.0800 210.2200 39.4600 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.231 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.312 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.1693 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 374.151 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 78.8600 210.2200 79.2400 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0161 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.7908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 20.7088 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 110.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 77.5000 210.2200 77.8800 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.5969 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.699 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 75.8000 210.2200 76.1800 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.148 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.8901 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.0559 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 74.4400 210.2200 74.8200 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.4994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 50.5959 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 268.548 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 73.0800 210.2200 73.4600 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.605 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 205.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 60.3164 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.896 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 71.3800 210.2200 71.7600 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.454 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1181 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.196 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 70.0200 210.2200 70.4000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.8348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 45.2766 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 236.668 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 68.6600 210.2200 69.0400 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.08 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.74492 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.33 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 66.9600 210.2200 67.3400 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.44 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.9732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.6552 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 335.417 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 65.6000 210.2200 65.9800 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.219 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8972 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.5521 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 305.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 64.2400 210.2200 64.6200 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.0297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4227 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 62.5400 210.2200 62.9200 ;
    END
  END W6END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2522 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 4.53963 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 23.4106 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 88.8200 0.0000 89.2000 0.7200 ;
    END
  END UserCLK
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.8858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.328 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 39.6544 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 196.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.891943 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 64.6836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 347.312 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 63.5458 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 329.177 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.891943 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 209.4200 0.7200 209.8000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.639 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met2  ;
    ANTENNAMAXAREACAR 21.8752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.382662 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.23 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 29.6406 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 146.903 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.442053 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.5015 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.944 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 67.7383 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.048 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.653459 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 207.7200 0.7200 208.1000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.505 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 70.1376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 376.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 89.2429 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 453.84 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 206.0200 0.7200 206.4000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.3522 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 66.5266 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.257 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 204.3200 0.7200 204.7000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.408 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 26.922 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.277 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.3128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 31.7706 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.101 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.941719 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.8776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.288 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 48.5923 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 242.389 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.941719 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 202.6200 0.7200 203.0000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.4163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.746 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7865 LAYER met2  ;
    ANTENNAMAXAREACAR 25.725 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.192 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.50956 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.3796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.632 LAYER met3  ;
    ANTENNAGATEAREA 3.2175 LAYER met3  ;
    ANTENNAMAXAREACAR 41.9823 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 204.765 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 200.9200 0.7200 201.3000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3615 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met2  ;
    ANTENNAMAXAREACAR 8.62684 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.733 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.524171 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 10.6551 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49.243 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.583562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.4726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.128 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 41.3344 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 204.633 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.666038 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 198.8800 0.7200 199.2600 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4545 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met2  ;
    ANTENNAMAXAREACAR 24.4133 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 115.856 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.665681 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 25.9292 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 124.634 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.725072 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.6044 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 57.968 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 40.6995 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 205.018 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.01824 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 197.1800 0.7200 197.5600 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2611 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.0265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 67.4962 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 332.28 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.9314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.096 LAYER met3  ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 71.1835 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 352.526 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.625157 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.1932 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.912 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 79.6352 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 398.187 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 195.4800 0.7200 195.8600 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.696 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 41.7497 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 202.802 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.6248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 47.6457 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.23 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.0942 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.776 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 60.7286 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.022 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 193.7800 0.7200 194.1600 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.23 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.7555 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 75.5309 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 382.324 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 192.0800 0.7200 192.4600 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.5665 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.138 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5815 LAYER met2  ;
    ANTENNAMAXAREACAR 60.5204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 297.045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.637279 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.42947 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met3  ;
    ANTENNAGATEAREA 2.7405 LAYER met3  ;
    ANTENNAMAXAREACAR 62.1367 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 305.995 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.651875 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 63.791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 314.972 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 190.0400 0.7200 190.4200 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.769 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 79.791 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 430.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 63.5431 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.468 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 188.3400 0.7200 188.7200 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.501 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 36.9984 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 180.892 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 186.6400 0.7200 187.0200 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.2048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.52 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 101.563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 534.529 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 184.9400 0.7200 185.3200 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.294 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met2  ;
    ANTENNAMAXAREACAR 61.9523 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 302.937 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.843895 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5215 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.696 LAYER met3  ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 62.5787 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 307.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.939991 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.439 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.88 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 77.1084 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.48 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.939991 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 183.2400 0.7200 183.6200 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.5246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 45.2725 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.041 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.528173 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 181.2000 0.7200 181.5800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.1808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.6673 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 66.3389 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 338.614 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.41342 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 179.5000 0.7200 179.8800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.3979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.4372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 52.9567 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.965 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.616771 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.1365 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.016 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 65.7527 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.285 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 177.8000 0.7200 178.1800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 75.2163 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 407.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 100.711 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 526.108 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 176.1000 0.7200 176.4800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.4568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6275 LAYER met3  ;
    ANTENNAMAXAREACAR 48.0373 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 241.45 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.538513 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.0806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.704 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 49.3714 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.874 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.662194 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 174.4000 0.7200 174.7800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.0138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 56.8031 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.745 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.839493 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 172.3600 0.7200 172.7400 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.507 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.1996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 89.7201 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 465.526 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 170.6600 0.7200 171.0400 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.1068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.2821 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 40.1146 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 200.9 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.855607 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 168.9600 0.7200 169.3400 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.3638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 60.6025 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.018 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.943842 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.0691 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 207.264 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 73.0495 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 380.784 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 167.2600 0.7200 167.6400 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0205 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met2  ;
    ANTENNAMAXAREACAR 54.106 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 265.554 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.577297 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 55.2311 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 272.868 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.689815 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.0872 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.032 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 70.2997 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 354.618 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 165.5600 0.7200 165.9400 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.4196 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 55.9182 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.729 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.757473 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 163.5200 0.7200 163.9000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 93.464 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met2  ;
    ANTENNAMAXAREACAR 34.0365 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 164.868 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.524171 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 34.6304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 168.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.583562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.1144 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.688 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 48.3404 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.645 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 161.8200 0.7200 162.2000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.239 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 92.877 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 498.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 95.96 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 489.716 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.19033 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 160.1200 0.7200 160.5000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.212 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.2307 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 67.3773 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.119 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.10943 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 158.4200 0.7200 158.8000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.1986 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 93.321 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 501.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 97.2652 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 511.847 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.10943 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 156.7200 0.7200 157.1000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.5519 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 84.7975 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 431.822 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.3687 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 262.656 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 100.612 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 517.699 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 155.0200 0.7200 155.4000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 209.4200 210.2200 209.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.5198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.576 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 207.7200 210.2200 208.1000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.1422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.367 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 206.0200 210.2200 206.4000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.8918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.233 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 204.3200 210.2200 204.7000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.56 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.802 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 202.6200 210.2200 203.0000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.1078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.712 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 200.9200 210.2200 201.3000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 198.8800 210.2200 199.2600 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0852 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 197.1800 210.2200 197.5600 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1397 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.322 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.072 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 195.4800 210.2200 195.8600 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.7878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.672 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 193.7800 210.2200 194.1600 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.9886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.88 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 192.0800 210.2200 192.4600 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.9976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 190.0400 210.2200 190.4200 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.4858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 188.3400 210.2200 188.7200 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.14 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 186.6400 210.2200 187.0200 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 184.9400 210.2200 185.3200 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.8538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.808 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 183.2400 210.2200 183.6200 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.6285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.592 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.9938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.104 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 181.2000 210.2200 181.5800 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.621 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 179.5000 210.2200 179.8800 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.441 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.9052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 177.8000 210.2200 178.1800 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 176.1000 210.2200 176.4800 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0372 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 174.4000 210.2200 174.7800 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.3618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 194.4 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 172.3600 210.2200 172.7400 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.9528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 170.6600 210.2200 171.0400 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 168.9600 210.2200 169.3400 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.0445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.6764 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.352 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 167.2600 210.2200 167.6400 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 250.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 165.5600 210.2200 165.9400 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 163.5200 210.2200 163.9000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.1326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 305.648 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 161.8200 210.2200 162.2000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.4552 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 160.1200 210.2200 160.5000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.571 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 158.4200 210.2200 158.8000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.5798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4674 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.904 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 156.7200 210.2200 157.1000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4346 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 155.0200 210.2200 155.4000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.9778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.1263 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 367.301 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 199.2200 0.0000 199.6000 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.103 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5112 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.0412 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 197.3800 0.0000 197.7600 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.873 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 100.317 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met2  ;
    ANTENNAMAXAREACAR 17.341 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.3795 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 195.0800 0.0000 195.4600 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 21.611 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 102.51 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.780525 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 192.7800 0.0000 193.1600 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.7655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.1715 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2472 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.6551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.757388 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.344 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 15.5621 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.4233 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.757388 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 190.4800 0.0000 190.8600 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.0832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 102.179 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.8075 LAYER met2  ;
    ANTENNAMAXAREACAR 11.9251 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.7446 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.654861 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 12.1043 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 53.7892 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.654861 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 188.1800 0.0000 188.5600 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3601 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.3644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 39.2882 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 197.195 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.792453 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 185.4200 0.0000 185.8000 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.7723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.3465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 63.3368 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 305.178 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.913836 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.0049 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.488 LAYER met3  ;
    ANTENNAGATEAREA 1.1505 LAYER met3  ;
    ANTENNAMAXAREACAR 84.2015 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 416.858 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.948604 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 84.4318 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.175 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.948604 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 184.0400 0.0000 184.4200 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.9422 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 31.8125 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 154.622 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.88232 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 181.2800 0.0000 181.6600 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 33.8879 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 164.907 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.833984 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 179.4400 0.0000 179.8200 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.0548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 29.5849 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.375 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.62172 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 174.8400 0.0000 175.2200 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 60.1317 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 325.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 42.2221 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 217.376 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 172.5400 0.0000 172.9200 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.599 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 38.4948 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.272 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 170.2400 0.0000 170.6200 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.127 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.5754 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 49.2555 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.502 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.762937 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 168.4000 0.0000 168.7800 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.29 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 13.3522 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.3931 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.3158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.288 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 26.4274 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 131.601 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.9712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.728 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 46.4591 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.629 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.871908 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 166.1000 0.0000 166.4800 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.4774 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 24.6796 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 119.962 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.819497 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 163.8000 0.0000 164.1800 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.3307 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 33.1719 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.04 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 161.0400 0.0000 161.4200 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.3286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 38.9532 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.448 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.772009 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 159.2000 0.0000 159.5800 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.1339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 147.304 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0125 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6825 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.7852 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.474749 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAGATEAREA 4.0125 LAYER met3  ;
    ANTENNAMAXAREACAR 18.0746 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 86.9923 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.484718 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.1166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.896 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 36.2939 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.573 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 156.9000 0.0000 157.2800 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.3832 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 23.9194 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 115.206 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.639571 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 155.0600 0.0000 155.4400 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1594 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.689 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 199.2200 218.9200 199.6000 219.6400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 197.3800 218.9200 197.7600 219.6400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.8328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 343.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 194.6200 218.9200 195.0000 219.6400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.1214 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 192.7800 218.9200 193.1600 219.6400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.492 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 190.4800 218.9200 190.8600 219.6400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.8058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 188.1800 218.9200 188.5600 219.6400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.1068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 185.8800 218.9200 186.2600 219.6400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.7242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 184.0400 218.9200 184.4200 219.6400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5825 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.0918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 181.2800 218.9200 181.6600 219.6400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 179.4400 218.9200 179.8200 219.6400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.052 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.8400 218.9200 175.2200 219.6400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0158 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.853 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 172.5400 218.9200 172.9200 219.6400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.961 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 170.2400 218.9200 170.6200 219.6400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.137 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 168.4000 218.9200 168.7800 219.6400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.1000 218.9200 166.4800 219.6400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.033 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.8000 218.9200 164.1800 219.6400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2895 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.8558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.368 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 161.5000 218.9200 161.8800 219.6400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.8458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 322 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 159.2000 218.9200 159.5800 219.6400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.7208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 156.4400 218.9200 156.8200 219.6400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.3718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 155.0600 218.9200 155.4400 219.6400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 204.6600 8.4300 ;
        RECT 5.5600 210.5300 204.6600 213.5300 ;
        RECT 5.5600 12.3400 8.5600 12.8200 ;
        RECT 5.5600 23.2200 8.5600 23.7000 ;
        RECT 5.5600 17.7800 8.5600 18.2600 ;
        RECT 5.5600 39.5400 8.5600 40.0200 ;
        RECT 5.5600 28.6600 8.5600 29.1400 ;
        RECT 5.5600 34.1000 8.5600 34.5800 ;
        RECT 5.5600 50.4200 8.5600 50.9000 ;
        RECT 5.5600 44.9800 8.5600 45.4600 ;
        RECT 55.1200 12.3400 56.7200 12.8200 ;
        RECT 55.1200 17.7800 56.7200 18.2600 ;
        RECT 55.1200 23.2200 56.7200 23.7000 ;
        RECT 100.1200 12.3400 101.7200 12.8200 ;
        RECT 100.1200 17.7800 101.7200 18.2600 ;
        RECT 100.1200 23.2200 101.7200 23.7000 ;
        RECT 55.1200 39.5400 56.7200 40.0200 ;
        RECT 55.1200 34.1000 56.7200 34.5800 ;
        RECT 55.1200 28.6600 56.7200 29.1400 ;
        RECT 55.1200 50.4200 56.7200 50.9000 ;
        RECT 55.1200 44.9800 56.7200 45.4600 ;
        RECT 100.1200 39.5400 101.7200 40.0200 ;
        RECT 100.1200 34.1000 101.7200 34.5800 ;
        RECT 100.1200 28.6600 101.7200 29.1400 ;
        RECT 100.1200 50.4200 101.7200 50.9000 ;
        RECT 100.1200 44.9800 101.7200 45.4600 ;
        RECT 5.5600 66.7400 8.5600 67.2200 ;
        RECT 5.5600 55.8600 8.5600 56.3400 ;
        RECT 5.5600 61.3000 8.5600 61.7800 ;
        RECT 5.5600 77.6200 8.5600 78.1000 ;
        RECT 5.5600 72.1800 8.5600 72.6600 ;
        RECT 5.5600 93.9400 8.5600 94.4200 ;
        RECT 5.5600 83.0600 8.5600 83.5400 ;
        RECT 5.5600 88.5000 8.5600 88.9800 ;
        RECT 5.5600 104.8200 8.5600 105.3000 ;
        RECT 5.5600 99.3800 8.5600 99.8600 ;
        RECT 55.1200 66.7400 56.7200 67.2200 ;
        RECT 55.1200 61.3000 56.7200 61.7800 ;
        RECT 55.1200 55.8600 56.7200 56.3400 ;
        RECT 55.1200 77.6200 56.7200 78.1000 ;
        RECT 55.1200 72.1800 56.7200 72.6600 ;
        RECT 100.1200 66.7400 101.7200 67.2200 ;
        RECT 100.1200 61.3000 101.7200 61.7800 ;
        RECT 100.1200 55.8600 101.7200 56.3400 ;
        RECT 100.1200 77.6200 101.7200 78.1000 ;
        RECT 100.1200 72.1800 101.7200 72.6600 ;
        RECT 55.1200 93.9400 56.7200 94.4200 ;
        RECT 55.1200 88.5000 56.7200 88.9800 ;
        RECT 55.1200 83.0600 56.7200 83.5400 ;
        RECT 55.1200 104.8200 56.7200 105.3000 ;
        RECT 55.1200 99.3800 56.7200 99.8600 ;
        RECT 100.1200 93.9400 101.7200 94.4200 ;
        RECT 100.1200 88.5000 101.7200 88.9800 ;
        RECT 100.1200 83.0600 101.7200 83.5400 ;
        RECT 100.1200 104.8200 101.7200 105.3000 ;
        RECT 100.1200 99.3800 101.7200 99.8600 ;
        RECT 145.1200 12.3400 146.7200 12.8200 ;
        RECT 145.1200 23.2200 146.7200 23.7000 ;
        RECT 145.1200 17.7800 146.7200 18.2600 ;
        RECT 145.1200 39.5400 146.7200 40.0200 ;
        RECT 145.1200 34.1000 146.7200 34.5800 ;
        RECT 145.1200 28.6600 146.7200 29.1400 ;
        RECT 145.1200 50.4200 146.7200 50.9000 ;
        RECT 145.1200 44.9800 146.7200 45.4600 ;
        RECT 190.1200 12.3400 191.7200 12.8200 ;
        RECT 201.6600 12.3400 204.6600 12.8200 ;
        RECT 190.1200 23.2200 191.7200 23.7000 ;
        RECT 190.1200 17.7800 191.7200 18.2600 ;
        RECT 201.6600 23.2200 204.6600 23.7000 ;
        RECT 201.6600 17.7800 204.6600 18.2600 ;
        RECT 190.1200 39.5400 191.7200 40.0200 ;
        RECT 190.1200 34.1000 191.7200 34.5800 ;
        RECT 190.1200 28.6600 191.7200 29.1400 ;
        RECT 201.6600 39.5400 204.6600 40.0200 ;
        RECT 201.6600 34.1000 204.6600 34.5800 ;
        RECT 201.6600 28.6600 204.6600 29.1400 ;
        RECT 190.1200 50.4200 191.7200 50.9000 ;
        RECT 190.1200 44.9800 191.7200 45.4600 ;
        RECT 201.6600 50.4200 204.6600 50.9000 ;
        RECT 201.6600 44.9800 204.6600 45.4600 ;
        RECT 145.1200 66.7400 146.7200 67.2200 ;
        RECT 145.1200 61.3000 146.7200 61.7800 ;
        RECT 145.1200 55.8600 146.7200 56.3400 ;
        RECT 145.1200 77.6200 146.7200 78.1000 ;
        RECT 145.1200 72.1800 146.7200 72.6600 ;
        RECT 145.1200 93.9400 146.7200 94.4200 ;
        RECT 145.1200 88.5000 146.7200 88.9800 ;
        RECT 145.1200 83.0600 146.7200 83.5400 ;
        RECT 145.1200 104.8200 146.7200 105.3000 ;
        RECT 145.1200 99.3800 146.7200 99.8600 ;
        RECT 190.1200 66.7400 191.7200 67.2200 ;
        RECT 190.1200 61.3000 191.7200 61.7800 ;
        RECT 190.1200 55.8600 191.7200 56.3400 ;
        RECT 201.6600 66.7400 204.6600 67.2200 ;
        RECT 201.6600 61.3000 204.6600 61.7800 ;
        RECT 201.6600 55.8600 204.6600 56.3400 ;
        RECT 190.1200 77.6200 191.7200 78.1000 ;
        RECT 190.1200 72.1800 191.7200 72.6600 ;
        RECT 201.6600 77.6200 204.6600 78.1000 ;
        RECT 201.6600 72.1800 204.6600 72.6600 ;
        RECT 190.1200 93.9400 191.7200 94.4200 ;
        RECT 190.1200 88.5000 191.7200 88.9800 ;
        RECT 190.1200 83.0600 191.7200 83.5400 ;
        RECT 201.6600 93.9400 204.6600 94.4200 ;
        RECT 201.6600 88.5000 204.6600 88.9800 ;
        RECT 201.6600 83.0600 204.6600 83.5400 ;
        RECT 190.1200 104.8200 191.7200 105.3000 ;
        RECT 190.1200 99.3800 191.7200 99.8600 ;
        RECT 201.6600 104.8200 204.6600 105.3000 ;
        RECT 201.6600 99.3800 204.6600 99.8600 ;
        RECT 100.1200 164.6600 101.7200 165.1400 ;
        RECT 55.1200 164.6600 56.7200 165.1400 ;
        RECT 5.5600 164.6600 8.5600 165.1400 ;
        RECT 5.5600 121.1400 8.5600 121.6200 ;
        RECT 5.5600 110.2600 8.5600 110.7400 ;
        RECT 5.5600 115.7000 8.5600 116.1800 ;
        RECT 5.5600 132.0200 8.5600 132.5000 ;
        RECT 5.5600 126.5800 8.5600 127.0600 ;
        RECT 5.5600 148.3400 8.5600 148.8200 ;
        RECT 5.5600 137.4600 8.5600 137.9400 ;
        RECT 5.5600 142.9000 8.5600 143.3800 ;
        RECT 5.5600 159.2200 8.5600 159.7000 ;
        RECT 5.5600 153.7800 8.5600 154.2600 ;
        RECT 55.1200 121.1400 56.7200 121.6200 ;
        RECT 55.1200 115.7000 56.7200 116.1800 ;
        RECT 55.1200 110.2600 56.7200 110.7400 ;
        RECT 55.1200 132.0200 56.7200 132.5000 ;
        RECT 55.1200 126.5800 56.7200 127.0600 ;
        RECT 100.1200 121.1400 101.7200 121.6200 ;
        RECT 100.1200 115.7000 101.7200 116.1800 ;
        RECT 100.1200 110.2600 101.7200 110.7400 ;
        RECT 100.1200 132.0200 101.7200 132.5000 ;
        RECT 100.1200 126.5800 101.7200 127.0600 ;
        RECT 55.1200 148.3400 56.7200 148.8200 ;
        RECT 55.1200 142.9000 56.7200 143.3800 ;
        RECT 55.1200 137.4600 56.7200 137.9400 ;
        RECT 55.1200 159.2200 56.7200 159.7000 ;
        RECT 55.1200 153.7800 56.7200 154.2600 ;
        RECT 100.1200 148.3400 101.7200 148.8200 ;
        RECT 100.1200 142.9000 101.7200 143.3800 ;
        RECT 100.1200 137.4600 101.7200 137.9400 ;
        RECT 100.1200 159.2200 101.7200 159.7000 ;
        RECT 100.1200 153.7800 101.7200 154.2600 ;
        RECT 5.5600 191.8600 8.5600 192.3400 ;
        RECT 5.5600 170.1000 8.5600 170.5800 ;
        RECT 5.5600 175.5400 8.5600 176.0200 ;
        RECT 5.5600 180.9800 8.5600 181.4600 ;
        RECT 5.5600 186.4200 8.5600 186.9000 ;
        RECT 5.5600 197.3000 8.5600 197.7800 ;
        RECT 5.5600 202.7400 8.5600 203.2200 ;
        RECT 5.5600 208.1800 8.5600 208.6600 ;
        RECT 100.1200 191.8600 101.7200 192.3400 ;
        RECT 55.1200 191.8600 56.7200 192.3400 ;
        RECT 55.1200 175.5400 56.7200 176.0200 ;
        RECT 55.1200 170.1000 56.7200 170.5800 ;
        RECT 55.1200 186.4200 56.7200 186.9000 ;
        RECT 55.1200 180.9800 56.7200 181.4600 ;
        RECT 100.1200 175.5400 101.7200 176.0200 ;
        RECT 100.1200 170.1000 101.7200 170.5800 ;
        RECT 100.1200 186.4200 101.7200 186.9000 ;
        RECT 100.1200 180.9800 101.7200 181.4600 ;
        RECT 55.1200 208.1800 56.7200 208.6600 ;
        RECT 55.1200 202.7400 56.7200 203.2200 ;
        RECT 55.1200 197.3000 56.7200 197.7800 ;
        RECT 100.1200 208.1800 101.7200 208.6600 ;
        RECT 100.1200 202.7400 101.7200 203.2200 ;
        RECT 100.1200 197.3000 101.7200 197.7800 ;
        RECT 190.1200 164.6600 191.7200 165.1400 ;
        RECT 145.1200 164.6600 146.7200 165.1400 ;
        RECT 201.6600 164.6600 204.6600 165.1400 ;
        RECT 145.1200 121.1400 146.7200 121.6200 ;
        RECT 145.1200 115.7000 146.7200 116.1800 ;
        RECT 145.1200 110.2600 146.7200 110.7400 ;
        RECT 145.1200 132.0200 146.7200 132.5000 ;
        RECT 145.1200 126.5800 146.7200 127.0600 ;
        RECT 145.1200 148.3400 146.7200 148.8200 ;
        RECT 145.1200 142.9000 146.7200 143.3800 ;
        RECT 145.1200 137.4600 146.7200 137.9400 ;
        RECT 145.1200 159.2200 146.7200 159.7000 ;
        RECT 145.1200 153.7800 146.7200 154.2600 ;
        RECT 190.1200 121.1400 191.7200 121.6200 ;
        RECT 190.1200 115.7000 191.7200 116.1800 ;
        RECT 190.1200 110.2600 191.7200 110.7400 ;
        RECT 201.6600 121.1400 204.6600 121.6200 ;
        RECT 201.6600 115.7000 204.6600 116.1800 ;
        RECT 201.6600 110.2600 204.6600 110.7400 ;
        RECT 190.1200 132.0200 191.7200 132.5000 ;
        RECT 190.1200 126.5800 191.7200 127.0600 ;
        RECT 201.6600 132.0200 204.6600 132.5000 ;
        RECT 201.6600 126.5800 204.6600 127.0600 ;
        RECT 190.1200 148.3400 191.7200 148.8200 ;
        RECT 190.1200 142.9000 191.7200 143.3800 ;
        RECT 190.1200 137.4600 191.7200 137.9400 ;
        RECT 201.6600 148.3400 204.6600 148.8200 ;
        RECT 201.6600 142.9000 204.6600 143.3800 ;
        RECT 201.6600 137.4600 204.6600 137.9400 ;
        RECT 190.1200 159.2200 191.7200 159.7000 ;
        RECT 190.1200 153.7800 191.7200 154.2600 ;
        RECT 201.6600 159.2200 204.6600 159.7000 ;
        RECT 201.6600 153.7800 204.6600 154.2600 ;
        RECT 145.1200 191.8600 146.7200 192.3400 ;
        RECT 145.1200 170.1000 146.7200 170.5800 ;
        RECT 145.1200 175.5400 146.7200 176.0200 ;
        RECT 145.1200 186.4200 146.7200 186.9000 ;
        RECT 145.1200 180.9800 146.7200 181.4600 ;
        RECT 145.1200 208.1800 146.7200 208.6600 ;
        RECT 145.1200 202.7400 146.7200 203.2200 ;
        RECT 145.1200 197.3000 146.7200 197.7800 ;
        RECT 190.1200 191.8600 191.7200 192.3400 ;
        RECT 201.6600 191.8600 204.6600 192.3400 ;
        RECT 190.1200 175.5400 191.7200 176.0200 ;
        RECT 190.1200 170.1000 191.7200 170.5800 ;
        RECT 201.6600 175.5400 204.6600 176.0200 ;
        RECT 201.6600 170.1000 204.6600 170.5800 ;
        RECT 190.1200 186.4200 191.7200 186.9000 ;
        RECT 190.1200 180.9800 191.7200 181.4600 ;
        RECT 201.6600 186.4200 204.6600 186.9000 ;
        RECT 201.6600 180.9800 204.6600 181.4600 ;
        RECT 190.1200 202.7400 191.7200 203.2200 ;
        RECT 190.1200 197.3000 191.7200 197.7800 ;
        RECT 201.6600 202.7400 204.6600 203.2200 ;
        RECT 201.6600 197.3000 204.6600 197.7800 ;
        RECT 190.1200 208.1800 191.7200 208.6600 ;
        RECT 201.6600 208.1800 204.6600 208.6600 ;
      LAYER met4 ;
        RECT 5.5600 5.4300 8.5600 213.5300 ;
        RECT 201.6600 5.4300 204.6600 213.5300 ;
        RECT 55.1200 5.4300 56.7200 213.5300 ;
        RECT 100.1200 5.4300 101.7200 213.5300 ;
        RECT 145.1200 5.4300 146.7200 213.5300 ;
        RECT 190.1200 5.4300 191.7200 213.5300 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 1.5600 1.4300 208.6600 4.4300 ;
        RECT 1.5600 214.5300 208.6600 217.5300 ;
        RECT 13.3200 9.6200 14.9200 10.1000 ;
        RECT 1.5600 9.6200 4.5600 10.1000 ;
        RECT 1.5600 25.9400 4.5600 26.4200 ;
        RECT 1.5600 20.5000 4.5600 20.9800 ;
        RECT 1.5600 15.0600 4.5600 15.5400 ;
        RECT 13.3200 25.9400 14.9200 26.4200 ;
        RECT 13.3200 20.5000 14.9200 20.9800 ;
        RECT 13.3200 15.0600 14.9200 15.5400 ;
        RECT 1.5600 36.8200 4.5600 37.3000 ;
        RECT 1.5600 31.3800 4.5600 31.8600 ;
        RECT 13.3200 36.8200 14.9200 37.3000 ;
        RECT 13.3200 31.3800 14.9200 31.8600 ;
        RECT 1.5600 53.1400 4.5600 53.6200 ;
        RECT 1.5600 47.7000 4.5600 48.1800 ;
        RECT 1.5600 42.2600 4.5600 42.7400 ;
        RECT 13.3200 53.1400 14.9200 53.6200 ;
        RECT 13.3200 47.7000 14.9200 48.1800 ;
        RECT 13.3200 42.2600 14.9200 42.7400 ;
        RECT 58.3200 9.6200 59.9200 10.1000 ;
        RECT 58.3200 25.9400 59.9200 26.4200 ;
        RECT 58.3200 20.5000 59.9200 20.9800 ;
        RECT 58.3200 15.0600 59.9200 15.5400 ;
        RECT 103.3200 9.6200 104.9200 10.1000 ;
        RECT 103.3200 25.9400 104.9200 26.4200 ;
        RECT 103.3200 20.5000 104.9200 20.9800 ;
        RECT 103.3200 15.0600 104.9200 15.5400 ;
        RECT 58.3200 36.8200 59.9200 37.3000 ;
        RECT 58.3200 31.3800 59.9200 31.8600 ;
        RECT 58.3200 53.1400 59.9200 53.6200 ;
        RECT 58.3200 47.7000 59.9200 48.1800 ;
        RECT 58.3200 42.2600 59.9200 42.7400 ;
        RECT 103.3200 36.8200 104.9200 37.3000 ;
        RECT 103.3200 31.3800 104.9200 31.8600 ;
        RECT 103.3200 53.1400 104.9200 53.6200 ;
        RECT 103.3200 47.7000 104.9200 48.1800 ;
        RECT 103.3200 42.2600 104.9200 42.7400 ;
        RECT 1.5600 64.0200 4.5600 64.5000 ;
        RECT 1.5600 58.5800 4.5600 59.0600 ;
        RECT 13.3200 64.0200 14.9200 64.5000 ;
        RECT 13.3200 58.5800 14.9200 59.0600 ;
        RECT 1.5600 80.3400 4.5600 80.8200 ;
        RECT 1.5600 74.9000 4.5600 75.3800 ;
        RECT 1.5600 69.4600 4.5600 69.9400 ;
        RECT 13.3200 80.3400 14.9200 80.8200 ;
        RECT 13.3200 74.9000 14.9200 75.3800 ;
        RECT 13.3200 69.4600 14.9200 69.9400 ;
        RECT 1.5600 91.2200 4.5600 91.7000 ;
        RECT 1.5600 85.7800 4.5600 86.2600 ;
        RECT 13.3200 91.2200 14.9200 91.7000 ;
        RECT 13.3200 85.7800 14.9200 86.2600 ;
        RECT 1.5600 107.5400 4.5600 108.0200 ;
        RECT 1.5600 102.1000 4.5600 102.5800 ;
        RECT 1.5600 96.6600 4.5600 97.1400 ;
        RECT 13.3200 107.5400 14.9200 108.0200 ;
        RECT 13.3200 102.1000 14.9200 102.5800 ;
        RECT 13.3200 96.6600 14.9200 97.1400 ;
        RECT 58.3200 64.0200 59.9200 64.5000 ;
        RECT 58.3200 58.5800 59.9200 59.0600 ;
        RECT 58.3200 80.3400 59.9200 80.8200 ;
        RECT 58.3200 74.9000 59.9200 75.3800 ;
        RECT 58.3200 69.4600 59.9200 69.9400 ;
        RECT 103.3200 64.0200 104.9200 64.5000 ;
        RECT 103.3200 58.5800 104.9200 59.0600 ;
        RECT 103.3200 80.3400 104.9200 80.8200 ;
        RECT 103.3200 74.9000 104.9200 75.3800 ;
        RECT 103.3200 69.4600 104.9200 69.9400 ;
        RECT 58.3200 91.2200 59.9200 91.7000 ;
        RECT 58.3200 85.7800 59.9200 86.2600 ;
        RECT 58.3200 107.5400 59.9200 108.0200 ;
        RECT 58.3200 102.1000 59.9200 102.5800 ;
        RECT 58.3200 96.6600 59.9200 97.1400 ;
        RECT 103.3200 91.2200 104.9200 91.7000 ;
        RECT 103.3200 85.7800 104.9200 86.2600 ;
        RECT 103.3200 107.5400 104.9200 108.0200 ;
        RECT 103.3200 102.1000 104.9200 102.5800 ;
        RECT 103.3200 96.6600 104.9200 97.1400 ;
        RECT 148.3200 9.6200 149.9200 10.1000 ;
        RECT 148.3200 25.9400 149.9200 26.4200 ;
        RECT 148.3200 20.5000 149.9200 20.9800 ;
        RECT 148.3200 15.0600 149.9200 15.5400 ;
        RECT 148.3200 36.8200 149.9200 37.3000 ;
        RECT 148.3200 31.3800 149.9200 31.8600 ;
        RECT 148.3200 53.1400 149.9200 53.6200 ;
        RECT 148.3200 47.7000 149.9200 48.1800 ;
        RECT 148.3200 42.2600 149.9200 42.7400 ;
        RECT 193.3200 9.6200 194.9200 10.1000 ;
        RECT 205.6600 9.6200 208.6600 10.1000 ;
        RECT 193.3200 25.9400 194.9200 26.4200 ;
        RECT 193.3200 20.5000 194.9200 20.9800 ;
        RECT 193.3200 15.0600 194.9200 15.5400 ;
        RECT 205.6600 25.9400 208.6600 26.4200 ;
        RECT 205.6600 20.5000 208.6600 20.9800 ;
        RECT 205.6600 15.0600 208.6600 15.5400 ;
        RECT 193.3200 36.8200 194.9200 37.3000 ;
        RECT 193.3200 31.3800 194.9200 31.8600 ;
        RECT 205.6600 36.8200 208.6600 37.3000 ;
        RECT 205.6600 31.3800 208.6600 31.8600 ;
        RECT 193.3200 53.1400 194.9200 53.6200 ;
        RECT 193.3200 47.7000 194.9200 48.1800 ;
        RECT 193.3200 42.2600 194.9200 42.7400 ;
        RECT 205.6600 53.1400 208.6600 53.6200 ;
        RECT 205.6600 47.7000 208.6600 48.1800 ;
        RECT 205.6600 42.2600 208.6600 42.7400 ;
        RECT 148.3200 64.0200 149.9200 64.5000 ;
        RECT 148.3200 58.5800 149.9200 59.0600 ;
        RECT 148.3200 80.3400 149.9200 80.8200 ;
        RECT 148.3200 74.9000 149.9200 75.3800 ;
        RECT 148.3200 69.4600 149.9200 69.9400 ;
        RECT 148.3200 91.2200 149.9200 91.7000 ;
        RECT 148.3200 85.7800 149.9200 86.2600 ;
        RECT 148.3200 107.5400 149.9200 108.0200 ;
        RECT 148.3200 102.1000 149.9200 102.5800 ;
        RECT 148.3200 96.6600 149.9200 97.1400 ;
        RECT 193.3200 64.0200 194.9200 64.5000 ;
        RECT 193.3200 58.5800 194.9200 59.0600 ;
        RECT 205.6600 64.0200 208.6600 64.5000 ;
        RECT 205.6600 58.5800 208.6600 59.0600 ;
        RECT 193.3200 80.3400 194.9200 80.8200 ;
        RECT 193.3200 74.9000 194.9200 75.3800 ;
        RECT 193.3200 69.4600 194.9200 69.9400 ;
        RECT 205.6600 80.3400 208.6600 80.8200 ;
        RECT 205.6600 74.9000 208.6600 75.3800 ;
        RECT 205.6600 69.4600 208.6600 69.9400 ;
        RECT 193.3200 91.2200 194.9200 91.7000 ;
        RECT 193.3200 85.7800 194.9200 86.2600 ;
        RECT 205.6600 91.2200 208.6600 91.7000 ;
        RECT 205.6600 85.7800 208.6600 86.2600 ;
        RECT 193.3200 107.5400 194.9200 108.0200 ;
        RECT 193.3200 102.1000 194.9200 102.5800 ;
        RECT 193.3200 96.6600 194.9200 97.1400 ;
        RECT 205.6600 107.5400 208.6600 108.0200 ;
        RECT 205.6600 102.1000 208.6600 102.5800 ;
        RECT 205.6600 96.6600 208.6600 97.1400 ;
        RECT 1.5600 118.4200 4.5600 118.9000 ;
        RECT 1.5600 112.9800 4.5600 113.4600 ;
        RECT 13.3200 118.4200 14.9200 118.9000 ;
        RECT 13.3200 112.9800 14.9200 113.4600 ;
        RECT 1.5600 134.7400 4.5600 135.2200 ;
        RECT 1.5600 129.3000 4.5600 129.7800 ;
        RECT 1.5600 123.8600 4.5600 124.3400 ;
        RECT 13.3200 134.7400 14.9200 135.2200 ;
        RECT 13.3200 129.3000 14.9200 129.7800 ;
        RECT 13.3200 123.8600 14.9200 124.3400 ;
        RECT 1.5600 145.6200 4.5600 146.1000 ;
        RECT 1.5600 140.1800 4.5600 140.6600 ;
        RECT 13.3200 145.6200 14.9200 146.1000 ;
        RECT 13.3200 140.1800 14.9200 140.6600 ;
        RECT 1.5600 161.9400 4.5600 162.4200 ;
        RECT 1.5600 156.5000 4.5600 156.9800 ;
        RECT 1.5600 151.0600 4.5600 151.5400 ;
        RECT 13.3200 161.9400 14.9200 162.4200 ;
        RECT 13.3200 156.5000 14.9200 156.9800 ;
        RECT 13.3200 151.0600 14.9200 151.5400 ;
        RECT 58.3200 118.4200 59.9200 118.9000 ;
        RECT 58.3200 112.9800 59.9200 113.4600 ;
        RECT 58.3200 134.7400 59.9200 135.2200 ;
        RECT 58.3200 129.3000 59.9200 129.7800 ;
        RECT 58.3200 123.8600 59.9200 124.3400 ;
        RECT 103.3200 118.4200 104.9200 118.9000 ;
        RECT 103.3200 112.9800 104.9200 113.4600 ;
        RECT 103.3200 134.7400 104.9200 135.2200 ;
        RECT 103.3200 129.3000 104.9200 129.7800 ;
        RECT 103.3200 123.8600 104.9200 124.3400 ;
        RECT 58.3200 145.6200 59.9200 146.1000 ;
        RECT 58.3200 140.1800 59.9200 140.6600 ;
        RECT 58.3200 161.9400 59.9200 162.4200 ;
        RECT 58.3200 156.5000 59.9200 156.9800 ;
        RECT 58.3200 151.0600 59.9200 151.5400 ;
        RECT 103.3200 145.6200 104.9200 146.1000 ;
        RECT 103.3200 140.1800 104.9200 140.6600 ;
        RECT 103.3200 161.9400 104.9200 162.4200 ;
        RECT 103.3200 156.5000 104.9200 156.9800 ;
        RECT 103.3200 151.0600 104.9200 151.5400 ;
        RECT 13.3200 178.2600 14.9200 178.7400 ;
        RECT 1.5600 178.2600 4.5600 178.7400 ;
        RECT 1.5600 167.3800 4.5600 167.8600 ;
        RECT 1.5600 172.8200 4.5600 173.3000 ;
        RECT 13.3200 172.8200 14.9200 173.3000 ;
        RECT 13.3200 167.3800 14.9200 167.8600 ;
        RECT 1.5600 183.7000 4.5600 184.1800 ;
        RECT 1.5600 189.1400 4.5600 189.6200 ;
        RECT 13.3200 189.1400 14.9200 189.6200 ;
        RECT 13.3200 183.7000 14.9200 184.1800 ;
        RECT 13.3200 205.4600 14.9200 205.9400 ;
        RECT 1.5600 205.4600 4.5600 205.9400 ;
        RECT 1.5600 194.5800 4.5600 195.0600 ;
        RECT 1.5600 200.0200 4.5600 200.5000 ;
        RECT 13.3200 200.0200 14.9200 200.5000 ;
        RECT 13.3200 194.5800 14.9200 195.0600 ;
        RECT 58.3200 178.2600 59.9200 178.7400 ;
        RECT 58.3200 172.8200 59.9200 173.3000 ;
        RECT 58.3200 167.3800 59.9200 167.8600 ;
        RECT 58.3200 189.1400 59.9200 189.6200 ;
        RECT 58.3200 183.7000 59.9200 184.1800 ;
        RECT 103.3200 178.2600 104.9200 178.7400 ;
        RECT 103.3200 172.8200 104.9200 173.3000 ;
        RECT 103.3200 167.3800 104.9200 167.8600 ;
        RECT 103.3200 189.1400 104.9200 189.6200 ;
        RECT 103.3200 183.7000 104.9200 184.1800 ;
        RECT 58.3200 205.4600 59.9200 205.9400 ;
        RECT 58.3200 200.0200 59.9200 200.5000 ;
        RECT 58.3200 194.5800 59.9200 195.0600 ;
        RECT 103.3200 205.4600 104.9200 205.9400 ;
        RECT 103.3200 200.0200 104.9200 200.5000 ;
        RECT 103.3200 194.5800 104.9200 195.0600 ;
        RECT 148.3200 118.4200 149.9200 118.9000 ;
        RECT 148.3200 112.9800 149.9200 113.4600 ;
        RECT 148.3200 134.7400 149.9200 135.2200 ;
        RECT 148.3200 129.3000 149.9200 129.7800 ;
        RECT 148.3200 123.8600 149.9200 124.3400 ;
        RECT 148.3200 145.6200 149.9200 146.1000 ;
        RECT 148.3200 140.1800 149.9200 140.6600 ;
        RECT 148.3200 161.9400 149.9200 162.4200 ;
        RECT 148.3200 156.5000 149.9200 156.9800 ;
        RECT 148.3200 151.0600 149.9200 151.5400 ;
        RECT 193.3200 118.4200 194.9200 118.9000 ;
        RECT 193.3200 112.9800 194.9200 113.4600 ;
        RECT 205.6600 118.4200 208.6600 118.9000 ;
        RECT 205.6600 112.9800 208.6600 113.4600 ;
        RECT 193.3200 134.7400 194.9200 135.2200 ;
        RECT 193.3200 129.3000 194.9200 129.7800 ;
        RECT 193.3200 123.8600 194.9200 124.3400 ;
        RECT 205.6600 134.7400 208.6600 135.2200 ;
        RECT 205.6600 129.3000 208.6600 129.7800 ;
        RECT 205.6600 123.8600 208.6600 124.3400 ;
        RECT 193.3200 145.6200 194.9200 146.1000 ;
        RECT 193.3200 140.1800 194.9200 140.6600 ;
        RECT 205.6600 145.6200 208.6600 146.1000 ;
        RECT 205.6600 140.1800 208.6600 140.6600 ;
        RECT 193.3200 161.9400 194.9200 162.4200 ;
        RECT 193.3200 156.5000 194.9200 156.9800 ;
        RECT 193.3200 151.0600 194.9200 151.5400 ;
        RECT 205.6600 161.9400 208.6600 162.4200 ;
        RECT 205.6600 156.5000 208.6600 156.9800 ;
        RECT 205.6600 151.0600 208.6600 151.5400 ;
        RECT 148.3200 178.2600 149.9200 178.7400 ;
        RECT 148.3200 172.8200 149.9200 173.3000 ;
        RECT 148.3200 167.3800 149.9200 167.8600 ;
        RECT 148.3200 189.1400 149.9200 189.6200 ;
        RECT 148.3200 183.7000 149.9200 184.1800 ;
        RECT 148.3200 205.4600 149.9200 205.9400 ;
        RECT 148.3200 200.0200 149.9200 200.5000 ;
        RECT 148.3200 194.5800 149.9200 195.0600 ;
        RECT 193.3200 178.2600 194.9200 178.7400 ;
        RECT 205.6600 178.2600 208.6600 178.7400 ;
        RECT 193.3200 172.8200 194.9200 173.3000 ;
        RECT 193.3200 167.3800 194.9200 167.8600 ;
        RECT 205.6600 172.8200 208.6600 173.3000 ;
        RECT 205.6600 167.3800 208.6600 167.8600 ;
        RECT 193.3200 189.1400 194.9200 189.6200 ;
        RECT 193.3200 183.7000 194.9200 184.1800 ;
        RECT 205.6600 189.1400 208.6600 189.6200 ;
        RECT 205.6600 183.7000 208.6600 184.1800 ;
        RECT 193.3200 205.4600 194.9200 205.9400 ;
        RECT 205.6600 205.4600 208.6600 205.9400 ;
        RECT 193.3200 200.0200 194.9200 200.5000 ;
        RECT 193.3200 194.5800 194.9200 195.0600 ;
        RECT 205.6600 200.0200 208.6600 200.5000 ;
        RECT 205.6600 194.5800 208.6600 195.0600 ;
      LAYER met4 ;
        RECT 1.5600 1.4300 4.5600 217.5300 ;
        RECT 205.6600 1.4300 208.6600 217.5300 ;
        RECT 13.3200 1.4300 14.9200 217.5300 ;
        RECT 58.3200 1.4300 59.9200 217.5300 ;
        RECT 103.3200 1.4300 104.9200 217.5300 ;
        RECT 148.3200 1.4300 149.9200 217.5300 ;
        RECT 193.3200 1.4300 194.9200 217.5300 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.6300 218.7500 210.2200 219.6400 ;
      RECT 148.7100 218.7500 148.9100 219.6400 ;
      RECT 147.3300 218.7500 147.9900 219.6400 ;
      RECT 145.9500 218.7500 146.6100 219.6400 ;
      RECT 144.5700 218.7500 145.2300 219.6400 ;
      RECT 143.1900 218.7500 143.8500 219.6400 ;
      RECT 141.8100 218.7500 142.4700 219.6400 ;
      RECT 140.4300 218.7500 141.0900 219.6400 ;
      RECT 139.0500 218.7500 139.7100 219.6400 ;
      RECT 137.6700 218.7500 138.3300 219.6400 ;
      RECT 136.2900 218.7500 136.9500 219.6400 ;
      RECT 134.9100 218.7500 135.5700 219.6400 ;
      RECT 133.5300 218.7500 134.1900 219.6400 ;
      RECT 132.1500 218.7500 132.8100 219.6400 ;
      RECT 130.7700 218.7500 131.4300 219.6400 ;
      RECT 129.3900 218.7500 130.0500 219.6400 ;
      RECT 128.0100 218.7500 128.6700 219.6400 ;
      RECT 126.6300 218.7500 127.2900 219.6400 ;
      RECT 125.7100 218.7500 125.9100 219.6400 ;
      RECT 124.3300 218.7500 124.9900 219.6400 ;
      RECT 122.9500 218.7500 123.6100 219.6400 ;
      RECT 121.5700 218.7500 122.2300 219.6400 ;
      RECT 120.1900 218.7500 120.8500 219.6400 ;
      RECT 118.8100 218.7500 119.4700 219.6400 ;
      RECT 117.4300 218.7500 118.0900 219.6400 ;
      RECT 116.0500 218.7500 116.7100 219.6400 ;
      RECT 114.6700 218.7500 115.3300 219.6400 ;
      RECT 113.2900 218.7500 113.9500 219.6400 ;
      RECT 111.9100 218.7500 112.5700 219.6400 ;
      RECT 110.5300 218.7500 111.1900 219.6400 ;
      RECT 109.1500 218.7500 109.8100 219.6400 ;
      RECT 107.7700 218.7500 108.4300 219.6400 ;
      RECT 106.3900 218.7500 107.0500 219.6400 ;
      RECT 105.0100 218.7500 105.6700 219.6400 ;
      RECT 103.6300 218.7500 104.2900 219.6400 ;
      RECT 102.7100 218.7500 102.9100 219.6400 ;
      RECT 101.3300 218.7500 101.9900 219.6400 ;
      RECT 99.9500 218.7500 100.6100 219.6400 ;
      RECT 98.5700 218.7500 99.2300 219.6400 ;
      RECT 97.1900 218.7500 97.8500 219.6400 ;
      RECT 95.8100 218.7500 96.4700 219.6400 ;
      RECT 94.4300 218.7500 95.0900 219.6400 ;
      RECT 93.0500 218.7500 93.7100 219.6400 ;
      RECT 91.6700 218.7500 92.3300 219.6400 ;
      RECT 90.2900 218.7500 90.9500 219.6400 ;
      RECT 88.9100 218.7500 89.5700 219.6400 ;
      RECT 87.5300 218.7500 88.1900 219.6400 ;
      RECT 86.1500 218.7500 86.8100 219.6400 ;
      RECT 84.7700 218.7500 85.4300 219.6400 ;
      RECT 83.3900 218.7500 84.0500 219.6400 ;
      RECT 82.0100 218.7500 82.6700 219.6400 ;
      RECT 80.6300 218.7500 81.2900 219.6400 ;
      RECT 79.7100 218.7500 79.9100 219.6400 ;
      RECT 78.3300 218.7500 78.9900 219.6400 ;
      RECT 76.9500 218.7500 77.6100 219.6400 ;
      RECT 75.5700 218.7500 76.2300 219.6400 ;
      RECT 74.1900 218.7500 74.8500 219.6400 ;
      RECT 72.8100 218.7500 73.4700 219.6400 ;
      RECT 71.4300 218.7500 72.0900 219.6400 ;
      RECT 70.0500 218.7500 70.7100 219.6400 ;
      RECT 68.6700 218.7500 69.3300 219.6400 ;
      RECT 67.2900 218.7500 67.9500 219.6400 ;
      RECT 65.9100 218.7500 66.5700 219.6400 ;
      RECT 64.5300 218.7500 65.1900 219.6400 ;
      RECT 63.1500 218.7500 63.8100 219.6400 ;
      RECT 61.7700 218.7500 62.4300 219.6400 ;
      RECT 60.3900 218.7500 61.0500 219.6400 ;
      RECT 59.0100 218.7500 59.6700 219.6400 ;
      RECT 57.6300 218.7500 58.2900 219.6400 ;
      RECT 56.7100 218.7500 56.9100 219.6400 ;
      RECT 55.3300 218.7500 55.9900 219.6400 ;
      RECT 53.9500 218.7500 54.6100 219.6400 ;
      RECT 52.5700 218.7500 53.2300 219.6400 ;
      RECT 51.1900 218.7500 51.8500 219.6400 ;
      RECT 49.8100 218.7500 50.4700 219.6400 ;
      RECT 48.4300 218.7500 49.0900 219.6400 ;
      RECT 47.0500 218.7500 47.7100 219.6400 ;
      RECT 45.6700 218.7500 46.3300 219.6400 ;
      RECT 44.2900 218.7500 44.9500 219.6400 ;
      RECT 42.9100 218.7500 43.5700 219.6400 ;
      RECT 41.5300 218.7500 42.1900 219.6400 ;
      RECT 40.1500 218.7500 40.8100 219.6400 ;
      RECT 38.7700 218.7500 39.4300 219.6400 ;
      RECT 37.3900 218.7500 38.0500 219.6400 ;
      RECT 36.0100 218.7500 36.6700 219.6400 ;
      RECT 34.6300 218.7500 35.2900 219.6400 ;
      RECT 33.7100 218.7500 33.9100 219.6400 ;
      RECT 32.3300 218.7500 32.9900 219.6400 ;
      RECT 30.9500 218.7500 31.6100 219.6400 ;
      RECT 29.5700 218.7500 30.2300 219.6400 ;
      RECT 28.1900 218.7500 28.8500 219.6400 ;
      RECT 26.8100 218.7500 27.4700 219.6400 ;
      RECT 25.4300 218.7500 26.0900 219.6400 ;
      RECT 24.0500 218.7500 24.7100 219.6400 ;
      RECT 22.6700 218.7500 23.3300 219.6400 ;
      RECT 21.2900 218.7500 21.9500 219.6400 ;
      RECT 19.9100 218.7500 20.5700 219.6400 ;
      RECT 18.5300 218.7500 19.1900 219.6400 ;
      RECT 17.1500 218.7500 17.8100 219.6400 ;
      RECT 15.7700 218.7500 16.4300 219.6400 ;
      RECT 14.3900 218.7500 15.0500 219.6400 ;
      RECT 13.0100 218.7500 13.6700 219.6400 ;
      RECT 11.6300 218.7500 12.2900 219.6400 ;
      RECT 10.7100 218.7500 10.9100 219.6400 ;
      RECT 0.0000 218.7500 9.9900 219.6400 ;
      RECT 0.0000 0.8900 210.2200 218.7500 ;
      RECT 149.6300 0.0000 210.2200 0.8900 ;
      RECT 148.7100 0.0000 148.9100 0.8900 ;
      RECT 147.3300 0.0000 147.9900 0.8900 ;
      RECT 145.9500 0.0000 146.6100 0.8900 ;
      RECT 144.5700 0.0000 145.2300 0.8900 ;
      RECT 143.1900 0.0000 143.8500 0.8900 ;
      RECT 141.8100 0.0000 142.4700 0.8900 ;
      RECT 140.4300 0.0000 141.0900 0.8900 ;
      RECT 139.0500 0.0000 139.7100 0.8900 ;
      RECT 137.6700 0.0000 138.3300 0.8900 ;
      RECT 136.2900 0.0000 136.9500 0.8900 ;
      RECT 134.9100 0.0000 135.5700 0.8900 ;
      RECT 133.5300 0.0000 134.1900 0.8900 ;
      RECT 132.1500 0.0000 132.8100 0.8900 ;
      RECT 130.7700 0.0000 131.4300 0.8900 ;
      RECT 129.3900 0.0000 130.0500 0.8900 ;
      RECT 128.0100 0.0000 128.6700 0.8900 ;
      RECT 126.6300 0.0000 127.2900 0.8900 ;
      RECT 125.7100 0.0000 125.9100 0.8900 ;
      RECT 124.3300 0.0000 124.9900 0.8900 ;
      RECT 122.9500 0.0000 123.6100 0.8900 ;
      RECT 121.5700 0.0000 122.2300 0.8900 ;
      RECT 120.1900 0.0000 120.8500 0.8900 ;
      RECT 118.8100 0.0000 119.4700 0.8900 ;
      RECT 117.4300 0.0000 118.0900 0.8900 ;
      RECT 116.0500 0.0000 116.7100 0.8900 ;
      RECT 114.6700 0.0000 115.3300 0.8900 ;
      RECT 113.2900 0.0000 113.9500 0.8900 ;
      RECT 111.9100 0.0000 112.5700 0.8900 ;
      RECT 110.5300 0.0000 111.1900 0.8900 ;
      RECT 109.1500 0.0000 109.8100 0.8900 ;
      RECT 107.7700 0.0000 108.4300 0.8900 ;
      RECT 106.3900 0.0000 107.0500 0.8900 ;
      RECT 105.0100 0.0000 105.6700 0.8900 ;
      RECT 103.6300 0.0000 104.2900 0.8900 ;
      RECT 102.7100 0.0000 102.9100 0.8900 ;
      RECT 101.3300 0.0000 101.9900 0.8900 ;
      RECT 99.9500 0.0000 100.6100 0.8900 ;
      RECT 98.5700 0.0000 99.2300 0.8900 ;
      RECT 97.1900 0.0000 97.8500 0.8900 ;
      RECT 95.8100 0.0000 96.4700 0.8900 ;
      RECT 94.4300 0.0000 95.0900 0.8900 ;
      RECT 93.0500 0.0000 93.7100 0.8900 ;
      RECT 91.6700 0.0000 92.3300 0.8900 ;
      RECT 90.2900 0.0000 90.9500 0.8900 ;
      RECT 88.9100 0.0000 89.5700 0.8900 ;
      RECT 87.5300 0.0000 88.1900 0.8900 ;
      RECT 86.1500 0.0000 86.8100 0.8900 ;
      RECT 84.7700 0.0000 85.4300 0.8900 ;
      RECT 83.3900 0.0000 84.0500 0.8900 ;
      RECT 82.0100 0.0000 82.6700 0.8900 ;
      RECT 80.6300 0.0000 81.2900 0.8900 ;
      RECT 79.7100 0.0000 79.9100 0.8900 ;
      RECT 78.3300 0.0000 78.9900 0.8900 ;
      RECT 76.9500 0.0000 77.6100 0.8900 ;
      RECT 75.5700 0.0000 76.2300 0.8900 ;
      RECT 74.1900 0.0000 74.8500 0.8900 ;
      RECT 72.8100 0.0000 73.4700 0.8900 ;
      RECT 71.4300 0.0000 72.0900 0.8900 ;
      RECT 70.0500 0.0000 70.7100 0.8900 ;
      RECT 68.6700 0.0000 69.3300 0.8900 ;
      RECT 67.2900 0.0000 67.9500 0.8900 ;
      RECT 65.9100 0.0000 66.5700 0.8900 ;
      RECT 64.5300 0.0000 65.1900 0.8900 ;
      RECT 63.1500 0.0000 63.8100 0.8900 ;
      RECT 61.7700 0.0000 62.4300 0.8900 ;
      RECT 60.3900 0.0000 61.0500 0.8900 ;
      RECT 59.0100 0.0000 59.6700 0.8900 ;
      RECT 57.6300 0.0000 58.2900 0.8900 ;
      RECT 56.7100 0.0000 56.9100 0.8900 ;
      RECT 55.3300 0.0000 55.9900 0.8900 ;
      RECT 53.9500 0.0000 54.6100 0.8900 ;
      RECT 52.5700 0.0000 53.2300 0.8900 ;
      RECT 51.1900 0.0000 51.8500 0.8900 ;
      RECT 49.8100 0.0000 50.4700 0.8900 ;
      RECT 48.4300 0.0000 49.0900 0.8900 ;
      RECT 47.0500 0.0000 47.7100 0.8900 ;
      RECT 45.6700 0.0000 46.3300 0.8900 ;
      RECT 44.2900 0.0000 44.9500 0.8900 ;
      RECT 42.9100 0.0000 43.5700 0.8900 ;
      RECT 41.5300 0.0000 42.1900 0.8900 ;
      RECT 40.1500 0.0000 40.8100 0.8900 ;
      RECT 38.7700 0.0000 39.4300 0.8900 ;
      RECT 37.3900 0.0000 38.0500 0.8900 ;
      RECT 36.0100 0.0000 36.6700 0.8900 ;
      RECT 34.6300 0.0000 35.2900 0.8900 ;
      RECT 33.7100 0.0000 33.9100 0.8900 ;
      RECT 32.3300 0.0000 32.9900 0.8900 ;
      RECT 30.9500 0.0000 31.6100 0.8900 ;
      RECT 29.5700 0.0000 30.2300 0.8900 ;
      RECT 28.1900 0.0000 28.8500 0.8900 ;
      RECT 26.8100 0.0000 27.4700 0.8900 ;
      RECT 25.4300 0.0000 26.0900 0.8900 ;
      RECT 24.0500 0.0000 24.7100 0.8900 ;
      RECT 22.6700 0.0000 23.3300 0.8900 ;
      RECT 21.2900 0.0000 21.9500 0.8900 ;
      RECT 19.9100 0.0000 20.5700 0.8900 ;
      RECT 18.5300 0.0000 19.1900 0.8900 ;
      RECT 17.1500 0.0000 17.8100 0.8900 ;
      RECT 15.7700 0.0000 16.4300 0.8900 ;
      RECT 14.3900 0.0000 15.0500 0.8900 ;
      RECT 13.0100 0.0000 13.6700 0.8900 ;
      RECT 11.6300 0.0000 12.2900 0.8900 ;
      RECT 10.7100 0.0000 10.9100 0.8900 ;
      RECT 0.0000 0.0000 9.9900 0.8900 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 210.2200 219.6400 ;
    LAYER met2 ;
      RECT 199.7400 218.7800 210.2200 219.6400 ;
      RECT 197.9000 218.7800 199.0800 219.6400 ;
      RECT 195.1400 218.7800 197.2400 219.6400 ;
      RECT 193.3000 218.7800 194.4800 219.6400 ;
      RECT 191.0000 218.7800 192.6400 219.6400 ;
      RECT 188.7000 218.7800 190.3400 219.6400 ;
      RECT 186.4000 218.7800 188.0400 219.6400 ;
      RECT 184.5600 218.7800 185.7400 219.6400 ;
      RECT 181.8000 218.7800 183.9000 219.6400 ;
      RECT 179.9600 218.7800 181.1400 219.6400 ;
      RECT 177.6600 218.7800 179.3000 219.6400 ;
      RECT 175.3600 218.7800 177.0000 219.6400 ;
      RECT 173.0600 218.7800 174.7000 219.6400 ;
      RECT 170.7600 218.7800 172.4000 219.6400 ;
      RECT 168.9200 218.7800 170.1000 219.6400 ;
      RECT 166.6200 218.7800 168.2600 219.6400 ;
      RECT 164.3200 218.7800 165.9600 219.6400 ;
      RECT 162.0200 218.7800 163.6600 219.6400 ;
      RECT 159.7200 218.7800 161.3600 219.6400 ;
      RECT 156.9600 218.7800 159.0600 219.6400 ;
      RECT 155.5800 218.7800 156.3000 219.6400 ;
      RECT 0.0000 218.7800 154.9200 219.6400 ;
      RECT 0.0000 209.9400 210.2200 218.7800 ;
      RECT 0.8600 209.2800 209.3600 209.9400 ;
      RECT 0.0000 208.2400 210.2200 209.2800 ;
      RECT 0.8600 207.5800 209.3600 208.2400 ;
      RECT 0.0000 206.5400 210.2200 207.5800 ;
      RECT 0.8600 205.8800 209.3600 206.5400 ;
      RECT 0.0000 204.8400 210.2200 205.8800 ;
      RECT 0.8600 204.1800 209.3600 204.8400 ;
      RECT 0.0000 203.1400 210.2200 204.1800 ;
      RECT 0.8600 202.4800 209.3600 203.1400 ;
      RECT 0.0000 201.4400 210.2200 202.4800 ;
      RECT 0.8600 200.7800 209.3600 201.4400 ;
      RECT 0.0000 199.4000 210.2200 200.7800 ;
      RECT 0.8600 198.7400 209.3600 199.4000 ;
      RECT 0.0000 197.7000 210.2200 198.7400 ;
      RECT 0.8600 197.0400 209.3600 197.7000 ;
      RECT 0.0000 196.0000 210.2200 197.0400 ;
      RECT 0.8600 195.3400 209.3600 196.0000 ;
      RECT 0.0000 194.3000 210.2200 195.3400 ;
      RECT 0.8600 193.6400 209.3600 194.3000 ;
      RECT 0.0000 192.6000 210.2200 193.6400 ;
      RECT 0.8600 191.9400 209.3600 192.6000 ;
      RECT 0.0000 190.5600 210.2200 191.9400 ;
      RECT 0.8600 189.9000 209.3600 190.5600 ;
      RECT 0.0000 188.8600 210.2200 189.9000 ;
      RECT 0.8600 188.2000 209.3600 188.8600 ;
      RECT 0.0000 187.1600 210.2200 188.2000 ;
      RECT 0.8600 186.5000 209.3600 187.1600 ;
      RECT 0.0000 185.4600 210.2200 186.5000 ;
      RECT 0.8600 184.8000 209.3600 185.4600 ;
      RECT 0.0000 183.7600 210.2200 184.8000 ;
      RECT 0.8600 183.1000 209.3600 183.7600 ;
      RECT 0.0000 181.7200 210.2200 183.1000 ;
      RECT 0.8600 181.0600 209.3600 181.7200 ;
      RECT 0.0000 180.0200 210.2200 181.0600 ;
      RECT 0.8600 179.3600 209.3600 180.0200 ;
      RECT 0.0000 178.3200 210.2200 179.3600 ;
      RECT 0.8600 177.6600 209.3600 178.3200 ;
      RECT 0.0000 176.6200 210.2200 177.6600 ;
      RECT 0.8600 175.9600 209.3600 176.6200 ;
      RECT 0.0000 174.9200 210.2200 175.9600 ;
      RECT 0.8600 174.2600 209.3600 174.9200 ;
      RECT 0.0000 172.8800 210.2200 174.2600 ;
      RECT 0.8600 172.2200 209.3600 172.8800 ;
      RECT 0.0000 171.1800 210.2200 172.2200 ;
      RECT 0.8600 170.5200 209.3600 171.1800 ;
      RECT 0.0000 169.4800 210.2200 170.5200 ;
      RECT 0.8600 168.8200 209.3600 169.4800 ;
      RECT 0.0000 167.7800 210.2200 168.8200 ;
      RECT 0.8600 167.1200 209.3600 167.7800 ;
      RECT 0.0000 166.0800 210.2200 167.1200 ;
      RECT 0.8600 165.4200 209.3600 166.0800 ;
      RECT 0.0000 164.0400 210.2200 165.4200 ;
      RECT 0.8600 163.3800 209.3600 164.0400 ;
      RECT 0.0000 162.3400 210.2200 163.3800 ;
      RECT 0.8600 161.6800 209.3600 162.3400 ;
      RECT 0.0000 160.6400 210.2200 161.6800 ;
      RECT 0.8600 159.9800 209.3600 160.6400 ;
      RECT 0.0000 158.9400 210.2200 159.9800 ;
      RECT 0.8600 158.2800 209.3600 158.9400 ;
      RECT 0.0000 157.2400 210.2200 158.2800 ;
      RECT 0.8600 156.5800 209.3600 157.2400 ;
      RECT 0.0000 155.5400 210.2200 156.5800 ;
      RECT 0.8600 154.8800 209.3600 155.5400 ;
      RECT 0.0000 150.1000 210.2200 154.8800 ;
      RECT 0.8600 149.4400 209.3600 150.1000 ;
      RECT 0.0000 148.4000 210.2200 149.4400 ;
      RECT 0.8600 147.7400 209.3600 148.4000 ;
      RECT 0.0000 147.0400 210.2200 147.7400 ;
      RECT 0.8600 146.3800 209.3600 147.0400 ;
      RECT 0.0000 145.6800 210.2200 146.3800 ;
      RECT 0.8600 145.0200 209.3600 145.6800 ;
      RECT 0.0000 143.9800 210.2200 145.0200 ;
      RECT 0.8600 143.3200 209.3600 143.9800 ;
      RECT 0.0000 142.6200 210.2200 143.3200 ;
      RECT 0.8600 141.9600 209.3600 142.6200 ;
      RECT 0.0000 141.2600 210.2200 141.9600 ;
      RECT 0.8600 140.6000 209.3600 141.2600 ;
      RECT 0.0000 139.5600 210.2200 140.6000 ;
      RECT 0.8600 138.9000 209.3600 139.5600 ;
      RECT 0.0000 138.2000 210.2200 138.9000 ;
      RECT 0.8600 137.5400 209.3600 138.2000 ;
      RECT 0.0000 136.8400 210.2200 137.5400 ;
      RECT 0.8600 136.1800 209.3600 136.8400 ;
      RECT 0.0000 135.1400 210.2200 136.1800 ;
      RECT 0.8600 134.4800 209.3600 135.1400 ;
      RECT 0.0000 133.7800 210.2200 134.4800 ;
      RECT 0.8600 133.1200 209.3600 133.7800 ;
      RECT 0.0000 132.4200 210.2200 133.1200 ;
      RECT 0.8600 131.7600 209.3600 132.4200 ;
      RECT 0.0000 130.7200 210.2200 131.7600 ;
      RECT 0.8600 130.0600 209.3600 130.7200 ;
      RECT 0.0000 129.3600 210.2200 130.0600 ;
      RECT 0.8600 128.7000 209.3600 129.3600 ;
      RECT 0.0000 128.0000 210.2200 128.7000 ;
      RECT 0.8600 127.3400 209.3600 128.0000 ;
      RECT 0.0000 126.3000 210.2200 127.3400 ;
      RECT 0.8600 125.6400 209.3600 126.3000 ;
      RECT 0.0000 124.9400 210.2200 125.6400 ;
      RECT 0.8600 124.2800 209.3600 124.9400 ;
      RECT 0.0000 123.5800 210.2200 124.2800 ;
      RECT 0.8600 122.9200 209.3600 123.5800 ;
      RECT 0.0000 121.8800 210.2200 122.9200 ;
      RECT 0.8600 121.2200 209.3600 121.8800 ;
      RECT 0.0000 120.5200 210.2200 121.2200 ;
      RECT 0.8600 119.8600 209.3600 120.5200 ;
      RECT 0.0000 119.1600 210.2200 119.8600 ;
      RECT 0.8600 118.5000 209.3600 119.1600 ;
      RECT 0.0000 117.4600 210.2200 118.5000 ;
      RECT 0.8600 116.8000 209.3600 117.4600 ;
      RECT 0.0000 116.1000 210.2200 116.8000 ;
      RECT 0.8600 115.4400 209.3600 116.1000 ;
      RECT 0.0000 114.7400 210.2200 115.4400 ;
      RECT 0.8600 114.0800 209.3600 114.7400 ;
      RECT 0.0000 113.0400 210.2200 114.0800 ;
      RECT 0.8600 112.3800 209.3600 113.0400 ;
      RECT 0.0000 111.6800 210.2200 112.3800 ;
      RECT 0.8600 111.0200 209.3600 111.6800 ;
      RECT 0.0000 110.3200 210.2200 111.0200 ;
      RECT 0.8600 109.6600 209.3600 110.3200 ;
      RECT 0.0000 108.6200 210.2200 109.6600 ;
      RECT 0.8600 107.9600 209.3600 108.6200 ;
      RECT 0.0000 107.2600 210.2200 107.9600 ;
      RECT 0.8600 106.6000 209.3600 107.2600 ;
      RECT 0.0000 105.9000 210.2200 106.6000 ;
      RECT 0.8600 105.2400 209.3600 105.9000 ;
      RECT 0.0000 104.2000 210.2200 105.2400 ;
      RECT 0.8600 103.5400 209.3600 104.2000 ;
      RECT 0.0000 102.8400 210.2200 103.5400 ;
      RECT 0.8600 102.1800 209.3600 102.8400 ;
      RECT 0.0000 101.4800 210.2200 102.1800 ;
      RECT 0.8600 100.8200 209.3600 101.4800 ;
      RECT 0.0000 99.7800 210.2200 100.8200 ;
      RECT 0.8600 99.1200 209.3600 99.7800 ;
      RECT 0.0000 98.4200 210.2200 99.1200 ;
      RECT 0.8600 97.7600 209.3600 98.4200 ;
      RECT 0.0000 97.0600 210.2200 97.7600 ;
      RECT 0.8600 96.4000 209.3600 97.0600 ;
      RECT 0.0000 95.3600 210.2200 96.4000 ;
      RECT 0.8600 94.7000 209.3600 95.3600 ;
      RECT 0.0000 94.0000 210.2200 94.7000 ;
      RECT 0.8600 93.3400 209.3600 94.0000 ;
      RECT 0.0000 92.6400 210.2200 93.3400 ;
      RECT 0.8600 91.9800 209.3600 92.6400 ;
      RECT 0.0000 90.9400 210.2200 91.9800 ;
      RECT 0.8600 90.2800 209.3600 90.9400 ;
      RECT 0.0000 89.5800 210.2200 90.2800 ;
      RECT 0.8600 88.9200 209.3600 89.5800 ;
      RECT 0.0000 88.2200 210.2200 88.9200 ;
      RECT 0.8600 87.5600 209.3600 88.2200 ;
      RECT 0.0000 86.5200 210.2200 87.5600 ;
      RECT 0.8600 85.8600 209.3600 86.5200 ;
      RECT 0.0000 85.1600 210.2200 85.8600 ;
      RECT 0.8600 84.5000 209.3600 85.1600 ;
      RECT 0.0000 83.8000 210.2200 84.5000 ;
      RECT 0.8600 83.1400 209.3600 83.8000 ;
      RECT 0.0000 82.1000 210.2200 83.1400 ;
      RECT 0.8600 81.4400 209.3600 82.1000 ;
      RECT 0.0000 80.7400 210.2200 81.4400 ;
      RECT 0.8600 80.0800 209.3600 80.7400 ;
      RECT 0.0000 79.3800 210.2200 80.0800 ;
      RECT 0.8600 78.7200 209.3600 79.3800 ;
      RECT 0.0000 78.0200 210.2200 78.7200 ;
      RECT 0.8600 77.3600 209.3600 78.0200 ;
      RECT 0.0000 76.3200 210.2200 77.3600 ;
      RECT 0.8600 75.6600 209.3600 76.3200 ;
      RECT 0.0000 74.9600 210.2200 75.6600 ;
      RECT 0.8600 74.3000 209.3600 74.9600 ;
      RECT 0.0000 73.6000 210.2200 74.3000 ;
      RECT 0.8600 72.9400 209.3600 73.6000 ;
      RECT 0.0000 71.9000 210.2200 72.9400 ;
      RECT 0.8600 71.2400 209.3600 71.9000 ;
      RECT 0.0000 70.5400 210.2200 71.2400 ;
      RECT 0.8600 69.8800 209.3600 70.5400 ;
      RECT 0.0000 69.1800 210.2200 69.8800 ;
      RECT 0.8600 68.5200 209.3600 69.1800 ;
      RECT 0.0000 67.4800 210.2200 68.5200 ;
      RECT 0.8600 66.8200 209.3600 67.4800 ;
      RECT 0.0000 66.1200 210.2200 66.8200 ;
      RECT 0.8600 65.4600 209.3600 66.1200 ;
      RECT 0.0000 64.7600 210.2200 65.4600 ;
      RECT 0.8600 64.1000 209.3600 64.7600 ;
      RECT 0.0000 63.0600 210.2200 64.1000 ;
      RECT 0.8600 62.4000 209.3600 63.0600 ;
      RECT 0.0000 61.7000 210.2200 62.4000 ;
      RECT 0.8600 61.0400 209.3600 61.7000 ;
      RECT 0.0000 60.3400 210.2200 61.0400 ;
      RECT 0.8600 59.6800 209.3600 60.3400 ;
      RECT 0.0000 58.6400 210.2200 59.6800 ;
      RECT 0.8600 57.9800 209.3600 58.6400 ;
      RECT 0.0000 57.2800 210.2200 57.9800 ;
      RECT 0.8600 56.6200 209.3600 57.2800 ;
      RECT 0.0000 55.9200 210.2200 56.6200 ;
      RECT 0.8600 55.2600 209.3600 55.9200 ;
      RECT 0.0000 54.2200 210.2200 55.2600 ;
      RECT 0.8600 53.5600 209.3600 54.2200 ;
      RECT 0.0000 52.8600 210.2200 53.5600 ;
      RECT 0.8600 52.2000 209.3600 52.8600 ;
      RECT 0.0000 51.5000 210.2200 52.2000 ;
      RECT 0.8600 50.8400 209.3600 51.5000 ;
      RECT 0.0000 49.8000 210.2200 50.8400 ;
      RECT 0.8600 49.1400 209.3600 49.8000 ;
      RECT 0.0000 48.4400 210.2200 49.1400 ;
      RECT 0.8600 47.7800 209.3600 48.4400 ;
      RECT 0.0000 47.0800 210.2200 47.7800 ;
      RECT 0.8600 46.4200 209.3600 47.0800 ;
      RECT 0.0000 45.3800 210.2200 46.4200 ;
      RECT 0.8600 44.7200 209.3600 45.3800 ;
      RECT 0.0000 44.0200 210.2200 44.7200 ;
      RECT 0.8600 43.3600 209.3600 44.0200 ;
      RECT 0.0000 42.6600 210.2200 43.3600 ;
      RECT 0.8600 42.0000 209.3600 42.6600 ;
      RECT 0.0000 40.9600 210.2200 42.0000 ;
      RECT 0.8600 40.3000 209.3600 40.9600 ;
      RECT 0.0000 39.6000 210.2200 40.3000 ;
      RECT 0.8600 38.9400 209.3600 39.6000 ;
      RECT 0.0000 38.2400 210.2200 38.9400 ;
      RECT 0.8600 37.5800 209.3600 38.2400 ;
      RECT 0.0000 36.5400 210.2200 37.5800 ;
      RECT 0.8600 35.8800 209.3600 36.5400 ;
      RECT 0.0000 35.1800 210.2200 35.8800 ;
      RECT 0.8600 34.5200 209.3600 35.1800 ;
      RECT 0.0000 33.8200 210.2200 34.5200 ;
      RECT 0.8600 33.1600 209.3600 33.8200 ;
      RECT 0.0000 32.1200 210.2200 33.1600 ;
      RECT 0.8600 31.4600 209.3600 32.1200 ;
      RECT 0.0000 30.7600 210.2200 31.4600 ;
      RECT 0.8600 30.1000 209.3600 30.7600 ;
      RECT 0.0000 29.4000 210.2200 30.1000 ;
      RECT 0.8600 28.7400 209.3600 29.4000 ;
      RECT 0.0000 27.7000 210.2200 28.7400 ;
      RECT 0.8600 27.0400 209.3600 27.7000 ;
      RECT 0.0000 26.3400 210.2200 27.0400 ;
      RECT 0.8600 25.6800 209.3600 26.3400 ;
      RECT 0.0000 24.9800 210.2200 25.6800 ;
      RECT 0.8600 24.3200 209.3600 24.9800 ;
      RECT 0.0000 23.2800 210.2200 24.3200 ;
      RECT 0.8600 22.6200 209.3600 23.2800 ;
      RECT 0.0000 21.9200 210.2200 22.6200 ;
      RECT 0.8600 21.2600 209.3600 21.9200 ;
      RECT 0.0000 20.5600 210.2200 21.2600 ;
      RECT 0.8600 19.9000 209.3600 20.5600 ;
      RECT 0.0000 18.8600 210.2200 19.9000 ;
      RECT 0.8600 18.2000 209.3600 18.8600 ;
      RECT 0.0000 17.5000 210.2200 18.2000 ;
      RECT 0.8600 16.8400 209.3600 17.5000 ;
      RECT 0.0000 16.1400 210.2200 16.8400 ;
      RECT 0.8600 15.4800 209.3600 16.1400 ;
      RECT 0.0000 14.4400 210.2200 15.4800 ;
      RECT 0.8600 13.7800 209.3600 14.4400 ;
      RECT 0.0000 13.0800 210.2200 13.7800 ;
      RECT 0.8600 12.4200 209.3600 13.0800 ;
      RECT 0.0000 11.7200 210.2200 12.4200 ;
      RECT 0.8600 11.0600 209.3600 11.7200 ;
      RECT 0.0000 10.3600 210.2200 11.0600 ;
      RECT 0.8600 9.7000 209.3600 10.3600 ;
      RECT 0.0000 0.8600 210.2200 9.7000 ;
      RECT 199.7400 0.0000 210.2200 0.8600 ;
      RECT 197.9000 0.0000 199.0800 0.8600 ;
      RECT 195.6000 0.0000 197.2400 0.8600 ;
      RECT 193.3000 0.0000 194.9400 0.8600 ;
      RECT 191.0000 0.0000 192.6400 0.8600 ;
      RECT 188.7000 0.0000 190.3400 0.8600 ;
      RECT 185.9400 0.0000 188.0400 0.8600 ;
      RECT 184.5600 0.0000 185.2800 0.8600 ;
      RECT 181.8000 0.0000 183.9000 0.8600 ;
      RECT 179.9600 0.0000 181.1400 0.8600 ;
      RECT 177.6600 0.0000 179.3000 0.8600 ;
      RECT 175.3600 0.0000 177.0000 0.8600 ;
      RECT 173.0600 0.0000 174.7000 0.8600 ;
      RECT 170.7600 0.0000 172.4000 0.8600 ;
      RECT 168.9200 0.0000 170.1000 0.8600 ;
      RECT 166.6200 0.0000 168.2600 0.8600 ;
      RECT 164.3200 0.0000 165.9600 0.8600 ;
      RECT 161.5600 0.0000 163.6600 0.8600 ;
      RECT 159.7200 0.0000 160.9000 0.8600 ;
      RECT 157.4200 0.0000 159.0600 0.8600 ;
      RECT 155.5800 0.0000 156.7600 0.8600 ;
      RECT 0.0000 0.0000 154.9200 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 217.8300 210.2200 219.6400 ;
      RECT 208.9600 214.2300 210.2200 217.8300 ;
      RECT 0.0000 214.2300 1.2600 217.8300 ;
      RECT 0.0000 213.8300 210.2200 214.2300 ;
      RECT 204.9600 210.2300 210.2200 213.8300 ;
      RECT 0.0000 210.2300 5.2600 213.8300 ;
      RECT 0.0000 208.9600 210.2200 210.2300 ;
      RECT 204.9600 207.8800 210.2200 208.9600 ;
      RECT 192.0200 207.8800 201.3600 208.9600 ;
      RECT 147.0200 207.8800 189.8200 208.9600 ;
      RECT 102.0200 207.8800 144.8200 208.9600 ;
      RECT 57.0200 207.8800 99.8200 208.9600 ;
      RECT 8.8600 207.8800 54.8200 208.9600 ;
      RECT 0.0000 207.8800 5.2600 208.9600 ;
      RECT 0.0000 206.2400 210.2200 207.8800 ;
      RECT 208.9600 205.1600 210.2200 206.2400 ;
      RECT 195.2200 205.1600 205.3600 206.2400 ;
      RECT 150.2200 205.1600 193.0200 206.2400 ;
      RECT 105.2200 205.1600 148.0200 206.2400 ;
      RECT 60.2200 205.1600 103.0200 206.2400 ;
      RECT 15.2200 205.1600 58.0200 206.2400 ;
      RECT 4.8600 205.1600 13.0200 206.2400 ;
      RECT 0.0000 205.1600 1.2600 206.2400 ;
      RECT 0.0000 203.5200 210.2200 205.1600 ;
      RECT 204.9600 202.4400 210.2200 203.5200 ;
      RECT 192.0200 202.4400 201.3600 203.5200 ;
      RECT 147.0200 202.4400 189.8200 203.5200 ;
      RECT 102.0200 202.4400 144.8200 203.5200 ;
      RECT 57.0200 202.4400 99.8200 203.5200 ;
      RECT 8.8600 202.4400 54.8200 203.5200 ;
      RECT 0.0000 202.4400 5.2600 203.5200 ;
      RECT 0.0000 200.8000 210.2200 202.4400 ;
      RECT 208.9600 199.7200 210.2200 200.8000 ;
      RECT 195.2200 199.7200 205.3600 200.8000 ;
      RECT 150.2200 199.7200 193.0200 200.8000 ;
      RECT 105.2200 199.7200 148.0200 200.8000 ;
      RECT 60.2200 199.7200 103.0200 200.8000 ;
      RECT 15.2200 199.7200 58.0200 200.8000 ;
      RECT 4.8600 199.7200 13.0200 200.8000 ;
      RECT 0.0000 199.7200 1.2600 200.8000 ;
      RECT 0.0000 198.0800 210.2200 199.7200 ;
      RECT 204.9600 197.0000 210.2200 198.0800 ;
      RECT 192.0200 197.0000 201.3600 198.0800 ;
      RECT 147.0200 197.0000 189.8200 198.0800 ;
      RECT 102.0200 197.0000 144.8200 198.0800 ;
      RECT 57.0200 197.0000 99.8200 198.0800 ;
      RECT 8.8600 197.0000 54.8200 198.0800 ;
      RECT 0.0000 197.0000 5.2600 198.0800 ;
      RECT 0.0000 195.3600 210.2200 197.0000 ;
      RECT 208.9600 194.2800 210.2200 195.3600 ;
      RECT 195.2200 194.2800 205.3600 195.3600 ;
      RECT 150.2200 194.2800 193.0200 195.3600 ;
      RECT 105.2200 194.2800 148.0200 195.3600 ;
      RECT 60.2200 194.2800 103.0200 195.3600 ;
      RECT 15.2200 194.2800 58.0200 195.3600 ;
      RECT 4.8600 194.2800 13.0200 195.3600 ;
      RECT 0.0000 194.2800 1.2600 195.3600 ;
      RECT 0.0000 192.6400 210.2200 194.2800 ;
      RECT 204.9600 191.5600 210.2200 192.6400 ;
      RECT 192.0200 191.5600 201.3600 192.6400 ;
      RECT 147.0200 191.5600 189.8200 192.6400 ;
      RECT 102.0200 191.5600 144.8200 192.6400 ;
      RECT 57.0200 191.5600 99.8200 192.6400 ;
      RECT 8.8600 191.5600 54.8200 192.6400 ;
      RECT 0.0000 191.5600 5.2600 192.6400 ;
      RECT 0.0000 189.9200 210.2200 191.5600 ;
      RECT 208.9600 188.8400 210.2200 189.9200 ;
      RECT 195.2200 188.8400 205.3600 189.9200 ;
      RECT 150.2200 188.8400 193.0200 189.9200 ;
      RECT 105.2200 188.8400 148.0200 189.9200 ;
      RECT 60.2200 188.8400 103.0200 189.9200 ;
      RECT 15.2200 188.8400 58.0200 189.9200 ;
      RECT 4.8600 188.8400 13.0200 189.9200 ;
      RECT 0.0000 188.8400 1.2600 189.9200 ;
      RECT 0.0000 187.2000 210.2200 188.8400 ;
      RECT 204.9600 186.1200 210.2200 187.2000 ;
      RECT 192.0200 186.1200 201.3600 187.2000 ;
      RECT 147.0200 186.1200 189.8200 187.2000 ;
      RECT 102.0200 186.1200 144.8200 187.2000 ;
      RECT 57.0200 186.1200 99.8200 187.2000 ;
      RECT 8.8600 186.1200 54.8200 187.2000 ;
      RECT 0.0000 186.1200 5.2600 187.2000 ;
      RECT 0.0000 184.4800 210.2200 186.1200 ;
      RECT 208.9600 183.4000 210.2200 184.4800 ;
      RECT 195.2200 183.4000 205.3600 184.4800 ;
      RECT 150.2200 183.4000 193.0200 184.4800 ;
      RECT 105.2200 183.4000 148.0200 184.4800 ;
      RECT 60.2200 183.4000 103.0200 184.4800 ;
      RECT 15.2200 183.4000 58.0200 184.4800 ;
      RECT 4.8600 183.4000 13.0200 184.4800 ;
      RECT 0.0000 183.4000 1.2600 184.4800 ;
      RECT 0.0000 181.7600 210.2200 183.4000 ;
      RECT 204.9600 180.6800 210.2200 181.7600 ;
      RECT 192.0200 180.6800 201.3600 181.7600 ;
      RECT 147.0200 180.6800 189.8200 181.7600 ;
      RECT 102.0200 180.6800 144.8200 181.7600 ;
      RECT 57.0200 180.6800 99.8200 181.7600 ;
      RECT 8.8600 180.6800 54.8200 181.7600 ;
      RECT 0.0000 180.6800 5.2600 181.7600 ;
      RECT 0.0000 179.0400 210.2200 180.6800 ;
      RECT 208.9600 177.9600 210.2200 179.0400 ;
      RECT 195.2200 177.9600 205.3600 179.0400 ;
      RECT 150.2200 177.9600 193.0200 179.0400 ;
      RECT 105.2200 177.9600 148.0200 179.0400 ;
      RECT 60.2200 177.9600 103.0200 179.0400 ;
      RECT 15.2200 177.9600 58.0200 179.0400 ;
      RECT 4.8600 177.9600 13.0200 179.0400 ;
      RECT 0.0000 177.9600 1.2600 179.0400 ;
      RECT 0.0000 176.3200 210.2200 177.9600 ;
      RECT 204.9600 175.2400 210.2200 176.3200 ;
      RECT 192.0200 175.2400 201.3600 176.3200 ;
      RECT 147.0200 175.2400 189.8200 176.3200 ;
      RECT 102.0200 175.2400 144.8200 176.3200 ;
      RECT 57.0200 175.2400 99.8200 176.3200 ;
      RECT 8.8600 175.2400 54.8200 176.3200 ;
      RECT 0.0000 175.2400 5.2600 176.3200 ;
      RECT 0.0000 173.6000 210.2200 175.2400 ;
      RECT 208.9600 172.5200 210.2200 173.6000 ;
      RECT 195.2200 172.5200 205.3600 173.6000 ;
      RECT 150.2200 172.5200 193.0200 173.6000 ;
      RECT 105.2200 172.5200 148.0200 173.6000 ;
      RECT 60.2200 172.5200 103.0200 173.6000 ;
      RECT 15.2200 172.5200 58.0200 173.6000 ;
      RECT 4.8600 172.5200 13.0200 173.6000 ;
      RECT 0.0000 172.5200 1.2600 173.6000 ;
      RECT 0.0000 170.8800 210.2200 172.5200 ;
      RECT 204.9600 169.8000 210.2200 170.8800 ;
      RECT 192.0200 169.8000 201.3600 170.8800 ;
      RECT 147.0200 169.8000 189.8200 170.8800 ;
      RECT 102.0200 169.8000 144.8200 170.8800 ;
      RECT 57.0200 169.8000 99.8200 170.8800 ;
      RECT 8.8600 169.8000 54.8200 170.8800 ;
      RECT 0.0000 169.8000 5.2600 170.8800 ;
      RECT 0.0000 168.1600 210.2200 169.8000 ;
      RECT 208.9600 167.0800 210.2200 168.1600 ;
      RECT 195.2200 167.0800 205.3600 168.1600 ;
      RECT 150.2200 167.0800 193.0200 168.1600 ;
      RECT 105.2200 167.0800 148.0200 168.1600 ;
      RECT 60.2200 167.0800 103.0200 168.1600 ;
      RECT 15.2200 167.0800 58.0200 168.1600 ;
      RECT 4.8600 167.0800 13.0200 168.1600 ;
      RECT 0.0000 167.0800 1.2600 168.1600 ;
      RECT 0.0000 165.4400 210.2200 167.0800 ;
      RECT 204.9600 164.3600 210.2200 165.4400 ;
      RECT 192.0200 164.3600 201.3600 165.4400 ;
      RECT 147.0200 164.3600 189.8200 165.4400 ;
      RECT 102.0200 164.3600 144.8200 165.4400 ;
      RECT 57.0200 164.3600 99.8200 165.4400 ;
      RECT 8.8600 164.3600 54.8200 165.4400 ;
      RECT 0.0000 164.3600 5.2600 165.4400 ;
      RECT 0.0000 162.7200 210.2200 164.3600 ;
      RECT 208.9600 161.6400 210.2200 162.7200 ;
      RECT 195.2200 161.6400 205.3600 162.7200 ;
      RECT 150.2200 161.6400 193.0200 162.7200 ;
      RECT 105.2200 161.6400 148.0200 162.7200 ;
      RECT 60.2200 161.6400 103.0200 162.7200 ;
      RECT 15.2200 161.6400 58.0200 162.7200 ;
      RECT 4.8600 161.6400 13.0200 162.7200 ;
      RECT 0.0000 161.6400 1.2600 162.7200 ;
      RECT 0.0000 160.0000 210.2200 161.6400 ;
      RECT 204.9600 158.9200 210.2200 160.0000 ;
      RECT 192.0200 158.9200 201.3600 160.0000 ;
      RECT 147.0200 158.9200 189.8200 160.0000 ;
      RECT 102.0200 158.9200 144.8200 160.0000 ;
      RECT 57.0200 158.9200 99.8200 160.0000 ;
      RECT 8.8600 158.9200 54.8200 160.0000 ;
      RECT 0.0000 158.9200 5.2600 160.0000 ;
      RECT 0.0000 157.2800 210.2200 158.9200 ;
      RECT 208.9600 156.2000 210.2200 157.2800 ;
      RECT 195.2200 156.2000 205.3600 157.2800 ;
      RECT 150.2200 156.2000 193.0200 157.2800 ;
      RECT 105.2200 156.2000 148.0200 157.2800 ;
      RECT 60.2200 156.2000 103.0200 157.2800 ;
      RECT 15.2200 156.2000 58.0200 157.2800 ;
      RECT 4.8600 156.2000 13.0200 157.2800 ;
      RECT 0.0000 156.2000 1.2600 157.2800 ;
      RECT 0.0000 154.5600 210.2200 156.2000 ;
      RECT 204.9600 153.4800 210.2200 154.5600 ;
      RECT 192.0200 153.4800 201.3600 154.5600 ;
      RECT 147.0200 153.4800 189.8200 154.5600 ;
      RECT 102.0200 153.4800 144.8200 154.5600 ;
      RECT 57.0200 153.4800 99.8200 154.5600 ;
      RECT 8.8600 153.4800 54.8200 154.5600 ;
      RECT 0.0000 153.4800 5.2600 154.5600 ;
      RECT 0.0000 151.8400 210.2200 153.4800 ;
      RECT 208.9600 150.7600 210.2200 151.8400 ;
      RECT 195.2200 150.7600 205.3600 151.8400 ;
      RECT 150.2200 150.7600 193.0200 151.8400 ;
      RECT 105.2200 150.7600 148.0200 151.8400 ;
      RECT 60.2200 150.7600 103.0200 151.8400 ;
      RECT 15.2200 150.7600 58.0200 151.8400 ;
      RECT 4.8600 150.7600 13.0200 151.8400 ;
      RECT 0.0000 150.7600 1.2600 151.8400 ;
      RECT 0.0000 149.1200 210.2200 150.7600 ;
      RECT 204.9600 148.0400 210.2200 149.1200 ;
      RECT 192.0200 148.0400 201.3600 149.1200 ;
      RECT 147.0200 148.0400 189.8200 149.1200 ;
      RECT 102.0200 148.0400 144.8200 149.1200 ;
      RECT 57.0200 148.0400 99.8200 149.1200 ;
      RECT 8.8600 148.0400 54.8200 149.1200 ;
      RECT 0.0000 148.0400 5.2600 149.1200 ;
      RECT 0.0000 146.4000 210.2200 148.0400 ;
      RECT 208.9600 145.3200 210.2200 146.4000 ;
      RECT 195.2200 145.3200 205.3600 146.4000 ;
      RECT 150.2200 145.3200 193.0200 146.4000 ;
      RECT 105.2200 145.3200 148.0200 146.4000 ;
      RECT 60.2200 145.3200 103.0200 146.4000 ;
      RECT 15.2200 145.3200 58.0200 146.4000 ;
      RECT 4.8600 145.3200 13.0200 146.4000 ;
      RECT 0.0000 145.3200 1.2600 146.4000 ;
      RECT 0.0000 143.6800 210.2200 145.3200 ;
      RECT 204.9600 142.6000 210.2200 143.6800 ;
      RECT 192.0200 142.6000 201.3600 143.6800 ;
      RECT 147.0200 142.6000 189.8200 143.6800 ;
      RECT 102.0200 142.6000 144.8200 143.6800 ;
      RECT 57.0200 142.6000 99.8200 143.6800 ;
      RECT 8.8600 142.6000 54.8200 143.6800 ;
      RECT 0.0000 142.6000 5.2600 143.6800 ;
      RECT 0.0000 140.9600 210.2200 142.6000 ;
      RECT 208.9600 139.8800 210.2200 140.9600 ;
      RECT 195.2200 139.8800 205.3600 140.9600 ;
      RECT 150.2200 139.8800 193.0200 140.9600 ;
      RECT 105.2200 139.8800 148.0200 140.9600 ;
      RECT 60.2200 139.8800 103.0200 140.9600 ;
      RECT 15.2200 139.8800 58.0200 140.9600 ;
      RECT 4.8600 139.8800 13.0200 140.9600 ;
      RECT 0.0000 139.8800 1.2600 140.9600 ;
      RECT 0.0000 138.2400 210.2200 139.8800 ;
      RECT 204.9600 137.1600 210.2200 138.2400 ;
      RECT 192.0200 137.1600 201.3600 138.2400 ;
      RECT 147.0200 137.1600 189.8200 138.2400 ;
      RECT 102.0200 137.1600 144.8200 138.2400 ;
      RECT 57.0200 137.1600 99.8200 138.2400 ;
      RECT 8.8600 137.1600 54.8200 138.2400 ;
      RECT 0.0000 137.1600 5.2600 138.2400 ;
      RECT 0.0000 135.5200 210.2200 137.1600 ;
      RECT 208.9600 134.4400 210.2200 135.5200 ;
      RECT 195.2200 134.4400 205.3600 135.5200 ;
      RECT 150.2200 134.4400 193.0200 135.5200 ;
      RECT 105.2200 134.4400 148.0200 135.5200 ;
      RECT 60.2200 134.4400 103.0200 135.5200 ;
      RECT 15.2200 134.4400 58.0200 135.5200 ;
      RECT 4.8600 134.4400 13.0200 135.5200 ;
      RECT 0.0000 134.4400 1.2600 135.5200 ;
      RECT 0.0000 132.8000 210.2200 134.4400 ;
      RECT 204.9600 131.7200 210.2200 132.8000 ;
      RECT 192.0200 131.7200 201.3600 132.8000 ;
      RECT 147.0200 131.7200 189.8200 132.8000 ;
      RECT 102.0200 131.7200 144.8200 132.8000 ;
      RECT 57.0200 131.7200 99.8200 132.8000 ;
      RECT 8.8600 131.7200 54.8200 132.8000 ;
      RECT 0.0000 131.7200 5.2600 132.8000 ;
      RECT 0.0000 130.0800 210.2200 131.7200 ;
      RECT 208.9600 129.0000 210.2200 130.0800 ;
      RECT 195.2200 129.0000 205.3600 130.0800 ;
      RECT 150.2200 129.0000 193.0200 130.0800 ;
      RECT 105.2200 129.0000 148.0200 130.0800 ;
      RECT 60.2200 129.0000 103.0200 130.0800 ;
      RECT 15.2200 129.0000 58.0200 130.0800 ;
      RECT 4.8600 129.0000 13.0200 130.0800 ;
      RECT 0.0000 129.0000 1.2600 130.0800 ;
      RECT 0.0000 127.3600 210.2200 129.0000 ;
      RECT 204.9600 126.2800 210.2200 127.3600 ;
      RECT 192.0200 126.2800 201.3600 127.3600 ;
      RECT 147.0200 126.2800 189.8200 127.3600 ;
      RECT 102.0200 126.2800 144.8200 127.3600 ;
      RECT 57.0200 126.2800 99.8200 127.3600 ;
      RECT 8.8600 126.2800 54.8200 127.3600 ;
      RECT 0.0000 126.2800 5.2600 127.3600 ;
      RECT 0.0000 124.6400 210.2200 126.2800 ;
      RECT 208.9600 123.5600 210.2200 124.6400 ;
      RECT 195.2200 123.5600 205.3600 124.6400 ;
      RECT 150.2200 123.5600 193.0200 124.6400 ;
      RECT 105.2200 123.5600 148.0200 124.6400 ;
      RECT 60.2200 123.5600 103.0200 124.6400 ;
      RECT 15.2200 123.5600 58.0200 124.6400 ;
      RECT 4.8600 123.5600 13.0200 124.6400 ;
      RECT 0.0000 123.5600 1.2600 124.6400 ;
      RECT 0.0000 121.9200 210.2200 123.5600 ;
      RECT 204.9600 120.8400 210.2200 121.9200 ;
      RECT 192.0200 120.8400 201.3600 121.9200 ;
      RECT 147.0200 120.8400 189.8200 121.9200 ;
      RECT 102.0200 120.8400 144.8200 121.9200 ;
      RECT 57.0200 120.8400 99.8200 121.9200 ;
      RECT 8.8600 120.8400 54.8200 121.9200 ;
      RECT 0.0000 120.8400 5.2600 121.9200 ;
      RECT 0.0000 119.2000 210.2200 120.8400 ;
      RECT 208.9600 118.1200 210.2200 119.2000 ;
      RECT 195.2200 118.1200 205.3600 119.2000 ;
      RECT 150.2200 118.1200 193.0200 119.2000 ;
      RECT 105.2200 118.1200 148.0200 119.2000 ;
      RECT 60.2200 118.1200 103.0200 119.2000 ;
      RECT 15.2200 118.1200 58.0200 119.2000 ;
      RECT 4.8600 118.1200 13.0200 119.2000 ;
      RECT 0.0000 118.1200 1.2600 119.2000 ;
      RECT 0.0000 116.4800 210.2200 118.1200 ;
      RECT 204.9600 115.4000 210.2200 116.4800 ;
      RECT 192.0200 115.4000 201.3600 116.4800 ;
      RECT 147.0200 115.4000 189.8200 116.4800 ;
      RECT 102.0200 115.4000 144.8200 116.4800 ;
      RECT 57.0200 115.4000 99.8200 116.4800 ;
      RECT 8.8600 115.4000 54.8200 116.4800 ;
      RECT 0.0000 115.4000 5.2600 116.4800 ;
      RECT 0.0000 113.7600 210.2200 115.4000 ;
      RECT 208.9600 112.6800 210.2200 113.7600 ;
      RECT 195.2200 112.6800 205.3600 113.7600 ;
      RECT 150.2200 112.6800 193.0200 113.7600 ;
      RECT 105.2200 112.6800 148.0200 113.7600 ;
      RECT 60.2200 112.6800 103.0200 113.7600 ;
      RECT 15.2200 112.6800 58.0200 113.7600 ;
      RECT 4.8600 112.6800 13.0200 113.7600 ;
      RECT 0.0000 112.6800 1.2600 113.7600 ;
      RECT 0.0000 111.0400 210.2200 112.6800 ;
      RECT 204.9600 109.9600 210.2200 111.0400 ;
      RECT 192.0200 109.9600 201.3600 111.0400 ;
      RECT 147.0200 109.9600 189.8200 111.0400 ;
      RECT 102.0200 109.9600 144.8200 111.0400 ;
      RECT 57.0200 109.9600 99.8200 111.0400 ;
      RECT 8.8600 109.9600 54.8200 111.0400 ;
      RECT 0.0000 109.9600 5.2600 111.0400 ;
      RECT 0.0000 108.3200 210.2200 109.9600 ;
      RECT 208.9600 107.2400 210.2200 108.3200 ;
      RECT 195.2200 107.2400 205.3600 108.3200 ;
      RECT 150.2200 107.2400 193.0200 108.3200 ;
      RECT 105.2200 107.2400 148.0200 108.3200 ;
      RECT 60.2200 107.2400 103.0200 108.3200 ;
      RECT 15.2200 107.2400 58.0200 108.3200 ;
      RECT 4.8600 107.2400 13.0200 108.3200 ;
      RECT 0.0000 107.2400 1.2600 108.3200 ;
      RECT 0.0000 105.6000 210.2200 107.2400 ;
      RECT 204.9600 104.5200 210.2200 105.6000 ;
      RECT 192.0200 104.5200 201.3600 105.6000 ;
      RECT 147.0200 104.5200 189.8200 105.6000 ;
      RECT 102.0200 104.5200 144.8200 105.6000 ;
      RECT 57.0200 104.5200 99.8200 105.6000 ;
      RECT 8.8600 104.5200 54.8200 105.6000 ;
      RECT 0.0000 104.5200 5.2600 105.6000 ;
      RECT 0.0000 102.8800 210.2200 104.5200 ;
      RECT 208.9600 101.8000 210.2200 102.8800 ;
      RECT 195.2200 101.8000 205.3600 102.8800 ;
      RECT 150.2200 101.8000 193.0200 102.8800 ;
      RECT 105.2200 101.8000 148.0200 102.8800 ;
      RECT 60.2200 101.8000 103.0200 102.8800 ;
      RECT 15.2200 101.8000 58.0200 102.8800 ;
      RECT 4.8600 101.8000 13.0200 102.8800 ;
      RECT 0.0000 101.8000 1.2600 102.8800 ;
      RECT 0.0000 100.1600 210.2200 101.8000 ;
      RECT 204.9600 99.0800 210.2200 100.1600 ;
      RECT 192.0200 99.0800 201.3600 100.1600 ;
      RECT 147.0200 99.0800 189.8200 100.1600 ;
      RECT 102.0200 99.0800 144.8200 100.1600 ;
      RECT 57.0200 99.0800 99.8200 100.1600 ;
      RECT 8.8600 99.0800 54.8200 100.1600 ;
      RECT 0.0000 99.0800 5.2600 100.1600 ;
      RECT 0.0000 97.4400 210.2200 99.0800 ;
      RECT 208.9600 96.3600 210.2200 97.4400 ;
      RECT 195.2200 96.3600 205.3600 97.4400 ;
      RECT 150.2200 96.3600 193.0200 97.4400 ;
      RECT 105.2200 96.3600 148.0200 97.4400 ;
      RECT 60.2200 96.3600 103.0200 97.4400 ;
      RECT 15.2200 96.3600 58.0200 97.4400 ;
      RECT 4.8600 96.3600 13.0200 97.4400 ;
      RECT 0.0000 96.3600 1.2600 97.4400 ;
      RECT 0.0000 94.7200 210.2200 96.3600 ;
      RECT 204.9600 93.6400 210.2200 94.7200 ;
      RECT 192.0200 93.6400 201.3600 94.7200 ;
      RECT 147.0200 93.6400 189.8200 94.7200 ;
      RECT 102.0200 93.6400 144.8200 94.7200 ;
      RECT 57.0200 93.6400 99.8200 94.7200 ;
      RECT 8.8600 93.6400 54.8200 94.7200 ;
      RECT 0.0000 93.6400 5.2600 94.7200 ;
      RECT 0.0000 92.0000 210.2200 93.6400 ;
      RECT 208.9600 90.9200 210.2200 92.0000 ;
      RECT 195.2200 90.9200 205.3600 92.0000 ;
      RECT 150.2200 90.9200 193.0200 92.0000 ;
      RECT 105.2200 90.9200 148.0200 92.0000 ;
      RECT 60.2200 90.9200 103.0200 92.0000 ;
      RECT 15.2200 90.9200 58.0200 92.0000 ;
      RECT 4.8600 90.9200 13.0200 92.0000 ;
      RECT 0.0000 90.9200 1.2600 92.0000 ;
      RECT 0.0000 89.2800 210.2200 90.9200 ;
      RECT 204.9600 88.2000 210.2200 89.2800 ;
      RECT 192.0200 88.2000 201.3600 89.2800 ;
      RECT 147.0200 88.2000 189.8200 89.2800 ;
      RECT 102.0200 88.2000 144.8200 89.2800 ;
      RECT 57.0200 88.2000 99.8200 89.2800 ;
      RECT 8.8600 88.2000 54.8200 89.2800 ;
      RECT 0.0000 88.2000 5.2600 89.2800 ;
      RECT 0.0000 86.5600 210.2200 88.2000 ;
      RECT 208.9600 85.4800 210.2200 86.5600 ;
      RECT 195.2200 85.4800 205.3600 86.5600 ;
      RECT 150.2200 85.4800 193.0200 86.5600 ;
      RECT 105.2200 85.4800 148.0200 86.5600 ;
      RECT 60.2200 85.4800 103.0200 86.5600 ;
      RECT 15.2200 85.4800 58.0200 86.5600 ;
      RECT 4.8600 85.4800 13.0200 86.5600 ;
      RECT 0.0000 85.4800 1.2600 86.5600 ;
      RECT 0.0000 83.8400 210.2200 85.4800 ;
      RECT 204.9600 82.7600 210.2200 83.8400 ;
      RECT 192.0200 82.7600 201.3600 83.8400 ;
      RECT 147.0200 82.7600 189.8200 83.8400 ;
      RECT 102.0200 82.7600 144.8200 83.8400 ;
      RECT 57.0200 82.7600 99.8200 83.8400 ;
      RECT 8.8600 82.7600 54.8200 83.8400 ;
      RECT 0.0000 82.7600 5.2600 83.8400 ;
      RECT 0.0000 81.1200 210.2200 82.7600 ;
      RECT 208.9600 80.0400 210.2200 81.1200 ;
      RECT 195.2200 80.0400 205.3600 81.1200 ;
      RECT 150.2200 80.0400 193.0200 81.1200 ;
      RECT 105.2200 80.0400 148.0200 81.1200 ;
      RECT 60.2200 80.0400 103.0200 81.1200 ;
      RECT 15.2200 80.0400 58.0200 81.1200 ;
      RECT 4.8600 80.0400 13.0200 81.1200 ;
      RECT 0.0000 80.0400 1.2600 81.1200 ;
      RECT 0.0000 78.4000 210.2200 80.0400 ;
      RECT 204.9600 77.3200 210.2200 78.4000 ;
      RECT 192.0200 77.3200 201.3600 78.4000 ;
      RECT 147.0200 77.3200 189.8200 78.4000 ;
      RECT 102.0200 77.3200 144.8200 78.4000 ;
      RECT 57.0200 77.3200 99.8200 78.4000 ;
      RECT 8.8600 77.3200 54.8200 78.4000 ;
      RECT 0.0000 77.3200 5.2600 78.4000 ;
      RECT 0.0000 75.6800 210.2200 77.3200 ;
      RECT 208.9600 74.6000 210.2200 75.6800 ;
      RECT 195.2200 74.6000 205.3600 75.6800 ;
      RECT 150.2200 74.6000 193.0200 75.6800 ;
      RECT 105.2200 74.6000 148.0200 75.6800 ;
      RECT 60.2200 74.6000 103.0200 75.6800 ;
      RECT 15.2200 74.6000 58.0200 75.6800 ;
      RECT 4.8600 74.6000 13.0200 75.6800 ;
      RECT 0.0000 74.6000 1.2600 75.6800 ;
      RECT 0.0000 72.9600 210.2200 74.6000 ;
      RECT 204.9600 71.8800 210.2200 72.9600 ;
      RECT 192.0200 71.8800 201.3600 72.9600 ;
      RECT 147.0200 71.8800 189.8200 72.9600 ;
      RECT 102.0200 71.8800 144.8200 72.9600 ;
      RECT 57.0200 71.8800 99.8200 72.9600 ;
      RECT 8.8600 71.8800 54.8200 72.9600 ;
      RECT 0.0000 71.8800 5.2600 72.9600 ;
      RECT 0.0000 70.2400 210.2200 71.8800 ;
      RECT 208.9600 69.1600 210.2200 70.2400 ;
      RECT 195.2200 69.1600 205.3600 70.2400 ;
      RECT 150.2200 69.1600 193.0200 70.2400 ;
      RECT 105.2200 69.1600 148.0200 70.2400 ;
      RECT 60.2200 69.1600 103.0200 70.2400 ;
      RECT 15.2200 69.1600 58.0200 70.2400 ;
      RECT 4.8600 69.1600 13.0200 70.2400 ;
      RECT 0.0000 69.1600 1.2600 70.2400 ;
      RECT 0.0000 67.5200 210.2200 69.1600 ;
      RECT 204.9600 66.4400 210.2200 67.5200 ;
      RECT 192.0200 66.4400 201.3600 67.5200 ;
      RECT 147.0200 66.4400 189.8200 67.5200 ;
      RECT 102.0200 66.4400 144.8200 67.5200 ;
      RECT 57.0200 66.4400 99.8200 67.5200 ;
      RECT 8.8600 66.4400 54.8200 67.5200 ;
      RECT 0.0000 66.4400 5.2600 67.5200 ;
      RECT 0.0000 64.8000 210.2200 66.4400 ;
      RECT 208.9600 63.7200 210.2200 64.8000 ;
      RECT 195.2200 63.7200 205.3600 64.8000 ;
      RECT 150.2200 63.7200 193.0200 64.8000 ;
      RECT 105.2200 63.7200 148.0200 64.8000 ;
      RECT 60.2200 63.7200 103.0200 64.8000 ;
      RECT 15.2200 63.7200 58.0200 64.8000 ;
      RECT 4.8600 63.7200 13.0200 64.8000 ;
      RECT 0.0000 63.7200 1.2600 64.8000 ;
      RECT 0.0000 62.0800 210.2200 63.7200 ;
      RECT 204.9600 61.0000 210.2200 62.0800 ;
      RECT 192.0200 61.0000 201.3600 62.0800 ;
      RECT 147.0200 61.0000 189.8200 62.0800 ;
      RECT 102.0200 61.0000 144.8200 62.0800 ;
      RECT 57.0200 61.0000 99.8200 62.0800 ;
      RECT 8.8600 61.0000 54.8200 62.0800 ;
      RECT 0.0000 61.0000 5.2600 62.0800 ;
      RECT 0.0000 59.3600 210.2200 61.0000 ;
      RECT 208.9600 58.2800 210.2200 59.3600 ;
      RECT 195.2200 58.2800 205.3600 59.3600 ;
      RECT 150.2200 58.2800 193.0200 59.3600 ;
      RECT 105.2200 58.2800 148.0200 59.3600 ;
      RECT 60.2200 58.2800 103.0200 59.3600 ;
      RECT 15.2200 58.2800 58.0200 59.3600 ;
      RECT 4.8600 58.2800 13.0200 59.3600 ;
      RECT 0.0000 58.2800 1.2600 59.3600 ;
      RECT 0.0000 56.6400 210.2200 58.2800 ;
      RECT 204.9600 55.5600 210.2200 56.6400 ;
      RECT 192.0200 55.5600 201.3600 56.6400 ;
      RECT 147.0200 55.5600 189.8200 56.6400 ;
      RECT 102.0200 55.5600 144.8200 56.6400 ;
      RECT 57.0200 55.5600 99.8200 56.6400 ;
      RECT 8.8600 55.5600 54.8200 56.6400 ;
      RECT 0.0000 55.5600 5.2600 56.6400 ;
      RECT 0.0000 53.9200 210.2200 55.5600 ;
      RECT 208.9600 52.8400 210.2200 53.9200 ;
      RECT 195.2200 52.8400 205.3600 53.9200 ;
      RECT 150.2200 52.8400 193.0200 53.9200 ;
      RECT 105.2200 52.8400 148.0200 53.9200 ;
      RECT 60.2200 52.8400 103.0200 53.9200 ;
      RECT 15.2200 52.8400 58.0200 53.9200 ;
      RECT 4.8600 52.8400 13.0200 53.9200 ;
      RECT 0.0000 52.8400 1.2600 53.9200 ;
      RECT 0.0000 51.2000 210.2200 52.8400 ;
      RECT 204.9600 50.1200 210.2200 51.2000 ;
      RECT 192.0200 50.1200 201.3600 51.2000 ;
      RECT 147.0200 50.1200 189.8200 51.2000 ;
      RECT 102.0200 50.1200 144.8200 51.2000 ;
      RECT 57.0200 50.1200 99.8200 51.2000 ;
      RECT 8.8600 50.1200 54.8200 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 210.2200 50.1200 ;
      RECT 208.9600 47.4000 210.2200 48.4800 ;
      RECT 195.2200 47.4000 205.3600 48.4800 ;
      RECT 150.2200 47.4000 193.0200 48.4800 ;
      RECT 105.2200 47.4000 148.0200 48.4800 ;
      RECT 60.2200 47.4000 103.0200 48.4800 ;
      RECT 15.2200 47.4000 58.0200 48.4800 ;
      RECT 4.8600 47.4000 13.0200 48.4800 ;
      RECT 0.0000 47.4000 1.2600 48.4800 ;
      RECT 0.0000 45.7600 210.2200 47.4000 ;
      RECT 204.9600 44.6800 210.2200 45.7600 ;
      RECT 192.0200 44.6800 201.3600 45.7600 ;
      RECT 147.0200 44.6800 189.8200 45.7600 ;
      RECT 102.0200 44.6800 144.8200 45.7600 ;
      RECT 57.0200 44.6800 99.8200 45.7600 ;
      RECT 8.8600 44.6800 54.8200 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 210.2200 44.6800 ;
      RECT 208.9600 41.9600 210.2200 43.0400 ;
      RECT 195.2200 41.9600 205.3600 43.0400 ;
      RECT 150.2200 41.9600 193.0200 43.0400 ;
      RECT 105.2200 41.9600 148.0200 43.0400 ;
      RECT 60.2200 41.9600 103.0200 43.0400 ;
      RECT 15.2200 41.9600 58.0200 43.0400 ;
      RECT 4.8600 41.9600 13.0200 43.0400 ;
      RECT 0.0000 41.9600 1.2600 43.0400 ;
      RECT 0.0000 40.3200 210.2200 41.9600 ;
      RECT 204.9600 39.2400 210.2200 40.3200 ;
      RECT 192.0200 39.2400 201.3600 40.3200 ;
      RECT 147.0200 39.2400 189.8200 40.3200 ;
      RECT 102.0200 39.2400 144.8200 40.3200 ;
      RECT 57.0200 39.2400 99.8200 40.3200 ;
      RECT 8.8600 39.2400 54.8200 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 210.2200 39.2400 ;
      RECT 208.9600 36.5200 210.2200 37.6000 ;
      RECT 195.2200 36.5200 205.3600 37.6000 ;
      RECT 150.2200 36.5200 193.0200 37.6000 ;
      RECT 105.2200 36.5200 148.0200 37.6000 ;
      RECT 60.2200 36.5200 103.0200 37.6000 ;
      RECT 15.2200 36.5200 58.0200 37.6000 ;
      RECT 4.8600 36.5200 13.0200 37.6000 ;
      RECT 0.0000 36.5200 1.2600 37.6000 ;
      RECT 0.0000 34.8800 210.2200 36.5200 ;
      RECT 204.9600 33.8000 210.2200 34.8800 ;
      RECT 192.0200 33.8000 201.3600 34.8800 ;
      RECT 147.0200 33.8000 189.8200 34.8800 ;
      RECT 102.0200 33.8000 144.8200 34.8800 ;
      RECT 57.0200 33.8000 99.8200 34.8800 ;
      RECT 8.8600 33.8000 54.8200 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 210.2200 33.8000 ;
      RECT 208.9600 31.0800 210.2200 32.1600 ;
      RECT 195.2200 31.0800 205.3600 32.1600 ;
      RECT 150.2200 31.0800 193.0200 32.1600 ;
      RECT 105.2200 31.0800 148.0200 32.1600 ;
      RECT 60.2200 31.0800 103.0200 32.1600 ;
      RECT 15.2200 31.0800 58.0200 32.1600 ;
      RECT 4.8600 31.0800 13.0200 32.1600 ;
      RECT 0.0000 31.0800 1.2600 32.1600 ;
      RECT 0.0000 29.4400 210.2200 31.0800 ;
      RECT 204.9600 28.3600 210.2200 29.4400 ;
      RECT 192.0200 28.3600 201.3600 29.4400 ;
      RECT 147.0200 28.3600 189.8200 29.4400 ;
      RECT 102.0200 28.3600 144.8200 29.4400 ;
      RECT 57.0200 28.3600 99.8200 29.4400 ;
      RECT 8.8600 28.3600 54.8200 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 210.2200 28.3600 ;
      RECT 208.9600 25.6400 210.2200 26.7200 ;
      RECT 195.2200 25.6400 205.3600 26.7200 ;
      RECT 150.2200 25.6400 193.0200 26.7200 ;
      RECT 105.2200 25.6400 148.0200 26.7200 ;
      RECT 60.2200 25.6400 103.0200 26.7200 ;
      RECT 15.2200 25.6400 58.0200 26.7200 ;
      RECT 4.8600 25.6400 13.0200 26.7200 ;
      RECT 0.0000 25.6400 1.2600 26.7200 ;
      RECT 0.0000 24.0000 210.2200 25.6400 ;
      RECT 204.9600 22.9200 210.2200 24.0000 ;
      RECT 192.0200 22.9200 201.3600 24.0000 ;
      RECT 147.0200 22.9200 189.8200 24.0000 ;
      RECT 102.0200 22.9200 144.8200 24.0000 ;
      RECT 57.0200 22.9200 99.8200 24.0000 ;
      RECT 8.8600 22.9200 54.8200 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 210.2200 22.9200 ;
      RECT 208.9600 20.2000 210.2200 21.2800 ;
      RECT 195.2200 20.2000 205.3600 21.2800 ;
      RECT 150.2200 20.2000 193.0200 21.2800 ;
      RECT 105.2200 20.2000 148.0200 21.2800 ;
      RECT 60.2200 20.2000 103.0200 21.2800 ;
      RECT 15.2200 20.2000 58.0200 21.2800 ;
      RECT 4.8600 20.2000 13.0200 21.2800 ;
      RECT 0.0000 20.2000 1.2600 21.2800 ;
      RECT 0.0000 18.5600 210.2200 20.2000 ;
      RECT 204.9600 17.4800 210.2200 18.5600 ;
      RECT 192.0200 17.4800 201.3600 18.5600 ;
      RECT 147.0200 17.4800 189.8200 18.5600 ;
      RECT 102.0200 17.4800 144.8200 18.5600 ;
      RECT 57.0200 17.4800 99.8200 18.5600 ;
      RECT 8.8600 17.4800 54.8200 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 210.2200 17.4800 ;
      RECT 208.9600 14.7600 210.2200 15.8400 ;
      RECT 195.2200 14.7600 205.3600 15.8400 ;
      RECT 150.2200 14.7600 193.0200 15.8400 ;
      RECT 105.2200 14.7600 148.0200 15.8400 ;
      RECT 60.2200 14.7600 103.0200 15.8400 ;
      RECT 15.2200 14.7600 58.0200 15.8400 ;
      RECT 4.8600 14.7600 13.0200 15.8400 ;
      RECT 0.0000 14.7600 1.2600 15.8400 ;
      RECT 0.0000 13.1200 210.2200 14.7600 ;
      RECT 204.9600 12.0400 210.2200 13.1200 ;
      RECT 192.0200 12.0400 201.3600 13.1200 ;
      RECT 147.0200 12.0400 189.8200 13.1200 ;
      RECT 102.0200 12.0400 144.8200 13.1200 ;
      RECT 57.0200 12.0400 99.8200 13.1200 ;
      RECT 8.8600 12.0400 54.8200 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 210.2200 12.0400 ;
      RECT 208.9600 9.3200 210.2200 10.4000 ;
      RECT 195.2200 9.3200 205.3600 10.4000 ;
      RECT 150.2200 9.3200 193.0200 10.4000 ;
      RECT 105.2200 9.3200 148.0200 10.4000 ;
      RECT 60.2200 9.3200 103.0200 10.4000 ;
      RECT 15.2200 9.3200 58.0200 10.4000 ;
      RECT 4.8600 9.3200 13.0200 10.4000 ;
      RECT 0.0000 9.3200 1.2600 10.4000 ;
      RECT 0.0000 8.7300 210.2200 9.3200 ;
      RECT 204.9600 5.1300 210.2200 8.7300 ;
      RECT 0.0000 5.1300 5.2600 8.7300 ;
      RECT 0.0000 4.7300 210.2200 5.1300 ;
      RECT 208.9600 1.1300 210.2200 4.7300 ;
      RECT 0.0000 1.1300 1.2600 4.7300 ;
      RECT 0.0000 0.0000 210.2200 1.1300 ;
    LAYER met4 ;
      RECT 0.0000 217.8300 210.2200 219.6400 ;
      RECT 195.2200 213.8300 205.3600 217.8300 ;
      RECT 150.2200 213.8300 193.0200 217.8300 ;
      RECT 105.2200 213.8300 148.0200 217.8300 ;
      RECT 60.2200 213.8300 103.0200 217.8300 ;
      RECT 15.2200 213.8300 58.0200 217.8300 ;
      RECT 4.8600 213.8300 13.0200 217.8300 ;
      RECT 204.9600 5.1300 205.3600 213.8300 ;
      RECT 195.2200 5.1300 201.3600 213.8300 ;
      RECT 192.0200 5.1300 193.0200 213.8300 ;
      RECT 150.2200 5.1300 189.8200 213.8300 ;
      RECT 147.0200 5.1300 148.0200 213.8300 ;
      RECT 105.2200 5.1300 144.8200 213.8300 ;
      RECT 102.0200 5.1300 103.0200 213.8300 ;
      RECT 60.2200 5.1300 99.8200 213.8300 ;
      RECT 57.0200 5.1300 58.0200 213.8300 ;
      RECT 15.2200 5.1300 54.8200 213.8300 ;
      RECT 8.8600 5.1300 13.0200 213.8300 ;
      RECT 4.8600 5.1300 5.2600 213.8300 ;
      RECT 208.9600 1.1300 210.2200 217.8300 ;
      RECT 195.2200 1.1300 205.3600 5.1300 ;
      RECT 150.2200 1.1300 193.0200 5.1300 ;
      RECT 105.2200 1.1300 148.0200 5.1300 ;
      RECT 60.2200 1.1300 103.0200 5.1300 ;
      RECT 15.2200 1.1300 58.0200 5.1300 ;
      RECT 4.8600 1.1300 13.0200 5.1300 ;
      RECT 0.0000 1.1300 1.2600 217.8300 ;
      RECT 0.0000 1.0200 210.2200 1.1300 ;
      RECT 89.5000 0.0000 210.2200 1.0200 ;
      RECT 0.0000 0.0000 88.5200 1.0200 ;
  END
END LUT4AB

END LIBRARY
