##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Sat Jun 19 03:30:33 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BlockRAM_1KB
  CLASS BLOCK ;
  SIZE 480.2400 BY 449.8200 ;
  FOREIGN BlockRAM_1KB 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 134.524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 718.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.406 LAYER met4  ;
    ANTENNAMAXAREACAR 60.7259 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 302.798 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.990122 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 9.4700 0.0000 9.8500 0.7200 ;
    END
  END clk
  PIN rd_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9582 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.683 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 48.2241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 240.831 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6969 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.192 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 97.5600 0.7200 97.9400 ;
    END
  END rd_addr[7]
  PIN rd_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6362 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.073 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 49.0221 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 244.822 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.0749 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.208 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 94.1600 0.7200 94.5400 ;
    END
  END rd_addr[6]
  PIN rd_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2032 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.908 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 49.3861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 246.642 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.48 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 90.7600 0.7200 91.1400 ;
    END
  END rd_addr[5]
  PIN rd_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.332 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.552 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 49.3441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 246.432 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6552 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.96 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 87.7000 0.7200 88.0800 ;
    END
  END rd_addr[4]
  PIN rd_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.765 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.717 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 50.0973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 250.198 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.5969 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.992 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 84.3000 0.7200 84.6800 ;
    END
  END rd_addr[3]
  PIN rd_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3426 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.568 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 48.3669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 241.546 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.0089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.856 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 81.2400 0.7200 81.6200 ;
    END
  END rd_addr[2]
  PIN rd_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2498 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 50.9849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 254.635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.2089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.256 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 77.8400 0.7200 78.2200 ;
    END
  END rd_addr[1]
  PIN rd_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6372 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.078 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 45.2031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 225.844 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.888 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 74.7800 0.7200 75.1600 ;
    END
  END rd_addr[0]
  PIN rd_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5002 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.393 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 38.0099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 189.878 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.4108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.328 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 291.0200 0.7200 291.4000 ;
    END
  END rd_data[31]
  PIN rd_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.985 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.817 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 36.5371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 182.514 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.6668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.36 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 287.6200 0.7200 288.0000 ;
    END
  END rd_data[30]
  PIN rd_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7578 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.681 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 34.7773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 173.715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.3768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.48 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 284.2200 0.7200 284.6000 ;
    END
  END rd_data[29]
  PIN rd_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4698 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.241 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 37.1502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 185.633 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 280.8200 0.7200 281.2000 ;
    END
  END rd_data[28]
  PIN rd_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.3178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 66.444 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 277.4200 0.7200 277.8000 ;
    END
  END rd_data[27]
  PIN rd_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.1844 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.885 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 274.0200 0.7200 274.4000 ;
    END
  END rd_data[26]
  PIN rd_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7274 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.529 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 36.4152 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 181.958 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 270.6200 0.7200 271.0000 ;
    END
  END rd_data[25]
  PIN rd_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.389 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8405 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 267.2200 0.7200 267.6000 ;
    END
  END rd_data[24]
  PIN rd_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.62 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 31.6987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 158.322 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.464 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 263.8200 0.7200 264.2000 ;
    END
  END rd_data[23]
  PIN rd_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1782 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.783 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 33.7721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 168.689 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.4 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 260.4200 0.7200 260.8000 ;
    END
  END rd_data[22]
  PIN rd_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0118 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.951 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 34.4254 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 171.773 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 257.0200 0.7200 257.4000 ;
    END
  END rd_data[21]
  PIN rd_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9546 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 33.5774 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 167.769 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 253.6200 0.7200 254.0000 ;
    END
  END rd_data[20]
  PIN rd_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.663 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.207 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 32.5135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 162.396 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.856 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 250.2200 0.7200 250.6000 ;
    END
  END rd_data[19]
  PIN rd_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9252 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.518 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 31.1428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 155.596 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 246.8200 0.7200 247.2000 ;
    END
  END rd_data[18]
  PIN rd_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4572 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.178 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 32.624 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 163.002 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 243.4200 0.7200 243.8000 ;
    END
  END rd_data[17]
  PIN rd_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.629 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.037 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 30.6668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.216 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 240.0200 0.7200 240.4000 ;
    END
  END rd_data[16]
  PIN rd_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 71.015 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.74 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 58.4600 0.7200 58.8400 ;
    END
  END rd_data[15]
  PIN rd_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8518 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 74.151 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8988 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.376 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 55.0600 0.7200 55.4400 ;
    END
  END rd_data[14]
  PIN rd_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7062 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.28 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 52.0000 0.7200 52.3800 ;
    END
  END rd_data[13]
  PIN rd_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.243 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.107 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.376 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 48.6000 0.7200 48.9800 ;
    END
  END rd_data[12]
  PIN rd_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7282 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.533 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.4428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.832 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 45.5400 0.7200 45.9200 ;
    END
  END rd_data[11]
  PIN rd_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.549 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.0668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.16 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 42.1400 0.7200 42.5200 ;
    END
  END rd_data[10]
  PIN rd_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5078 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.431 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0486 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.125 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 39.0800 0.7200 39.4600 ;
    END
  END rd_data[9]
  PIN rd_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.087 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.327 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.8478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.992 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 35.6800 0.7200 36.0600 ;
    END
  END rd_data[8]
  PIN rd_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6974 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.379 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.3248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.536 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 32.2800 0.7200 32.6600 ;
    END
  END rd_data[7]
  PIN rd_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.5188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.904 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 29.2200 0.7200 29.6000 ;
    END
  END rd_data[6]
  PIN rd_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.8188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.504 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 25.8200 0.7200 26.2000 ;
    END
  END rd_data[5]
  PIN rd_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7006 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3793 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.3888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.544 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 22.7600 0.7200 23.1400 ;
    END
  END rd_data[4]
  PIN rd_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0226 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.7148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.616 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 19.3600 0.7200 19.7400 ;
    END
  END rd_data[3]
  PIN rd_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.333 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.5975 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 16.3000 0.7200 16.6800 ;
    END
  END rd_data[2]
  PIN rd_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.8088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.9765 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 12.9000 0.7200 13.2800 ;
    END
  END rd_data[1]
  PIN rd_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6702 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.243 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.37 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 9.8400 0.7200 10.2200 ;
    END
  END rd_data[0]
  PIN wr_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2086 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.935 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 37.0481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 185.07 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.552 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 325.0200 0.7200 325.4000 ;
    END
  END wr_addr[7]
  PIN wr_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4546 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 36.5721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 182.689 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 321.6200 0.7200 322.0000 ;
    END
  END wr_addr[6]
  PIN wr_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3338 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.561 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 36.0667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 180.162 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 318.2200 0.7200 318.6000 ;
    END
  END wr_addr[5]
  PIN wr_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.199 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.887 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 35.5935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 177.796 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.552 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 314.8200 0.7200 315.2000 ;
    END
  END wr_addr[4]
  PIN wr_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4948 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.366 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 35.0893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 175.158 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.9684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.64 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 311.4200 0.7200 311.8000 ;
    END
  END wr_addr[3]
  PIN wr_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.771 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.988 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.648 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 308.0200 0.7200 308.4000 ;
    END
  END wr_addr[2]
  PIN wr_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1926 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.818 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.1861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 304.6200 0.7200 305.0000 ;
    END
  END wr_addr[1]
  PIN wr_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.908 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.432 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 29.6279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 147.85 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.697 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.840075 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.936 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 301.2200 0.7200 301.6000 ;
    END
  END wr_addr[0]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.2878 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 296.331 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 50.5091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 252.374 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 35.727 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.643 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 379.4200 0.7200 379.8000 ;
    END
  END wr_data[31]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.7698 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 293.741 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 49.9701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 249.68 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.37 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2222 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 151.123 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 376.0200 0.7200 376.4000 ;
    END
  END wr_data[30]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.4334 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 297.059 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 48.2215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 240.936 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 44.5778 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.262 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 372.6200 0.7200 373.0000 ;
    END
  END wr_data[29]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.7518 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 308.651 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 45.0209 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 224.816 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 9.10873 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.5794 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 369.2200 0.7200 369.6000 ;
    END
  END wr_data[28]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.6982 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 278.383 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 46.7268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 233.345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 9.81032 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.5516 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 365.8200 0.7200 366.2000 ;
    END
  END wr_data[27]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.0792 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 295.288 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 48.6653 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 243.156 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.0888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 79.6968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 407.663 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 362.4200 0.7200 362.8000 ;
    END
  END wr_data[26]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.2028 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 85.869 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.798 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 24.0325 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.552 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 359.0200 0.7200 359.4000 ;
    END
  END wr_data[25]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3964 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.837 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.3065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.1255 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 61.2619 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 285.302 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 63.9238 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 301.365 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 355.6200 0.7200 356.0000 ;
    END
  END wr_data[24]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 62.581 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 312.76 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 122.073 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 634.369 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 352.2200 0.7200 352.6000 ;
    END
  END wr_data[23]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 62.3598 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 311.654 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.802 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 69.4865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 328.718 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 348.8200 0.7200 349.2000 ;
    END
  END wr_data[22]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 62.2184 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 310.947 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.3908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.836 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 81.8643 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 390.607 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 345.4200 0.7200 345.8000 ;
    END
  END wr_data[21]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6064 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.887 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.7148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.22 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 39.2335 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 177.82 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 342.0200 0.7200 342.4000 ;
    END
  END wr_data[20]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 63.0612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 315.161 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.46 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 57.3754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 268.163 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 338.6200 0.7200 339.0000 ;
    END
  END wr_data[19]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 62.7952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 313.831 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.82 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.982 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 67.0087 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 316.329 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 335.2200 0.7200 335.6000 ;
    END
  END wr_data[18]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 309.645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.77 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.737 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2664 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.6608 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 331.8200 0.7200 332.2000 ;
    END
  END wr_data[17]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.425 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 301.98 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.2424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.642 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.494 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1876 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.9217 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 328.4200 0.7200 328.8000 ;
    END
  END wr_data[16]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 63.5064 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 317.387 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.252 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 37.0786 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 166.718 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 149.2400 0.7200 149.6200 ;
    END
  END wr_data[15]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.0058 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 319.921 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.184 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 74.4341 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 353.496 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 146.1800 0.7200 146.5600 ;
    END
  END wr_data[14]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.7554 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 298.669 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.9815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.7365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 44.8496 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.522 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 142.7800 0.7200 143.1600 ;
    END
  END wr_data[13]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.1428 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 305.606 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.954 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 59.4008 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 278.329 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 139.7200 0.7200 140.1000 ;
    END
  END wr_data[12]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.9968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 309.876 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.5524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.536 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 61.0675 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 286.663 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 136.3200 0.7200 136.7000 ;
    END
  END wr_data[11]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 63.2876 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 316.33 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 15.6328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.938 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 67.8897 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 320.774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 133.2600 0.7200 133.6400 ;
    END
  END wr_data[10]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.6444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 303.114 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 14.1236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.392 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 61.9008 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 290.829 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 129.8600 0.7200 130.2400 ;
    END
  END wr_data[9]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.768 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 228.732 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.7444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.541 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.1844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 16.2317 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 69.1905 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 126.8000 0.7200 127.1800 ;
    END
  END wr_data[8]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.509 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 322.329 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNAPARTIALMETALAREA 21.1492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 105.007 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.5854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 18.9504 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 95.4246 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0029 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.824 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 22.9302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 118.536 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 123.4000 0.7200 123.7800 ;
    END
  END wr_data[7]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.6038 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 327.803 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.9555 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 80.3294 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 389.05 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 81.369 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 396.446 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2019 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.552 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 105.98 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 529.589 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 120.0000 0.7200 120.3800 ;
    END
  END wr_data[6]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 63.9698 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 319.704 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.2261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.5745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 90.7944 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 440.744 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 93.2032 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 455.442 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1589 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.656 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 97.802 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 481.855 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 116.9400 0.7200 117.3200 ;
    END
  END wr_data[5]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.9356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 304.57 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 14.5417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.0755 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 69.0659 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 330.939 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 71.4746 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 345.637 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0539 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.096 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 75.6567 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 369.827 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 113.5400 0.7200 113.9200 ;
    END
  END wr_data[4]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.6822 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 328.195 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.9077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.0135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 70.369 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 337.883 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 71.6825 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 346.74 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.0589 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.456 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 103.662 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 519.185 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 110.4800 0.7200 110.8600 ;
    END
  END wr_data[3]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 63.7496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 318.64 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.81 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.6 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9797 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 45.0619 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 224.54 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0269 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.952 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 49.1369 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.159 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884127 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 107.0800 0.7200 107.4600 ;
    END
  END wr_data[2]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.413 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 306.957 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 14.1711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 63.8937 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 306.911 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.477381 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 66.3024 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 321.609 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.636111 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1049 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.368 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 70.6869 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.879 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.636111 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 104.0200 0.7200 104.4000 ;
    END
  END wr_data[1]
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.1966 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 280.875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.2839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.8945 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 58.773 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 280.439 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 61.1817 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 295.137 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1829 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.784 LAYER met4  ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 65.8758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.058 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 100.6200 0.7200 101.0000 ;
    END
  END wr_data[0]
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.968 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.254 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.611 LAYER met2  ;
    ANTENNAMAXAREACAR 52.6425 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 261.667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.265597 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 61.5200 0.7200 61.9000 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.6932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 78.358 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.3716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.622 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met2  ;
    ANTENNAMAXAREACAR 83.0117 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 408.321 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.265597 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 64.9200 0.7200 65.3000 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.713 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 58.457 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.9404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.466 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2655 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.1152 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.149293 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 68.3200 0.7200 68.7000 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6114 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 67.949 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.7374 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.451 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7048 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.3171 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 71.3800 0.7200 71.7600 ;
    END
  END C3
  PIN C4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.4394 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 87.052 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.4316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.922 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4319 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.5798 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 294.4200 0.7200 294.8000 ;
    END
  END C4
  PIN C5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.994 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 51.1648 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 253.652 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.064 LAYER met2  ;
    ANTENNAMAXAREACAR 21.3603 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.2664 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.293254 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 297.8200 0.7200 298.2000 ;
    END
  END C5
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 474.6800 6.9300 ;
        RECT 5.5600 442.7200 474.6800 444.2200 ;
        RECT 466.1650 250.9400 474.6800 252.4400 ;
        RECT 5.5600 12.3400 7.0600 12.8200 ;
        RECT 5.5600 17.7800 7.0600 18.2600 ;
        RECT 5.5600 28.6600 7.0600 29.1400 ;
        RECT 5.5600 23.2200 7.0600 23.7000 ;
        RECT 5.5600 34.1000 7.0600 34.5800 ;
        RECT 5.5600 39.5400 7.0600 40.0200 ;
        RECT 5.5600 44.9800 7.0600 45.4600 ;
        RECT 5.5600 50.4200 7.0600 50.9000 ;
        RECT 473.1800 12.3400 474.6800 12.8200 ;
        RECT 473.1800 17.7800 474.6800 18.2600 ;
        RECT 473.1800 28.6600 474.6800 29.1400 ;
        RECT 473.1800 23.2200 474.6800 23.7000 ;
        RECT 473.1800 34.1000 474.6800 34.5800 ;
        RECT 473.1800 39.5400 474.6800 40.0200 ;
        RECT 473.1800 44.9800 474.6800 45.4600 ;
        RECT 473.1800 50.4200 474.6800 50.9000 ;
      LAYER met4 ;
        RECT 473.1800 5.4300 474.6800 444.2200 ;
        RECT 5.5600 5.4300 7.0600 444.2200 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 3.0600 2.9300 477.1800 4.4300 ;
        RECT 3.0600 445.2200 477.1800 446.7200 ;
        RECT 3.0600 433.5200 20.7650 435.0200 ;
        RECT 3.0600 9.6200 4.5600 10.1000 ;
        RECT 3.0600 15.0600 4.5600 15.5400 ;
        RECT 3.0600 20.5000 4.5600 20.9800 ;
        RECT 3.0600 25.9400 4.5600 26.4200 ;
        RECT 3.0600 31.3800 4.5600 31.8600 ;
        RECT 3.0600 36.8200 4.5600 37.3000 ;
        RECT 3.0600 42.2600 4.5600 42.7400 ;
        RECT 3.0600 47.7000 4.5600 48.1800 ;
        RECT 3.0600 53.1400 4.5600 53.6200 ;
        RECT 475.6800 9.6200 477.1800 10.1000 ;
        RECT 475.6800 15.0600 477.1800 15.5400 ;
        RECT 475.6800 20.5000 477.1800 20.9800 ;
        RECT 475.6800 25.9400 477.1800 26.4200 ;
        RECT 475.6800 31.3800 477.1800 31.8600 ;
        RECT 475.6800 36.8200 477.1800 37.3000 ;
        RECT 475.6800 42.2600 477.1800 42.7400 ;
        RECT 475.6800 47.7000 477.1800 48.1800 ;
        RECT 475.6800 53.1400 477.1800 53.6200 ;
      LAYER met4 ;
        RECT 475.6800 2.9300 477.1800 446.7200 ;
        RECT 3.0600 2.9300 4.5600 446.7200 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 480.2400 449.8200 ;
    LAYER met1 ;
      RECT 0.0000 379.9400 480.2400 449.8200 ;
      RECT 0.8600 379.2800 480.2400 379.9400 ;
      RECT 0.0000 376.5400 480.2400 379.2800 ;
      RECT 0.8600 375.8800 480.2400 376.5400 ;
      RECT 0.0000 373.1400 480.2400 375.8800 ;
      RECT 0.8600 372.4800 480.2400 373.1400 ;
      RECT 0.0000 369.7400 480.2400 372.4800 ;
      RECT 0.8600 369.0800 480.2400 369.7400 ;
      RECT 0.0000 366.3400 480.2400 369.0800 ;
      RECT 0.8600 365.6800 480.2400 366.3400 ;
      RECT 0.0000 362.9400 480.2400 365.6800 ;
      RECT 0.8600 362.2800 480.2400 362.9400 ;
      RECT 0.0000 359.5400 480.2400 362.2800 ;
      RECT 0.8600 358.8800 480.2400 359.5400 ;
      RECT 0.0000 356.1400 480.2400 358.8800 ;
      RECT 0.8600 355.4800 480.2400 356.1400 ;
      RECT 0.0000 352.7400 480.2400 355.4800 ;
      RECT 0.8600 352.0800 480.2400 352.7400 ;
      RECT 0.0000 349.3400 480.2400 352.0800 ;
      RECT 0.8600 348.6800 480.2400 349.3400 ;
      RECT 0.0000 345.9400 480.2400 348.6800 ;
      RECT 0.8600 345.2800 480.2400 345.9400 ;
      RECT 0.0000 342.5400 480.2400 345.2800 ;
      RECT 0.8600 341.8800 480.2400 342.5400 ;
      RECT 0.0000 339.1400 480.2400 341.8800 ;
      RECT 0.8600 338.4800 480.2400 339.1400 ;
      RECT 0.0000 335.7400 480.2400 338.4800 ;
      RECT 0.8600 335.0800 480.2400 335.7400 ;
      RECT 0.0000 332.3400 480.2400 335.0800 ;
      RECT 0.8600 331.6800 480.2400 332.3400 ;
      RECT 0.0000 328.9400 480.2400 331.6800 ;
      RECT 0.8600 328.2800 480.2400 328.9400 ;
      RECT 0.0000 325.5400 480.2400 328.2800 ;
      RECT 0.8600 324.8800 480.2400 325.5400 ;
      RECT 0.0000 322.1400 480.2400 324.8800 ;
      RECT 0.8600 321.4800 480.2400 322.1400 ;
      RECT 0.0000 318.7400 480.2400 321.4800 ;
      RECT 0.8600 318.0800 480.2400 318.7400 ;
      RECT 0.0000 315.3400 480.2400 318.0800 ;
      RECT 0.8600 314.6800 480.2400 315.3400 ;
      RECT 0.0000 311.9400 480.2400 314.6800 ;
      RECT 0.8600 311.2800 480.2400 311.9400 ;
      RECT 0.0000 308.5400 480.2400 311.2800 ;
      RECT 0.8600 307.8800 480.2400 308.5400 ;
      RECT 0.0000 305.1400 480.2400 307.8800 ;
      RECT 0.8600 304.4800 480.2400 305.1400 ;
      RECT 0.0000 301.7400 480.2400 304.4800 ;
      RECT 0.8600 301.0800 480.2400 301.7400 ;
      RECT 0.0000 298.3400 480.2400 301.0800 ;
      RECT 0.8600 297.6800 480.2400 298.3400 ;
      RECT 0.0000 294.9400 480.2400 297.6800 ;
      RECT 0.8600 294.2800 480.2400 294.9400 ;
      RECT 0.0000 291.5400 480.2400 294.2800 ;
      RECT 0.8600 290.8800 480.2400 291.5400 ;
      RECT 0.0000 288.1400 480.2400 290.8800 ;
      RECT 0.8600 287.4800 480.2400 288.1400 ;
      RECT 0.0000 284.7400 480.2400 287.4800 ;
      RECT 0.8600 284.0800 480.2400 284.7400 ;
      RECT 0.0000 281.3400 480.2400 284.0800 ;
      RECT 0.8600 280.6800 480.2400 281.3400 ;
      RECT 0.0000 277.9400 480.2400 280.6800 ;
      RECT 0.8600 277.2800 480.2400 277.9400 ;
      RECT 0.0000 274.5400 480.2400 277.2800 ;
      RECT 0.8600 273.8800 480.2400 274.5400 ;
      RECT 0.0000 271.1400 480.2400 273.8800 ;
      RECT 0.8600 270.4800 480.2400 271.1400 ;
      RECT 0.0000 267.7400 480.2400 270.4800 ;
      RECT 0.8600 267.0800 480.2400 267.7400 ;
      RECT 0.0000 264.3400 480.2400 267.0800 ;
      RECT 0.8600 263.6800 480.2400 264.3400 ;
      RECT 0.0000 260.9400 480.2400 263.6800 ;
      RECT 0.8600 260.2800 480.2400 260.9400 ;
      RECT 0.0000 257.5400 480.2400 260.2800 ;
      RECT 0.8600 256.8800 480.2400 257.5400 ;
      RECT 0.0000 254.1400 480.2400 256.8800 ;
      RECT 0.8600 253.4800 480.2400 254.1400 ;
      RECT 0.0000 250.7400 480.2400 253.4800 ;
      RECT 0.8600 250.0800 480.2400 250.7400 ;
      RECT 0.0000 247.3400 480.2400 250.0800 ;
      RECT 0.8600 246.6800 480.2400 247.3400 ;
      RECT 0.0000 243.9400 480.2400 246.6800 ;
      RECT 0.8600 243.2800 480.2400 243.9400 ;
      RECT 0.0000 240.5400 480.2400 243.2800 ;
      RECT 0.8600 239.8800 480.2400 240.5400 ;
      RECT 0.0000 149.7600 480.2400 239.8800 ;
      RECT 0.8600 149.1000 480.2400 149.7600 ;
      RECT 0.0000 146.7000 480.2400 149.1000 ;
      RECT 0.8600 146.0400 480.2400 146.7000 ;
      RECT 0.0000 143.3000 480.2400 146.0400 ;
      RECT 0.8600 142.6400 480.2400 143.3000 ;
      RECT 0.0000 140.2400 480.2400 142.6400 ;
      RECT 0.8600 139.5800 480.2400 140.2400 ;
      RECT 0.0000 136.8400 480.2400 139.5800 ;
      RECT 0.8600 136.1800 480.2400 136.8400 ;
      RECT 0.0000 133.7800 480.2400 136.1800 ;
      RECT 0.8600 133.1200 480.2400 133.7800 ;
      RECT 0.0000 130.3800 480.2400 133.1200 ;
      RECT 0.8600 129.7200 480.2400 130.3800 ;
      RECT 0.0000 127.3200 480.2400 129.7200 ;
      RECT 0.8600 126.6600 480.2400 127.3200 ;
      RECT 0.0000 123.9200 480.2400 126.6600 ;
      RECT 0.8600 123.2600 480.2400 123.9200 ;
      RECT 0.0000 120.5200 480.2400 123.2600 ;
      RECT 0.8600 119.8600 480.2400 120.5200 ;
      RECT 0.0000 117.4600 480.2400 119.8600 ;
      RECT 0.8600 116.8000 480.2400 117.4600 ;
      RECT 0.0000 114.0600 480.2400 116.8000 ;
      RECT 0.8600 113.4000 480.2400 114.0600 ;
      RECT 0.0000 111.0000 480.2400 113.4000 ;
      RECT 0.8600 110.3400 480.2400 111.0000 ;
      RECT 0.0000 107.6000 480.2400 110.3400 ;
      RECT 0.8600 106.9400 480.2400 107.6000 ;
      RECT 0.0000 104.5400 480.2400 106.9400 ;
      RECT 0.8600 103.8800 480.2400 104.5400 ;
      RECT 0.0000 101.1400 480.2400 103.8800 ;
      RECT 0.8600 100.4800 480.2400 101.1400 ;
      RECT 0.0000 98.0800 480.2400 100.4800 ;
      RECT 0.8600 97.4200 480.2400 98.0800 ;
      RECT 0.0000 94.6800 480.2400 97.4200 ;
      RECT 0.8600 94.0200 480.2400 94.6800 ;
      RECT 0.0000 91.2800 480.2400 94.0200 ;
      RECT 0.8600 90.6200 480.2400 91.2800 ;
      RECT 0.0000 88.2200 480.2400 90.6200 ;
      RECT 0.8600 87.5600 480.2400 88.2200 ;
      RECT 0.0000 84.8200 480.2400 87.5600 ;
      RECT 0.8600 84.1600 480.2400 84.8200 ;
      RECT 0.0000 81.7600 480.2400 84.1600 ;
      RECT 0.8600 81.1000 480.2400 81.7600 ;
      RECT 0.0000 78.3600 480.2400 81.1000 ;
      RECT 0.8600 77.7000 480.2400 78.3600 ;
      RECT 0.0000 75.3000 480.2400 77.7000 ;
      RECT 0.8600 74.6400 480.2400 75.3000 ;
      RECT 0.0000 71.9000 480.2400 74.6400 ;
      RECT 0.8600 71.2400 480.2400 71.9000 ;
      RECT 0.0000 68.8400 480.2400 71.2400 ;
      RECT 0.8600 68.1800 480.2400 68.8400 ;
      RECT 0.0000 65.4400 480.2400 68.1800 ;
      RECT 0.8600 64.7800 480.2400 65.4400 ;
      RECT 0.0000 62.0400 480.2400 64.7800 ;
      RECT 0.8600 61.3800 480.2400 62.0400 ;
      RECT 0.0000 58.9800 480.2400 61.3800 ;
      RECT 0.8600 58.3200 480.2400 58.9800 ;
      RECT 0.0000 55.5800 480.2400 58.3200 ;
      RECT 0.8600 54.9200 480.2400 55.5800 ;
      RECT 0.0000 52.5200 480.2400 54.9200 ;
      RECT 0.8600 51.8600 480.2400 52.5200 ;
      RECT 0.0000 49.1200 480.2400 51.8600 ;
      RECT 0.8600 48.4600 480.2400 49.1200 ;
      RECT 0.0000 46.0600 480.2400 48.4600 ;
      RECT 0.8600 45.4000 480.2400 46.0600 ;
      RECT 0.0000 42.6600 480.2400 45.4000 ;
      RECT 0.8600 42.0000 480.2400 42.6600 ;
      RECT 0.0000 39.6000 480.2400 42.0000 ;
      RECT 0.8600 38.9400 480.2400 39.6000 ;
      RECT 0.0000 36.2000 480.2400 38.9400 ;
      RECT 0.8600 35.5400 480.2400 36.2000 ;
      RECT 0.0000 32.8000 480.2400 35.5400 ;
      RECT 0.8600 32.1400 480.2400 32.8000 ;
      RECT 0.0000 29.7400 480.2400 32.1400 ;
      RECT 0.8600 29.0800 480.2400 29.7400 ;
      RECT 0.0000 26.3400 480.2400 29.0800 ;
      RECT 0.8600 25.6800 480.2400 26.3400 ;
      RECT 0.0000 23.2800 480.2400 25.6800 ;
      RECT 0.8600 22.6200 480.2400 23.2800 ;
      RECT 0.0000 19.8800 480.2400 22.6200 ;
      RECT 0.8600 19.2200 480.2400 19.8800 ;
      RECT 0.0000 16.8200 480.2400 19.2200 ;
      RECT 0.8600 16.1600 480.2400 16.8200 ;
      RECT 0.0000 13.4200 480.2400 16.1600 ;
      RECT 0.8600 12.7600 480.2400 13.4200 ;
      RECT 0.0000 10.3600 480.2400 12.7600 ;
      RECT 0.8600 9.7000 480.2400 10.3600 ;
      RECT 0.0000 0.0000 480.2400 9.7000 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 480.2400 449.8200 ;
    LAYER met3 ;
      RECT 0.0000 447.0200 480.2400 449.8200 ;
      RECT 477.4800 444.9200 480.2400 447.0200 ;
      RECT 0.0000 444.9200 2.7600 447.0200 ;
      RECT 0.0000 444.5200 480.2400 444.9200 ;
      RECT 474.9800 442.4200 480.2400 444.5200 ;
      RECT 0.0000 442.4200 5.2600 444.5200 ;
      RECT 0.0000 435.3200 480.2400 442.4200 ;
      RECT 21.0650 433.2200 480.2400 435.3200 ;
      RECT 0.0000 433.2200 2.7600 435.3200 ;
      RECT 0.0000 252.7400 480.2400 433.2200 ;
      RECT 474.9800 250.6400 480.2400 252.7400 ;
      RECT 0.0000 250.6400 465.8650 252.7400 ;
      RECT 0.0000 53.9200 480.2400 250.6400 ;
      RECT 477.4800 52.8400 480.2400 53.9200 ;
      RECT 4.8600 52.8400 475.3800 53.9200 ;
      RECT 0.0000 52.8400 2.7600 53.9200 ;
      RECT 0.0000 51.2000 480.2400 52.8400 ;
      RECT 474.9800 50.1200 480.2400 51.2000 ;
      RECT 7.3600 50.1200 472.8800 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 480.2400 50.1200 ;
      RECT 477.4800 47.4000 480.2400 48.4800 ;
      RECT 4.8600 47.4000 475.3800 48.4800 ;
      RECT 0.0000 47.4000 2.7600 48.4800 ;
      RECT 0.0000 45.7600 480.2400 47.4000 ;
      RECT 474.9800 44.6800 480.2400 45.7600 ;
      RECT 7.3600 44.6800 472.8800 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 480.2400 44.6800 ;
      RECT 477.4800 41.9600 480.2400 43.0400 ;
      RECT 4.8600 41.9600 475.3800 43.0400 ;
      RECT 0.0000 41.9600 2.7600 43.0400 ;
      RECT 0.0000 40.3200 480.2400 41.9600 ;
      RECT 474.9800 39.2400 480.2400 40.3200 ;
      RECT 7.3600 39.2400 472.8800 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 480.2400 39.2400 ;
      RECT 477.4800 36.5200 480.2400 37.6000 ;
      RECT 4.8600 36.5200 475.3800 37.6000 ;
      RECT 0.0000 36.5200 2.7600 37.6000 ;
      RECT 0.0000 34.8800 480.2400 36.5200 ;
      RECT 474.9800 33.8000 480.2400 34.8800 ;
      RECT 7.3600 33.8000 472.8800 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 480.2400 33.8000 ;
      RECT 477.4800 31.0800 480.2400 32.1600 ;
      RECT 4.8600 31.0800 475.3800 32.1600 ;
      RECT 0.0000 31.0800 2.7600 32.1600 ;
      RECT 0.0000 29.4400 480.2400 31.0800 ;
      RECT 474.9800 28.3600 480.2400 29.4400 ;
      RECT 7.3600 28.3600 472.8800 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 480.2400 28.3600 ;
      RECT 477.4800 25.6400 480.2400 26.7200 ;
      RECT 4.8600 25.6400 475.3800 26.7200 ;
      RECT 0.0000 25.6400 2.7600 26.7200 ;
      RECT 0.0000 24.0000 480.2400 25.6400 ;
      RECT 474.9800 22.9200 480.2400 24.0000 ;
      RECT 7.3600 22.9200 472.8800 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 480.2400 22.9200 ;
      RECT 477.4800 20.2000 480.2400 21.2800 ;
      RECT 4.8600 20.2000 475.3800 21.2800 ;
      RECT 0.0000 20.2000 2.7600 21.2800 ;
      RECT 0.0000 18.5600 480.2400 20.2000 ;
      RECT 474.9800 17.4800 480.2400 18.5600 ;
      RECT 7.3600 17.4800 472.8800 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 480.2400 17.4800 ;
      RECT 477.4800 14.7600 480.2400 15.8400 ;
      RECT 4.8600 14.7600 475.3800 15.8400 ;
      RECT 0.0000 14.7600 2.7600 15.8400 ;
      RECT 0.0000 13.1200 480.2400 14.7600 ;
      RECT 474.9800 12.0400 480.2400 13.1200 ;
      RECT 7.3600 12.0400 472.8800 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 480.2400 12.0400 ;
      RECT 477.4800 9.3200 480.2400 10.4000 ;
      RECT 4.8600 9.3200 475.3800 10.4000 ;
      RECT 0.0000 9.3200 2.7600 10.4000 ;
      RECT 0.0000 7.2300 480.2400 9.3200 ;
      RECT 474.9800 5.1300 480.2400 7.2300 ;
      RECT 0.0000 5.1300 5.2600 7.2300 ;
      RECT 0.0000 4.7300 480.2400 5.1300 ;
      RECT 477.4800 2.6300 480.2400 4.7300 ;
      RECT 0.0000 2.6300 2.7600 4.7300 ;
      RECT 0.0000 0.0000 480.2400 2.6300 ;
    LAYER met4 ;
      RECT 0.0000 447.0200 480.2400 449.8200 ;
      RECT 4.8600 444.5200 475.3800 447.0200 ;
      RECT 474.9800 5.1300 475.3800 444.5200 ;
      RECT 7.3600 5.1300 472.8800 444.5200 ;
      RECT 4.8600 5.1300 5.2600 444.5200 ;
      RECT 477.4800 2.6300 480.2400 447.0200 ;
      RECT 4.8600 2.6300 475.3800 5.1300 ;
      RECT 0.0000 2.6300 2.7600 447.0200 ;
      RECT 0.0000 1.0200 480.2400 2.6300 ;
      RECT 10.1500 0.0000 480.2400 1.0200 ;
      RECT 0.0000 0.0000 9.1700 1.0200 ;
  END
END BlockRAM_1KB

END LIBRARY
