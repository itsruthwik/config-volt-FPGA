magic
tech sky130A
magscale 1 2
timestamp 1762063560
<< viali >>
rect 7021 22729 7055 22763
rect 8217 22729 8251 22763
rect 2789 22661 2823 22695
rect 9505 22661 9539 22695
rect 16221 22661 16255 22695
rect 18797 22661 18831 22695
rect 21005 22661 21039 22695
rect 5549 22593 5583 22627
rect 7113 22593 7147 22627
rect 8125 22593 8159 22627
rect 8401 22593 8435 22627
rect 9321 22593 9355 22627
rect 11805 22593 11839 22627
rect 13185 22593 13219 22627
rect 16124 22593 16158 22627
rect 16313 22593 16347 22627
rect 16497 22593 16531 22627
rect 17417 22593 17451 22627
rect 18653 22593 18687 22627
rect 18889 22593 18923 22627
rect 19073 22593 19107 22627
rect 19257 22593 19291 22627
rect 20729 22593 20763 22627
rect 20821 22593 20855 22627
rect 21097 22593 21131 22627
rect 21194 22593 21228 22627
rect 2697 22525 2731 22559
rect 2881 22525 2915 22559
rect 4813 22525 4847 22559
rect 7021 22525 7055 22559
rect 9597 22525 9631 22559
rect 16681 22525 16715 22559
rect 17969 22525 18003 22559
rect 19809 22525 19843 22559
rect 20177 22525 20211 22559
rect 6561 22457 6595 22491
rect 2329 22389 2363 22423
rect 5457 22389 5491 22423
rect 5733 22389 5767 22423
rect 8677 22389 8711 22423
rect 9045 22389 9079 22423
rect 11621 22389 11655 22423
rect 13001 22389 13035 22423
rect 15945 22389 15979 22423
rect 17325 22389 17359 22423
rect 18521 22389 18555 22423
rect 21373 22389 21407 22423
rect 7113 22185 7147 22219
rect 14197 22185 14231 22219
rect 7389 22117 7423 22151
rect 17785 22117 17819 22151
rect 5365 22049 5399 22083
rect 5733 22049 5767 22083
rect 9321 22049 9355 22083
rect 16405 22049 16439 22083
rect 18521 22049 18555 22083
rect 2053 21981 2087 22015
rect 2145 21981 2179 22015
rect 5641 21981 5675 22015
rect 5989 21981 6023 22015
rect 8769 21981 8803 22015
rect 9137 21981 9171 22015
rect 11109 21981 11143 22015
rect 11529 21981 11563 22015
rect 11621 21981 11655 22015
rect 12173 21981 12207 22015
rect 12449 21981 12483 22015
rect 12716 21981 12750 22015
rect 14749 21981 14783 22015
rect 15945 21981 15979 22015
rect 16672 21981 16706 22015
rect 19809 21981 19843 22015
rect 2412 21913 2446 21947
rect 5120 21913 5154 21947
rect 8524 21913 8558 21947
rect 9566 21913 9600 21947
rect 11253 21913 11287 21947
rect 11345 21913 11379 21947
rect 14473 21913 14507 21947
rect 15301 21913 15335 21947
rect 15577 21913 15611 21947
rect 18521 21913 18555 21947
rect 18613 21913 18647 21947
rect 20076 21913 20110 21947
rect 1869 21845 1903 21879
rect 3525 21845 3559 21879
rect 3985 21845 4019 21879
rect 5457 21845 5491 21879
rect 8953 21845 8987 21879
rect 10701 21845 10735 21879
rect 10960 21845 10994 21879
rect 13829 21845 13863 21879
rect 14657 21845 14691 21879
rect 15015 21845 15049 21879
rect 15485 21845 15519 21879
rect 15761 21845 15795 21879
rect 18051 21845 18085 21879
rect 21189 21845 21223 21879
rect 2973 21641 3007 21675
rect 3985 21641 4019 21675
rect 5733 21641 5767 21675
rect 9597 21641 9631 21675
rect 11253 21641 11287 21675
rect 12081 21641 12115 21675
rect 16773 21641 16807 21675
rect 19625 21641 19659 21675
rect 6469 21573 6503 21607
rect 7389 21573 7423 21607
rect 7573 21573 7607 21607
rect 10140 21573 10174 21607
rect 12173 21573 12207 21607
rect 20076 21573 20110 21607
rect 1409 21505 1443 21539
rect 1676 21505 1710 21539
rect 3157 21505 3191 21539
rect 4353 21505 4387 21539
rect 4620 21505 4654 21539
rect 6009 21505 6043 21539
rect 8217 21505 8251 21539
rect 8484 21505 8518 21539
rect 9873 21505 9907 21539
rect 11897 21505 11931 21539
rect 12725 21505 12759 21539
rect 13001 21505 13035 21539
rect 13257 21505 13291 21539
rect 14565 21505 14599 21539
rect 14832 21505 14866 21539
rect 16129 21505 16163 21539
rect 17886 21505 17920 21539
rect 18153 21505 18187 21539
rect 18245 21505 18279 21539
rect 18512 21505 18546 21539
rect 3893 21437 3927 21471
rect 4077 21437 4111 21471
rect 7665 21437 7699 21471
rect 19809 21437 19843 21471
rect 2789 21369 2823 21403
rect 3525 21369 3559 21403
rect 7113 21369 7147 21403
rect 11621 21369 11655 21403
rect 12909 21369 12943 21403
rect 16313 21369 16347 21403
rect 6193 21301 6227 21335
rect 6745 21301 6779 21335
rect 14381 21301 14415 21335
rect 15945 21301 15979 21335
rect 21189 21301 21223 21335
rect 3893 21097 3927 21131
rect 5273 21097 5307 21131
rect 6009 21097 6043 21131
rect 8953 21097 8987 21131
rect 9413 21097 9447 21131
rect 11897 21097 11931 21131
rect 14197 21097 14231 21131
rect 14933 21097 14967 21131
rect 16681 21097 16715 21131
rect 18613 21097 18647 21131
rect 2145 21029 2179 21063
rect 2973 21029 3007 21063
rect 7849 21029 7883 21063
rect 12541 21029 12575 21063
rect 2605 20961 2639 20995
rect 3433 20961 3467 20995
rect 4813 20961 4847 20995
rect 10517 20961 10551 20995
rect 13921 20961 13955 20995
rect 15301 20961 15335 20995
rect 4169 20893 4203 20927
rect 5457 20893 5491 20927
rect 5641 20893 5675 20927
rect 5733 20893 5767 20927
rect 5877 20893 5911 20927
rect 6193 20893 6227 20927
rect 6469 20893 6503 20927
rect 6725 20893 6759 20927
rect 9137 20893 9171 20927
rect 9597 20893 9631 20927
rect 9763 20893 9797 20927
rect 10057 20893 10091 20927
rect 10784 20893 10818 20927
rect 14473 20893 14507 20927
rect 15117 20893 15151 20927
rect 17233 20893 17267 20927
rect 18889 20893 18923 20927
rect 19257 20893 19291 20927
rect 21557 20893 21591 20927
rect 2697 20825 2731 20859
rect 3433 20825 3467 20859
rect 3525 20825 3559 20859
rect 4445 20825 4479 20859
rect 4721 20825 4755 20859
rect 8309 20825 8343 20859
rect 10333 20825 10367 20859
rect 13654 20825 13688 20859
rect 14657 20825 14691 20859
rect 14749 20825 14783 20859
rect 15568 20825 15602 20859
rect 17500 20825 17534 20859
rect 19502 20825 19536 20859
rect 2605 20757 2639 20791
rect 4353 20757 4387 20791
rect 4813 20757 4847 20791
rect 6377 20757 6411 20791
rect 8401 20757 8435 20791
rect 10241 20757 10275 20791
rect 19073 20757 19107 20791
rect 20637 20757 20671 20791
rect 21005 20757 21039 20791
rect 5917 20553 5951 20587
rect 6653 20553 6687 20587
rect 8677 20553 8711 20587
rect 9689 20553 9723 20587
rect 11345 20553 11379 20587
rect 14197 20553 14231 20587
rect 17509 20553 17543 20587
rect 18429 20553 18463 20587
rect 3525 20485 3559 20519
rect 3709 20485 3743 20519
rect 3801 20485 3835 20519
rect 4721 20485 4755 20519
rect 5365 20485 5399 20519
rect 5457 20485 5491 20519
rect 5825 20485 5859 20519
rect 8493 20485 8527 20519
rect 9505 20485 9539 20519
rect 12173 20485 12207 20519
rect 13185 20485 13219 20519
rect 14381 20485 14415 20519
rect 16129 20485 16163 20519
rect 16313 20485 16347 20519
rect 17049 20485 17083 20519
rect 17141 20485 17175 20519
rect 18613 20485 18647 20519
rect 1409 20417 1443 20451
rect 1676 20417 1710 20451
rect 5268 20417 5302 20451
rect 5641 20417 5675 20451
rect 7766 20417 7800 20451
rect 8033 20417 8067 20451
rect 10793 20417 10827 20451
rect 11989 20417 12023 20451
rect 12449 20417 12483 20451
rect 12909 20417 12943 20451
rect 13093 20417 13127 20451
rect 13282 20417 13316 20451
rect 16952 20417 16986 20451
rect 17325 20417 17359 20451
rect 17693 20417 17727 20451
rect 19073 20417 19107 20451
rect 20085 20417 20119 20451
rect 21045 20417 21079 20451
rect 21189 20417 21223 20451
rect 21281 20417 21315 20451
rect 21465 20417 21499 20451
rect 4629 20349 4663 20383
rect 4813 20349 4847 20383
rect 8769 20349 8803 20383
rect 9781 20349 9815 20383
rect 12265 20349 12299 20383
rect 14105 20349 14139 20383
rect 16405 20349 16439 20383
rect 18337 20349 18371 20383
rect 19809 20349 19843 20383
rect 2789 20281 2823 20315
rect 9229 20281 9263 20315
rect 11713 20281 11747 20315
rect 13461 20281 13495 20315
rect 14657 20281 14691 20315
rect 15853 20281 15887 20315
rect 16773 20281 16807 20315
rect 18889 20281 18923 20315
rect 3249 20213 3283 20247
rect 4261 20213 4295 20247
rect 5089 20213 5123 20247
rect 8217 20213 8251 20247
rect 12633 20213 12667 20247
rect 20729 20213 20763 20247
rect 20913 20213 20947 20247
rect 1777 20009 1811 20043
rect 3433 20009 3467 20043
rect 5917 20009 5951 20043
rect 7757 20009 7791 20043
rect 11713 20009 11747 20043
rect 13277 20009 13311 20043
rect 18981 20009 19015 20043
rect 21557 20009 21591 20043
rect 5733 19941 5767 19975
rect 9045 19941 9079 19975
rect 14197 19941 14231 19975
rect 16497 19941 16531 19975
rect 17877 19941 17911 19975
rect 6469 19873 6503 19907
rect 9505 19873 9539 19907
rect 13093 19873 13127 19907
rect 1961 19805 1995 19839
rect 2053 19805 2087 19839
rect 3985 19805 4019 19839
rect 4353 19805 4387 19839
rect 7941 19805 7975 19839
rect 9597 19805 9631 19839
rect 11253 19805 11287 19839
rect 12826 19805 12860 19839
rect 14473 19805 14507 19839
rect 15117 19805 15151 19839
rect 16129 19805 16163 19839
rect 18061 19805 18095 19839
rect 18521 19805 18555 19839
rect 18613 19805 18647 19839
rect 18797 19805 18831 19839
rect 20177 19805 20211 19839
rect 20444 19805 20478 19839
rect 2320 19737 2354 19771
rect 4620 19737 4654 19771
rect 7297 19737 7331 19771
rect 7573 19737 7607 19771
rect 10609 19737 10643 19771
rect 13553 19737 13587 19771
rect 13737 19737 13771 19771
rect 13829 19737 13863 19771
rect 14749 19737 14783 19771
rect 16773 19737 16807 19771
rect 16957 19737 16991 19771
rect 17049 19737 17083 19771
rect 17325 19737 17359 19771
rect 17601 19737 17635 19771
rect 19441 19737 19475 19771
rect 19533 19737 19567 19771
rect 19717 19737 19751 19771
rect 3801 19669 3835 19703
rect 7003 19669 7037 19703
rect 7481 19669 7515 19703
rect 9505 19669 9539 19703
rect 10885 19669 10919 19703
rect 11437 19669 11471 19703
rect 14657 19669 14691 19703
rect 14933 19669 14967 19703
rect 16313 19669 16347 19703
rect 17417 19669 17451 19703
rect 18245 19669 18279 19703
rect 20011 19669 20045 19703
rect 2237 19465 2271 19499
rect 4721 19465 4755 19499
rect 6009 19465 6043 19499
rect 7839 19465 7873 19499
rect 8309 19465 8343 19499
rect 9873 19465 9907 19499
rect 12909 19465 12943 19499
rect 14657 19465 14691 19499
rect 16221 19465 16255 19499
rect 18061 19465 18095 19499
rect 19625 19465 19659 19499
rect 21189 19465 21223 19499
rect 21373 19465 21407 19499
rect 2513 19397 2547 19431
rect 3608 19397 3642 19431
rect 5825 19397 5859 19431
rect 6101 19397 6135 19431
rect 7481 19397 7515 19431
rect 7573 19397 7607 19431
rect 15108 19397 15142 19431
rect 20076 19397 20110 19431
rect 2053 19329 2087 19363
rect 3249 19329 3283 19363
rect 3341 19329 3375 19363
rect 6469 19329 6503 19363
rect 8125 19329 8159 19363
rect 8401 19329 8435 19363
rect 8585 19329 8619 19363
rect 10986 19329 11020 19363
rect 11253 19329 11287 19363
rect 11529 19329 11563 19363
rect 11785 19329 11819 19363
rect 13277 19329 13311 19363
rect 13544 19329 13578 19363
rect 14841 19329 14875 19363
rect 16681 19329 16715 19363
rect 16948 19329 16982 19363
rect 18245 19329 18279 19363
rect 18501 19329 18535 19363
rect 19809 19329 19843 19363
rect 21557 19329 21591 19363
rect 7481 19261 7515 19295
rect 9321 19261 9355 19295
rect 5549 19125 5583 19159
rect 6745 19125 6779 19159
rect 7021 19125 7055 19159
rect 2789 18921 2823 18955
rect 4721 18921 4755 18955
rect 7941 18921 7975 18955
rect 10701 18921 10735 18955
rect 13737 18921 13771 18955
rect 15209 18921 15243 18955
rect 17601 18921 17635 18955
rect 18245 18921 18279 18955
rect 20637 18921 20671 18955
rect 3893 18853 3927 18887
rect 10977 18853 11011 18887
rect 16129 18853 16163 18887
rect 21373 18853 21407 18887
rect 3065 18785 3099 18819
rect 4353 18785 4387 18819
rect 6101 18785 6135 18819
rect 6561 18785 6595 18819
rect 8953 18785 8987 18819
rect 12357 18785 12391 18819
rect 14197 18785 14231 18819
rect 16221 18785 16255 18819
rect 18705 18785 18739 18819
rect 1409 18717 1443 18751
rect 3617 18717 3651 18751
rect 6285 18717 6319 18751
rect 8309 18717 8343 18751
rect 8585 18717 8619 18751
rect 10517 18717 10551 18751
rect 11253 18717 11287 18751
rect 15485 18717 15519 18751
rect 15945 18717 15979 18751
rect 17785 18717 17819 18751
rect 19257 18717 19291 18751
rect 20821 18717 20855 18751
rect 21097 18717 21131 18751
rect 21241 18717 21275 18751
rect 1654 18649 1688 18683
rect 4445 18649 4479 18683
rect 5856 18649 5890 18683
rect 6806 18649 6840 18683
rect 9198 18649 9232 18683
rect 11529 18649 11563 18683
rect 12624 18649 12658 18683
rect 15025 18649 15059 18683
rect 15761 18649 15795 18683
rect 16466 18649 16500 18683
rect 18797 18649 18831 18683
rect 19524 18649 19558 18683
rect 21005 18649 21039 18683
rect 4353 18581 4387 18615
rect 6469 18581 6503 18615
rect 8493 18581 8527 18615
rect 8769 18581 8803 18615
rect 10333 18581 10367 18615
rect 11437 18581 11471 18615
rect 15669 18581 15703 18615
rect 17969 18581 18003 18615
rect 18705 18581 18739 18615
rect 1501 18377 1535 18411
rect 2697 18377 2731 18411
rect 4353 18377 4387 18411
rect 6193 18377 6227 18411
rect 7757 18377 7791 18411
rect 9873 18377 9907 18411
rect 10609 18377 10643 18411
rect 12725 18377 12759 18411
rect 13461 18377 13495 18411
rect 14657 18377 14691 18411
rect 17233 18377 17267 18411
rect 2329 18309 2363 18343
rect 6622 18309 6656 18343
rect 10425 18309 10459 18343
rect 12081 18309 12115 18343
rect 13921 18309 13955 18343
rect 14473 18309 14507 18343
rect 17049 18309 17083 18343
rect 18153 18309 18187 18343
rect 18245 18309 18279 18343
rect 1685 18241 1719 18275
rect 2145 18241 2179 18275
rect 3821 18241 3855 18275
rect 4077 18241 4111 18275
rect 5477 18241 5511 18275
rect 6009 18241 6043 18275
rect 8493 18241 8527 18275
rect 8749 18241 8783 18275
rect 10701 18241 10735 18275
rect 12173 18241 12207 18275
rect 12541 18241 12575 18275
rect 13001 18241 13035 18275
rect 13277 18241 13311 18275
rect 14749 18241 14783 18275
rect 15117 18241 15151 18275
rect 17969 18241 18003 18275
rect 18389 18241 18423 18275
rect 18705 18241 18739 18275
rect 2421 18173 2455 18207
rect 5733 18173 5767 18207
rect 6377 18173 6411 18207
rect 12081 18173 12115 18207
rect 17325 18173 17359 18207
rect 19441 18173 19475 18207
rect 20361 18173 20395 18207
rect 21005 18173 21039 18207
rect 1869 18105 1903 18139
rect 10149 18105 10183 18139
rect 11621 18105 11655 18139
rect 14197 18105 14231 18139
rect 16773 18105 16807 18139
rect 18521 18105 18555 18139
rect 12817 18037 12851 18071
rect 13645 18037 13679 18071
rect 14933 18037 14967 18071
rect 19717 18037 19751 18071
rect 21649 18037 21683 18071
rect 3249 17833 3283 17867
rect 3617 17833 3651 17867
rect 6101 17833 6135 17867
rect 6285 17833 6319 17867
rect 9689 17833 9723 17867
rect 12357 17833 12391 17867
rect 13185 17833 13219 17867
rect 17693 17833 17727 17867
rect 21557 17833 21591 17867
rect 3893 17765 3927 17799
rect 6653 17765 6687 17799
rect 8493 17765 8527 17799
rect 10885 17765 10919 17799
rect 15209 17765 15243 17799
rect 17325 17765 17359 17799
rect 18521 17765 18555 17799
rect 4353 17697 4387 17731
rect 7205 17697 7239 17731
rect 8125 17697 8159 17731
rect 11345 17697 11379 17731
rect 11437 17697 11471 17731
rect 13737 17697 13771 17731
rect 18337 17697 18371 17731
rect 19441 17697 19475 17731
rect 20177 17697 20211 17731
rect 1869 17629 1903 17663
rect 3433 17629 3467 17663
rect 4813 17629 4847 17663
rect 5549 17629 5583 17663
rect 5733 17629 5767 17663
rect 5825 17629 5859 17663
rect 5922 17629 5956 17663
rect 6469 17629 6503 17663
rect 7941 17629 7975 17663
rect 9965 17629 9999 17663
rect 10701 17629 10735 17663
rect 14197 17629 14231 17663
rect 15388 17629 15422 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 16405 17629 16439 17663
rect 16773 17629 16807 17663
rect 16865 17629 16899 17663
rect 17141 17629 17175 17663
rect 18653 17629 18687 17663
rect 18797 17629 18831 17663
rect 19073 17629 19107 17663
rect 19717 17629 19751 17663
rect 2114 17561 2148 17595
rect 4353 17561 4387 17595
rect 4445 17561 4479 17595
rect 6929 17561 6963 17595
rect 10241 17561 10275 17595
rect 11345 17561 11379 17595
rect 12633 17561 12667 17595
rect 12909 17561 12943 17595
rect 13461 17561 13495 17595
rect 15025 17561 15059 17595
rect 15485 17561 15519 17595
rect 15577 17561 15611 17595
rect 18889 17561 18923 17595
rect 20444 17561 20478 17595
rect 5457 17493 5491 17527
rect 7113 17493 7147 17527
rect 8033 17493 8067 17527
rect 10149 17493 10183 17527
rect 10517 17493 10551 17527
rect 12817 17493 12851 17527
rect 13645 17493 13679 17527
rect 16589 17493 16623 17527
rect 17049 17493 17083 17527
rect 19533 17493 19567 17527
rect 20011 17493 20045 17527
rect 5199 17289 5233 17323
rect 7095 17289 7129 17323
rect 11253 17289 11287 17323
rect 14087 17289 14121 17323
rect 16313 17289 16347 17323
rect 19441 17289 19475 17323
rect 21557 17289 21591 17323
rect 2789 17221 2823 17255
rect 3065 17221 3099 17255
rect 3801 17221 3835 17255
rect 4721 17221 4755 17255
rect 5641 17221 5675 17255
rect 7573 17221 7607 17255
rect 8033 17221 8067 17255
rect 10140 17221 10174 17255
rect 12081 17221 12115 17255
rect 12716 17221 12750 17255
rect 14565 17221 14599 17255
rect 15200 17221 15234 17255
rect 17233 17221 17267 17255
rect 2145 17153 2179 17187
rect 2605 17153 2639 17187
rect 5365 17153 5399 17187
rect 5549 17153 5583 17187
rect 5785 17153 5819 17187
rect 6561 17153 6595 17187
rect 6745 17153 6779 17187
rect 11897 17153 11931 17187
rect 14933 17153 14967 17187
rect 17325 17153 17359 17187
rect 17877 17153 17911 17187
rect 18061 17153 18095 17187
rect 18328 17153 18362 17187
rect 19809 17153 19843 17187
rect 20085 17153 20119 17187
rect 20444 17153 20478 17187
rect 2881 17085 2915 17119
rect 4629 17085 4663 17119
rect 4813 17085 4847 17119
rect 7573 17085 7607 17119
rect 7665 17085 7699 17119
rect 8861 17085 8895 17119
rect 9873 17085 9907 17119
rect 12173 17085 12207 17119
rect 12449 17085 12483 17119
rect 14565 17085 14599 17119
rect 14657 17085 14691 17119
rect 17141 17085 17175 17119
rect 20177 17085 20211 17119
rect 1961 17017 1995 17051
rect 2329 17017 2363 17051
rect 13829 17017 13863 17051
rect 5917 16949 5951 16983
rect 6377 16949 6411 16983
rect 6929 16949 6963 16983
rect 11621 16949 11655 16983
rect 16773 16949 16807 16983
rect 17693 16949 17727 16983
rect 19625 16949 19659 16983
rect 19901 16949 19935 16983
rect 5365 16745 5399 16779
rect 10057 16745 10091 16779
rect 11805 16745 11839 16779
rect 13829 16745 13863 16779
rect 20637 16745 20671 16779
rect 21465 16745 21499 16779
rect 8217 16677 8251 16711
rect 9229 16677 9263 16711
rect 15485 16677 15519 16711
rect 4353 16609 4387 16643
rect 6745 16609 6779 16643
rect 6837 16609 6871 16643
rect 10425 16609 10459 16643
rect 14105 16609 14139 16643
rect 15853 16609 15887 16643
rect 17417 16609 17451 16643
rect 19257 16609 19291 16643
rect 21005 16609 21039 16643
rect 1409 16541 1443 16575
rect 3157 16541 3191 16575
rect 3617 16541 3651 16575
rect 4445 16541 4479 16575
rect 6478 16541 6512 16575
rect 7093 16541 7127 16575
rect 8493 16541 8527 16575
rect 9045 16541 9079 16575
rect 9597 16541 9631 16575
rect 10681 16541 10715 16575
rect 12173 16541 12207 16575
rect 12449 16541 12483 16575
rect 14372 16541 14406 16575
rect 16120 16541 16154 16575
rect 17684 16541 17718 16575
rect 20913 16541 20947 16575
rect 1676 16473 1710 16507
rect 9965 16473 9999 16507
rect 12694 16473 12728 16507
rect 19524 16473 19558 16507
rect 2789 16405 2823 16439
rect 2973 16405 3007 16439
rect 3433 16405 3467 16439
rect 3875 16405 3909 16439
rect 4353 16405 4387 16439
rect 8677 16405 8711 16439
rect 9781 16405 9815 16439
rect 12357 16405 12391 16439
rect 17233 16405 17267 16439
rect 18797 16405 18831 16439
rect 21005 16405 21039 16439
rect 1685 16201 1719 16235
rect 2513 16201 2547 16235
rect 4169 16201 4203 16235
rect 7757 16201 7791 16235
rect 8493 16201 8527 16235
rect 10333 16201 10367 16235
rect 12081 16201 12115 16235
rect 12817 16201 12851 16235
rect 20821 16201 20855 16235
rect 3056 16133 3090 16167
rect 5558 16133 5592 16167
rect 8309 16133 8343 16167
rect 11253 16133 11287 16167
rect 12173 16133 12207 16167
rect 13461 16133 13495 16167
rect 13982 16133 14016 16167
rect 15853 16133 15887 16167
rect 15945 16133 15979 16167
rect 16129 16133 16163 16167
rect 18613 16133 18647 16167
rect 18797 16133 18831 16167
rect 21373 16133 21407 16167
rect 1869 16065 1903 16099
rect 2329 16065 2363 16099
rect 5825 16065 5859 16099
rect 5917 16065 5951 16099
rect 6377 16065 6411 16099
rect 6633 16065 6667 16099
rect 8953 16065 8987 16099
rect 9209 16065 9243 16099
rect 11897 16065 11931 16099
rect 12633 16065 12667 16099
rect 13553 16065 13587 16099
rect 15485 16065 15519 16099
rect 16681 16065 16715 16099
rect 16948 16065 16982 16099
rect 19441 16065 19475 16099
rect 19708 16065 19742 16099
rect 21229 16065 21263 16099
rect 21465 16065 21499 16099
rect 21649 16065 21683 16099
rect 2605 15997 2639 16031
rect 2789 15997 2823 16031
rect 8585 15997 8619 16031
rect 13461 15997 13495 16031
rect 13737 15997 13771 16031
rect 18889 15997 18923 16031
rect 2053 15929 2087 15963
rect 6101 15929 6135 15963
rect 8033 15929 8067 15963
rect 11621 15929 11655 15963
rect 13001 15929 13035 15963
rect 15117 15929 15151 15963
rect 16405 15929 16439 15963
rect 18337 15929 18371 15963
rect 21097 15929 21131 15963
rect 4445 15861 4479 15895
rect 11161 15861 11195 15895
rect 15669 15861 15703 15895
rect 18061 15861 18095 15895
rect 3893 15657 3927 15691
rect 6101 15657 6135 15691
rect 7297 15657 7331 15691
rect 10057 15657 10091 15691
rect 10241 15657 10275 15691
rect 11069 15657 11103 15691
rect 13185 15657 13219 15691
rect 15025 15657 15059 15691
rect 16589 15657 16623 15691
rect 3525 15589 3559 15623
rect 9597 15589 9631 15623
rect 20729 15589 20763 15623
rect 4261 15521 4295 15555
rect 4445 15521 4479 15555
rect 5549 15521 5583 15555
rect 13645 15521 13679 15555
rect 14473 15521 14507 15555
rect 14565 15521 14599 15555
rect 17049 15521 17083 15555
rect 17141 15521 17175 15555
rect 21189 15521 21223 15555
rect 2145 15453 2179 15487
rect 5825 15453 5859 15487
rect 7481 15453 7515 15487
rect 8953 15453 8987 15487
rect 10701 15453 10735 15487
rect 11345 15453 11379 15487
rect 11621 15453 11655 15487
rect 13737 15453 13771 15487
rect 15945 15453 15979 15487
rect 17877 15453 17911 15487
rect 2412 15385 2446 15419
rect 4353 15385 4387 15419
rect 5641 15385 5675 15419
rect 9781 15385 9815 15419
rect 10609 15385 10643 15419
rect 14565 15385 14599 15419
rect 21281 15385 21315 15419
rect 9045 15317 9079 15351
rect 10232 15317 10266 15351
rect 11078 15317 11112 15351
rect 11437 15317 11471 15351
rect 13645 15317 13679 15351
rect 16129 15317 16163 15351
rect 17049 15317 17083 15351
rect 17693 15317 17727 15351
rect 21189 15317 21223 15351
rect 3709 15113 3743 15147
rect 10701 15113 10735 15147
rect 20085 15113 20119 15147
rect 3525 15045 3559 15079
rect 10333 15045 10367 15079
rect 10517 15045 10551 15079
rect 10885 15045 10919 15079
rect 11253 15045 11287 15079
rect 12081 15045 12115 15079
rect 13461 15045 13495 15079
rect 16313 15045 16347 15079
rect 20422 15045 20456 15079
rect 3065 14977 3099 15011
rect 8125 14977 8159 15011
rect 11897 14977 11931 15011
rect 13185 14977 13219 15011
rect 15485 14977 15519 15011
rect 16129 14977 16163 15011
rect 17233 14977 17267 15011
rect 17489 14977 17523 15011
rect 19625 14977 19659 15011
rect 19901 14977 19935 15011
rect 3801 14909 3835 14943
rect 8401 14909 8435 14943
rect 12173 14909 12207 14943
rect 13369 14909 13403 14943
rect 16405 14909 16439 14943
rect 20177 14909 20211 14943
rect 3249 14841 3283 14875
rect 11621 14841 11655 14875
rect 15853 14841 15887 14875
rect 2973 14773 3007 14807
rect 9873 14773 9907 14807
rect 10517 14773 10551 14807
rect 13001 14773 13035 14807
rect 13461 14773 13495 14807
rect 15301 14773 15335 14807
rect 18613 14773 18647 14807
rect 19441 14773 19475 14807
rect 21557 14773 21591 14807
rect 5825 14569 5859 14603
rect 10057 14569 10091 14603
rect 11989 14569 12023 14603
rect 17969 14569 18003 14603
rect 18245 14569 18279 14603
rect 20913 14569 20947 14603
rect 9045 14501 9079 14535
rect 20637 14501 20671 14535
rect 1593 14433 1627 14467
rect 5365 14433 5399 14467
rect 7757 14433 7791 14467
rect 8493 14433 8527 14467
rect 10609 14433 10643 14467
rect 15025 14433 15059 14467
rect 18797 14433 18831 14467
rect 21373 14433 21407 14467
rect 21465 14433 21499 14467
rect 3985 14365 4019 14399
rect 4169 14365 4203 14399
rect 4445 14365 4479 14399
rect 4537 14365 4571 14399
rect 4905 14365 4939 14399
rect 5089 14365 5123 14399
rect 5641 14365 5675 14399
rect 6469 14365 6503 14399
rect 6653 14365 6687 14399
rect 7389 14365 7423 14399
rect 9781 14365 9815 14399
rect 10876 14365 10910 14399
rect 12173 14365 12207 14399
rect 13737 14365 13771 14399
rect 14749 14365 14783 14399
rect 15292 14365 15326 14399
rect 16589 14365 16623 14399
rect 18521 14365 18555 14399
rect 19257 14365 19291 14399
rect 1869 14297 1903 14331
rect 3801 14297 3835 14331
rect 4813 14297 4847 14331
rect 9321 14297 9355 14331
rect 9597 14297 9631 14331
rect 10057 14297 10091 14331
rect 10241 14297 10275 14331
rect 12440 14297 12474 14331
rect 16834 14297 16868 14331
rect 19524 14297 19558 14331
rect 3341 14229 3375 14263
rect 6285 14229 6319 14263
rect 6745 14229 6779 14263
rect 7573 14229 7607 14263
rect 9505 14229 9539 14263
rect 13553 14229 13587 14263
rect 13921 14229 13955 14263
rect 14933 14229 14967 14263
rect 16405 14229 16439 14263
rect 18705 14229 18739 14263
rect 21373 14229 21407 14263
rect 1593 14025 1627 14059
rect 5825 14025 5859 14059
rect 6561 14025 6595 14059
rect 11805 14025 11839 14059
rect 17233 14025 17267 14059
rect 18705 14025 18739 14059
rect 21281 14025 21315 14059
rect 2053 13957 2087 13991
rect 3249 13957 3283 13991
rect 5365 13957 5399 13991
rect 5641 13957 5675 13991
rect 7849 13957 7883 13991
rect 10425 13957 10459 13991
rect 12449 13957 12483 13991
rect 13930 13957 13964 13991
rect 14657 13957 14691 13991
rect 14841 13957 14875 13991
rect 15853 13957 15887 13991
rect 16037 13957 16071 13991
rect 17592 13957 17626 13991
rect 20637 13957 20671 13991
rect 20821 13957 20855 13991
rect 1685 13889 1719 13923
rect 2789 13889 2823 13923
rect 2973 13889 3007 13923
rect 5181 13889 5215 13923
rect 6193 13889 6227 13923
rect 6561 13889 6595 13923
rect 7113 13889 7147 13923
rect 7389 13889 7423 13923
rect 7573 13889 7607 13923
rect 9781 13889 9815 13923
rect 9965 13889 9999 13923
rect 10333 13889 10367 13923
rect 10701 13889 10735 13923
rect 10793 13889 10827 13923
rect 11069 13889 11103 13923
rect 11253 13889 11287 13923
rect 11621 13889 11655 13923
rect 11971 13889 12005 13923
rect 12265 13889 12299 13923
rect 14933 13889 14967 13923
rect 17049 13889 17083 13923
rect 17325 13889 17359 13923
rect 18889 13889 18923 13923
rect 19145 13889 19179 13923
rect 21465 13889 21499 13923
rect 4721 13821 4755 13855
rect 4905 13821 4939 13855
rect 5273 13821 5307 13855
rect 6101 13821 6135 13855
rect 6377 13821 6411 13855
rect 6929 13821 6963 13855
rect 7481 13821 7515 13855
rect 9321 13821 9355 13855
rect 12541 13821 12575 13855
rect 14197 13821 14231 13855
rect 16129 13821 16163 13855
rect 20545 13821 20579 13855
rect 15577 13753 15611 13787
rect 21097 13753 21131 13787
rect 6009 13685 6043 13719
rect 9597 13685 9631 13719
rect 12817 13685 12851 13719
rect 14381 13685 14415 13719
rect 20269 13685 20303 13719
rect 3525 13481 3559 13515
rect 4537 13481 4571 13515
rect 4905 13481 4939 13515
rect 5181 13481 5215 13515
rect 5273 13481 5307 13515
rect 7757 13481 7791 13515
rect 8585 13481 8619 13515
rect 9137 13481 9171 13515
rect 10793 13481 10827 13515
rect 12173 13481 12207 13515
rect 13645 13481 13679 13515
rect 17785 13481 17819 13515
rect 19257 13481 19291 13515
rect 21373 13481 21407 13515
rect 16773 13413 16807 13447
rect 1777 13345 1811 13379
rect 4353 13345 4387 13379
rect 5365 13345 5399 13379
rect 5641 13345 5675 13379
rect 5733 13345 5767 13379
rect 6009 13345 6043 13379
rect 7481 13345 7515 13379
rect 7941 13345 7975 13379
rect 8125 13345 8159 13379
rect 9689 13345 9723 13379
rect 9873 13345 9907 13379
rect 10425 13345 10459 13379
rect 12265 13345 12299 13379
rect 15945 13345 15979 13379
rect 18245 13345 18279 13379
rect 19993 13345 20027 13379
rect 3801 13277 3835 13311
rect 3985 13277 4019 13311
rect 4629 13277 4663 13311
rect 8217 13277 8251 13311
rect 8493 13277 8527 13311
rect 9230 13277 9264 13311
rect 9597 13277 9631 13311
rect 9781 13277 9815 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 10609 13277 10643 13311
rect 11989 13277 12023 13311
rect 15669 13277 15703 13311
rect 19441 13277 19475 13311
rect 20260 13277 20294 13311
rect 2053 13209 2087 13243
rect 12510 13209 12544 13243
rect 15853 13209 15887 13243
rect 16221 13209 16255 13243
rect 16313 13209 16347 13243
rect 16497 13209 16531 13243
rect 18337 13209 18371 13243
rect 3985 13141 4019 13175
rect 5549 13141 5583 13175
rect 15375 13141 15409 13175
rect 18245 13141 18279 13175
rect 3065 12937 3099 12971
rect 4169 12937 4203 12971
rect 4353 12937 4387 12971
rect 5457 12937 5491 12971
rect 6469 12937 6503 12971
rect 11897 12937 11931 12971
rect 14749 12937 14783 12971
rect 16221 12937 16255 12971
rect 18061 12937 18095 12971
rect 20269 12937 20303 12971
rect 4537 12869 4571 12903
rect 6193 12869 6227 12903
rect 7297 12869 7331 12903
rect 7389 12869 7423 12903
rect 10333 12869 10367 12903
rect 13185 12869 13219 12903
rect 13277 12869 13311 12903
rect 15086 12869 15120 12903
rect 18153 12869 18187 12903
rect 18889 12869 18923 12903
rect 20453 12869 20487 12903
rect 3157 12801 3191 12835
rect 5089 12801 5123 12835
rect 5365 12801 5399 12835
rect 5917 12801 5951 12835
rect 6101 12801 6135 12835
rect 6653 12801 6687 12835
rect 7757 12801 7791 12835
rect 8125 12801 8159 12835
rect 8401 12801 8435 12835
rect 8585 12801 8619 12835
rect 8953 12801 8987 12835
rect 9137 12801 9171 12835
rect 10057 12801 10091 12835
rect 10517 12801 10551 12835
rect 10701 12801 10735 12835
rect 12173 12801 12207 12835
rect 12541 12801 12575 12835
rect 14565 12801 14599 12835
rect 16865 12801 16899 12835
rect 18705 12801 18739 12835
rect 20177 12801 20211 12835
rect 7297 12733 7331 12767
rect 7941 12733 7975 12767
rect 8493 12733 8527 12767
rect 9781 12733 9815 12767
rect 9873 12733 9907 12767
rect 9965 12733 9999 12767
rect 12357 12733 12391 12767
rect 13277 12733 13311 12767
rect 14841 12733 14875 12767
rect 18061 12733 18095 12767
rect 18981 12733 19015 12767
rect 7665 12665 7699 12699
rect 8677 12665 8711 12699
rect 12265 12665 12299 12699
rect 13737 12665 13771 12699
rect 20729 12665 20763 12699
rect 4353 12597 4387 12631
rect 4905 12597 4939 12631
rect 5733 12597 5767 12631
rect 6837 12597 6871 12631
rect 10241 12597 10275 12631
rect 12449 12597 12483 12631
rect 16681 12597 16715 12631
rect 17601 12597 17635 12631
rect 18429 12597 18463 12631
rect 6745 12393 6779 12427
rect 11161 12393 11195 12427
rect 13737 12393 13771 12427
rect 16313 12393 16347 12427
rect 2421 12325 2455 12359
rect 9045 12325 9079 12359
rect 10793 12325 10827 12359
rect 18521 12325 18555 12359
rect 21189 12325 21223 12359
rect 2881 12257 2915 12291
rect 4997 12257 5031 12291
rect 5273 12257 5307 12291
rect 7941 12257 7975 12291
rect 10609 12257 10643 12291
rect 13277 12257 13311 12291
rect 20269 12257 20303 12291
rect 2145 12189 2179 12223
rect 4353 12189 4387 12223
rect 7665 12189 7699 12223
rect 8493 12189 8527 12223
rect 8585 12189 8619 12223
rect 8677 12189 8711 12223
rect 9413 12189 9447 12223
rect 9781 12189 9815 12223
rect 10057 12189 10091 12223
rect 10149 12189 10183 12223
rect 10425 12189 10459 12223
rect 10977 12189 11011 12223
rect 11437 12189 11471 12223
rect 11529 12189 11563 12223
rect 13369 12189 13403 12223
rect 13829 12189 13863 12223
rect 14933 12189 14967 12223
rect 16589 12189 16623 12223
rect 16865 12189 16899 12223
rect 17141 12189 17175 12223
rect 20637 12189 20671 12223
rect 2973 12121 3007 12155
rect 4629 12121 4663 12155
rect 10517 12121 10551 12155
rect 15200 12121 15234 12155
rect 17386 12121 17420 12155
rect 20361 12121 20395 12155
rect 20913 12121 20947 12155
rect 1961 12053 1995 12087
rect 2881 12053 2915 12087
rect 4059 12053 4093 12087
rect 4537 12053 4571 12087
rect 7757 12053 7791 12087
rect 8125 12053 8159 12087
rect 9965 12053 9999 12087
rect 11253 12053 11287 12087
rect 13553 12053 13587 12087
rect 16773 12053 16807 12087
rect 17049 12053 17083 12087
rect 19791 12053 19825 12087
rect 20269 12053 20303 12087
rect 20729 12053 20763 12087
rect 3525 11849 3559 11883
rect 9321 11849 9355 11883
rect 10149 11849 10183 11883
rect 11713 11849 11747 11883
rect 15301 11849 15335 11883
rect 18521 11849 18555 11883
rect 19441 11849 19475 11883
rect 20913 11849 20947 11883
rect 3862 11781 3896 11815
rect 10241 11781 10275 11815
rect 11161 11781 11195 11815
rect 11253 11781 11287 11815
rect 16037 11781 16071 11815
rect 17386 11781 17420 11815
rect 19778 11781 19812 11815
rect 1593 11713 1627 11747
rect 1860 11713 1894 11747
rect 3341 11713 3375 11747
rect 5365 11713 5399 11747
rect 10057 11713 10091 11747
rect 11529 11713 11563 11747
rect 11897 11713 11931 11747
rect 12173 11713 12207 11747
rect 13470 11713 13504 11747
rect 13829 11713 13863 11747
rect 15117 11713 15151 11747
rect 15853 11713 15887 11747
rect 16497 11713 16531 11747
rect 17141 11713 17175 11747
rect 19257 11713 19291 11747
rect 21281 11713 21315 11747
rect 3617 11645 3651 11679
rect 7573 11645 7607 11679
rect 7849 11645 7883 11679
rect 9505 11645 9539 11679
rect 9689 11645 9723 11679
rect 11161 11645 11195 11679
rect 13737 11645 13771 11679
rect 16129 11645 16163 11679
rect 19533 11645 19567 11679
rect 4997 11577 5031 11611
rect 10701 11577 10735 11611
rect 12357 11577 12391 11611
rect 2973 11509 3007 11543
rect 5181 11509 5215 11543
rect 11897 11509 11931 11543
rect 14013 11509 14047 11543
rect 15577 11509 15611 11543
rect 16313 11509 16347 11543
rect 21097 11509 21131 11543
rect 4353 11305 4387 11339
rect 9781 11305 9815 11339
rect 10609 11305 10643 11339
rect 12357 11305 12391 11339
rect 13277 11305 13311 11339
rect 13737 11305 13771 11339
rect 14197 11305 14231 11339
rect 16773 11305 16807 11339
rect 21373 11305 21407 11339
rect 1685 11237 1719 11271
rect 6653 11237 6687 11271
rect 7297 11237 7331 11271
rect 17693 11237 17727 11271
rect 9387 11169 9421 11203
rect 10241 11169 10275 11203
rect 14565 11169 14599 11203
rect 17233 11169 17267 11203
rect 18245 11169 18279 11203
rect 19993 11169 20027 11203
rect 1501 11101 1535 11135
rect 1777 11101 1811 11135
rect 2033 11101 2067 11135
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 4221 11101 4255 11135
rect 4537 11101 4571 11135
rect 4804 11101 4838 11135
rect 6101 11101 6135 11135
rect 6521 11101 6555 11135
rect 8677 11101 8711 11135
rect 9229 11101 9263 11135
rect 9597 11101 9631 11135
rect 10057 11101 10091 11135
rect 10425 11101 10459 11135
rect 10977 11101 11011 11135
rect 11244 11101 11278 11135
rect 13645 11101 13679 11135
rect 15117 11101 15151 11135
rect 15384 11101 15418 11135
rect 19717 11101 19751 11135
rect 20260 11101 20294 11135
rect 4077 11033 4111 11067
rect 6285 11033 6319 11067
rect 6377 11033 6411 11067
rect 6929 11033 6963 11067
rect 7113 11033 7147 11067
rect 8125 11033 8159 11067
rect 12725 11033 12759 11067
rect 13001 11033 13035 11067
rect 13461 11033 13495 11067
rect 14749 11033 14783 11067
rect 17325 11033 17359 11067
rect 17969 11033 18003 11067
rect 3157 10965 3191 10999
rect 5917 10965 5951 10999
rect 7849 10965 7883 10999
rect 8401 10965 8435 10999
rect 9873 10965 9907 10999
rect 12817 10965 12851 10999
rect 14657 10965 14691 10999
rect 16497 10965 16531 10999
rect 17233 10965 17267 10999
rect 18153 10965 18187 10999
rect 19901 10965 19935 10999
rect 3801 10761 3835 10795
rect 5549 10761 5583 10795
rect 12909 10761 12943 10795
rect 16405 10761 16439 10795
rect 19165 10761 19199 10795
rect 20637 10761 20671 10795
rect 3617 10693 3651 10727
rect 4353 10693 4387 10727
rect 5365 10693 5399 10727
rect 7481 10693 7515 10727
rect 10149 10693 10183 10727
rect 14390 10693 14424 10727
rect 19502 10693 19536 10727
rect 21005 10693 21039 10727
rect 1952 10625 1986 10659
rect 4629 10625 4663 10659
rect 7665 10625 7699 10659
rect 8125 10625 8159 10659
rect 8493 10625 8527 10659
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 9873 10625 9907 10659
rect 10609 10625 10643 10659
rect 10793 10625 10827 10659
rect 10977 10625 11011 10659
rect 11161 10625 11195 10659
rect 11785 10625 11819 10659
rect 14657 10625 14691 10659
rect 15025 10625 15059 10659
rect 15292 10625 15326 10659
rect 18357 10625 18391 10659
rect 18613 10625 18647 10659
rect 18889 10625 18923 10659
rect 18981 10625 19015 10659
rect 1685 10557 1719 10591
rect 3893 10557 3927 10591
rect 4537 10557 4571 10591
rect 5641 10557 5675 10591
rect 10425 10557 10459 10591
rect 11529 10557 11563 10591
rect 19257 10557 19291 10591
rect 20913 10557 20947 10591
rect 21005 10557 21039 10591
rect 3341 10489 3375 10523
rect 5089 10489 5123 10523
rect 13277 10489 13311 10523
rect 18705 10489 18739 10523
rect 21465 10489 21499 10523
rect 3065 10421 3099 10455
rect 4629 10421 4663 10455
rect 4813 10421 4847 10455
rect 7389 10421 7423 10455
rect 7757 10421 7791 10455
rect 11069 10421 11103 10455
rect 17233 10421 17267 10455
rect 2053 10217 2087 10251
rect 6561 10217 6595 10251
rect 8125 10217 8159 10251
rect 10885 10217 10919 10251
rect 13001 10217 13035 10251
rect 15393 10217 15427 10251
rect 15761 10217 15795 10251
rect 16957 10217 16991 10251
rect 18521 10217 18555 10251
rect 2421 10149 2455 10183
rect 3525 10149 3559 10183
rect 6377 10149 6411 10183
rect 8033 10149 8067 10183
rect 8217 10149 8251 10183
rect 11529 10149 11563 10183
rect 6653 10081 6687 10115
rect 10241 10081 10275 10115
rect 11989 10081 12023 10115
rect 12909 10081 12943 10115
rect 17141 10081 17175 10115
rect 2237 10013 2271 10047
rect 3249 10013 3283 10047
rect 3985 10013 4019 10047
rect 4261 10013 4295 10047
rect 5825 10013 5859 10047
rect 6009 10013 6043 10047
rect 6101 10013 6135 10047
rect 6245 10013 6279 10047
rect 6561 10013 6595 10047
rect 6837 10013 6871 10047
rect 7941 10013 7975 10047
rect 8309 10013 8343 10047
rect 8953 10013 8987 10047
rect 9321 10013 9355 10047
rect 9965 10013 9999 10047
rect 10057 10013 10091 10047
rect 10701 10013 10735 10047
rect 12081 10013 12115 10047
rect 13093 10013 13127 10047
rect 14289 10013 14323 10047
rect 14473 10013 14507 10047
rect 15577 10013 15611 10047
rect 19809 10013 19843 10047
rect 20065 10013 20099 10047
rect 21557 10013 21591 10047
rect 2697 9945 2731 9979
rect 2973 9945 3007 9979
rect 4506 9945 4540 9979
rect 12817 9945 12851 9979
rect 14657 9945 14691 9979
rect 16037 9945 16071 9979
rect 16681 9945 16715 9979
rect 17408 9945 17442 9979
rect 2881 9877 2915 9911
rect 4169 9877 4203 9911
rect 5641 9877 5675 9911
rect 7021 9877 7055 9911
rect 7665 9877 7699 9911
rect 11989 9877 12023 9911
rect 13277 9877 13311 9911
rect 21189 9877 21223 9911
rect 21373 9877 21407 9911
rect 6009 9673 6043 9707
rect 8309 9673 8343 9707
rect 8953 9673 8987 9707
rect 17417 9673 17451 9707
rect 17969 9673 18003 9707
rect 21373 9673 21407 9707
rect 2605 9605 2639 9639
rect 2789 9605 2823 9639
rect 5089 9605 5123 9639
rect 5273 9605 5307 9639
rect 5825 9605 5859 9639
rect 10057 9605 10091 9639
rect 13185 9605 13219 9639
rect 13277 9605 13311 9639
rect 14381 9605 14415 9639
rect 14473 9605 14507 9639
rect 16313 9605 16347 9639
rect 19717 9605 19751 9639
rect 20177 9605 20211 9639
rect 21465 9605 21499 9639
rect 2145 9537 2179 9571
rect 3341 9537 3375 9571
rect 3801 9537 3835 9571
rect 3985 9537 4019 9571
rect 4077 9537 4111 9571
rect 4221 9537 4255 9571
rect 5963 9537 5997 9571
rect 6193 9537 6227 9571
rect 6469 9537 6503 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 7196 9537 7230 9571
rect 8769 9537 8803 9571
rect 9045 9537 9079 9571
rect 9413 9537 9447 9571
rect 9873 9537 9907 9571
rect 12541 9537 12575 9571
rect 13553 9537 13587 9571
rect 16129 9537 16163 9571
rect 17601 9537 17635 9571
rect 18981 9537 19015 9571
rect 20361 9537 20395 9571
rect 2881 9469 2915 9503
rect 3617 9469 3651 9503
rect 5365 9469 5399 9503
rect 6837 9469 6871 9503
rect 9597 9469 9631 9503
rect 13185 9469 13219 9503
rect 14381 9469 14415 9503
rect 16405 9469 16439 9503
rect 17877 9469 17911 9503
rect 18061 9469 18095 9503
rect 20085 9469 20119 9503
rect 21373 9469 21407 9503
rect 2329 9401 2363 9435
rect 4353 9401 4387 9435
rect 4813 9401 4847 9435
rect 5641 9401 5675 9435
rect 8585 9401 8619 9435
rect 12725 9401 12759 9435
rect 13921 9401 13955 9435
rect 18429 9401 18463 9435
rect 20637 9401 20671 9435
rect 20913 9401 20947 9435
rect 1961 9333 1995 9367
rect 9229 9333 9263 9367
rect 9781 9333 9815 9367
rect 12357 9333 12391 9367
rect 13737 9333 13771 9367
rect 15853 9333 15887 9367
rect 7389 9129 7423 9163
rect 17049 9129 17083 9163
rect 18613 9129 18647 9163
rect 7573 9061 7607 9095
rect 8309 9061 8343 9095
rect 10977 9061 11011 9095
rect 13277 9061 13311 9095
rect 10517 8993 10551 9027
rect 11897 8993 11931 9027
rect 14105 8993 14139 9027
rect 17233 8993 17267 9027
rect 20177 8993 20211 9027
rect 1685 8925 1719 8959
rect 1952 8925 1986 8959
rect 3433 8925 3467 8959
rect 4905 8925 4939 8959
rect 5325 8925 5359 8959
rect 6009 8925 6043 8959
rect 7757 8925 7791 8959
rect 7895 8925 7929 8959
rect 8493 8925 8527 8959
rect 8769 8925 8803 8959
rect 10793 8925 10827 8959
rect 13645 8925 13679 8959
rect 14361 8925 14395 8959
rect 15669 8925 15703 8959
rect 18981 8925 19015 8959
rect 19331 8925 19365 8959
rect 19901 8925 19935 8959
rect 3801 8857 3835 8891
rect 4629 8857 4663 8891
rect 5089 8857 5123 8891
rect 5181 8857 5215 8891
rect 6254 8857 6288 8891
rect 8125 8857 8159 8891
rect 8677 8857 8711 8891
rect 10250 8857 10284 8891
rect 11253 8857 11287 8891
rect 11529 8857 11563 8891
rect 12164 8857 12198 8891
rect 15936 8857 15970 8891
rect 17478 8857 17512 8891
rect 19625 8857 19659 8891
rect 20444 8857 20478 8891
rect 3065 8789 3099 8823
rect 3617 8789 3651 8823
rect 5474 8789 5508 8823
rect 7941 8789 7975 8823
rect 9137 8789 9171 8823
rect 10609 8789 10643 8823
rect 11437 8789 11471 8823
rect 13461 8789 13495 8823
rect 15485 8789 15519 8823
rect 18797 8789 18831 8823
rect 19809 8789 19843 8823
rect 21557 8789 21591 8823
rect 5457 8585 5491 8619
rect 7297 8585 7331 8619
rect 7849 8585 7883 8619
rect 7941 8585 7975 8619
rect 14289 8585 14323 8619
rect 18061 8585 18095 8619
rect 21373 8585 21407 8619
rect 6929 8517 6963 8551
rect 7389 8517 7423 8551
rect 7573 8517 7607 8551
rect 8462 8517 8496 8551
rect 12633 8517 12667 8551
rect 13176 8517 13210 8551
rect 15209 8517 15243 8551
rect 15853 8517 15887 8551
rect 15945 8517 15979 8551
rect 17233 8517 17267 8551
rect 18153 8517 18187 8551
rect 20260 8517 20294 8551
rect 1777 8449 1811 8483
rect 2053 8449 2087 8483
rect 2309 8449 2343 8483
rect 4077 8449 4111 8483
rect 4333 8449 4367 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 5917 8449 5951 8483
rect 7113 8449 7147 8483
rect 7757 8449 7791 8483
rect 8125 8449 8159 8483
rect 9873 8449 9907 8483
rect 10140 8449 10174 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 12909 8449 12943 8483
rect 14473 8449 14507 8483
rect 18337 8449 18371 8483
rect 18604 8449 18638 8483
rect 19993 8449 20027 8483
rect 8217 8381 8251 8415
rect 12633 8381 12667 8415
rect 12725 8381 12759 8415
rect 15945 8381 15979 8415
rect 17141 8381 17175 8415
rect 17325 8381 17359 8415
rect 18061 8381 18095 8415
rect 1961 8313 1995 8347
rect 11253 8313 11287 8347
rect 12173 8313 12207 8347
rect 16405 8313 16439 8347
rect 3433 8245 3467 8279
rect 5641 8245 5675 8279
rect 6101 8245 6135 8279
rect 9597 8245 9631 8279
rect 11529 8245 11563 8279
rect 11989 8245 12023 8279
rect 16773 8245 16807 8279
rect 17601 8245 17635 8279
rect 19717 8245 19751 8279
rect 4353 8041 4387 8075
rect 7297 8041 7331 8075
rect 10149 8041 10183 8075
rect 13369 8041 13403 8075
rect 15117 8041 15151 8075
rect 16957 8041 16991 8075
rect 20637 8041 20671 8075
rect 4629 7973 4663 8007
rect 15393 7973 15427 8007
rect 16497 7973 16531 8007
rect 20913 7973 20947 8007
rect 5181 7905 5215 7939
rect 9781 7905 9815 7939
rect 10241 7905 10275 7939
rect 11989 7905 12023 7939
rect 18337 7905 18371 7939
rect 19257 7905 19291 7939
rect 21373 7905 21407 7939
rect 1869 7837 1903 7871
rect 3801 7837 3835 7871
rect 4077 7837 4111 7871
rect 4174 7837 4208 7871
rect 5917 7837 5951 7871
rect 7757 7837 7791 7871
rect 7849 7837 7883 7871
rect 8309 7837 8343 7871
rect 9965 7837 9999 7871
rect 10508 7837 10542 7871
rect 12245 7837 12279 7871
rect 14841 7837 14875 7871
rect 15669 7837 15703 7871
rect 18613 7837 18647 7871
rect 18889 7837 18923 7871
rect 21465 7837 21499 7871
rect 2136 7769 2170 7803
rect 3985 7769 4019 7803
rect 4905 7769 4939 7803
rect 5089 7769 5123 7803
rect 6184 7769 6218 7803
rect 8125 7769 8159 7803
rect 8493 7769 8527 7803
rect 8953 7769 8987 7803
rect 14565 7769 14599 7803
rect 15853 7769 15887 7803
rect 15945 7769 15979 7803
rect 16221 7769 16255 7803
rect 18092 7769 18126 7803
rect 19524 7769 19558 7803
rect 21373 7769 21407 7803
rect 3249 7701 3283 7735
rect 7573 7701 7607 7735
rect 11621 7701 11655 7735
rect 14657 7701 14691 7735
rect 18429 7701 18463 7735
rect 18705 7701 18739 7735
rect 2237 7497 2271 7531
rect 6561 7497 6595 7531
rect 6745 7497 6779 7531
rect 6837 7497 6871 7531
rect 7757 7497 7791 7531
rect 8493 7497 8527 7531
rect 9597 7497 9631 7531
rect 15945 7497 15979 7531
rect 16129 7497 16163 7531
rect 16865 7497 16899 7531
rect 17049 7497 17083 7531
rect 19901 7497 19935 7531
rect 21005 7497 21039 7531
rect 3525 7429 3559 7463
rect 3985 7429 4019 7463
rect 6653 7429 6687 7463
rect 7021 7429 7055 7463
rect 7849 7429 7883 7463
rect 8953 7429 8987 7463
rect 9505 7429 9539 7463
rect 9781 7429 9815 7463
rect 11897 7429 11931 7463
rect 12081 7429 12115 7463
rect 12909 7429 12943 7463
rect 14810 7429 14844 7463
rect 18184 7429 18218 7463
rect 19073 7429 19107 7463
rect 19165 7429 19199 7463
rect 20545 7429 20579 7463
rect 20729 7429 20763 7463
rect 20821 7429 20855 7463
rect 2421 7361 2455 7395
rect 2789 7361 2823 7395
rect 3801 7361 3835 7395
rect 4077 7361 4111 7395
rect 4174 7361 4208 7395
rect 4905 7361 4939 7395
rect 5181 7361 5215 7395
rect 7573 7361 7607 7395
rect 8309 7361 8343 7395
rect 8447 7361 8481 7395
rect 8677 7361 8711 7395
rect 9137 7361 9171 7395
rect 12725 7361 12759 7395
rect 14013 7361 14047 7395
rect 14289 7361 14323 7395
rect 14565 7361 14599 7395
rect 16313 7361 16347 7395
rect 16681 7361 16715 7395
rect 18889 7361 18923 7395
rect 19717 7361 19751 7395
rect 21189 7361 21223 7395
rect 4997 7293 5031 7327
rect 7389 7293 7423 7327
rect 9321 7293 9355 7327
rect 12173 7293 12207 7327
rect 13001 7293 13035 7327
rect 18429 7293 18463 7327
rect 19993 7293 20027 7327
rect 4353 7225 4387 7259
rect 5365 7225 5399 7259
rect 8125 7225 8159 7259
rect 10057 7225 10091 7259
rect 11621 7225 11655 7259
rect 14473 7225 14507 7259
rect 19441 7225 19475 7259
rect 4997 7157 5031 7191
rect 12449 7157 12483 7191
rect 14197 7157 14231 7191
rect 18613 7157 18647 7191
rect 20269 7157 20303 7191
rect 1869 6953 1903 6987
rect 5181 6953 5215 6987
rect 7389 6953 7423 6987
rect 17969 6953 18003 6987
rect 20729 6953 20763 6987
rect 2697 6885 2731 6919
rect 3249 6817 3283 6851
rect 4353 6817 4387 6851
rect 7205 6817 7239 6851
rect 8769 6817 8803 6851
rect 10057 6817 10091 6851
rect 13001 6817 13035 6851
rect 17509 6817 17543 6851
rect 21557 6817 21591 6851
rect 2145 6749 2179 6783
rect 2421 6749 2455 6783
rect 3617 6749 3651 6783
rect 3875 6749 3909 6783
rect 4445 6749 4479 6783
rect 4629 6749 4663 6783
rect 5049 6749 5083 6783
rect 5365 6749 5399 6783
rect 6561 6749 6595 6783
rect 7021 6749 7055 6783
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 9505 6749 9539 6783
rect 9689 6749 9723 6783
rect 9873 6749 9907 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 12357 6749 12391 6783
rect 14565 6749 14599 6783
rect 14832 6749 14866 6783
rect 16405 6749 16439 6783
rect 16773 6749 16807 6783
rect 17417 6749 17451 6783
rect 18153 6749 18187 6783
rect 19349 6749 19383 6783
rect 2973 6681 3007 6715
rect 3157 6681 3191 6715
rect 4813 6681 4847 6715
rect 4905 6681 4939 6715
rect 5549 6681 5583 6715
rect 5917 6681 5951 6715
rect 6837 6681 6871 6715
rect 8502 6681 8536 6715
rect 10517 6681 10551 6715
rect 13001 6681 13035 6715
rect 13093 6681 13127 6715
rect 18981 6681 19015 6715
rect 19594 6681 19628 6715
rect 20987 6681 21021 6715
rect 21281 6681 21315 6715
rect 2329 6613 2363 6647
rect 3433 6613 3467 6647
rect 4353 6613 4387 6647
rect 5641 6613 5675 6647
rect 5733 6613 5767 6647
rect 6009 6613 6043 6647
rect 9045 6613 9079 6647
rect 12173 6613 12207 6647
rect 12523 6613 12557 6647
rect 15945 6613 15979 6647
rect 17509 6613 17543 6647
rect 21465 6613 21499 6647
rect 2237 6409 2271 6443
rect 4169 6409 4203 6443
rect 6101 6409 6135 6443
rect 7757 6409 7791 6443
rect 9413 6409 9447 6443
rect 10057 6409 10091 6443
rect 13185 6409 13219 6443
rect 19349 6409 19383 6443
rect 19441 6409 19475 6443
rect 2053 6341 2087 6375
rect 8300 6341 8334 6375
rect 10517 6341 10551 6375
rect 10609 6341 10643 6375
rect 12072 6341 12106 6375
rect 13461 6341 13495 6375
rect 15117 6341 15151 6375
rect 19962 6341 19996 6375
rect 2513 6273 2547 6307
rect 2789 6273 2823 6307
rect 3056 6273 3090 6307
rect 4721 6273 4755 6307
rect 4988 6273 5022 6307
rect 6377 6273 6411 6307
rect 6633 6273 6667 6307
rect 8033 6273 8067 6307
rect 9597 6273 9631 6307
rect 9873 6273 9907 6307
rect 10793 6273 10827 6307
rect 11529 6273 11563 6307
rect 11805 6273 11839 6307
rect 15577 6273 15611 6307
rect 17049 6273 17083 6307
rect 17325 6273 17359 6307
rect 17581 6273 17615 6307
rect 18889 6273 18923 6307
rect 19165 6273 19199 6307
rect 19625 6273 19659 6307
rect 2329 6205 2363 6239
rect 9781 6205 9815 6239
rect 14197 6205 14231 6239
rect 15117 6205 15151 6239
rect 15209 6205 15243 6239
rect 19717 6205 19751 6239
rect 1777 6137 1811 6171
rect 21097 6137 21131 6171
rect 2697 6069 2731 6103
rect 9781 6069 9815 6103
rect 11069 6069 11103 6103
rect 11713 6069 11747 6103
rect 14657 6069 14691 6103
rect 15393 6069 15427 6103
rect 17233 6069 17267 6103
rect 18705 6069 18739 6103
rect 19073 6069 19107 6103
rect 1593 5865 1627 5899
rect 4997 5865 5031 5899
rect 5181 5865 5215 5899
rect 5365 5865 5399 5899
rect 6285 5865 6319 5899
rect 7941 5865 7975 5899
rect 13277 5865 13311 5899
rect 15485 5865 15519 5899
rect 15761 5865 15795 5899
rect 19349 5865 19383 5899
rect 4537 5797 4571 5831
rect 7665 5797 7699 5831
rect 8309 5797 8343 5831
rect 11437 5797 11471 5831
rect 17141 5797 17175 5831
rect 18613 5797 18647 5831
rect 20177 5797 20211 5831
rect 21557 5797 21591 5831
rect 4813 5729 4847 5763
rect 5808 5729 5842 5763
rect 6009 5729 6043 5763
rect 9045 5729 9079 5763
rect 10057 5729 10091 5763
rect 16313 5729 16347 5763
rect 19809 5729 19843 5763
rect 20729 5729 20763 5763
rect 2706 5661 2740 5695
rect 2973 5661 3007 5695
rect 3985 5661 4019 5695
rect 4358 5661 4392 5695
rect 4721 5661 4755 5695
rect 4997 5661 5031 5695
rect 6101 5661 6135 5695
rect 6469 5661 6503 5695
rect 7481 5661 7515 5695
rect 8125 5661 8159 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 11805 5661 11839 5695
rect 11897 5661 11931 5695
rect 12164 5661 12198 5695
rect 13737 5661 13771 5695
rect 14105 5661 14139 5695
rect 16957 5661 16991 5695
rect 17233 5661 17267 5695
rect 20453 5661 20487 5695
rect 4169 5593 4203 5627
rect 4261 5593 4295 5627
rect 5549 5593 5583 5627
rect 6745 5593 6779 5627
rect 7205 5593 7239 5627
rect 9873 5593 9907 5627
rect 10302 5593 10336 5627
rect 14350 5593 14384 5627
rect 16037 5593 16071 5627
rect 16221 5593 16255 5627
rect 17478 5593 17512 5627
rect 19809 5593 19843 5627
rect 19901 5593 19935 5627
rect 21005 5593 21039 5627
rect 21281 5593 21315 5627
rect 5917 5525 5951 5559
rect 6653 5525 6687 5559
rect 7297 5525 7331 5559
rect 11621 5525 11655 5559
rect 13921 5525 13955 5559
rect 20637 5525 20671 5559
rect 21097 5525 21131 5559
rect 3341 5321 3375 5355
rect 9781 5321 9815 5355
rect 11253 5321 11287 5355
rect 12081 5321 12115 5355
rect 19717 5321 19751 5355
rect 21189 5321 21223 5355
rect 4353 5253 4387 5287
rect 6929 5253 6963 5287
rect 8493 5253 8527 5287
rect 8861 5253 8895 5287
rect 10140 5253 10174 5287
rect 12909 5253 12943 5287
rect 13093 5253 13127 5287
rect 13921 5253 13955 5287
rect 14013 5253 14047 5287
rect 14464 5253 14498 5287
rect 18613 5253 18647 5287
rect 18797 5253 18831 5287
rect 18889 5253 18923 5287
rect 20054 5253 20088 5287
rect 1685 5185 1719 5219
rect 1961 5185 1995 5219
rect 2217 5185 2251 5219
rect 3985 5185 4019 5219
rect 4078 5185 4112 5219
rect 4261 5185 4295 5219
rect 4491 5185 4525 5219
rect 5825 5185 5859 5219
rect 7849 5185 7883 5219
rect 8033 5185 8067 5219
rect 8125 5185 8159 5219
rect 8251 5185 8285 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 9005 5185 9039 5219
rect 9597 5185 9631 5219
rect 9873 5185 9907 5219
rect 11897 5185 11931 5219
rect 12173 5185 12207 5219
rect 13737 5185 13771 5219
rect 16313 5185 16347 5219
rect 16681 5185 16715 5219
rect 16937 5185 16971 5219
rect 19533 5185 19567 5219
rect 21557 5185 21591 5219
rect 6837 5117 6871 5151
rect 7021 5117 7055 5151
rect 13185 5117 13219 5151
rect 14197 5117 14231 5151
rect 19809 5117 19843 5151
rect 1869 5049 1903 5083
rect 4629 5049 4663 5083
rect 6469 5049 6503 5083
rect 9137 5049 9171 5083
rect 11621 5049 11655 5083
rect 13461 5049 13495 5083
rect 16497 5049 16531 5083
rect 18337 5049 18371 5083
rect 5641 4981 5675 5015
rect 12633 4981 12667 5015
rect 15577 4981 15611 5015
rect 18061 4981 18095 5015
rect 21373 4981 21407 5015
rect 3893 4777 3927 4811
rect 4721 4777 4755 4811
rect 6745 4777 6779 4811
rect 7665 4777 7699 4811
rect 13461 4777 13495 4811
rect 21557 4777 21591 4811
rect 8125 4709 8159 4743
rect 8585 4641 8619 4675
rect 1869 4573 1903 4607
rect 2145 4573 2179 4607
rect 4169 4573 4203 4607
rect 4900 4573 4934 4607
rect 5089 4573 5123 4607
rect 5273 4573 5307 4607
rect 5365 4573 5399 4607
rect 5632 4573 5666 4607
rect 7113 4573 7147 4607
rect 7533 4573 7567 4607
rect 8953 4573 8987 4607
rect 11529 4573 11563 4607
rect 11805 4573 11839 4607
rect 12081 4573 12115 4607
rect 16313 4573 16347 4607
rect 16589 4573 16623 4607
rect 20177 4573 20211 4607
rect 20444 4573 20478 4607
rect 2390 4505 2424 4539
rect 4445 4505 4479 4539
rect 4997 4505 5031 4539
rect 7297 4505 7331 4539
rect 7389 4505 7423 4539
rect 8677 4505 8711 4539
rect 9198 4505 9232 4539
rect 12326 4505 12360 4539
rect 16834 4505 16868 4539
rect 2053 4437 2087 4471
rect 3525 4437 3559 4471
rect 4353 4437 4387 4471
rect 8585 4437 8619 4471
rect 10333 4437 10367 4471
rect 11713 4437 11747 4471
rect 11989 4437 12023 4471
rect 16497 4437 16531 4471
rect 17969 4437 18003 4471
rect 4537 4233 4571 4267
rect 8401 4233 8435 4267
rect 13461 4233 13495 4267
rect 17693 4233 17727 4267
rect 2237 4165 2271 4199
rect 3065 4165 3099 4199
rect 5365 4165 5399 4199
rect 6929 4165 6963 4199
rect 7389 4165 7423 4199
rect 11161 4165 11195 4199
rect 12326 4165 12360 4199
rect 14749 4165 14783 4199
rect 14841 4165 14875 4199
rect 18521 4165 18555 4199
rect 20085 4165 20119 4199
rect 1409 4097 1443 4131
rect 2881 4097 2915 4131
rect 4353 4097 4387 4131
rect 5181 4097 5215 4131
rect 6745 4097 6779 4131
rect 7021 4097 7055 4131
rect 7205 4097 7239 4131
rect 7481 4097 7515 4131
rect 7578 4097 7612 4131
rect 7941 4097 7975 4131
rect 8217 4097 8251 4131
rect 8493 4097 8527 4131
rect 8677 4097 8711 4131
rect 8769 4097 8803 4131
rect 8913 4097 8947 4131
rect 10517 4097 10551 4131
rect 11253 4097 11287 4131
rect 14105 4097 14139 4131
rect 15292 4097 15326 4131
rect 17509 4097 17543 4131
rect 18981 4097 19015 4131
rect 19257 4097 19291 4131
rect 19607 4097 19641 4131
rect 20177 4097 20211 4131
rect 2237 4029 2271 4063
rect 2329 4029 2363 4063
rect 3157 4029 3191 4063
rect 4629 4029 4663 4063
rect 5457 4029 5491 4063
rect 11069 4029 11103 4063
rect 12081 4029 12115 4063
rect 14271 4029 14305 4063
rect 14749 4029 14783 4063
rect 15025 4029 15059 4063
rect 17785 4029 17819 4063
rect 18521 4029 18555 4063
rect 18613 4029 18647 4063
rect 19993 4029 20027 4063
rect 1777 3961 1811 3995
rect 7757 3961 7791 3995
rect 9045 3961 9079 3995
rect 10701 3961 10735 3995
rect 17233 3961 17267 3995
rect 19441 3961 19475 3995
rect 1593 3893 1627 3927
rect 2605 3893 2639 3927
rect 4077 3893 4111 3927
rect 4905 3893 4939 3927
rect 6469 3893 6503 3927
rect 8125 3893 8159 3927
rect 10333 3893 10367 3927
rect 13921 3893 13955 3927
rect 16405 3893 16439 3927
rect 18061 3893 18095 3927
rect 19165 3893 19199 3927
rect 5181 3689 5215 3723
rect 6837 3689 6871 3723
rect 9045 3689 9079 3723
rect 15485 3689 15519 3723
rect 20637 3689 20671 3723
rect 20913 3689 20947 3723
rect 8125 3621 8159 3655
rect 12081 3621 12115 3655
rect 13461 3621 13495 3655
rect 17877 3621 17911 3655
rect 18705 3621 18739 3655
rect 3801 3553 3835 3587
rect 5457 3553 5491 3587
rect 9597 3553 9631 3587
rect 9873 3553 9907 3587
rect 12541 3553 12575 3587
rect 14105 3553 14139 3587
rect 17417 3553 17451 3587
rect 18153 3553 18187 3587
rect 21373 3553 21407 3587
rect 1593 3485 1627 3519
rect 3157 3485 3191 3519
rect 3433 3485 3467 3519
rect 7389 3485 7423 3519
rect 8677 3485 8711 3519
rect 9321 3485 9355 3519
rect 10140 3485 10174 3519
rect 11621 3485 11655 3519
rect 11897 3485 11931 3519
rect 13737 3485 13771 3519
rect 15669 3485 15703 3519
rect 18429 3485 18463 3519
rect 19073 3485 19107 3519
rect 19257 3485 19291 3519
rect 21465 3485 21499 3519
rect 1860 3417 1894 3451
rect 4046 3417 4080 3451
rect 5724 3417 5758 3451
rect 7095 3417 7129 3451
rect 7573 3417 7607 3451
rect 7665 3417 7699 3451
rect 8401 3417 8435 3451
rect 9505 3417 9539 3451
rect 12633 3417 12667 3451
rect 12909 3417 12943 3451
rect 13185 3417 13219 3451
rect 14350 3417 14384 3451
rect 15914 3417 15948 3451
rect 17325 3417 17359 3451
rect 19524 3417 19558 3451
rect 2973 3349 3007 3383
rect 3341 3349 3375 3383
rect 3617 3349 3651 3383
rect 8585 3349 8619 3383
rect 11253 3349 11287 3383
rect 11437 3349 11471 3383
rect 11713 3349 11747 3383
rect 12541 3349 12575 3383
rect 13001 3349 13035 3383
rect 13921 3349 13955 3383
rect 17049 3349 17083 3383
rect 17417 3349 17451 3383
rect 18245 3349 18279 3383
rect 18889 3349 18923 3383
rect 21373 3349 21407 3383
rect 2973 3145 3007 3179
rect 5089 3145 5123 3179
rect 5733 3145 5767 3179
rect 7757 3145 7791 3179
rect 9413 3145 9447 3179
rect 11161 3145 11195 3179
rect 13185 3145 13219 3179
rect 15577 3145 15611 3179
rect 16221 3145 16255 3179
rect 17325 3145 17359 3179
rect 20361 3145 20395 3179
rect 1838 3077 1872 3111
rect 3954 3077 3988 3111
rect 8300 3077 8334 3111
rect 10048 3077 10082 3111
rect 11888 3077 11922 3111
rect 14074 3077 14108 3111
rect 16037 3077 16071 3111
rect 18460 3077 18494 3111
rect 19226 3077 19260 3111
rect 1593 3009 1627 3043
rect 3709 3009 3743 3043
rect 5917 3009 5951 3043
rect 6009 3009 6043 3043
rect 6377 3009 6411 3043
rect 6633 3009 6667 3043
rect 8033 3009 8067 3043
rect 9781 3009 9815 3043
rect 13369 3009 13403 3043
rect 13829 3009 13863 3043
rect 15393 3009 15427 3043
rect 16313 3009 16347 3043
rect 16957 3009 16991 3043
rect 11621 2941 11655 2975
rect 18705 2941 18739 2975
rect 18981 2941 19015 2975
rect 6193 2873 6227 2907
rect 13001 2873 13035 2907
rect 15761 2873 15795 2907
rect 15209 2805 15243 2839
rect 17141 2805 17175 2839
rect 1961 2601 1995 2635
rect 4353 2601 4387 2635
rect 8677 2601 8711 2635
rect 10977 2601 11011 2635
rect 12909 2601 12943 2635
rect 14565 2601 14599 2635
rect 15393 2601 15427 2635
rect 2421 2533 2455 2567
rect 2789 2465 2823 2499
rect 2973 2465 3007 2499
rect 7297 2465 7331 2499
rect 10425 2465 10459 2499
rect 11529 2465 11563 2499
rect 15025 2465 15059 2499
rect 2145 2397 2179 2431
rect 3801 2397 3835 2431
rect 3985 2397 4019 2431
rect 4077 2397 4111 2431
rect 4221 2397 4255 2431
rect 7021 2397 7055 2431
rect 10701 2397 10735 2431
rect 11796 2397 11830 2431
rect 15117 2397 15151 2431
rect 15577 2397 15611 2431
rect 17233 2397 17267 2431
rect 2881 2329 2915 2363
rect 7542 2329 7576 2363
rect 15025 2329 15059 2363
rect 17478 2329 17512 2363
rect 7205 2261 7239 2295
rect 10517 2261 10551 2295
rect 18613 2261 18647 2295
<< metal1 >>
rect 1104 22874 21988 22896
rect 1104 22822 4220 22874
rect 4272 22822 4284 22874
rect 4336 22822 4348 22874
rect 4400 22822 4412 22874
rect 4464 22822 4476 22874
rect 4528 22822 9441 22874
rect 9493 22822 9505 22874
rect 9557 22822 9569 22874
rect 9621 22822 9633 22874
rect 9685 22822 9697 22874
rect 9749 22822 14662 22874
rect 14714 22822 14726 22874
rect 14778 22822 14790 22874
rect 14842 22822 14854 22874
rect 14906 22822 14918 22874
rect 14970 22822 19883 22874
rect 19935 22822 19947 22874
rect 19999 22822 20011 22874
rect 20063 22822 20075 22874
rect 20127 22822 20139 22874
rect 20191 22822 21988 22874
rect 1104 22800 21988 22822
rect 7009 22763 7067 22769
rect 7009 22729 7021 22763
rect 7055 22760 7067 22763
rect 7098 22760 7104 22772
rect 7055 22732 7104 22760
rect 7055 22729 7067 22732
rect 7009 22723 7067 22729
rect 7098 22720 7104 22732
rect 7156 22720 7162 22772
rect 7374 22720 7380 22772
rect 7432 22760 7438 22772
rect 8205 22763 8263 22769
rect 8205 22760 8217 22763
rect 7432 22732 8217 22760
rect 7432 22720 7438 22732
rect 8205 22729 8217 22732
rect 8251 22760 8263 22763
rect 9030 22760 9036 22772
rect 8251 22732 9036 22760
rect 8251 22729 8263 22732
rect 8205 22723 8263 22729
rect 9030 22720 9036 22732
rect 9088 22720 9094 22772
rect 16127 22732 18082 22760
rect 2777 22695 2835 22701
rect 2777 22661 2789 22695
rect 2823 22692 2835 22695
rect 3050 22692 3056 22704
rect 2823 22664 3056 22692
rect 2823 22661 2835 22664
rect 2777 22655 2835 22661
rect 3050 22652 3056 22664
rect 3108 22652 3114 22704
rect 8570 22652 8576 22704
rect 8628 22692 8634 22704
rect 9493 22695 9551 22701
rect 9493 22692 9505 22695
rect 8628 22664 9505 22692
rect 8628 22652 8634 22664
rect 9493 22661 9505 22664
rect 9539 22661 9551 22695
rect 9493 22655 9551 22661
rect 5537 22627 5595 22633
rect 5537 22593 5549 22627
rect 5583 22624 5595 22627
rect 5583 22596 6592 22624
rect 5583 22593 5595 22596
rect 5537 22587 5595 22593
rect 2685 22559 2743 22565
rect 2685 22525 2697 22559
rect 2731 22556 2743 22559
rect 2774 22556 2780 22568
rect 2731 22528 2780 22556
rect 2731 22525 2743 22528
rect 2685 22519 2743 22525
rect 2774 22516 2780 22528
rect 2832 22516 2838 22568
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22525 2927 22559
rect 2869 22519 2927 22525
rect 2038 22380 2044 22432
rect 2096 22420 2102 22432
rect 2317 22423 2375 22429
rect 2317 22420 2329 22423
rect 2096 22392 2329 22420
rect 2096 22380 2102 22392
rect 2317 22389 2329 22392
rect 2363 22389 2375 22423
rect 2317 22383 2375 22389
rect 2774 22380 2780 22432
rect 2832 22420 2838 22432
rect 2884 22420 2912 22519
rect 4798 22516 4804 22568
rect 4856 22516 4862 22568
rect 6564 22497 6592 22596
rect 6914 22584 6920 22636
rect 6972 22624 6978 22636
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 6972 22596 7113 22624
rect 6972 22584 6978 22596
rect 7101 22593 7113 22596
rect 7147 22624 7159 22627
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 7147 22596 8125 22624
rect 7147 22593 7159 22596
rect 7101 22587 7159 22593
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 8386 22584 8392 22636
rect 8444 22584 8450 22636
rect 9214 22584 9220 22636
rect 9272 22624 9278 22636
rect 9309 22627 9367 22633
rect 9309 22624 9321 22627
rect 9272 22596 9321 22624
rect 9272 22584 9278 22596
rect 9309 22593 9321 22596
rect 9355 22593 9367 22627
rect 9309 22587 9367 22593
rect 11606 22584 11612 22636
rect 11664 22624 11670 22636
rect 11793 22627 11851 22633
rect 11793 22624 11805 22627
rect 11664 22596 11805 22624
rect 11664 22584 11670 22596
rect 11793 22593 11805 22596
rect 11839 22593 11851 22627
rect 11793 22587 11851 22593
rect 13173 22627 13231 22633
rect 13173 22593 13185 22627
rect 13219 22624 13231 22627
rect 13814 22624 13820 22636
rect 13219 22596 13820 22624
rect 13219 22593 13231 22596
rect 13173 22587 13231 22593
rect 13814 22584 13820 22596
rect 13872 22584 13878 22636
rect 16127 22633 16155 22732
rect 16209 22695 16267 22701
rect 16209 22661 16221 22695
rect 16255 22692 16267 22695
rect 17862 22692 17868 22704
rect 16255 22664 17868 22692
rect 16255 22661 16267 22664
rect 16209 22655 16267 22661
rect 17862 22652 17868 22664
rect 17920 22652 17926 22704
rect 16112 22627 16170 22633
rect 16112 22593 16124 22627
rect 16158 22593 16170 22627
rect 16112 22587 16170 22593
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22624 16359 22627
rect 16390 22624 16396 22636
rect 16347 22596 16396 22624
rect 16347 22593 16359 22596
rect 16301 22587 16359 22593
rect 16390 22584 16396 22596
rect 16448 22584 16454 22636
rect 16485 22627 16543 22633
rect 16485 22593 16497 22627
rect 16531 22624 16543 22627
rect 17405 22627 17463 22633
rect 17405 22624 17417 22627
rect 16531 22596 17417 22624
rect 16531 22593 16543 22596
rect 16485 22587 16543 22593
rect 17405 22593 17417 22596
rect 17451 22593 17463 22627
rect 18054 22624 18082 22732
rect 18785 22695 18843 22701
rect 18785 22661 18797 22695
rect 18831 22692 18843 22695
rect 19334 22692 19340 22704
rect 18831 22664 19340 22692
rect 18831 22661 18843 22664
rect 18785 22655 18843 22661
rect 19334 22652 19340 22664
rect 19392 22692 19398 22704
rect 19610 22692 19616 22704
rect 19392 22664 19616 22692
rect 19392 22652 19398 22664
rect 19610 22652 19616 22664
rect 19668 22652 19674 22704
rect 20993 22695 21051 22701
rect 20993 22692 21005 22695
rect 19996 22664 21005 22692
rect 18690 22633 18696 22636
rect 18641 22627 18696 22633
rect 18641 22624 18653 22627
rect 18054 22596 18653 22624
rect 17405 22587 17463 22593
rect 18641 22593 18653 22596
rect 18687 22593 18696 22627
rect 18641 22587 18696 22593
rect 18690 22584 18696 22587
rect 18748 22584 18754 22636
rect 18877 22627 18935 22633
rect 18877 22593 18889 22627
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 19061 22627 19119 22633
rect 19061 22593 19073 22627
rect 19107 22624 19119 22627
rect 19245 22627 19303 22633
rect 19245 22624 19257 22627
rect 19107 22596 19257 22624
rect 19107 22593 19119 22596
rect 19061 22587 19119 22593
rect 19245 22593 19257 22596
rect 19291 22593 19303 22627
rect 19996 22624 20024 22664
rect 20993 22661 21005 22664
rect 21039 22692 21051 22695
rect 21358 22692 21364 22704
rect 21039 22664 21364 22692
rect 21039 22661 21051 22664
rect 20993 22655 21051 22661
rect 21358 22652 21364 22664
rect 21416 22652 21422 22704
rect 19245 22587 19303 22593
rect 19352 22596 20024 22624
rect 20717 22627 20775 22633
rect 7006 22516 7012 22568
rect 7064 22516 7070 22568
rect 9582 22516 9588 22568
rect 9640 22516 9646 22568
rect 16022 22516 16028 22568
rect 16080 22556 16086 22568
rect 16669 22559 16727 22565
rect 16669 22556 16681 22559
rect 16080 22528 16681 22556
rect 16080 22516 16086 22528
rect 16669 22525 16681 22528
rect 16715 22525 16727 22559
rect 16669 22519 16727 22525
rect 16850 22516 16856 22568
rect 16908 22556 16914 22568
rect 17957 22559 18015 22565
rect 17957 22556 17969 22559
rect 16908 22528 17969 22556
rect 16908 22516 16914 22528
rect 17957 22525 17969 22528
rect 18003 22525 18015 22559
rect 18892 22556 18920 22587
rect 19352 22556 19380 22596
rect 20717 22593 20729 22627
rect 20763 22624 20775 22627
rect 20809 22627 20867 22633
rect 20809 22624 20821 22627
rect 20763 22596 20821 22624
rect 20763 22593 20775 22596
rect 20717 22587 20775 22593
rect 20809 22593 20821 22596
rect 20855 22593 20867 22627
rect 20809 22587 20867 22593
rect 21082 22584 21088 22636
rect 21140 22584 21146 22636
rect 21182 22627 21240 22633
rect 21182 22593 21194 22627
rect 21228 22593 21240 22627
rect 21182 22587 21240 22593
rect 17957 22519 18015 22525
rect 18708 22528 19380 22556
rect 6549 22491 6607 22497
rect 6549 22457 6561 22491
rect 6595 22457 6607 22491
rect 6549 22451 6607 22457
rect 16390 22448 16396 22500
rect 16448 22488 16454 22500
rect 18708 22488 18736 22528
rect 19702 22516 19708 22568
rect 19760 22556 19766 22568
rect 19797 22559 19855 22565
rect 19797 22556 19809 22559
rect 19760 22528 19809 22556
rect 19760 22516 19766 22528
rect 19797 22525 19809 22528
rect 19843 22525 19855 22559
rect 19797 22519 19855 22525
rect 20165 22559 20223 22565
rect 20165 22525 20177 22559
rect 20211 22556 20223 22559
rect 20530 22556 20536 22568
rect 20211 22528 20536 22556
rect 20211 22525 20223 22528
rect 20165 22519 20223 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 20990 22516 20996 22568
rect 21048 22556 21054 22568
rect 21192 22556 21220 22587
rect 21048 22528 21220 22556
rect 21048 22516 21054 22528
rect 16448 22460 18736 22488
rect 16448 22448 16454 22460
rect 18782 22448 18788 22500
rect 18840 22488 18846 22500
rect 21008 22488 21036 22516
rect 18840 22460 21036 22488
rect 18840 22448 18846 22460
rect 2832 22392 2912 22420
rect 2832 22380 2838 22392
rect 5442 22380 5448 22432
rect 5500 22380 5506 22432
rect 5721 22423 5779 22429
rect 5721 22389 5733 22423
rect 5767 22420 5779 22423
rect 5810 22420 5816 22432
rect 5767 22392 5816 22420
rect 5767 22389 5779 22392
rect 5721 22383 5779 22389
rect 5810 22380 5816 22392
rect 5868 22380 5874 22432
rect 8662 22380 8668 22432
rect 8720 22380 8726 22432
rect 9033 22423 9091 22429
rect 9033 22389 9045 22423
rect 9079 22420 9091 22423
rect 9122 22420 9128 22432
rect 9079 22392 9128 22420
rect 9079 22389 9091 22392
rect 9033 22383 9091 22389
rect 9122 22380 9128 22392
rect 9180 22380 9186 22432
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 11609 22423 11667 22429
rect 11609 22420 11621 22423
rect 11112 22392 11621 22420
rect 11112 22380 11118 22392
rect 11609 22389 11621 22392
rect 11655 22389 11667 22423
rect 11609 22383 11667 22389
rect 12986 22380 12992 22432
rect 13044 22380 13050 22432
rect 15933 22423 15991 22429
rect 15933 22389 15945 22423
rect 15979 22420 15991 22423
rect 16666 22420 16672 22432
rect 15979 22392 16672 22420
rect 15979 22389 15991 22392
rect 15933 22383 15991 22389
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 17310 22380 17316 22432
rect 17368 22380 17374 22432
rect 18506 22380 18512 22432
rect 18564 22380 18570 22432
rect 20622 22380 20628 22432
rect 20680 22420 20686 22432
rect 21361 22423 21419 22429
rect 21361 22420 21373 22423
rect 20680 22392 21373 22420
rect 20680 22380 20686 22392
rect 21361 22389 21373 22392
rect 21407 22389 21419 22423
rect 21361 22383 21419 22389
rect 1104 22330 21988 22352
rect 1104 22278 3560 22330
rect 3612 22278 3624 22330
rect 3676 22278 3688 22330
rect 3740 22278 3752 22330
rect 3804 22278 3816 22330
rect 3868 22278 8781 22330
rect 8833 22278 8845 22330
rect 8897 22278 8909 22330
rect 8961 22278 8973 22330
rect 9025 22278 9037 22330
rect 9089 22278 14002 22330
rect 14054 22278 14066 22330
rect 14118 22278 14130 22330
rect 14182 22278 14194 22330
rect 14246 22278 14258 22330
rect 14310 22278 19223 22330
rect 19275 22278 19287 22330
rect 19339 22278 19351 22330
rect 19403 22278 19415 22330
rect 19467 22278 19479 22330
rect 19531 22278 21988 22330
rect 1104 22256 21988 22278
rect 4172 22188 6914 22216
rect 3970 22040 3976 22092
rect 4028 22080 4034 22092
rect 4172 22080 4200 22188
rect 6886 22148 6914 22188
rect 7098 22176 7104 22228
rect 7156 22176 7162 22228
rect 9582 22216 9588 22228
rect 7300 22188 9588 22216
rect 7300 22148 7328 22188
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 13814 22176 13820 22228
rect 13872 22216 13878 22228
rect 14185 22219 14243 22225
rect 14185 22216 14197 22219
rect 13872 22188 14197 22216
rect 13872 22176 13878 22188
rect 14185 22185 14197 22188
rect 14231 22185 14243 22219
rect 14185 22179 14243 22185
rect 6886 22120 7328 22148
rect 7374 22108 7380 22160
rect 7432 22108 7438 22160
rect 8938 22108 8944 22160
rect 8996 22148 9002 22160
rect 9214 22148 9220 22160
rect 8996 22120 9220 22148
rect 8996 22108 9002 22120
rect 9214 22108 9220 22120
rect 9272 22108 9278 22160
rect 17773 22151 17831 22157
rect 10888 22120 11284 22148
rect 4028 22052 4200 22080
rect 5353 22083 5411 22089
rect 4028 22040 4034 22052
rect 5353 22049 5365 22083
rect 5399 22080 5411 22083
rect 5721 22083 5779 22089
rect 5721 22080 5733 22083
rect 5399 22052 5733 22080
rect 5399 22049 5411 22052
rect 5353 22043 5411 22049
rect 5721 22049 5733 22052
rect 5767 22049 5779 22083
rect 9306 22080 9312 22092
rect 5721 22043 5779 22049
rect 8772 22052 9312 22080
rect 2038 21972 2044 22024
rect 2096 21972 2102 22024
rect 2133 22015 2191 22021
rect 2133 21981 2145 22015
rect 2179 22012 2191 22015
rect 2774 22012 2780 22024
rect 2179 21984 2780 22012
rect 2179 21981 2191 21984
rect 2133 21975 2191 21981
rect 2774 21972 2780 21984
rect 2832 21972 2838 22024
rect 4062 21972 4068 22024
rect 4120 22012 4126 22024
rect 5368 22012 5396 22043
rect 4120 21984 5396 22012
rect 4120 21972 4126 21984
rect 5626 21972 5632 22024
rect 5684 21972 5690 22024
rect 5810 21972 5816 22024
rect 5868 22012 5874 22024
rect 8772 22021 8800 22052
rect 9306 22040 9312 22052
rect 9364 22040 9370 22092
rect 10888 22024 10916 22120
rect 11256 22080 11284 22120
rect 17773 22117 17785 22151
rect 17819 22117 17831 22151
rect 17773 22111 17831 22117
rect 11256 22052 12296 22080
rect 5977 22015 6035 22021
rect 5977 22012 5989 22015
rect 5868 21984 5989 22012
rect 5868 21972 5874 21984
rect 5977 21981 5989 21984
rect 6023 21981 6035 22015
rect 8757 22015 8815 22021
rect 8757 22012 8769 22015
rect 5977 21975 6035 21981
rect 8312 21984 8769 22012
rect 8312 21956 8340 21984
rect 8757 21981 8769 21984
rect 8803 21981 8815 22015
rect 8757 21975 8815 21981
rect 8846 21972 8852 22024
rect 8904 22012 8910 22024
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 8904 21984 9137 22012
rect 8904 21972 8910 21984
rect 9125 21981 9137 21984
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 10870 21972 10876 22024
rect 10928 22012 10934 22024
rect 11097 22015 11155 22021
rect 11097 22012 11109 22015
rect 10928 21984 11109 22012
rect 10928 21972 10934 21984
rect 11097 21981 11109 21984
rect 11143 21981 11155 22015
rect 11097 21975 11155 21981
rect 11517 22015 11575 22021
rect 11517 21981 11529 22015
rect 11563 22012 11575 22015
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 11563 21984 11621 22012
rect 11563 21981 11575 21984
rect 11517 21975 11575 21981
rect 11609 21981 11621 21984
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 2400 21947 2458 21953
rect 2400 21913 2412 21947
rect 2446 21944 2458 21947
rect 2958 21944 2964 21956
rect 2446 21916 2964 21944
rect 2446 21913 2458 21916
rect 2400 21907 2458 21913
rect 2958 21904 2964 21916
rect 3016 21904 3022 21956
rect 5108 21947 5166 21953
rect 5108 21913 5120 21947
rect 5154 21944 5166 21947
rect 5154 21916 5488 21944
rect 5154 21913 5166 21916
rect 5108 21907 5166 21913
rect 1670 21836 1676 21888
rect 1728 21876 1734 21888
rect 1857 21879 1915 21885
rect 1857 21876 1869 21879
rect 1728 21848 1869 21876
rect 1728 21836 1734 21848
rect 1857 21845 1869 21848
rect 1903 21845 1915 21879
rect 1857 21839 1915 21845
rect 3513 21879 3571 21885
rect 3513 21845 3525 21879
rect 3559 21876 3571 21879
rect 3878 21876 3884 21888
rect 3559 21848 3884 21876
rect 3559 21845 3571 21848
rect 3513 21839 3571 21845
rect 3878 21836 3884 21848
rect 3936 21836 3942 21888
rect 3973 21879 4031 21885
rect 3973 21845 3985 21879
rect 4019 21876 4031 21879
rect 4614 21876 4620 21888
rect 4019 21848 4620 21876
rect 4019 21845 4031 21848
rect 3973 21839 4031 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 5460 21885 5488 21916
rect 8294 21904 8300 21956
rect 8352 21904 8358 21956
rect 8512 21947 8570 21953
rect 8512 21913 8524 21947
rect 8558 21944 8570 21947
rect 8558 21916 8800 21944
rect 8558 21913 8570 21916
rect 8512 21907 8570 21913
rect 5445 21879 5503 21885
rect 5445 21845 5457 21879
rect 5491 21845 5503 21879
rect 8772 21876 8800 21916
rect 9214 21904 9220 21956
rect 9272 21944 9278 21956
rect 9554 21947 9612 21953
rect 9554 21944 9566 21947
rect 9272 21916 9566 21944
rect 9272 21904 9278 21916
rect 9554 21913 9566 21916
rect 9600 21913 9612 21947
rect 9554 21907 9612 21913
rect 10704 21916 11100 21944
rect 8941 21879 8999 21885
rect 8941 21876 8953 21879
rect 8772 21848 8953 21876
rect 5445 21839 5503 21845
rect 8941 21845 8953 21848
rect 8987 21845 8999 21879
rect 8941 21839 8999 21845
rect 10042 21836 10048 21888
rect 10100 21876 10106 21888
rect 10704 21885 10732 21916
rect 10689 21879 10747 21885
rect 10689 21876 10701 21879
rect 10100 21848 10701 21876
rect 10100 21836 10106 21848
rect 10689 21845 10701 21848
rect 10735 21845 10747 21879
rect 10689 21839 10747 21845
rect 10778 21836 10784 21888
rect 10836 21876 10842 21888
rect 10948 21879 11006 21885
rect 10948 21876 10960 21879
rect 10836 21848 10960 21876
rect 10836 21836 10842 21848
rect 10948 21845 10960 21848
rect 10994 21845 11006 21879
rect 11072 21876 11100 21916
rect 11238 21904 11244 21956
rect 11296 21904 11302 21956
rect 11330 21904 11336 21956
rect 11388 21904 11394 21956
rect 12176 21876 12204 21975
rect 12268 21944 12296 22052
rect 15102 22040 15108 22092
rect 15160 22080 15166 22092
rect 16393 22083 16451 22089
rect 16393 22080 16405 22083
rect 15160 22052 16405 22080
rect 15160 22040 15166 22052
rect 16393 22049 16405 22052
rect 16439 22049 16451 22083
rect 17788 22080 17816 22111
rect 18046 22080 18052 22092
rect 17788 22052 18052 22080
rect 16393 22043 16451 22049
rect 18046 22040 18052 22052
rect 18104 22040 18110 22092
rect 18509 22083 18567 22089
rect 18509 22049 18521 22083
rect 18555 22080 18567 22083
rect 19702 22080 19708 22092
rect 18555 22052 19708 22080
rect 18555 22049 18567 22052
rect 18509 22043 18567 22049
rect 19702 22040 19708 22052
rect 19760 22040 19766 22092
rect 12434 21972 12440 22024
rect 12492 21972 12498 22024
rect 12704 22015 12762 22021
rect 12704 21981 12716 22015
rect 12750 22012 12762 22015
rect 12986 22012 12992 22024
rect 12750 21984 12992 22012
rect 12750 21981 12762 21984
rect 12704 21975 12762 21981
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 14737 22015 14795 22021
rect 14737 22012 14749 22015
rect 13648 21984 14749 22012
rect 13262 21944 13268 21956
rect 12268 21916 13268 21944
rect 13262 21904 13268 21916
rect 13320 21904 13326 21956
rect 11072 21848 12204 21876
rect 10948 21839 11006 21845
rect 12342 21836 12348 21888
rect 12400 21876 12406 21888
rect 13648 21876 13676 21984
rect 14737 21981 14749 21984
rect 14783 21981 14795 22015
rect 14737 21975 14795 21981
rect 15930 21972 15936 22024
rect 15988 21972 15994 22024
rect 16666 22021 16672 22024
rect 16660 21975 16672 22021
rect 16666 21972 16672 21975
rect 16724 21972 16730 22024
rect 19794 21972 19800 22024
rect 19852 21972 19858 22024
rect 14461 21947 14519 21953
rect 14461 21913 14473 21947
rect 14507 21944 14519 21947
rect 14550 21944 14556 21956
rect 14507 21916 14556 21944
rect 14507 21913 14519 21916
rect 14461 21907 14519 21913
rect 14550 21904 14556 21916
rect 14608 21904 14614 21956
rect 15286 21904 15292 21956
rect 15344 21904 15350 21956
rect 15562 21904 15568 21956
rect 15620 21904 15626 21956
rect 17954 21904 17960 21956
rect 18012 21944 18018 21956
rect 18509 21947 18567 21953
rect 18509 21944 18521 21947
rect 18012 21916 18521 21944
rect 18012 21904 18018 21916
rect 18509 21913 18521 21916
rect 18555 21913 18567 21947
rect 18509 21907 18567 21913
rect 18601 21947 18659 21953
rect 18601 21913 18613 21947
rect 18647 21944 18659 21947
rect 18966 21944 18972 21956
rect 18647 21916 18972 21944
rect 18647 21913 18659 21916
rect 18601 21907 18659 21913
rect 18966 21904 18972 21916
rect 19024 21904 19030 21956
rect 20064 21947 20122 21953
rect 20064 21913 20076 21947
rect 20110 21944 20122 21947
rect 20346 21944 20352 21956
rect 20110 21916 20352 21944
rect 20110 21913 20122 21916
rect 20064 21907 20122 21913
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 13722 21876 13728 21888
rect 12400 21848 13728 21876
rect 12400 21836 12406 21848
rect 13722 21836 13728 21848
rect 13780 21836 13786 21888
rect 13817 21879 13875 21885
rect 13817 21845 13829 21879
rect 13863 21876 13875 21879
rect 13906 21876 13912 21888
rect 13863 21848 13912 21876
rect 13863 21845 13875 21848
rect 13817 21839 13875 21845
rect 13906 21836 13912 21848
rect 13964 21876 13970 21888
rect 15010 21885 15016 21888
rect 14645 21879 14703 21885
rect 14645 21876 14657 21879
rect 13964 21848 14657 21876
rect 13964 21836 13970 21848
rect 14645 21845 14657 21848
rect 14691 21845 14703 21879
rect 14645 21839 14703 21845
rect 15003 21879 15016 21885
rect 15003 21845 15015 21879
rect 15003 21839 15016 21845
rect 15010 21836 15016 21839
rect 15068 21836 15074 21888
rect 15378 21836 15384 21888
rect 15436 21876 15442 21888
rect 15473 21879 15531 21885
rect 15473 21876 15485 21879
rect 15436 21848 15485 21876
rect 15436 21836 15442 21848
rect 15473 21845 15485 21848
rect 15519 21845 15531 21879
rect 15473 21839 15531 21845
rect 15746 21836 15752 21888
rect 15804 21836 15810 21888
rect 18046 21885 18052 21888
rect 18039 21879 18052 21885
rect 18039 21845 18051 21879
rect 18039 21839 18052 21845
rect 18046 21836 18052 21839
rect 18104 21836 18110 21888
rect 21082 21836 21088 21888
rect 21140 21876 21146 21888
rect 21177 21879 21235 21885
rect 21177 21876 21189 21879
rect 21140 21848 21189 21876
rect 21140 21836 21146 21848
rect 21177 21845 21189 21848
rect 21223 21845 21235 21879
rect 21177 21839 21235 21845
rect 1104 21786 21988 21808
rect 1104 21734 4220 21786
rect 4272 21734 4284 21786
rect 4336 21734 4348 21786
rect 4400 21734 4412 21786
rect 4464 21734 4476 21786
rect 4528 21734 9441 21786
rect 9493 21734 9505 21786
rect 9557 21734 9569 21786
rect 9621 21734 9633 21786
rect 9685 21734 9697 21786
rect 9749 21734 14662 21786
rect 14714 21734 14726 21786
rect 14778 21734 14790 21786
rect 14842 21734 14854 21786
rect 14906 21734 14918 21786
rect 14970 21734 19883 21786
rect 19935 21734 19947 21786
rect 19999 21734 20011 21786
rect 20063 21734 20075 21786
rect 20127 21734 20139 21786
rect 20191 21734 21988 21786
rect 1104 21712 21988 21734
rect 2958 21632 2964 21684
rect 3016 21632 3022 21684
rect 3973 21675 4031 21681
rect 3973 21641 3985 21675
rect 4019 21672 4031 21675
rect 5258 21672 5264 21684
rect 4019 21644 5264 21672
rect 4019 21641 4031 21644
rect 3973 21635 4031 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 5718 21632 5724 21684
rect 5776 21632 5782 21684
rect 5994 21632 6000 21684
rect 6052 21672 6058 21684
rect 6052 21644 8524 21672
rect 6052 21632 6058 21644
rect 2774 21604 2780 21616
rect 1412 21576 2780 21604
rect 1412 21545 1440 21576
rect 2774 21564 2780 21576
rect 2832 21604 2838 21616
rect 2832 21576 3648 21604
rect 2832 21564 2838 21576
rect 1670 21545 1676 21548
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21505 1455 21539
rect 1664 21536 1676 21545
rect 1631 21508 1676 21536
rect 1397 21499 1455 21505
rect 1664 21499 1676 21508
rect 1670 21496 1676 21499
rect 1728 21496 1734 21548
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21536 3203 21539
rect 3620 21536 3648 21576
rect 4062 21564 4068 21616
rect 4120 21564 4126 21616
rect 4798 21564 4804 21616
rect 4856 21604 4862 21616
rect 5350 21604 5356 21616
rect 4856 21576 5356 21604
rect 4856 21564 4862 21576
rect 5350 21564 5356 21576
rect 5408 21564 5414 21616
rect 5534 21564 5540 21616
rect 5592 21604 5598 21616
rect 6457 21607 6515 21613
rect 6457 21604 6469 21607
rect 5592 21576 6469 21604
rect 5592 21564 5598 21576
rect 6457 21573 6469 21576
rect 6503 21573 6515 21607
rect 6457 21567 6515 21573
rect 6638 21564 6644 21616
rect 6696 21604 6702 21616
rect 7377 21607 7435 21613
rect 7377 21604 7389 21607
rect 6696 21576 7389 21604
rect 6696 21564 6702 21576
rect 7377 21573 7389 21576
rect 7423 21573 7435 21607
rect 7377 21567 7435 21573
rect 7561 21607 7619 21613
rect 7561 21573 7573 21607
rect 7607 21604 7619 21607
rect 8386 21604 8392 21616
rect 7607 21576 8392 21604
rect 7607 21573 7619 21576
rect 7561 21567 7619 21573
rect 8386 21564 8392 21576
rect 8444 21564 8450 21616
rect 8496 21604 8524 21644
rect 8938 21632 8944 21684
rect 8996 21672 9002 21684
rect 9398 21672 9404 21684
rect 8996 21644 9404 21672
rect 8996 21632 9002 21644
rect 9398 21632 9404 21644
rect 9456 21672 9462 21684
rect 9585 21675 9643 21681
rect 9585 21672 9597 21675
rect 9456 21644 9597 21672
rect 9456 21632 9462 21644
rect 9585 21641 9597 21644
rect 9631 21641 9643 21675
rect 9585 21635 9643 21641
rect 10962 21632 10968 21684
rect 11020 21672 11026 21684
rect 11238 21672 11244 21684
rect 11020 21644 11244 21672
rect 11020 21632 11026 21644
rect 11238 21632 11244 21644
rect 11296 21632 11302 21684
rect 12069 21675 12127 21681
rect 12069 21641 12081 21675
rect 12115 21672 12127 21675
rect 12250 21672 12256 21684
rect 12115 21644 12256 21672
rect 12115 21641 12127 21644
rect 12069 21635 12127 21641
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 13078 21632 13084 21684
rect 13136 21672 13142 21684
rect 13136 21644 15700 21672
rect 13136 21632 13142 21644
rect 10128 21607 10186 21613
rect 8496 21576 9996 21604
rect 4080 21536 4108 21564
rect 4341 21539 4399 21545
rect 4341 21536 4353 21539
rect 3191 21508 3556 21536
rect 3620 21508 4353 21536
rect 3191 21505 3203 21508
rect 3145 21499 3203 21505
rect 2777 21403 2835 21409
rect 2777 21369 2789 21403
rect 2823 21400 2835 21403
rect 3050 21400 3056 21412
rect 2823 21372 3056 21400
rect 2823 21369 2835 21372
rect 2777 21363 2835 21369
rect 3050 21360 3056 21372
rect 3108 21360 3114 21412
rect 3528 21409 3556 21508
rect 4341 21505 4353 21508
rect 4387 21505 4399 21539
rect 4341 21499 4399 21505
rect 4608 21539 4666 21545
rect 4608 21505 4620 21539
rect 4654 21536 4666 21539
rect 5810 21536 5816 21548
rect 4654 21508 5816 21536
rect 4654 21505 4666 21508
rect 4608 21499 4666 21505
rect 5810 21496 5816 21508
rect 5868 21496 5874 21548
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 3878 21428 3884 21480
rect 3936 21428 3942 21480
rect 3970 21428 3976 21480
rect 4028 21468 4034 21480
rect 4065 21471 4123 21477
rect 4065 21468 4077 21471
rect 4028 21440 4077 21468
rect 4028 21428 4034 21440
rect 4065 21437 4077 21440
rect 4111 21437 4123 21471
rect 6012 21468 6040 21499
rect 6546 21496 6552 21548
rect 6604 21536 6610 21548
rect 8205 21539 8263 21545
rect 6604 21508 7512 21536
rect 6604 21496 6610 21508
rect 7374 21468 7380 21480
rect 6012 21440 7380 21468
rect 4065 21431 4123 21437
rect 7374 21428 7380 21440
rect 7432 21428 7438 21480
rect 3513 21403 3571 21409
rect 3513 21369 3525 21403
rect 3559 21369 3571 21403
rect 3513 21363 3571 21369
rect 5350 21360 5356 21412
rect 5408 21400 5414 21412
rect 6822 21400 6828 21412
rect 5408 21372 6828 21400
rect 5408 21360 5414 21372
rect 6822 21360 6828 21372
rect 6880 21360 6886 21412
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 7101 21403 7159 21409
rect 7101 21400 7113 21403
rect 7064 21372 7113 21400
rect 7064 21360 7070 21372
rect 7101 21369 7113 21372
rect 7147 21369 7159 21403
rect 7484 21400 7512 21508
rect 8205 21505 8217 21539
rect 8251 21536 8263 21539
rect 8294 21536 8300 21548
rect 8251 21508 8300 21536
rect 8251 21505 8263 21508
rect 8205 21499 8263 21505
rect 8294 21496 8300 21508
rect 8352 21496 8358 21548
rect 8478 21545 8484 21548
rect 8472 21499 8484 21545
rect 8478 21496 8484 21499
rect 8536 21496 8542 21548
rect 9306 21496 9312 21548
rect 9364 21536 9370 21548
rect 9861 21539 9919 21545
rect 9861 21536 9873 21539
rect 9364 21508 9873 21536
rect 9364 21496 9370 21508
rect 9861 21505 9873 21508
rect 9907 21505 9919 21539
rect 9968 21536 9996 21576
rect 10128 21573 10140 21607
rect 10174 21604 10186 21607
rect 10778 21604 10784 21616
rect 10174 21576 10784 21604
rect 10174 21573 10186 21576
rect 10128 21567 10186 21573
rect 10778 21564 10784 21576
rect 10836 21564 10842 21616
rect 11146 21564 11152 21616
rect 11204 21604 11210 21616
rect 12161 21607 12219 21613
rect 12161 21604 12173 21607
rect 11204 21576 12173 21604
rect 11204 21564 11210 21576
rect 12161 21573 12173 21576
rect 12207 21604 12219 21607
rect 12342 21604 12348 21616
rect 12207 21576 12348 21604
rect 12207 21573 12219 21576
rect 12161 21567 12219 21573
rect 12342 21564 12348 21576
rect 12400 21564 12406 21616
rect 12434 21564 12440 21616
rect 12492 21604 12498 21616
rect 15102 21604 15108 21616
rect 12492 21576 15108 21604
rect 12492 21564 12498 21576
rect 11330 21536 11336 21548
rect 9968 21508 11336 21536
rect 9861 21499 9919 21505
rect 11330 21496 11336 21508
rect 11388 21496 11394 21548
rect 11698 21496 11704 21548
rect 11756 21536 11762 21548
rect 11885 21539 11943 21545
rect 11885 21536 11897 21539
rect 11756 21508 11897 21536
rect 11756 21496 11762 21508
rect 11885 21505 11897 21508
rect 11931 21505 11943 21539
rect 11885 21499 11943 21505
rect 12710 21496 12716 21548
rect 12768 21496 12774 21548
rect 13004 21545 13032 21576
rect 14568 21545 14596 21576
rect 15102 21564 15108 21576
rect 15160 21564 15166 21616
rect 15672 21548 15700 21644
rect 16114 21632 16120 21684
rect 16172 21672 16178 21684
rect 16761 21675 16819 21681
rect 16761 21672 16773 21675
rect 16172 21644 16773 21672
rect 16172 21632 16178 21644
rect 16761 21641 16773 21644
rect 16807 21672 16819 21675
rect 17034 21672 17040 21684
rect 16807 21644 17040 21672
rect 16807 21641 16819 21644
rect 16761 21635 16819 21641
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 19610 21632 19616 21684
rect 19668 21632 19674 21684
rect 19794 21604 19800 21616
rect 18248 21576 19800 21604
rect 14826 21545 14832 21548
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21505 13047 21539
rect 13245 21539 13303 21545
rect 13245 21536 13257 21539
rect 12989 21499 13047 21505
rect 13096 21508 13257 21536
rect 7653 21471 7711 21477
rect 7653 21437 7665 21471
rect 7699 21468 7711 21471
rect 8110 21468 8116 21480
rect 7699 21440 8116 21468
rect 7699 21437 7711 21440
rect 7653 21431 7711 21437
rect 8110 21428 8116 21440
rect 8168 21428 8174 21480
rect 13096 21468 13124 21508
rect 13245 21505 13257 21508
rect 13291 21505 13303 21539
rect 13245 21499 13303 21505
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21505 14611 21539
rect 14553 21499 14611 21505
rect 14820 21499 14832 21545
rect 14826 21496 14832 21499
rect 14884 21496 14890 21548
rect 15654 21496 15660 21548
rect 15712 21536 15718 21548
rect 16117 21539 16175 21545
rect 16117 21536 16129 21539
rect 15712 21508 16129 21536
rect 15712 21496 15718 21508
rect 16117 21505 16129 21508
rect 16163 21505 16175 21539
rect 16117 21499 16175 21505
rect 16758 21496 16764 21548
rect 16816 21536 16822 21548
rect 18248 21545 18276 21576
rect 19794 21564 19800 21576
rect 19852 21564 19858 21616
rect 20064 21607 20122 21613
rect 20064 21573 20076 21607
rect 20110 21604 20122 21607
rect 20622 21604 20628 21616
rect 20110 21576 20628 21604
rect 20110 21573 20122 21576
rect 20064 21567 20122 21573
rect 20622 21564 20628 21576
rect 20680 21564 20686 21616
rect 18506 21545 18512 21548
rect 17874 21539 17932 21545
rect 17874 21536 17886 21539
rect 16816 21508 17886 21536
rect 16816 21496 16822 21508
rect 17874 21505 17886 21508
rect 17920 21505 17932 21539
rect 17874 21499 17932 21505
rect 18141 21539 18199 21545
rect 18141 21505 18153 21539
rect 18187 21536 18199 21539
rect 18233 21539 18291 21545
rect 18233 21536 18245 21539
rect 18187 21508 18245 21536
rect 18187 21505 18199 21508
rect 18141 21499 18199 21505
rect 18233 21505 18245 21508
rect 18279 21505 18291 21539
rect 18500 21536 18512 21545
rect 18467 21508 18512 21536
rect 18233 21499 18291 21505
rect 18500 21499 18512 21508
rect 18506 21496 18512 21499
rect 18564 21496 18570 21548
rect 12912 21440 13124 21468
rect 7484 21372 8156 21400
rect 7101 21363 7159 21369
rect 5258 21292 5264 21344
rect 5316 21332 5322 21344
rect 6086 21332 6092 21344
rect 5316 21304 6092 21332
rect 5316 21292 5322 21304
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 6181 21335 6239 21341
rect 6181 21301 6193 21335
rect 6227 21332 6239 21335
rect 6362 21332 6368 21344
rect 6227 21304 6368 21332
rect 6227 21301 6239 21304
rect 6181 21295 6239 21301
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 6733 21335 6791 21341
rect 6733 21301 6745 21335
rect 6779 21332 6791 21335
rect 6914 21332 6920 21344
rect 6779 21304 6920 21332
rect 6779 21301 6791 21304
rect 6733 21295 6791 21301
rect 6914 21292 6920 21304
rect 6972 21332 6978 21344
rect 8018 21332 8024 21344
rect 6972 21304 8024 21332
rect 6972 21292 6978 21304
rect 8018 21292 8024 21304
rect 8076 21292 8082 21344
rect 8128 21332 8156 21372
rect 11606 21360 11612 21412
rect 11664 21360 11670 21412
rect 12912 21409 12940 21440
rect 19794 21428 19800 21480
rect 19852 21428 19858 21480
rect 12897 21403 12955 21409
rect 12897 21369 12909 21403
rect 12943 21369 12955 21403
rect 12897 21363 12955 21369
rect 16301 21403 16359 21409
rect 16301 21369 16313 21403
rect 16347 21400 16359 21403
rect 16390 21400 16396 21412
rect 16347 21372 16396 21400
rect 16347 21369 16359 21372
rect 16301 21363 16359 21369
rect 16390 21360 16396 21372
rect 16448 21360 16454 21412
rect 10870 21332 10876 21344
rect 8128 21304 10876 21332
rect 10870 21292 10876 21304
rect 10928 21292 10934 21344
rect 14369 21335 14427 21341
rect 14369 21301 14381 21335
rect 14415 21332 14427 21335
rect 14458 21332 14464 21344
rect 14415 21304 14464 21332
rect 14415 21301 14427 21304
rect 14369 21295 14427 21301
rect 14458 21292 14464 21304
rect 14516 21292 14522 21344
rect 15286 21292 15292 21344
rect 15344 21332 15350 21344
rect 15933 21335 15991 21341
rect 15933 21332 15945 21335
rect 15344 21304 15945 21332
rect 15344 21292 15350 21304
rect 15933 21301 15945 21304
rect 15979 21332 15991 21335
rect 16022 21332 16028 21344
rect 15979 21304 16028 21332
rect 15979 21301 15991 21304
rect 15933 21295 15991 21301
rect 16022 21292 16028 21304
rect 16080 21292 16086 21344
rect 21174 21292 21180 21344
rect 21232 21292 21238 21344
rect 1104 21242 21988 21264
rect 1104 21190 3560 21242
rect 3612 21190 3624 21242
rect 3676 21190 3688 21242
rect 3740 21190 3752 21242
rect 3804 21190 3816 21242
rect 3868 21190 8781 21242
rect 8833 21190 8845 21242
rect 8897 21190 8909 21242
rect 8961 21190 8973 21242
rect 9025 21190 9037 21242
rect 9089 21190 14002 21242
rect 14054 21190 14066 21242
rect 14118 21190 14130 21242
rect 14182 21190 14194 21242
rect 14246 21190 14258 21242
rect 14310 21190 19223 21242
rect 19275 21190 19287 21242
rect 19339 21190 19351 21242
rect 19403 21190 19415 21242
rect 19467 21190 19479 21242
rect 19531 21190 21988 21242
rect 1104 21168 21988 21190
rect 3881 21131 3939 21137
rect 3881 21128 3893 21131
rect 2746 21100 3893 21128
rect 1946 21020 1952 21072
rect 2004 21060 2010 21072
rect 2133 21063 2191 21069
rect 2133 21060 2145 21063
rect 2004 21032 2145 21060
rect 2004 21020 2010 21032
rect 2133 21029 2145 21032
rect 2179 21029 2191 21063
rect 2746 21060 2774 21100
rect 3881 21097 3893 21100
rect 3927 21097 3939 21131
rect 3881 21091 3939 21097
rect 5261 21131 5319 21137
rect 5261 21097 5273 21131
rect 5307 21128 5319 21131
rect 5626 21128 5632 21140
rect 5307 21100 5632 21128
rect 5307 21097 5319 21100
rect 5261 21091 5319 21097
rect 5626 21088 5632 21100
rect 5684 21088 5690 21140
rect 5810 21088 5816 21140
rect 5868 21128 5874 21140
rect 5997 21131 6055 21137
rect 5997 21128 6009 21131
rect 5868 21100 6009 21128
rect 5868 21088 5874 21100
rect 5997 21097 6009 21100
rect 6043 21097 6055 21131
rect 6638 21128 6644 21140
rect 5997 21091 6055 21097
rect 6288 21100 6644 21128
rect 2133 21023 2191 21029
rect 2608 21032 2774 21060
rect 2608 21001 2636 21032
rect 2866 21020 2872 21072
rect 2924 21060 2930 21072
rect 2961 21063 3019 21069
rect 2961 21060 2973 21063
rect 2924 21032 2973 21060
rect 2924 21020 2930 21032
rect 2961 21029 2973 21032
rect 3007 21029 3019 21063
rect 5534 21060 5540 21072
rect 2961 21023 3019 21029
rect 3344 21032 5540 21060
rect 2593 20995 2651 21001
rect 2593 20961 2605 20995
rect 2639 20961 2651 20995
rect 3344 20992 3372 21032
rect 5534 21020 5540 21032
rect 5592 21020 5598 21072
rect 2593 20955 2651 20961
rect 2746 20964 3372 20992
rect 3421 20995 3479 21001
rect 2746 20868 2774 20964
rect 3421 20961 3433 20995
rect 3467 20992 3479 20995
rect 4614 20992 4620 21004
rect 3467 20964 4620 20992
rect 3467 20961 3479 20964
rect 3421 20955 3479 20961
rect 4614 20952 4620 20964
rect 4672 20992 4678 21004
rect 4801 20995 4859 21001
rect 4801 20992 4813 20995
rect 4672 20964 4813 20992
rect 4672 20952 4678 20964
rect 4801 20961 4813 20964
rect 4847 20961 4859 20995
rect 5994 20992 6000 21004
rect 4801 20955 4859 20961
rect 5644 20964 6000 20992
rect 5644 20936 5672 20964
rect 5994 20952 6000 20964
rect 6052 20952 6058 21004
rect 3878 20924 3884 20936
rect 2406 20816 2412 20868
rect 2464 20856 2470 20868
rect 2682 20856 2688 20868
rect 2464 20828 2688 20856
rect 2464 20816 2470 20828
rect 2682 20816 2688 20828
rect 2740 20828 2774 20868
rect 3436 20896 3884 20924
rect 3436 20865 3464 20896
rect 3878 20884 3884 20896
rect 3936 20884 3942 20936
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 4890 20924 4896 20936
rect 4203 20896 4896 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 4890 20884 4896 20896
rect 4948 20884 4954 20936
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 5626 20884 5632 20936
rect 5684 20884 5690 20936
rect 5718 20884 5724 20936
rect 5776 20884 5782 20936
rect 5902 20933 5908 20936
rect 5865 20927 5908 20933
rect 5865 20893 5877 20927
rect 5865 20887 5908 20893
rect 5902 20884 5908 20887
rect 5960 20884 5966 20936
rect 6181 20927 6239 20933
rect 6181 20924 6193 20927
rect 6012 20896 6193 20924
rect 3421 20859 3479 20865
rect 2740 20816 2746 20828
rect 3421 20825 3433 20859
rect 3467 20825 3479 20859
rect 3421 20819 3479 20825
rect 3513 20859 3571 20865
rect 3513 20825 3525 20859
rect 3559 20856 3571 20859
rect 4433 20859 4491 20865
rect 4433 20856 4445 20859
rect 3559 20828 4445 20856
rect 3559 20825 3571 20828
rect 3513 20819 3571 20825
rect 4433 20825 4445 20828
rect 4479 20856 4491 20859
rect 4522 20856 4528 20868
rect 4479 20828 4528 20856
rect 4479 20825 4491 20828
rect 4433 20819 4491 20825
rect 4522 20816 4528 20828
rect 4580 20816 4586 20868
rect 4709 20859 4767 20865
rect 4709 20825 4721 20859
rect 4755 20856 4767 20859
rect 4982 20856 4988 20868
rect 4755 20828 4988 20856
rect 4755 20825 4767 20828
rect 4709 20819 4767 20825
rect 4982 20816 4988 20828
rect 5040 20816 5046 20868
rect 2590 20748 2596 20800
rect 2648 20748 2654 20800
rect 4341 20791 4399 20797
rect 4341 20757 4353 20791
rect 4387 20788 4399 20791
rect 4614 20788 4620 20800
rect 4387 20760 4620 20788
rect 4387 20757 4399 20760
rect 4341 20751 4399 20757
rect 4614 20748 4620 20760
rect 4672 20748 4678 20800
rect 4801 20791 4859 20797
rect 4801 20757 4813 20791
rect 4847 20788 4859 20791
rect 6012 20788 6040 20896
rect 6181 20893 6193 20896
rect 6227 20924 6239 20927
rect 6288 20924 6316 21100
rect 6638 21088 6644 21100
rect 6696 21088 6702 21140
rect 8478 21088 8484 21140
rect 8536 21128 8542 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8536 21100 8953 21128
rect 8536 21088 8542 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 8941 21091 8999 21097
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 9401 21131 9459 21137
rect 9401 21128 9413 21131
rect 9272 21100 9413 21128
rect 9272 21088 9278 21100
rect 9401 21097 9413 21100
rect 9447 21097 9459 21131
rect 9401 21091 9459 21097
rect 11885 21131 11943 21137
rect 11885 21097 11897 21131
rect 11931 21128 11943 21131
rect 12250 21128 12256 21140
rect 11931 21100 12256 21128
rect 11931 21097 11943 21100
rect 11885 21091 11943 21097
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 12710 21088 12716 21140
rect 12768 21128 12774 21140
rect 14185 21131 14243 21137
rect 14185 21128 14197 21131
rect 12768 21100 14197 21128
rect 12768 21088 12774 21100
rect 14185 21097 14197 21100
rect 14231 21097 14243 21131
rect 14185 21091 14243 21097
rect 14826 21088 14832 21140
rect 14884 21128 14890 21140
rect 14921 21131 14979 21137
rect 14921 21128 14933 21131
rect 14884 21100 14933 21128
rect 14884 21088 14890 21100
rect 14921 21097 14933 21100
rect 14967 21097 14979 21131
rect 14921 21091 14979 21097
rect 16669 21131 16727 21137
rect 16669 21097 16681 21131
rect 16715 21128 16727 21131
rect 16850 21128 16856 21140
rect 16715 21100 16856 21128
rect 16715 21097 16727 21100
rect 16669 21091 16727 21097
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 18601 21131 18659 21137
rect 18601 21097 18613 21131
rect 18647 21128 18659 21131
rect 19610 21128 19616 21140
rect 18647 21100 19616 21128
rect 18647 21097 18659 21100
rect 18601 21091 18659 21097
rect 19610 21088 19616 21100
rect 19668 21088 19674 21140
rect 7837 21063 7895 21069
rect 7837 21029 7849 21063
rect 7883 21060 7895 21063
rect 8386 21060 8392 21072
rect 7883 21032 8392 21060
rect 7883 21029 7895 21032
rect 7837 21023 7895 21029
rect 8386 21020 8392 21032
rect 8444 21020 8450 21072
rect 12529 21063 12587 21069
rect 12529 21029 12541 21063
rect 12575 21060 12587 21063
rect 12894 21060 12900 21072
rect 12575 21032 12900 21060
rect 12575 21029 12587 21032
rect 12529 21023 12587 21029
rect 12894 21020 12900 21032
rect 12952 21020 12958 21072
rect 15102 21020 15108 21072
rect 15160 21020 15166 21072
rect 6362 20952 6368 21004
rect 6420 20992 6426 21004
rect 6420 20964 6592 20992
rect 6420 20952 6426 20964
rect 6227 20896 6316 20924
rect 6457 20927 6515 20933
rect 6227 20893 6239 20896
rect 6181 20887 6239 20893
rect 6457 20893 6469 20927
rect 6503 20893 6515 20927
rect 6564 20924 6592 20964
rect 9306 20952 9312 21004
rect 9364 20992 9370 21004
rect 10505 20995 10563 21001
rect 10505 20992 10517 20995
rect 9364 20964 10517 20992
rect 9364 20952 9370 20964
rect 10505 20961 10517 20964
rect 10551 20961 10563 20995
rect 10505 20955 10563 20961
rect 13906 20952 13912 21004
rect 13964 20992 13970 21004
rect 15120 20992 15148 21020
rect 15289 20995 15347 21001
rect 15289 20992 15301 20995
rect 13964 20964 15301 20992
rect 13964 20952 13970 20964
rect 15289 20961 15301 20964
rect 15335 20961 15347 20995
rect 15289 20955 15347 20961
rect 6713 20927 6771 20933
rect 6713 20924 6725 20927
rect 6564 20896 6725 20924
rect 6457 20887 6515 20893
rect 6713 20893 6725 20896
rect 6759 20893 6771 20927
rect 6713 20887 6771 20893
rect 6086 20816 6092 20868
rect 6144 20856 6150 20868
rect 6472 20856 6500 20887
rect 9122 20884 9128 20936
rect 9180 20884 9186 20936
rect 9585 20927 9643 20933
rect 9585 20893 9597 20927
rect 9631 20924 9643 20927
rect 9751 20927 9809 20933
rect 9751 20924 9763 20927
rect 9631 20896 9763 20924
rect 9631 20893 9643 20896
rect 9585 20887 9643 20893
rect 9751 20893 9763 20896
rect 9797 20893 9809 20927
rect 9751 20887 9809 20893
rect 10042 20884 10048 20936
rect 10100 20884 10106 20936
rect 10772 20927 10830 20933
rect 10772 20893 10784 20927
rect 10818 20924 10830 20927
rect 11054 20924 11060 20936
rect 10818 20896 11060 20924
rect 10818 20893 10830 20896
rect 10772 20887 10830 20893
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 11330 20884 11336 20936
rect 11388 20924 11394 20936
rect 13078 20924 13084 20936
rect 11388 20896 13084 20924
rect 11388 20884 11394 20896
rect 13078 20884 13084 20896
rect 13136 20884 13142 20936
rect 14458 20884 14464 20936
rect 14516 20884 14522 20936
rect 14660 20896 14872 20924
rect 6144 20828 6500 20856
rect 6144 20816 6150 20828
rect 6822 20816 6828 20868
rect 6880 20856 6886 20868
rect 8297 20859 8355 20865
rect 8297 20856 8309 20859
rect 6880 20828 8309 20856
rect 6880 20816 6886 20828
rect 8297 20825 8309 20828
rect 8343 20856 8355 20859
rect 9858 20856 9864 20868
rect 8343 20828 9864 20856
rect 8343 20825 8355 20828
rect 8297 20819 8355 20825
rect 9858 20816 9864 20828
rect 9916 20816 9922 20868
rect 10321 20859 10379 20865
rect 10321 20825 10333 20859
rect 10367 20825 10379 20859
rect 10321 20819 10379 20825
rect 4847 20760 6040 20788
rect 4847 20757 4859 20760
rect 4801 20751 4859 20757
rect 6178 20748 6184 20800
rect 6236 20788 6242 20800
rect 6365 20791 6423 20797
rect 6365 20788 6377 20791
rect 6236 20760 6377 20788
rect 6236 20748 6242 20760
rect 6365 20757 6377 20760
rect 6411 20757 6423 20791
rect 6365 20751 6423 20757
rect 8110 20748 8116 20800
rect 8168 20788 8174 20800
rect 8389 20791 8447 20797
rect 8389 20788 8401 20791
rect 8168 20760 8401 20788
rect 8168 20748 8174 20760
rect 8389 20757 8401 20760
rect 8435 20757 8447 20791
rect 8389 20751 8447 20757
rect 10226 20748 10232 20800
rect 10284 20748 10290 20800
rect 10336 20788 10364 20819
rect 13446 20816 13452 20868
rect 13504 20856 13510 20868
rect 14660 20865 14688 20896
rect 13642 20859 13700 20865
rect 13642 20856 13654 20859
rect 13504 20828 13654 20856
rect 13504 20816 13510 20828
rect 13642 20825 13654 20828
rect 13688 20825 13700 20859
rect 13642 20819 13700 20825
rect 14645 20859 14703 20865
rect 14645 20825 14657 20859
rect 14691 20825 14703 20859
rect 14645 20819 14703 20825
rect 14737 20859 14795 20865
rect 14737 20825 14749 20859
rect 14783 20825 14795 20859
rect 14844 20856 14872 20896
rect 15010 20884 15016 20936
rect 15068 20924 15074 20936
rect 15105 20927 15163 20933
rect 15105 20924 15117 20927
rect 15068 20896 15117 20924
rect 15068 20884 15074 20896
rect 15105 20893 15117 20896
rect 15151 20893 15163 20927
rect 15105 20887 15163 20893
rect 17221 20927 17279 20933
rect 17221 20893 17233 20927
rect 17267 20924 17279 20927
rect 17267 20896 18828 20924
rect 17267 20893 17279 20896
rect 17221 20887 17279 20893
rect 15378 20856 15384 20868
rect 14844 20828 15384 20856
rect 14737 20819 14795 20825
rect 10962 20788 10968 20800
rect 10336 20760 10968 20788
rect 10962 20748 10968 20760
rect 11020 20788 11026 20800
rect 13814 20788 13820 20800
rect 11020 20760 13820 20788
rect 11020 20748 11026 20760
rect 13814 20748 13820 20760
rect 13872 20748 13878 20800
rect 14752 20788 14780 20819
rect 15378 20816 15384 20828
rect 15436 20856 15442 20868
rect 15556 20859 15614 20865
rect 15436 20828 15516 20856
rect 15436 20816 15442 20828
rect 15010 20788 15016 20800
rect 14752 20760 15016 20788
rect 15010 20748 15016 20760
rect 15068 20748 15074 20800
rect 15488 20788 15516 20828
rect 15556 20825 15568 20859
rect 15602 20856 15614 20859
rect 15746 20856 15752 20868
rect 15602 20828 15752 20856
rect 15602 20825 15614 20828
rect 15556 20819 15614 20825
rect 15746 20816 15752 20828
rect 15804 20816 15810 20868
rect 17494 20865 17500 20868
rect 17488 20819 17500 20865
rect 17494 20816 17500 20819
rect 17552 20816 17558 20868
rect 18800 20856 18828 20896
rect 18874 20884 18880 20936
rect 18932 20884 18938 20936
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 19794 20924 19800 20936
rect 19291 20896 19800 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 19260 20856 19288 20887
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 21266 20884 21272 20936
rect 21324 20924 21330 20936
rect 21545 20927 21603 20933
rect 21545 20924 21557 20927
rect 21324 20896 21557 20924
rect 21324 20884 21330 20896
rect 21545 20893 21557 20896
rect 21591 20893 21603 20927
rect 21545 20887 21603 20893
rect 19490 20859 19548 20865
rect 19490 20856 19502 20859
rect 18800 20828 19288 20856
rect 19352 20828 19502 20856
rect 17862 20788 17868 20800
rect 15488 20760 17868 20788
rect 17862 20748 17868 20760
rect 17920 20748 17926 20800
rect 19061 20791 19119 20797
rect 19061 20757 19073 20791
rect 19107 20788 19119 20791
rect 19352 20788 19380 20828
rect 19490 20825 19502 20828
rect 19536 20825 19548 20859
rect 19490 20819 19548 20825
rect 19107 20760 19380 20788
rect 19107 20757 19119 20760
rect 19061 20751 19119 20757
rect 20622 20748 20628 20800
rect 20680 20748 20686 20800
rect 20993 20791 21051 20797
rect 20993 20757 21005 20791
rect 21039 20788 21051 20791
rect 21450 20788 21456 20800
rect 21039 20760 21456 20788
rect 21039 20757 21051 20760
rect 20993 20751 21051 20757
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 1104 20698 21988 20720
rect 1104 20646 4220 20698
rect 4272 20646 4284 20698
rect 4336 20646 4348 20698
rect 4400 20646 4412 20698
rect 4464 20646 4476 20698
rect 4528 20646 9441 20698
rect 9493 20646 9505 20698
rect 9557 20646 9569 20698
rect 9621 20646 9633 20698
rect 9685 20646 9697 20698
rect 9749 20646 14662 20698
rect 14714 20646 14726 20698
rect 14778 20646 14790 20698
rect 14842 20646 14854 20698
rect 14906 20646 14918 20698
rect 14970 20646 19883 20698
rect 19935 20646 19947 20698
rect 19999 20646 20011 20698
rect 20063 20646 20075 20698
rect 20127 20646 20139 20698
rect 20191 20646 21988 20698
rect 1104 20624 21988 20646
rect 4154 20584 4160 20596
rect 3528 20556 4160 20584
rect 2774 20516 2780 20528
rect 1412 20488 2780 20516
rect 1412 20457 1440 20488
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 3528 20525 3556 20556
rect 4154 20544 4160 20556
rect 4212 20584 4218 20596
rect 4614 20584 4620 20596
rect 4212 20556 4620 20584
rect 4212 20544 4218 20556
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 5166 20544 5172 20596
rect 5224 20584 5230 20596
rect 5626 20584 5632 20596
rect 5224 20556 5396 20584
rect 5224 20544 5230 20556
rect 5368 20528 5396 20556
rect 5460 20556 5632 20584
rect 3513 20519 3571 20525
rect 3513 20485 3525 20519
rect 3559 20485 3571 20519
rect 3513 20479 3571 20485
rect 3697 20519 3755 20525
rect 3697 20485 3709 20519
rect 3743 20485 3755 20519
rect 3697 20479 3755 20485
rect 3789 20519 3847 20525
rect 3789 20485 3801 20519
rect 3835 20516 3847 20519
rect 3970 20516 3976 20528
rect 3835 20488 3976 20516
rect 3835 20485 3847 20488
rect 3789 20479 3847 20485
rect 1670 20457 1676 20460
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20417 1455 20451
rect 1397 20411 1455 20417
rect 1664 20411 1676 20457
rect 1670 20408 1676 20411
rect 1728 20408 1734 20460
rect 3712 20448 3740 20479
rect 3970 20476 3976 20488
rect 4028 20476 4034 20528
rect 4706 20476 4712 20528
rect 4764 20476 4770 20528
rect 5350 20476 5356 20528
rect 5408 20476 5414 20528
rect 5460 20525 5488 20556
rect 5626 20544 5632 20556
rect 5684 20544 5690 20596
rect 5902 20544 5908 20596
rect 5960 20584 5966 20596
rect 6546 20584 6552 20596
rect 5960 20556 6552 20584
rect 5960 20544 5966 20556
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 6638 20544 6644 20596
rect 6696 20544 6702 20596
rect 8662 20544 8668 20596
rect 8720 20544 8726 20596
rect 9306 20544 9312 20596
rect 9364 20584 9370 20596
rect 9677 20587 9735 20593
rect 9677 20584 9689 20587
rect 9364 20556 9689 20584
rect 9364 20544 9370 20556
rect 9677 20553 9689 20556
rect 9723 20553 9735 20587
rect 9677 20547 9735 20553
rect 11333 20587 11391 20593
rect 11333 20553 11345 20587
rect 11379 20584 11391 20587
rect 14185 20587 14243 20593
rect 11379 20556 12940 20584
rect 11379 20553 11391 20556
rect 11333 20547 11391 20553
rect 5445 20519 5503 20525
rect 5445 20485 5457 20519
rect 5491 20485 5503 20519
rect 5445 20479 5503 20485
rect 5534 20476 5540 20528
rect 5592 20516 5598 20528
rect 5813 20519 5871 20525
rect 5813 20516 5825 20519
rect 5592 20488 5825 20516
rect 5592 20476 5598 20488
rect 5813 20485 5825 20488
rect 5859 20485 5871 20519
rect 5813 20479 5871 20485
rect 6086 20476 6092 20528
rect 6144 20516 6150 20528
rect 8294 20516 8300 20528
rect 6144 20488 8300 20516
rect 6144 20476 6150 20488
rect 4890 20448 4896 20460
rect 3712 20420 3832 20448
rect 2682 20272 2688 20324
rect 2740 20312 2746 20324
rect 2777 20315 2835 20321
rect 2777 20312 2789 20315
rect 2740 20284 2789 20312
rect 2740 20272 2746 20284
rect 2777 20281 2789 20284
rect 2823 20281 2835 20315
rect 3804 20312 3832 20420
rect 4632 20420 4896 20448
rect 4632 20392 4660 20420
rect 4890 20408 4896 20420
rect 4948 20408 4954 20460
rect 5256 20451 5314 20457
rect 5256 20417 5268 20451
rect 5302 20448 5314 20451
rect 5302 20420 5580 20448
rect 5302 20417 5314 20420
rect 5256 20411 5314 20417
rect 4614 20340 4620 20392
rect 4672 20340 4678 20392
rect 4801 20383 4859 20389
rect 4801 20349 4813 20383
rect 4847 20380 4859 20383
rect 4982 20380 4988 20392
rect 4847 20352 4988 20380
rect 4847 20349 4859 20352
rect 4801 20343 4859 20349
rect 4982 20340 4988 20352
rect 5040 20340 5046 20392
rect 5552 20380 5580 20420
rect 5626 20408 5632 20460
rect 5684 20408 5690 20460
rect 7742 20408 7748 20460
rect 7800 20457 7806 20460
rect 8036 20457 8064 20488
rect 8294 20476 8300 20488
rect 8352 20476 8358 20528
rect 8386 20476 8392 20528
rect 8444 20516 8450 20528
rect 8481 20519 8539 20525
rect 8481 20516 8493 20519
rect 8444 20488 8493 20516
rect 8444 20476 8450 20488
rect 8481 20485 8493 20488
rect 8527 20485 8539 20519
rect 8481 20479 8539 20485
rect 9493 20519 9551 20525
rect 9493 20485 9505 20519
rect 9539 20516 9551 20519
rect 10042 20516 10048 20528
rect 9539 20488 10048 20516
rect 9539 20485 9551 20488
rect 9493 20479 9551 20485
rect 10042 20476 10048 20488
rect 10100 20476 10106 20528
rect 12066 20476 12072 20528
rect 12124 20516 12130 20528
rect 12161 20519 12219 20525
rect 12161 20516 12173 20519
rect 12124 20488 12173 20516
rect 12124 20476 12130 20488
rect 12161 20485 12173 20488
rect 12207 20485 12219 20519
rect 12161 20479 12219 20485
rect 7800 20411 7812 20457
rect 8021 20451 8079 20457
rect 8021 20417 8033 20451
rect 8067 20417 8079 20451
rect 8021 20411 8079 20417
rect 7800 20408 7806 20411
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 10781 20451 10839 20457
rect 8720 20420 9904 20448
rect 8720 20408 8726 20420
rect 5902 20380 5908 20392
rect 5552 20352 5908 20380
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 8202 20340 8208 20392
rect 8260 20380 8266 20392
rect 8757 20383 8815 20389
rect 8757 20380 8769 20383
rect 8260 20352 8769 20380
rect 8260 20340 8266 20352
rect 8757 20349 8769 20352
rect 8803 20349 8815 20383
rect 8757 20343 8815 20349
rect 9769 20383 9827 20389
rect 9769 20349 9781 20383
rect 9815 20349 9827 20383
rect 9876 20380 9904 20420
rect 10781 20417 10793 20451
rect 10827 20448 10839 20451
rect 11790 20448 11796 20460
rect 10827 20420 11796 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 11790 20408 11796 20420
rect 11848 20448 11854 20460
rect 11977 20451 12035 20457
rect 11977 20448 11989 20451
rect 11848 20420 11989 20448
rect 11848 20408 11854 20420
rect 11977 20417 11989 20420
rect 12023 20417 12035 20451
rect 11977 20411 12035 20417
rect 12434 20408 12440 20460
rect 12492 20408 12498 20460
rect 12912 20457 12940 20556
rect 14185 20553 14197 20587
rect 14231 20584 14243 20587
rect 14458 20584 14464 20596
rect 14231 20556 14464 20584
rect 14231 20553 14243 20556
rect 14185 20547 14243 20553
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 16850 20584 16856 20596
rect 16132 20556 16856 20584
rect 12986 20476 12992 20528
rect 13044 20516 13050 20528
rect 13173 20519 13231 20525
rect 13173 20516 13185 20519
rect 13044 20488 13185 20516
rect 13044 20476 13050 20488
rect 13173 20485 13185 20488
rect 13219 20485 13231 20519
rect 13173 20479 13231 20485
rect 14369 20519 14427 20525
rect 14369 20485 14381 20519
rect 14415 20516 14427 20519
rect 15286 20516 15292 20528
rect 14415 20488 15292 20516
rect 14415 20485 14427 20488
rect 14369 20479 14427 20485
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 16132 20525 16160 20556
rect 16850 20544 16856 20556
rect 16908 20544 16914 20596
rect 16960 20556 17172 20584
rect 16117 20519 16175 20525
rect 16117 20485 16129 20519
rect 16163 20485 16175 20519
rect 16117 20479 16175 20485
rect 16301 20519 16359 20525
rect 16301 20485 16313 20519
rect 16347 20485 16359 20519
rect 16301 20479 16359 20485
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 13078 20408 13084 20460
rect 13136 20408 13142 20460
rect 13262 20408 13268 20460
rect 13320 20457 13326 20460
rect 13320 20448 13328 20457
rect 16022 20448 16028 20460
rect 13320 20420 13365 20448
rect 14016 20420 16028 20448
rect 13320 20411 13328 20420
rect 13320 20408 13326 20411
rect 9876 20352 11836 20380
rect 9769 20343 9827 20349
rect 6822 20312 6828 20324
rect 3804 20284 6828 20312
rect 2777 20275 2835 20281
rect 6822 20272 6828 20284
rect 6880 20272 6886 20324
rect 8570 20272 8576 20324
rect 8628 20312 8634 20324
rect 9217 20315 9275 20321
rect 9217 20312 9229 20315
rect 8628 20284 9229 20312
rect 8628 20272 8634 20284
rect 9217 20281 9229 20284
rect 9263 20281 9275 20315
rect 9217 20275 9275 20281
rect 2038 20204 2044 20256
rect 2096 20244 2102 20256
rect 3237 20247 3295 20253
rect 3237 20244 3249 20247
rect 2096 20216 3249 20244
rect 2096 20204 2102 20216
rect 3237 20213 3249 20216
rect 3283 20213 3295 20247
rect 3237 20207 3295 20213
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 4249 20247 4307 20253
rect 4249 20244 4261 20247
rect 4028 20216 4261 20244
rect 4028 20204 4034 20216
rect 4249 20213 4261 20216
rect 4295 20213 4307 20247
rect 4249 20207 4307 20213
rect 5074 20204 5080 20256
rect 5132 20204 5138 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 8205 20247 8263 20253
rect 8205 20244 8217 20247
rect 7432 20216 8217 20244
rect 7432 20204 7438 20216
rect 8205 20213 8217 20216
rect 8251 20213 8263 20247
rect 9784 20244 9812 20343
rect 11698 20272 11704 20324
rect 11756 20272 11762 20324
rect 11808 20312 11836 20352
rect 12250 20340 12256 20392
rect 12308 20340 12314 20392
rect 14016 20380 14044 20420
rect 16022 20408 16028 20420
rect 16080 20448 16086 20460
rect 16316 20448 16344 20479
rect 16390 20476 16396 20528
rect 16448 20516 16454 20528
rect 16960 20516 16988 20556
rect 16448 20488 16988 20516
rect 16448 20476 16454 20488
rect 17034 20476 17040 20528
rect 17092 20476 17098 20528
rect 17144 20525 17172 20556
rect 17494 20544 17500 20596
rect 17552 20544 17558 20596
rect 18414 20544 18420 20596
rect 18472 20584 18478 20596
rect 20530 20584 20536 20596
rect 18472 20556 20536 20584
rect 18472 20544 18478 20556
rect 20530 20544 20536 20556
rect 20588 20544 20594 20596
rect 17129 20519 17187 20525
rect 17129 20485 17141 20519
rect 17175 20516 17187 20519
rect 18322 20516 18328 20528
rect 17175 20488 18328 20516
rect 17175 20485 17187 20488
rect 17129 20479 17187 20485
rect 18322 20476 18328 20488
rect 18380 20476 18386 20528
rect 18601 20519 18659 20525
rect 18601 20485 18613 20519
rect 18647 20516 18659 20519
rect 20622 20516 20628 20528
rect 18647 20488 20628 20516
rect 18647 20485 18659 20488
rect 18601 20479 18659 20485
rect 20622 20476 20628 20488
rect 20680 20476 20686 20528
rect 16080 20420 16344 20448
rect 16940 20451 16998 20457
rect 16080 20408 16086 20420
rect 16940 20417 16952 20451
rect 16986 20417 16998 20451
rect 16940 20411 16998 20417
rect 12406 20352 14044 20380
rect 14093 20383 14151 20389
rect 12406 20312 12434 20352
rect 14093 20349 14105 20383
rect 14139 20380 14151 20383
rect 14734 20380 14740 20392
rect 14139 20352 14740 20380
rect 14139 20349 14151 20352
rect 14093 20343 14151 20349
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 16393 20383 16451 20389
rect 16393 20349 16405 20383
rect 16439 20380 16451 20383
rect 16850 20380 16856 20392
rect 16439 20352 16856 20380
rect 16439 20349 16451 20352
rect 16393 20343 16451 20349
rect 16850 20340 16856 20352
rect 16908 20340 16914 20392
rect 11808 20284 12434 20312
rect 13446 20272 13452 20324
rect 13504 20272 13510 20324
rect 14550 20272 14556 20324
rect 14608 20312 14614 20324
rect 14645 20315 14703 20321
rect 14645 20312 14657 20315
rect 14608 20284 14657 20312
rect 14608 20272 14614 20284
rect 14645 20281 14657 20284
rect 14691 20281 14703 20315
rect 14645 20275 14703 20281
rect 15841 20315 15899 20321
rect 15841 20281 15853 20315
rect 15887 20312 15899 20315
rect 15930 20312 15936 20324
rect 15887 20284 15936 20312
rect 15887 20281 15899 20284
rect 15841 20275 15899 20281
rect 15930 20272 15936 20284
rect 15988 20272 15994 20324
rect 16758 20272 16764 20324
rect 16816 20272 16822 20324
rect 16955 20312 16983 20411
rect 17310 20408 17316 20460
rect 17368 20408 17374 20460
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20448 17739 20451
rect 18046 20448 18052 20460
rect 17727 20420 18052 20448
rect 17727 20417 17739 20420
rect 17681 20411 17739 20417
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 19061 20451 19119 20457
rect 19061 20448 19073 20451
rect 18748 20420 19073 20448
rect 18748 20408 18754 20420
rect 19061 20417 19073 20420
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 20073 20451 20131 20457
rect 20073 20448 20085 20451
rect 19668 20420 20085 20448
rect 19668 20408 19674 20420
rect 20073 20417 20085 20420
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 20990 20408 20996 20460
rect 21048 20457 21054 20460
rect 21048 20451 21091 20457
rect 21079 20417 21091 20451
rect 21048 20411 21091 20417
rect 21048 20408 21054 20411
rect 21174 20408 21180 20460
rect 21232 20408 21238 20460
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 21358 20448 21364 20460
rect 21315 20420 21364 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 21450 20408 21456 20460
rect 21508 20408 21514 20460
rect 17126 20340 17132 20392
rect 17184 20380 17190 20392
rect 18325 20383 18383 20389
rect 18325 20380 18337 20383
rect 17184 20352 18337 20380
rect 17184 20340 17190 20352
rect 18325 20349 18337 20352
rect 18371 20380 18383 20383
rect 18966 20380 18972 20392
rect 18371 20352 18972 20380
rect 18371 20349 18383 20352
rect 18325 20343 18383 20349
rect 18966 20340 18972 20352
rect 19024 20340 19030 20392
rect 19794 20340 19800 20392
rect 19852 20340 19858 20392
rect 18506 20312 18512 20324
rect 16955 20284 18512 20312
rect 18506 20272 18512 20284
rect 18564 20272 18570 20324
rect 18874 20272 18880 20324
rect 18932 20272 18938 20324
rect 9858 20244 9864 20256
rect 9784 20216 9864 20244
rect 8205 20207 8263 20213
rect 9858 20204 9864 20216
rect 9916 20244 9922 20256
rect 12250 20244 12256 20256
rect 9916 20216 12256 20244
rect 9916 20204 9922 20216
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 12621 20247 12679 20253
rect 12621 20213 12633 20247
rect 12667 20244 12679 20247
rect 12802 20244 12808 20256
rect 12667 20216 12808 20244
rect 12667 20213 12679 20216
rect 12621 20207 12679 20213
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 13262 20204 13268 20256
rect 13320 20244 13326 20256
rect 17218 20244 17224 20256
rect 13320 20216 17224 20244
rect 13320 20204 13326 20216
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 20717 20247 20775 20253
rect 20717 20213 20729 20247
rect 20763 20244 20775 20247
rect 20806 20244 20812 20256
rect 20763 20216 20812 20244
rect 20763 20213 20775 20216
rect 20717 20207 20775 20213
rect 20806 20204 20812 20216
rect 20864 20204 20870 20256
rect 20898 20204 20904 20256
rect 20956 20204 20962 20256
rect 1104 20154 21988 20176
rect 1104 20102 3560 20154
rect 3612 20102 3624 20154
rect 3676 20102 3688 20154
rect 3740 20102 3752 20154
rect 3804 20102 3816 20154
rect 3868 20102 8781 20154
rect 8833 20102 8845 20154
rect 8897 20102 8909 20154
rect 8961 20102 8973 20154
rect 9025 20102 9037 20154
rect 9089 20102 14002 20154
rect 14054 20102 14066 20154
rect 14118 20102 14130 20154
rect 14182 20102 14194 20154
rect 14246 20102 14258 20154
rect 14310 20102 19223 20154
rect 19275 20102 19287 20154
rect 19339 20102 19351 20154
rect 19403 20102 19415 20154
rect 19467 20102 19479 20154
rect 19531 20102 21988 20154
rect 1104 20080 21988 20102
rect 1670 20000 1676 20052
rect 1728 20040 1734 20052
rect 1765 20043 1823 20049
rect 1765 20040 1777 20043
rect 1728 20012 1777 20040
rect 1728 20000 1734 20012
rect 1765 20009 1777 20012
rect 1811 20009 1823 20043
rect 1765 20003 1823 20009
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20040 3479 20043
rect 4154 20040 4160 20052
rect 3467 20012 4160 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 4154 20000 4160 20012
rect 4212 20000 4218 20052
rect 5626 20000 5632 20052
rect 5684 20040 5690 20052
rect 5905 20043 5963 20049
rect 5905 20040 5917 20043
rect 5684 20012 5917 20040
rect 5684 20000 5690 20012
rect 5905 20009 5917 20012
rect 5951 20009 5963 20043
rect 5905 20003 5963 20009
rect 7742 20000 7748 20052
rect 7800 20000 7806 20052
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 10594 20040 10600 20052
rect 8260 20012 10600 20040
rect 8260 20000 8266 20012
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 11701 20043 11759 20049
rect 11701 20009 11713 20043
rect 11747 20040 11759 20043
rect 11790 20040 11796 20052
rect 11747 20012 11796 20040
rect 11747 20009 11759 20012
rect 11701 20003 11759 20009
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 12434 20000 12440 20052
rect 12492 20040 12498 20052
rect 13265 20043 13323 20049
rect 13265 20040 13277 20043
rect 12492 20012 13277 20040
rect 12492 20000 12498 20012
rect 13265 20009 13277 20012
rect 13311 20009 13323 20043
rect 13265 20003 13323 20009
rect 13446 20000 13452 20052
rect 13504 20040 13510 20052
rect 18414 20040 18420 20052
rect 13504 20012 18420 20040
rect 13504 20000 13510 20012
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 18969 20043 19027 20049
rect 18969 20009 18981 20043
rect 19015 20040 19027 20043
rect 20346 20040 20352 20052
rect 19015 20012 20352 20040
rect 19015 20009 19027 20012
rect 18969 20003 19027 20009
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 21545 20043 21603 20049
rect 21545 20040 21557 20043
rect 21232 20012 21557 20040
rect 21232 20000 21238 20012
rect 21545 20009 21557 20012
rect 21591 20009 21603 20043
rect 21545 20003 21603 20009
rect 5350 19932 5356 19984
rect 5408 19972 5414 19984
rect 5721 19975 5779 19981
rect 5721 19972 5733 19975
rect 5408 19944 5733 19972
rect 5408 19932 5414 19944
rect 5721 19941 5733 19944
rect 5767 19941 5779 19975
rect 5721 19935 5779 19941
rect 8386 19932 8392 19984
rect 8444 19972 8450 19984
rect 9033 19975 9091 19981
rect 9033 19972 9045 19975
rect 8444 19944 9045 19972
rect 8444 19932 8450 19944
rect 9033 19941 9045 19944
rect 9079 19941 9091 19975
rect 9033 19935 9091 19941
rect 14185 19975 14243 19981
rect 14185 19941 14197 19975
rect 14231 19972 14243 19975
rect 14458 19972 14464 19984
rect 14231 19944 14464 19972
rect 14231 19941 14243 19944
rect 14185 19935 14243 19941
rect 14458 19932 14464 19944
rect 14516 19932 14522 19984
rect 16485 19975 16543 19981
rect 16485 19941 16497 19975
rect 16531 19941 16543 19975
rect 16485 19935 16543 19941
rect 5442 19864 5448 19916
rect 5500 19904 5506 19916
rect 6457 19907 6515 19913
rect 6457 19904 6469 19907
rect 5500 19876 6469 19904
rect 5500 19864 5506 19876
rect 6457 19873 6469 19876
rect 6503 19873 6515 19907
rect 6457 19867 6515 19873
rect 9493 19907 9551 19913
rect 9493 19873 9505 19907
rect 9539 19904 9551 19907
rect 9766 19904 9772 19916
rect 9539 19876 9772 19904
rect 9539 19873 9551 19876
rect 9493 19867 9551 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 13081 19907 13139 19913
rect 13081 19873 13093 19907
rect 13127 19904 13139 19907
rect 13906 19904 13912 19916
rect 13127 19876 13912 19904
rect 13127 19873 13139 19876
rect 13081 19867 13139 19873
rect 13906 19864 13912 19876
rect 13964 19864 13970 19916
rect 15562 19904 15568 19916
rect 14568 19876 15568 19904
rect 1946 19796 1952 19848
rect 2004 19796 2010 19848
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19836 2099 19839
rect 2774 19836 2780 19848
rect 2087 19808 2780 19836
rect 2087 19805 2099 19808
rect 2041 19799 2099 19805
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 3970 19796 3976 19848
rect 4028 19796 4034 19848
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 6086 19836 6092 19848
rect 4387 19808 6092 19836
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 6086 19796 6092 19808
rect 6144 19796 6150 19848
rect 7926 19796 7932 19848
rect 7984 19796 7990 19848
rect 8018 19796 8024 19848
rect 8076 19836 8082 19848
rect 9585 19839 9643 19845
rect 9585 19836 9597 19839
rect 8076 19808 9597 19836
rect 8076 19796 8082 19808
rect 9585 19805 9597 19808
rect 9631 19836 9643 19839
rect 11146 19836 11152 19848
rect 9631 19808 11152 19836
rect 9631 19805 9643 19808
rect 9585 19799 9643 19805
rect 11146 19796 11152 19808
rect 11204 19796 11210 19848
rect 11238 19796 11244 19848
rect 11296 19796 11302 19848
rect 12802 19796 12808 19848
rect 12860 19845 12866 19848
rect 12860 19836 12872 19845
rect 14274 19836 14280 19848
rect 12860 19808 12905 19836
rect 13740 19808 14280 19836
rect 12860 19799 12872 19808
rect 12860 19796 12866 19799
rect 2314 19777 2320 19780
rect 2308 19731 2320 19777
rect 2314 19728 2320 19731
rect 2372 19728 2378 19780
rect 4608 19771 4666 19777
rect 4608 19737 4620 19771
rect 4654 19768 4666 19771
rect 5074 19768 5080 19780
rect 4654 19740 5080 19768
rect 4654 19737 4666 19740
rect 4608 19731 4666 19737
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 7282 19728 7288 19780
rect 7340 19728 7346 19780
rect 7561 19771 7619 19777
rect 7561 19737 7573 19771
rect 7607 19768 7619 19771
rect 8110 19768 8116 19780
rect 7607 19740 8116 19768
rect 7607 19737 7619 19740
rect 7561 19731 7619 19737
rect 8110 19728 8116 19740
rect 8168 19728 8174 19780
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 10226 19768 10232 19780
rect 9916 19740 10232 19768
rect 9916 19728 9922 19740
rect 10226 19728 10232 19740
rect 10284 19768 10290 19780
rect 10597 19771 10655 19777
rect 10597 19768 10609 19771
rect 10284 19740 10609 19768
rect 10284 19728 10290 19740
rect 10597 19737 10609 19740
rect 10643 19737 10655 19771
rect 13446 19768 13452 19780
rect 10597 19731 10655 19737
rect 10888 19740 13452 19768
rect 10888 19712 10916 19740
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 13740 19777 13768 19808
rect 14274 19796 14280 19808
rect 14332 19836 14338 19848
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 14332 19808 14473 19836
rect 14332 19796 14338 19808
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 13541 19771 13599 19777
rect 13541 19737 13553 19771
rect 13587 19737 13599 19771
rect 13541 19731 13599 19737
rect 13725 19771 13783 19777
rect 13725 19737 13737 19771
rect 13771 19737 13783 19771
rect 13725 19731 13783 19737
rect 3786 19660 3792 19712
rect 3844 19660 3850 19712
rect 5810 19660 5816 19712
rect 5868 19700 5874 19712
rect 6991 19703 7049 19709
rect 6991 19700 7003 19703
rect 5868 19672 7003 19700
rect 5868 19660 5874 19672
rect 6991 19669 7003 19672
rect 7037 19669 7049 19703
rect 6991 19663 7049 19669
rect 7466 19660 7472 19712
rect 7524 19660 7530 19712
rect 9493 19703 9551 19709
rect 9493 19669 9505 19703
rect 9539 19700 9551 19703
rect 9674 19700 9680 19712
rect 9539 19672 9680 19700
rect 9539 19669 9551 19672
rect 9493 19663 9551 19669
rect 9674 19660 9680 19672
rect 9732 19700 9738 19712
rect 9950 19700 9956 19712
rect 9732 19672 9956 19700
rect 9732 19660 9738 19672
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 10870 19660 10876 19712
rect 10928 19660 10934 19712
rect 11425 19703 11483 19709
rect 11425 19669 11437 19703
rect 11471 19700 11483 19703
rect 11606 19700 11612 19712
rect 11471 19672 11612 19700
rect 11471 19669 11483 19672
rect 11425 19663 11483 19669
rect 11606 19660 11612 19672
rect 11664 19660 11670 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 13556 19700 13584 19731
rect 13814 19728 13820 19780
rect 13872 19768 13878 19780
rect 14568 19768 14596 19876
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 15105 19839 15163 19845
rect 13872 19740 14596 19768
rect 14660 19808 15056 19836
rect 13872 19728 13878 19740
rect 14660 19709 14688 19808
rect 14734 19728 14740 19780
rect 14792 19728 14798 19780
rect 15028 19768 15056 19808
rect 15105 19805 15117 19839
rect 15151 19836 15163 19839
rect 15194 19836 15200 19848
rect 15151 19808 15200 19836
rect 15151 19805 15163 19808
rect 15105 19799 15163 19805
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19836 16175 19839
rect 16500 19836 16528 19935
rect 17034 19932 17040 19984
rect 17092 19972 17098 19984
rect 17865 19975 17923 19981
rect 17865 19972 17877 19975
rect 17092 19944 17877 19972
rect 17092 19932 17098 19944
rect 17865 19941 17877 19944
rect 17911 19941 17923 19975
rect 17865 19935 17923 19941
rect 18138 19864 18144 19916
rect 18196 19904 18202 19916
rect 18322 19904 18328 19916
rect 18196 19876 18328 19904
rect 18196 19864 18202 19876
rect 18322 19864 18328 19876
rect 18380 19904 18386 19916
rect 19702 19904 19708 19916
rect 18380 19876 18828 19904
rect 18380 19864 18386 19876
rect 17402 19836 17408 19848
rect 16163 19808 16528 19836
rect 16960 19808 17408 19836
rect 16163 19805 16175 19808
rect 16117 19799 16175 19805
rect 15470 19768 15476 19780
rect 15028 19740 15476 19768
rect 15470 19728 15476 19740
rect 15528 19768 15534 19780
rect 16206 19768 16212 19780
rect 15528 19740 16212 19768
rect 15528 19728 15534 19740
rect 16206 19728 16212 19740
rect 16264 19728 16270 19780
rect 16758 19728 16764 19780
rect 16816 19728 16822 19780
rect 16960 19777 16988 19808
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 18046 19796 18052 19848
rect 18104 19796 18110 19848
rect 18506 19796 18512 19848
rect 18564 19796 18570 19848
rect 18598 19796 18604 19848
rect 18656 19796 18662 19848
rect 18800 19845 18828 19876
rect 19536 19876 19708 19904
rect 18785 19839 18843 19845
rect 18785 19805 18797 19839
rect 18831 19805 18843 19839
rect 18785 19799 18843 19805
rect 16945 19771 17003 19777
rect 16945 19737 16957 19771
rect 16991 19737 17003 19771
rect 16945 19731 17003 19737
rect 17037 19771 17095 19777
rect 17037 19737 17049 19771
rect 17083 19737 17095 19771
rect 17037 19731 17095 19737
rect 11848 19672 13584 19700
rect 14645 19703 14703 19709
rect 11848 19660 11854 19672
rect 14645 19669 14657 19703
rect 14691 19669 14703 19703
rect 14645 19663 14703 19669
rect 14921 19703 14979 19709
rect 14921 19669 14933 19703
rect 14967 19700 14979 19703
rect 15102 19700 15108 19712
rect 14967 19672 15108 19700
rect 14967 19669 14979 19672
rect 14921 19663 14979 19669
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 16301 19703 16359 19709
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 16850 19700 16856 19712
rect 16347 19672 16856 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 17052 19700 17080 19731
rect 17126 19728 17132 19780
rect 17184 19768 17190 19780
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 17184 19740 17325 19768
rect 17184 19728 17190 19740
rect 17313 19737 17325 19740
rect 17359 19737 17371 19771
rect 17313 19731 17371 19737
rect 17586 19728 17592 19780
rect 17644 19728 17650 19780
rect 18966 19728 18972 19780
rect 19024 19768 19030 19780
rect 19536 19777 19564 19876
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 19852 19808 20177 19836
rect 19852 19796 19858 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 20432 19839 20490 19845
rect 20432 19805 20444 19839
rect 20478 19836 20490 19839
rect 20898 19836 20904 19848
rect 20478 19808 20904 19836
rect 20478 19805 20490 19808
rect 20432 19799 20490 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 19429 19771 19487 19777
rect 19429 19768 19441 19771
rect 19024 19740 19441 19768
rect 19024 19728 19030 19740
rect 19429 19737 19441 19740
rect 19475 19737 19487 19771
rect 19429 19731 19487 19737
rect 19521 19771 19579 19777
rect 19521 19737 19533 19771
rect 19567 19737 19579 19771
rect 19521 19731 19579 19737
rect 19705 19771 19763 19777
rect 19705 19737 19717 19771
rect 19751 19768 19763 19771
rect 21266 19768 21272 19780
rect 19751 19740 21272 19768
rect 19751 19737 19763 19740
rect 19705 19731 19763 19737
rect 21266 19728 21272 19740
rect 21324 19728 21330 19780
rect 17218 19700 17224 19712
rect 17052 19672 17224 19700
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 17405 19703 17463 19709
rect 17405 19669 17417 19703
rect 17451 19700 17463 19703
rect 17862 19700 17868 19712
rect 17451 19672 17868 19700
rect 17451 19669 17463 19672
rect 17405 19663 17463 19669
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 18233 19703 18291 19709
rect 18233 19669 18245 19703
rect 18279 19700 18291 19703
rect 18322 19700 18328 19712
rect 18279 19672 18328 19700
rect 18279 19669 18291 19672
rect 18233 19663 18291 19669
rect 18322 19660 18328 19672
rect 18380 19660 18386 19712
rect 19999 19703 20057 19709
rect 19999 19669 20011 19703
rect 20045 19700 20057 19703
rect 21450 19700 21456 19712
rect 20045 19672 21456 19700
rect 20045 19669 20057 19672
rect 19999 19663 20057 19669
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 1104 19610 21988 19632
rect 1104 19558 4220 19610
rect 4272 19558 4284 19610
rect 4336 19558 4348 19610
rect 4400 19558 4412 19610
rect 4464 19558 4476 19610
rect 4528 19558 9441 19610
rect 9493 19558 9505 19610
rect 9557 19558 9569 19610
rect 9621 19558 9633 19610
rect 9685 19558 9697 19610
rect 9749 19558 14662 19610
rect 14714 19558 14726 19610
rect 14778 19558 14790 19610
rect 14842 19558 14854 19610
rect 14906 19558 14918 19610
rect 14970 19558 19883 19610
rect 19935 19558 19947 19610
rect 19999 19558 20011 19610
rect 20063 19558 20075 19610
rect 20127 19558 20139 19610
rect 20191 19558 21988 19610
rect 1104 19536 21988 19558
rect 2225 19499 2283 19505
rect 2225 19465 2237 19499
rect 2271 19496 2283 19499
rect 2314 19496 2320 19508
rect 2271 19468 2320 19496
rect 2271 19465 2283 19468
rect 2225 19459 2283 19465
rect 2314 19456 2320 19468
rect 2372 19456 2378 19508
rect 4614 19456 4620 19508
rect 4672 19496 4678 19508
rect 4709 19499 4767 19505
rect 4709 19496 4721 19499
rect 4672 19468 4721 19496
rect 4672 19456 4678 19468
rect 4709 19465 4721 19468
rect 4755 19496 4767 19499
rect 5442 19496 5448 19508
rect 4755 19468 5448 19496
rect 4755 19465 4767 19468
rect 4709 19459 4767 19465
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 5997 19499 6055 19505
rect 5997 19465 6009 19499
rect 6043 19496 6055 19499
rect 7650 19496 7656 19508
rect 6043 19468 7656 19496
rect 6043 19465 6055 19468
rect 5997 19459 6055 19465
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 7827 19499 7885 19505
rect 7827 19465 7839 19499
rect 7873 19496 7885 19499
rect 7926 19496 7932 19508
rect 7873 19468 7932 19496
rect 7873 19465 7885 19468
rect 7827 19459 7885 19465
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8018 19456 8024 19508
rect 8076 19496 8082 19508
rect 8297 19499 8355 19505
rect 8297 19496 8309 19499
rect 8076 19468 8309 19496
rect 8076 19456 8082 19468
rect 8297 19465 8309 19468
rect 8343 19496 8355 19499
rect 8662 19496 8668 19508
rect 8343 19468 8668 19496
rect 8343 19465 8355 19468
rect 8297 19459 8355 19465
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 9674 19496 9680 19508
rect 9232 19468 9680 19496
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 2774 19428 2780 19440
rect 2547 19400 2780 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 2774 19388 2780 19400
rect 2832 19428 2838 19440
rect 3596 19431 3654 19437
rect 2832 19400 3372 19428
rect 2832 19388 2838 19400
rect 2038 19320 2044 19372
rect 2096 19320 2102 19372
rect 3050 19320 3056 19372
rect 3108 19360 3114 19372
rect 3344 19369 3372 19400
rect 3596 19397 3608 19431
rect 3642 19428 3654 19431
rect 3786 19428 3792 19440
rect 3642 19400 3792 19428
rect 3642 19397 3654 19400
rect 3596 19391 3654 19397
rect 3786 19388 3792 19400
rect 3844 19388 3850 19440
rect 5810 19388 5816 19440
rect 5868 19388 5874 19440
rect 6089 19431 6147 19437
rect 6089 19397 6101 19431
rect 6135 19428 6147 19431
rect 6914 19428 6920 19440
rect 6135 19400 6920 19428
rect 6135 19397 6147 19400
rect 6089 19391 6147 19397
rect 6914 19388 6920 19400
rect 6972 19388 6978 19440
rect 7469 19431 7527 19437
rect 7469 19428 7481 19431
rect 7392 19400 7481 19428
rect 3237 19363 3295 19369
rect 3237 19360 3249 19363
rect 3108 19332 3249 19360
rect 3108 19320 3114 19332
rect 3237 19329 3249 19332
rect 3283 19329 3295 19363
rect 3237 19323 3295 19329
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19329 3387 19363
rect 3329 19323 3387 19329
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 6457 19363 6515 19369
rect 6457 19360 6469 19363
rect 4764 19332 6469 19360
rect 4764 19320 4770 19332
rect 6457 19329 6469 19332
rect 6503 19360 6515 19363
rect 7282 19360 7288 19372
rect 6503 19332 7288 19360
rect 6503 19329 6515 19332
rect 6457 19323 6515 19329
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7392 19292 7420 19400
rect 7469 19397 7481 19400
rect 7515 19397 7527 19431
rect 7469 19391 7527 19397
rect 7561 19431 7619 19437
rect 7561 19397 7573 19431
rect 7607 19428 7619 19431
rect 8202 19428 8208 19440
rect 7607 19400 8208 19428
rect 7607 19397 7619 19400
rect 7561 19391 7619 19397
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 9122 19428 9128 19440
rect 8312 19400 9128 19428
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 8312 19360 8340 19400
rect 9122 19388 9128 19400
rect 9180 19428 9186 19440
rect 9232 19428 9260 19468
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 9858 19456 9864 19508
rect 9916 19456 9922 19508
rect 12066 19456 12072 19508
rect 12124 19496 12130 19508
rect 12897 19499 12955 19505
rect 12897 19496 12909 19499
rect 12124 19468 12909 19496
rect 12124 19456 12130 19468
rect 12897 19465 12909 19468
rect 12943 19465 12955 19499
rect 12897 19459 12955 19465
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 14645 19499 14703 19505
rect 14645 19496 14657 19499
rect 14608 19468 14657 19496
rect 14608 19456 14614 19468
rect 14645 19465 14657 19468
rect 14691 19465 14703 19499
rect 14645 19459 14703 19465
rect 16206 19456 16212 19508
rect 16264 19456 16270 19508
rect 17402 19456 17408 19508
rect 17460 19496 17466 19508
rect 18049 19499 18107 19505
rect 18049 19496 18061 19499
rect 17460 19468 18061 19496
rect 17460 19456 17466 19468
rect 18049 19465 18061 19468
rect 18095 19465 18107 19499
rect 18049 19459 18107 19465
rect 19610 19456 19616 19508
rect 19668 19456 19674 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 21266 19496 21272 19508
rect 21223 19468 21272 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 21361 19499 21419 19505
rect 21361 19465 21373 19499
rect 21407 19465 21419 19499
rect 21361 19459 21419 19465
rect 13906 19428 13912 19440
rect 9180 19400 9260 19428
rect 9324 19400 11284 19428
rect 9180 19388 9186 19400
rect 8159 19332 8340 19360
rect 8389 19363 8447 19369
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 8389 19329 8401 19363
rect 8435 19360 8447 19363
rect 8478 19360 8484 19372
rect 8435 19332 8484 19360
rect 8435 19329 8447 19332
rect 8389 19323 8447 19329
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 8570 19320 8576 19372
rect 8628 19320 8634 19372
rect 6840 19264 7420 19292
rect 6840 19168 6868 19264
rect 7466 19252 7472 19304
rect 7524 19252 7530 19304
rect 9324 19301 9352 19400
rect 10686 19320 10692 19372
rect 10744 19360 10750 19372
rect 11256 19369 11284 19400
rect 11532 19400 12434 19428
rect 11532 19369 11560 19400
rect 12406 19372 12434 19400
rect 10974 19363 11032 19369
rect 10974 19360 10986 19363
rect 10744 19332 10986 19360
rect 10744 19320 10750 19332
rect 10974 19329 10986 19332
rect 11020 19329 11032 19363
rect 10974 19323 11032 19329
rect 11241 19363 11299 19369
rect 11241 19329 11253 19363
rect 11287 19329 11299 19363
rect 11241 19323 11299 19329
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19329 11575 19363
rect 11517 19323 11575 19329
rect 11606 19320 11612 19372
rect 11664 19360 11670 19372
rect 11773 19363 11831 19369
rect 11773 19360 11785 19363
rect 11664 19332 11785 19360
rect 11664 19320 11670 19332
rect 11773 19329 11785 19332
rect 11819 19329 11831 19363
rect 11773 19323 11831 19329
rect 12342 19320 12348 19372
rect 12400 19360 12434 19372
rect 13280 19400 13912 19428
rect 13280 19369 13308 19400
rect 13906 19388 13912 19400
rect 13964 19388 13970 19440
rect 15102 19437 15108 19440
rect 15096 19428 15108 19437
rect 15063 19400 15108 19428
rect 15096 19391 15108 19400
rect 15102 19388 15108 19391
rect 15160 19388 15166 19440
rect 20064 19431 20122 19437
rect 16684 19400 19840 19428
rect 13538 19369 13544 19372
rect 13265 19363 13323 19369
rect 13265 19360 13277 19363
rect 12400 19332 13277 19360
rect 12400 19320 12406 19332
rect 13265 19329 13277 19332
rect 13311 19329 13323 19363
rect 13265 19323 13323 19329
rect 13532 19323 13544 19369
rect 13538 19320 13544 19323
rect 13596 19320 13602 19372
rect 13924 19360 13952 19388
rect 16684 19369 16712 19400
rect 16942 19369 16948 19372
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 13924 19332 14841 19360
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 14829 19323 14887 19329
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19329 16727 19363
rect 16936 19360 16948 19369
rect 16903 19332 16948 19360
rect 16669 19323 16727 19329
rect 16936 19323 16948 19332
rect 16942 19320 16948 19323
rect 17000 19320 17006 19372
rect 18248 19369 18276 19400
rect 19812 19372 19840 19400
rect 20064 19397 20076 19431
rect 20110 19428 20122 19431
rect 21376 19428 21404 19459
rect 20110 19400 21404 19428
rect 20110 19397 20122 19400
rect 20064 19391 20122 19397
rect 18233 19363 18291 19369
rect 18233 19329 18245 19363
rect 18279 19329 18291 19363
rect 18233 19323 18291 19329
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18489 19363 18547 19369
rect 18489 19360 18501 19363
rect 18380 19332 18501 19360
rect 18380 19320 18386 19332
rect 18489 19329 18501 19332
rect 18535 19329 18547 19363
rect 18489 19323 18547 19329
rect 19794 19320 19800 19372
rect 19852 19320 19858 19372
rect 21450 19320 21456 19372
rect 21508 19360 21514 19372
rect 21545 19363 21603 19369
rect 21545 19360 21557 19363
rect 21508 19332 21557 19360
rect 21508 19320 21514 19332
rect 21545 19329 21557 19332
rect 21591 19329 21603 19363
rect 21545 19323 21603 19329
rect 9309 19295 9367 19301
rect 9309 19261 9321 19295
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 9324 19224 9352 19255
rect 8352 19196 9352 19224
rect 8352 19184 8358 19196
rect 5537 19159 5595 19165
rect 5537 19125 5549 19159
rect 5583 19156 5595 19159
rect 5994 19156 6000 19168
rect 5583 19128 6000 19156
rect 5583 19125 5595 19128
rect 5537 19119 5595 19125
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 6733 19159 6791 19165
rect 6733 19125 6745 19159
rect 6779 19156 6791 19159
rect 6822 19156 6828 19168
rect 6779 19128 6828 19156
rect 6779 19125 6791 19128
rect 6733 19119 6791 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7009 19159 7067 19165
rect 7009 19125 7021 19159
rect 7055 19156 7067 19159
rect 7098 19156 7104 19168
rect 7055 19128 7104 19156
rect 7055 19125 7067 19128
rect 7009 19119 7067 19125
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 10870 19156 10876 19168
rect 9732 19128 10876 19156
rect 9732 19116 9738 19128
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 15010 19156 15016 19168
rect 11848 19128 15016 19156
rect 11848 19116 11854 19128
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 18506 19116 18512 19168
rect 18564 19156 18570 19168
rect 20990 19156 20996 19168
rect 18564 19128 20996 19156
rect 18564 19116 18570 19128
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 1104 19066 21988 19088
rect 1104 19014 3560 19066
rect 3612 19014 3624 19066
rect 3676 19014 3688 19066
rect 3740 19014 3752 19066
rect 3804 19014 3816 19066
rect 3868 19014 8781 19066
rect 8833 19014 8845 19066
rect 8897 19014 8909 19066
rect 8961 19014 8973 19066
rect 9025 19014 9037 19066
rect 9089 19014 14002 19066
rect 14054 19014 14066 19066
rect 14118 19014 14130 19066
rect 14182 19014 14194 19066
rect 14246 19014 14258 19066
rect 14310 19014 19223 19066
rect 19275 19014 19287 19066
rect 19339 19014 19351 19066
rect 19403 19014 19415 19066
rect 19467 19014 19479 19066
rect 19531 19014 21988 19066
rect 1104 18992 21988 19014
rect 1302 18912 1308 18964
rect 1360 18952 1366 18964
rect 2777 18955 2835 18961
rect 2777 18952 2789 18955
rect 1360 18924 2789 18952
rect 1360 18912 1366 18924
rect 2777 18921 2789 18924
rect 2823 18921 2835 18955
rect 2777 18915 2835 18921
rect 4706 18912 4712 18964
rect 4764 18912 4770 18964
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 7929 18955 7987 18961
rect 7929 18952 7941 18955
rect 7524 18924 7941 18952
rect 7524 18912 7530 18924
rect 7929 18921 7941 18924
rect 7975 18921 7987 18955
rect 7929 18915 7987 18921
rect 10686 18912 10692 18964
rect 10744 18912 10750 18964
rect 13725 18955 13783 18961
rect 13725 18921 13737 18955
rect 13771 18952 13783 18955
rect 14366 18952 14372 18964
rect 13771 18924 14372 18952
rect 13771 18921 13783 18924
rect 13725 18915 13783 18921
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 15194 18912 15200 18964
rect 15252 18912 15258 18964
rect 17586 18912 17592 18964
rect 17644 18912 17650 18964
rect 18046 18912 18052 18964
rect 18104 18952 18110 18964
rect 18233 18955 18291 18961
rect 18233 18952 18245 18955
rect 18104 18924 18245 18952
rect 18104 18912 18110 18924
rect 18233 18921 18245 18924
rect 18279 18921 18291 18955
rect 19610 18952 19616 18964
rect 18233 18915 18291 18921
rect 19260 18924 19616 18952
rect 2498 18844 2504 18896
rect 2556 18884 2562 18896
rect 3881 18887 3939 18893
rect 3881 18884 3893 18887
rect 2556 18856 3893 18884
rect 2556 18844 2562 18856
rect 3881 18853 3893 18856
rect 3927 18853 3939 18887
rect 3881 18847 3939 18853
rect 8294 18844 8300 18896
rect 8352 18844 8358 18896
rect 10965 18887 11023 18893
rect 10965 18853 10977 18887
rect 11011 18853 11023 18887
rect 10965 18847 11023 18853
rect 2682 18776 2688 18828
rect 2740 18816 2746 18828
rect 3053 18819 3111 18825
rect 3053 18816 3065 18819
rect 2740 18788 3065 18816
rect 2740 18776 2746 18788
rect 3053 18785 3065 18788
rect 3099 18816 3111 18819
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 3099 18788 4353 18816
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 4341 18785 4353 18788
rect 4387 18816 4399 18819
rect 4614 18816 4620 18828
rect 4387 18788 4620 18816
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 6086 18776 6092 18828
rect 6144 18816 6150 18828
rect 6549 18819 6607 18825
rect 6549 18816 6561 18819
rect 6144 18788 6561 18816
rect 6144 18776 6150 18788
rect 6549 18785 6561 18788
rect 6595 18785 6607 18819
rect 8312 18816 8340 18844
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 8312 18788 8953 18816
rect 6549 18779 6607 18785
rect 8941 18785 8953 18788
rect 8987 18785 8999 18819
rect 8941 18779 8999 18785
rect 1397 18751 1455 18757
rect 1397 18717 1409 18751
rect 1443 18748 1455 18751
rect 2774 18748 2780 18760
rect 1443 18720 2780 18748
rect 1443 18717 1455 18720
rect 1397 18711 1455 18717
rect 2774 18708 2780 18720
rect 2832 18708 2838 18760
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18748 3663 18751
rect 5534 18748 5540 18760
rect 3651 18720 5540 18748
rect 3651 18717 3663 18720
rect 3605 18711 3663 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 6273 18751 6331 18757
rect 6273 18717 6285 18751
rect 6319 18748 6331 18751
rect 7098 18748 7104 18760
rect 6319 18720 7104 18748
rect 6319 18717 6331 18720
rect 6273 18711 6331 18717
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 8386 18748 8392 18760
rect 8343 18720 8392 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18748 8631 18751
rect 10134 18748 10140 18760
rect 8619 18720 10140 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 10980 18748 11008 18847
rect 14274 18844 14280 18896
rect 14332 18884 14338 18896
rect 14734 18884 14740 18896
rect 14332 18856 14740 18884
rect 14332 18844 14338 18856
rect 14734 18844 14740 18856
rect 14792 18844 14798 18896
rect 16114 18844 16120 18896
rect 16172 18844 16178 18896
rect 12342 18776 12348 18828
rect 12400 18776 12406 18828
rect 13906 18776 13912 18828
rect 13964 18816 13970 18828
rect 14185 18819 14243 18825
rect 14185 18816 14197 18819
rect 13964 18788 14197 18816
rect 13964 18776 13970 18788
rect 14185 18785 14197 18788
rect 14231 18816 14243 18819
rect 16209 18819 16267 18825
rect 16209 18816 16221 18819
rect 14231 18788 16221 18816
rect 14231 18785 14243 18788
rect 14185 18779 14243 18785
rect 16209 18785 16221 18788
rect 16255 18785 16267 18819
rect 16209 18779 16267 18785
rect 18693 18819 18751 18825
rect 18693 18785 18705 18819
rect 18739 18816 18751 18819
rect 19260 18816 19288 18924
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 20622 18912 20628 18964
rect 20680 18912 20686 18964
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 21048 18924 21496 18952
rect 21048 18912 21054 18924
rect 21361 18887 21419 18893
rect 21361 18853 21373 18887
rect 21407 18853 21419 18887
rect 21361 18847 21419 18853
rect 21376 18816 21404 18847
rect 18739 18788 19288 18816
rect 20456 18788 21404 18816
rect 18739 18785 18751 18788
rect 18693 18779 18751 18785
rect 10551 18720 11008 18748
rect 11241 18751 11299 18757
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 11241 18717 11253 18751
rect 11287 18748 11299 18751
rect 11287 18720 12434 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 12406 18692 12434 18720
rect 15470 18708 15476 18760
rect 15528 18708 15534 18760
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 17034 18748 17040 18760
rect 15979 18720 17040 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 17034 18708 17040 18720
rect 17092 18708 17098 18760
rect 17773 18751 17831 18757
rect 17773 18717 17785 18751
rect 17819 18717 17831 18751
rect 17773 18711 17831 18717
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18748 19303 18751
rect 19794 18748 19800 18760
rect 19291 18720 19800 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 1486 18640 1492 18692
rect 1544 18680 1550 18692
rect 1642 18683 1700 18689
rect 1642 18680 1654 18683
rect 1544 18652 1654 18680
rect 1544 18640 1550 18652
rect 1642 18649 1654 18652
rect 1688 18649 1700 18683
rect 1642 18643 1700 18649
rect 4433 18683 4491 18689
rect 4433 18649 4445 18683
rect 4479 18680 4491 18683
rect 4890 18680 4896 18692
rect 4479 18652 4896 18680
rect 4479 18649 4491 18652
rect 4433 18643 4491 18649
rect 4890 18640 4896 18652
rect 4948 18680 4954 18692
rect 5074 18680 5080 18692
rect 4948 18652 5080 18680
rect 4948 18640 4954 18652
rect 5074 18640 5080 18652
rect 5132 18640 5138 18692
rect 5844 18683 5902 18689
rect 5844 18649 5856 18683
rect 5890 18680 5902 18683
rect 6178 18680 6184 18692
rect 5890 18652 6184 18680
rect 5890 18649 5902 18652
rect 5844 18643 5902 18649
rect 6178 18640 6184 18652
rect 6236 18640 6242 18692
rect 6794 18683 6852 18689
rect 6794 18680 6806 18683
rect 6472 18652 6806 18680
rect 3234 18572 3240 18624
rect 3292 18612 3298 18624
rect 6472 18621 6500 18652
rect 6794 18649 6806 18652
rect 6840 18649 6852 18683
rect 9186 18683 9244 18689
rect 9186 18680 9198 18683
rect 6794 18643 6852 18649
rect 8772 18652 9198 18680
rect 4341 18615 4399 18621
rect 4341 18612 4353 18615
rect 3292 18584 4353 18612
rect 3292 18572 3298 18584
rect 4341 18581 4353 18584
rect 4387 18581 4399 18615
rect 4341 18575 4399 18581
rect 6457 18615 6515 18621
rect 6457 18581 6469 18615
rect 6503 18581 6515 18615
rect 6457 18575 6515 18581
rect 8481 18615 8539 18621
rect 8481 18581 8493 18615
rect 8527 18612 8539 18615
rect 8570 18612 8576 18624
rect 8527 18584 8576 18612
rect 8527 18581 8539 18584
rect 8481 18575 8539 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8772 18621 8800 18652
rect 9186 18649 9198 18652
rect 9232 18649 9244 18683
rect 9186 18643 9244 18649
rect 11514 18640 11520 18692
rect 11572 18640 11578 18692
rect 12406 18652 12440 18692
rect 12434 18640 12440 18652
rect 12492 18640 12498 18692
rect 12612 18683 12670 18689
rect 12612 18649 12624 18683
rect 12658 18680 12670 18683
rect 12710 18680 12716 18692
rect 12658 18652 12716 18680
rect 12658 18649 12670 18652
rect 12612 18643 12670 18649
rect 12710 18640 12716 18652
rect 12768 18640 12774 18692
rect 15010 18640 15016 18692
rect 15068 18640 15074 18692
rect 15749 18683 15807 18689
rect 15749 18680 15761 18683
rect 15580 18652 15761 18680
rect 8757 18615 8815 18621
rect 8757 18581 8769 18615
rect 8803 18581 8815 18615
rect 8757 18575 8815 18581
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 11425 18615 11483 18621
rect 11425 18612 11437 18615
rect 11204 18584 11437 18612
rect 11204 18572 11210 18584
rect 11425 18581 11437 18584
rect 11471 18581 11483 18615
rect 11425 18575 11483 18581
rect 11606 18572 11612 18624
rect 11664 18612 11670 18624
rect 15580 18612 15608 18652
rect 15749 18649 15761 18652
rect 15795 18649 15807 18683
rect 15749 18643 15807 18649
rect 11664 18584 15608 18612
rect 11664 18572 11670 18584
rect 15654 18572 15660 18624
rect 15712 18572 15718 18624
rect 15764 18612 15792 18643
rect 16114 18640 16120 18692
rect 16172 18680 16178 18692
rect 16454 18683 16512 18689
rect 16454 18680 16466 18683
rect 16172 18652 16466 18680
rect 16172 18640 16178 18652
rect 16454 18649 16466 18652
rect 16500 18649 16512 18683
rect 16454 18643 16512 18649
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 17788 18680 17816 18711
rect 19794 18708 19800 18720
rect 19852 18708 19858 18760
rect 16724 18652 17816 18680
rect 18785 18683 18843 18689
rect 16724 18640 16730 18652
rect 18785 18649 18797 18683
rect 18831 18680 18843 18683
rect 18874 18680 18880 18692
rect 18831 18652 18880 18680
rect 18831 18649 18843 18652
rect 18785 18643 18843 18649
rect 18874 18640 18880 18652
rect 18932 18640 18938 18692
rect 19512 18683 19570 18689
rect 19512 18649 19524 18683
rect 19558 18680 19570 18683
rect 20456 18680 20484 18788
rect 20806 18708 20812 18760
rect 20864 18708 20870 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20916 18720 21097 18748
rect 19558 18652 20484 18680
rect 19558 18649 19570 18652
rect 19512 18643 19570 18649
rect 20622 18640 20628 18692
rect 20680 18680 20686 18692
rect 20916 18680 20944 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 21174 18708 21180 18760
rect 21232 18757 21238 18760
rect 21232 18751 21287 18757
rect 21232 18717 21241 18751
rect 21275 18748 21287 18751
rect 21468 18748 21496 18924
rect 21275 18720 21496 18748
rect 21275 18717 21287 18720
rect 21232 18711 21287 18717
rect 21232 18708 21238 18711
rect 20680 18652 20944 18680
rect 20993 18683 21051 18689
rect 20680 18640 20686 18652
rect 20993 18649 21005 18683
rect 21039 18680 21051 18683
rect 21358 18680 21364 18692
rect 21039 18652 21364 18680
rect 21039 18649 21051 18652
rect 20993 18643 21051 18649
rect 21358 18640 21364 18652
rect 21416 18640 21422 18692
rect 17126 18612 17132 18624
rect 15764 18584 17132 18612
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 17862 18572 17868 18624
rect 17920 18612 17926 18624
rect 17957 18615 18015 18621
rect 17957 18612 17969 18615
rect 17920 18584 17969 18612
rect 17920 18572 17926 18584
rect 17957 18581 17969 18584
rect 18003 18581 18015 18615
rect 17957 18575 18015 18581
rect 18414 18572 18420 18624
rect 18472 18612 18478 18624
rect 18693 18615 18751 18621
rect 18693 18612 18705 18615
rect 18472 18584 18705 18612
rect 18472 18572 18478 18584
rect 18693 18581 18705 18584
rect 18739 18581 18751 18615
rect 18693 18575 18751 18581
rect 1104 18522 21988 18544
rect 1104 18470 4220 18522
rect 4272 18470 4284 18522
rect 4336 18470 4348 18522
rect 4400 18470 4412 18522
rect 4464 18470 4476 18522
rect 4528 18470 9441 18522
rect 9493 18470 9505 18522
rect 9557 18470 9569 18522
rect 9621 18470 9633 18522
rect 9685 18470 9697 18522
rect 9749 18470 14662 18522
rect 14714 18470 14726 18522
rect 14778 18470 14790 18522
rect 14842 18470 14854 18522
rect 14906 18470 14918 18522
rect 14970 18470 19883 18522
rect 19935 18470 19947 18522
rect 19999 18470 20011 18522
rect 20063 18470 20075 18522
rect 20127 18470 20139 18522
rect 20191 18470 21988 18522
rect 1104 18448 21988 18470
rect 1486 18368 1492 18420
rect 1544 18368 1550 18420
rect 2682 18368 2688 18420
rect 2740 18368 2746 18420
rect 4338 18368 4344 18420
rect 4396 18368 4402 18420
rect 6181 18411 6239 18417
rect 6181 18377 6193 18411
rect 6227 18377 6239 18411
rect 6181 18371 6239 18377
rect 1302 18300 1308 18352
rect 1360 18340 1366 18352
rect 2317 18343 2375 18349
rect 2317 18340 2329 18343
rect 1360 18312 2329 18340
rect 1360 18300 1366 18312
rect 2317 18309 2329 18312
rect 2363 18309 2375 18343
rect 2317 18303 2375 18309
rect 2774 18300 2780 18352
rect 2832 18340 2838 18352
rect 6196 18340 6224 18371
rect 7650 18368 7656 18420
rect 7708 18408 7714 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7708 18380 7757 18408
rect 7708 18368 7714 18380
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 7745 18371 7803 18377
rect 9861 18411 9919 18417
rect 9861 18377 9873 18411
rect 9907 18408 9919 18411
rect 9950 18408 9956 18420
rect 9907 18380 9956 18408
rect 9907 18377 9919 18380
rect 9861 18371 9919 18377
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 10597 18411 10655 18417
rect 10597 18377 10609 18411
rect 10643 18408 10655 18411
rect 10870 18408 10876 18420
rect 10643 18380 10876 18408
rect 10643 18377 10655 18380
rect 10597 18371 10655 18377
rect 10870 18368 10876 18380
rect 10928 18408 10934 18420
rect 11146 18408 11152 18420
rect 10928 18380 11152 18408
rect 10928 18368 10934 18380
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 12710 18368 12716 18420
rect 12768 18368 12774 18420
rect 13449 18411 13507 18417
rect 13449 18377 13461 18411
rect 13495 18408 13507 18411
rect 13538 18408 13544 18420
rect 13495 18380 13544 18408
rect 13495 18377 13507 18380
rect 13449 18371 13507 18377
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 14550 18368 14556 18420
rect 14608 18408 14614 18420
rect 14645 18411 14703 18417
rect 14645 18408 14657 18411
rect 14608 18380 14657 18408
rect 14608 18368 14614 18380
rect 14645 18377 14657 18380
rect 14691 18377 14703 18411
rect 14645 18371 14703 18377
rect 15654 18368 15660 18420
rect 15712 18408 15718 18420
rect 17221 18411 17279 18417
rect 15712 18380 17172 18408
rect 15712 18368 15718 18380
rect 6610 18343 6668 18349
rect 6610 18340 6622 18343
rect 2832 18312 4108 18340
rect 6196 18312 6622 18340
rect 2832 18300 2838 18312
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 2133 18275 2191 18281
rect 1719 18244 1900 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1872 18145 1900 18244
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2498 18272 2504 18284
rect 2179 18244 2504 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2498 18232 2504 18244
rect 2556 18232 2562 18284
rect 3809 18275 3867 18281
rect 3809 18241 3821 18275
rect 3855 18272 3867 18275
rect 3970 18272 3976 18284
rect 3855 18244 3976 18272
rect 3855 18241 3867 18244
rect 3809 18235 3867 18241
rect 3970 18232 3976 18244
rect 4028 18232 4034 18284
rect 4080 18281 4108 18312
rect 6610 18309 6622 18312
rect 6656 18309 6668 18343
rect 6610 18303 6668 18309
rect 10318 18300 10324 18352
rect 10376 18340 10382 18352
rect 10413 18343 10471 18349
rect 10413 18340 10425 18343
rect 10376 18312 10425 18340
rect 10376 18300 10382 18312
rect 10413 18309 10425 18312
rect 10459 18309 10471 18343
rect 10413 18303 10471 18309
rect 12069 18343 12127 18349
rect 12069 18309 12081 18343
rect 12115 18340 12127 18343
rect 12434 18340 12440 18352
rect 12115 18312 12440 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 12434 18300 12440 18312
rect 12492 18340 12498 18352
rect 13170 18340 13176 18352
rect 12492 18312 13176 18340
rect 12492 18300 12498 18312
rect 13170 18300 13176 18312
rect 13228 18300 13234 18352
rect 13909 18343 13967 18349
rect 13909 18309 13921 18343
rect 13955 18340 13967 18343
rect 14366 18340 14372 18352
rect 13955 18312 14372 18340
rect 13955 18309 13967 18312
rect 13909 18303 13967 18309
rect 14366 18300 14372 18312
rect 14424 18300 14430 18352
rect 14458 18300 14464 18352
rect 14516 18300 14522 18352
rect 4065 18275 4123 18281
rect 4065 18241 4077 18275
rect 4111 18241 4123 18275
rect 4065 18235 4123 18241
rect 5465 18275 5523 18281
rect 5465 18241 5477 18275
rect 5511 18272 5523 18275
rect 5626 18272 5632 18284
rect 5511 18244 5632 18272
rect 5511 18241 5523 18244
rect 5465 18235 5523 18241
rect 5626 18232 5632 18244
rect 5684 18232 5690 18284
rect 5994 18232 6000 18284
rect 6052 18232 6058 18284
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 8352 18244 8493 18272
rect 8352 18232 8358 18244
rect 8481 18241 8493 18244
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 8570 18232 8576 18284
rect 8628 18272 8634 18284
rect 8737 18275 8795 18281
rect 8737 18272 8749 18275
rect 8628 18244 8749 18272
rect 8628 18232 8634 18244
rect 8737 18241 8749 18244
rect 8783 18241 8795 18275
rect 8737 18235 8795 18241
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 10689 18275 10747 18281
rect 10689 18272 10701 18275
rect 10652 18244 10701 18272
rect 10652 18232 10658 18244
rect 10689 18241 10701 18244
rect 10735 18272 10747 18275
rect 11606 18272 11612 18284
rect 10735 18244 11612 18272
rect 10735 18241 10747 18244
rect 10689 18235 10747 18241
rect 11606 18232 11612 18244
rect 11664 18232 11670 18284
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 11848 18244 12173 18272
rect 11848 18232 11854 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 12526 18232 12532 18284
rect 12584 18232 12590 18284
rect 12986 18232 12992 18284
rect 13044 18232 13050 18284
rect 13265 18275 13323 18281
rect 13265 18241 13277 18275
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 2406 18164 2412 18216
rect 2464 18164 2470 18216
rect 5721 18207 5779 18213
rect 5721 18173 5733 18207
rect 5767 18204 5779 18207
rect 6365 18207 6423 18213
rect 6365 18204 6377 18207
rect 5767 18176 6377 18204
rect 5767 18173 5779 18176
rect 5721 18167 5779 18173
rect 6365 18173 6377 18176
rect 6411 18173 6423 18207
rect 6365 18167 6423 18173
rect 1857 18139 1915 18145
rect 1857 18105 1869 18139
rect 1903 18105 1915 18139
rect 1857 18099 1915 18105
rect 6380 18068 6408 18167
rect 12066 18164 12072 18216
rect 12124 18164 12130 18216
rect 13280 18204 13308 18235
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14737 18275 14795 18281
rect 14737 18272 14749 18275
rect 13872 18244 14749 18272
rect 13872 18232 13878 18244
rect 14737 18241 14749 18244
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 15102 18232 15108 18284
rect 15160 18232 15166 18284
rect 15672 18204 15700 18368
rect 16666 18300 16672 18352
rect 16724 18340 16730 18352
rect 17037 18343 17095 18349
rect 17037 18340 17049 18343
rect 16724 18312 17049 18340
rect 16724 18300 16730 18312
rect 17037 18309 17049 18312
rect 17083 18309 17095 18343
rect 17144 18340 17172 18380
rect 17221 18377 17233 18411
rect 17267 18408 17279 18411
rect 17586 18408 17592 18420
rect 17267 18380 17592 18408
rect 17267 18377 17279 18380
rect 17221 18371 17279 18377
rect 17586 18368 17592 18380
rect 17644 18368 17650 18420
rect 19702 18408 19708 18420
rect 17696 18380 19708 18408
rect 17696 18340 17724 18380
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 17144 18312 17724 18340
rect 17037 18303 17095 18309
rect 18138 18300 18144 18352
rect 18196 18300 18202 18352
rect 18233 18343 18291 18349
rect 18233 18309 18245 18343
rect 18279 18340 18291 18343
rect 21266 18340 21272 18352
rect 18279 18312 21272 18340
rect 18279 18309 18291 18312
rect 18233 18303 18291 18309
rect 21266 18300 21272 18312
rect 21324 18300 21330 18352
rect 17954 18232 17960 18284
rect 18012 18232 18018 18284
rect 18377 18275 18435 18281
rect 18377 18241 18389 18275
rect 18423 18272 18435 18275
rect 18506 18272 18512 18284
rect 18423 18244 18512 18272
rect 18423 18241 18435 18244
rect 18377 18235 18435 18241
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 18690 18232 18696 18284
rect 18748 18232 18754 18284
rect 13280 18176 14228 18204
rect 10134 18096 10140 18148
rect 10192 18096 10198 18148
rect 11238 18096 11244 18148
rect 11296 18136 11302 18148
rect 14200 18145 14228 18176
rect 14292 18176 15700 18204
rect 11609 18139 11667 18145
rect 11609 18136 11621 18139
rect 11296 18108 11621 18136
rect 11296 18096 11302 18108
rect 11609 18105 11621 18108
rect 11655 18105 11667 18139
rect 11609 18099 11667 18105
rect 14185 18139 14243 18145
rect 14185 18105 14197 18139
rect 14231 18105 14243 18139
rect 14185 18099 14243 18105
rect 6730 18068 6736 18080
rect 6380 18040 6736 18068
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 12802 18028 12808 18080
rect 12860 18028 12866 18080
rect 13170 18028 13176 18080
rect 13228 18068 13234 18080
rect 13633 18071 13691 18077
rect 13633 18068 13645 18071
rect 13228 18040 13645 18068
rect 13228 18028 13234 18040
rect 13633 18037 13645 18040
rect 13679 18068 13691 18071
rect 14292 18068 14320 18176
rect 17310 18164 17316 18216
rect 17368 18164 17374 18216
rect 19058 18164 19064 18216
rect 19116 18204 19122 18216
rect 19429 18207 19487 18213
rect 19429 18204 19441 18207
rect 19116 18176 19441 18204
rect 19116 18164 19122 18176
rect 19429 18173 19441 18176
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 20346 18164 20352 18216
rect 20404 18164 20410 18216
rect 20990 18164 20996 18216
rect 21048 18164 21054 18216
rect 16758 18096 16764 18148
rect 16816 18096 16822 18148
rect 18509 18139 18567 18145
rect 18509 18105 18521 18139
rect 18555 18136 18567 18139
rect 20438 18136 20444 18148
rect 18555 18108 20444 18136
rect 18555 18105 18567 18108
rect 18509 18099 18567 18105
rect 20438 18096 20444 18108
rect 20496 18096 20502 18148
rect 13679 18040 14320 18068
rect 13679 18037 13691 18040
rect 13633 18031 13691 18037
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 14424 18040 14933 18068
rect 14424 18028 14430 18040
rect 14921 18037 14933 18040
rect 14967 18037 14979 18071
rect 14921 18031 14979 18037
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 19705 18071 19763 18077
rect 19705 18068 19717 18071
rect 19668 18040 19717 18068
rect 19668 18028 19674 18040
rect 19705 18037 19717 18040
rect 19751 18037 19763 18071
rect 19705 18031 19763 18037
rect 21634 18028 21640 18080
rect 21692 18028 21698 18080
rect 1104 17978 21988 18000
rect 1104 17926 3560 17978
rect 3612 17926 3624 17978
rect 3676 17926 3688 17978
rect 3740 17926 3752 17978
rect 3804 17926 3816 17978
rect 3868 17926 8781 17978
rect 8833 17926 8845 17978
rect 8897 17926 8909 17978
rect 8961 17926 8973 17978
rect 9025 17926 9037 17978
rect 9089 17926 14002 17978
rect 14054 17926 14066 17978
rect 14118 17926 14130 17978
rect 14182 17926 14194 17978
rect 14246 17926 14258 17978
rect 14310 17926 19223 17978
rect 19275 17926 19287 17978
rect 19339 17926 19351 17978
rect 19403 17926 19415 17978
rect 19467 17926 19479 17978
rect 19531 17926 21988 17978
rect 1104 17904 21988 17926
rect 3234 17824 3240 17876
rect 3292 17824 3298 17876
rect 3605 17867 3663 17873
rect 3605 17833 3617 17867
rect 3651 17864 3663 17867
rect 3970 17864 3976 17876
rect 3651 17836 3976 17864
rect 3651 17833 3663 17836
rect 3605 17827 3663 17833
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 4338 17824 4344 17876
rect 4396 17824 4402 17876
rect 5626 17824 5632 17876
rect 5684 17864 5690 17876
rect 6089 17867 6147 17873
rect 6089 17864 6101 17867
rect 5684 17836 6101 17864
rect 5684 17824 5690 17836
rect 6089 17833 6101 17836
rect 6135 17833 6147 17867
rect 6089 17827 6147 17833
rect 6178 17824 6184 17876
rect 6236 17864 6242 17876
rect 6273 17867 6331 17873
rect 6273 17864 6285 17867
rect 6236 17836 6285 17864
rect 6236 17824 6242 17836
rect 6273 17833 6285 17836
rect 6319 17833 6331 17867
rect 6273 17827 6331 17833
rect 9677 17867 9735 17873
rect 9677 17833 9689 17867
rect 9723 17864 9735 17867
rect 9766 17864 9772 17876
rect 9723 17836 9772 17864
rect 9723 17833 9735 17836
rect 9677 17827 9735 17833
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 12345 17867 12403 17873
rect 12345 17833 12357 17867
rect 12391 17864 12403 17867
rect 12526 17864 12532 17876
rect 12391 17836 12532 17864
rect 12391 17833 12403 17836
rect 12345 17827 12403 17833
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12986 17824 12992 17876
rect 13044 17864 13050 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 13044 17836 13185 17864
rect 13044 17824 13050 17836
rect 13173 17833 13185 17836
rect 13219 17833 13231 17867
rect 13173 17827 13231 17833
rect 17681 17867 17739 17873
rect 17681 17833 17693 17867
rect 17727 17864 17739 17867
rect 17954 17864 17960 17876
rect 17727 17836 17960 17864
rect 17727 17833 17739 17836
rect 17681 17827 17739 17833
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 20530 17864 20536 17876
rect 18340 17836 20536 17864
rect 3881 17799 3939 17805
rect 3881 17765 3893 17799
rect 3927 17765 3939 17799
rect 4356 17796 4384 17824
rect 5810 17796 5816 17808
rect 4356 17768 5816 17796
rect 3881 17759 3939 17765
rect 1854 17620 1860 17672
rect 1912 17620 1918 17672
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 3896 17660 3924 17759
rect 5810 17756 5816 17768
rect 5868 17756 5874 17808
rect 6546 17756 6552 17808
rect 6604 17796 6610 17808
rect 6641 17799 6699 17805
rect 6641 17796 6653 17799
rect 6604 17768 6653 17796
rect 6604 17756 6610 17768
rect 6641 17765 6653 17768
rect 6687 17765 6699 17799
rect 6641 17759 6699 17765
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 6880 17768 8156 17796
rect 6880 17756 6886 17768
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17728 4399 17731
rect 4614 17728 4620 17740
rect 4387 17700 4620 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 5994 17728 6000 17740
rect 4724 17700 6000 17728
rect 4724 17660 4752 17700
rect 5994 17688 6000 17700
rect 6052 17688 6058 17740
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 8128 17737 8156 17768
rect 8478 17756 8484 17808
rect 8536 17756 8542 17808
rect 10873 17799 10931 17805
rect 10873 17765 10885 17799
rect 10919 17765 10931 17799
rect 10873 17759 10931 17765
rect 7193 17731 7251 17737
rect 7193 17728 7205 17731
rect 6972 17700 7205 17728
rect 6972 17688 6978 17700
rect 7193 17697 7205 17700
rect 7239 17697 7251 17731
rect 7193 17691 7251 17697
rect 8113 17731 8171 17737
rect 8113 17697 8125 17731
rect 8159 17728 8171 17731
rect 10778 17728 10784 17740
rect 8159 17700 10784 17728
rect 8159 17697 8171 17700
rect 8113 17691 8171 17697
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 3467 17632 3924 17660
rect 4356 17632 4752 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 1946 17552 1952 17604
rect 2004 17592 2010 17604
rect 2102 17595 2160 17601
rect 2102 17592 2114 17595
rect 2004 17564 2114 17592
rect 2004 17552 2010 17564
rect 2102 17561 2114 17564
rect 2148 17561 2160 17595
rect 2102 17555 2160 17561
rect 2866 17552 2872 17604
rect 2924 17592 2930 17604
rect 4356 17601 4384 17632
rect 4798 17620 4804 17672
rect 4856 17620 4862 17672
rect 5534 17620 5540 17672
rect 5592 17620 5598 17672
rect 5718 17620 5724 17672
rect 5776 17620 5782 17672
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 5902 17620 5908 17672
rect 5960 17669 5966 17672
rect 5960 17660 5968 17669
rect 5960 17632 6005 17660
rect 5960 17623 5968 17632
rect 5960 17620 5966 17623
rect 6454 17620 6460 17672
rect 6512 17620 6518 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 6564 17632 7941 17660
rect 4341 17595 4399 17601
rect 4341 17592 4353 17595
rect 2924 17564 4353 17592
rect 2924 17552 2930 17564
rect 4341 17561 4353 17564
rect 4387 17561 4399 17595
rect 4341 17555 4399 17561
rect 4433 17595 4491 17601
rect 4433 17561 4445 17595
rect 4479 17592 4491 17595
rect 4982 17592 4988 17604
rect 4479 17564 4988 17592
rect 4479 17561 4491 17564
rect 4433 17555 4491 17561
rect 4982 17552 4988 17564
rect 5040 17552 5046 17604
rect 6564 17592 6592 17632
rect 7929 17629 7941 17632
rect 7975 17660 7987 17663
rect 8662 17660 8668 17672
rect 7975 17632 8668 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 9858 17620 9864 17672
rect 9916 17660 9922 17672
rect 9953 17663 10011 17669
rect 9953 17660 9965 17663
rect 9916 17632 9965 17660
rect 9916 17620 9922 17632
rect 9953 17629 9965 17632
rect 9999 17629 10011 17663
rect 9953 17623 10011 17629
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17660 10747 17663
rect 10888 17660 10916 17759
rect 11514 17756 11520 17808
rect 11572 17796 11578 17808
rect 13078 17796 13084 17808
rect 11572 17768 13084 17796
rect 11572 17756 11578 17768
rect 13078 17756 13084 17768
rect 13136 17756 13142 17808
rect 15194 17756 15200 17808
rect 15252 17756 15258 17808
rect 15838 17756 15844 17808
rect 15896 17756 15902 17808
rect 17313 17799 17371 17805
rect 17313 17765 17325 17799
rect 17359 17765 17371 17799
rect 17313 17759 17371 17765
rect 11330 17688 11336 17740
rect 11388 17688 11394 17740
rect 11425 17731 11483 17737
rect 11425 17697 11437 17731
rect 11471 17728 11483 17731
rect 13725 17731 13783 17737
rect 13725 17728 13737 17731
rect 11471 17700 13737 17728
rect 11471 17697 11483 17700
rect 11425 17691 11483 17697
rect 13725 17697 13737 17700
rect 13771 17728 13783 17731
rect 13814 17728 13820 17740
rect 13771 17700 13820 17728
rect 13771 17697 13783 17700
rect 13725 17691 13783 17697
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 15856 17728 15884 17756
rect 15396 17700 17172 17728
rect 10735 17632 10916 17660
rect 10735 17629 10747 17632
rect 10689 17623 10747 17629
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 15396 17669 15424 17700
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13688 17632 14197 17660
rect 13688 17620 13694 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 15376 17663 15434 17669
rect 15376 17629 15388 17663
rect 15422 17629 15434 17663
rect 15376 17623 15434 17629
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17660 15807 17663
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15795 17632 15853 17660
rect 15795 17629 15807 17632
rect 15749 17623 15807 17629
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 5276 17564 6592 17592
rect 4706 17484 4712 17536
rect 4764 17524 4770 17536
rect 5276 17524 5304 17564
rect 6914 17552 6920 17604
rect 6972 17552 6978 17604
rect 8202 17592 8208 17604
rect 8036 17564 8208 17592
rect 4764 17496 5304 17524
rect 4764 17484 4770 17496
rect 5350 17484 5356 17536
rect 5408 17524 5414 17536
rect 5445 17527 5503 17533
rect 5445 17524 5457 17527
rect 5408 17496 5457 17524
rect 5408 17484 5414 17496
rect 5445 17493 5457 17496
rect 5491 17493 5503 17527
rect 5445 17487 5503 17493
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 8036 17533 8064 17564
rect 8202 17552 8208 17564
rect 8260 17552 8266 17604
rect 10229 17595 10287 17601
rect 10229 17592 10241 17595
rect 8312 17564 10241 17592
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 5592 17496 7113 17524
rect 5592 17484 5598 17496
rect 7101 17493 7113 17496
rect 7147 17493 7159 17527
rect 7101 17487 7159 17493
rect 8021 17527 8079 17533
rect 8021 17493 8033 17527
rect 8067 17493 8079 17527
rect 8021 17487 8079 17493
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 8312 17524 8340 17564
rect 10229 17561 10241 17564
rect 10275 17592 10287 17595
rect 11333 17595 11391 17601
rect 10275 17564 10640 17592
rect 10275 17561 10287 17564
rect 10229 17555 10287 17561
rect 8168 17496 8340 17524
rect 10137 17527 10195 17533
rect 8168 17484 8174 17496
rect 10137 17493 10149 17527
rect 10183 17524 10195 17527
rect 10318 17524 10324 17536
rect 10183 17496 10324 17524
rect 10183 17493 10195 17496
rect 10137 17487 10195 17493
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 10502 17484 10508 17536
rect 10560 17484 10566 17536
rect 10612 17524 10640 17564
rect 11333 17561 11345 17595
rect 11379 17592 11391 17595
rect 11422 17592 11428 17604
rect 11379 17564 11428 17592
rect 11379 17561 11391 17564
rect 11333 17555 11391 17561
rect 11422 17552 11428 17564
rect 11480 17552 11486 17604
rect 12621 17595 12679 17601
rect 12621 17561 12633 17595
rect 12667 17592 12679 17595
rect 12710 17592 12716 17604
rect 12667 17564 12716 17592
rect 12667 17561 12679 17564
rect 12621 17555 12679 17561
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 12897 17595 12955 17601
rect 12897 17561 12909 17595
rect 12943 17592 12955 17595
rect 13078 17592 13084 17604
rect 12943 17564 13084 17592
rect 12943 17561 12955 17564
rect 12897 17555 12955 17561
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 13446 17552 13452 17604
rect 13504 17552 13510 17604
rect 15010 17552 15016 17604
rect 15068 17552 15074 17604
rect 15470 17552 15476 17604
rect 15528 17552 15534 17604
rect 15562 17552 15568 17604
rect 15620 17552 15626 17604
rect 15654 17552 15660 17604
rect 15712 17592 15718 17604
rect 16408 17592 16436 17623
rect 16666 17620 16672 17672
rect 16724 17660 16730 17672
rect 16761 17663 16819 17669
rect 16761 17660 16773 17663
rect 16724 17632 16773 17660
rect 16724 17620 16730 17632
rect 16761 17629 16773 17632
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 16850 17620 16856 17672
rect 16908 17620 16914 17672
rect 17144 17669 17172 17700
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17660 17187 17663
rect 17218 17660 17224 17672
rect 17175 17632 17224 17660
rect 17175 17629 17187 17632
rect 17129 17623 17187 17629
rect 17218 17620 17224 17632
rect 17276 17620 17282 17672
rect 17328 17660 17356 17759
rect 18340 17737 18368 17836
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 21542 17824 21548 17876
rect 21600 17824 21606 17876
rect 18509 17799 18567 17805
rect 18509 17765 18521 17799
rect 18555 17796 18567 17799
rect 18598 17796 18604 17808
rect 18555 17768 18604 17796
rect 18555 17765 18567 17768
rect 18509 17759 18567 17765
rect 18598 17756 18604 17768
rect 18656 17756 18662 17808
rect 18325 17731 18383 17737
rect 18325 17697 18337 17731
rect 18371 17697 18383 17731
rect 18325 17691 18383 17697
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 19429 17731 19487 17737
rect 19429 17728 19441 17731
rect 18932 17700 19441 17728
rect 18932 17688 18938 17700
rect 19429 17697 19441 17700
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 20165 17731 20223 17737
rect 20165 17728 20177 17731
rect 19852 17700 20177 17728
rect 19852 17688 19858 17700
rect 20165 17697 20177 17700
rect 20211 17697 20223 17731
rect 20165 17691 20223 17697
rect 18506 17660 18512 17672
rect 17328 17632 18512 17660
rect 18506 17620 18512 17632
rect 18564 17660 18570 17672
rect 18641 17663 18699 17669
rect 18641 17660 18653 17663
rect 18564 17632 18653 17660
rect 18564 17620 18570 17632
rect 18641 17629 18653 17632
rect 18687 17629 18699 17663
rect 18641 17623 18699 17629
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17660 18843 17663
rect 18966 17660 18972 17672
rect 18831 17632 18972 17660
rect 18831 17629 18843 17632
rect 18785 17623 18843 17629
rect 18966 17620 18972 17632
rect 19024 17620 19030 17672
rect 19061 17663 19119 17669
rect 19061 17629 19073 17663
rect 19107 17660 19119 17663
rect 19610 17660 19616 17672
rect 19107 17632 19616 17660
rect 19107 17629 19119 17632
rect 19061 17623 19119 17629
rect 19610 17620 19616 17632
rect 19668 17620 19674 17672
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 20990 17660 20996 17672
rect 19751 17632 20996 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 20990 17620 20996 17632
rect 21048 17620 21054 17672
rect 15712 17564 16436 17592
rect 16500 17564 17264 17592
rect 15712 17552 15718 17564
rect 12250 17524 12256 17536
rect 10612 17496 12256 17524
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 12584 17496 12817 17524
rect 12584 17484 12590 17496
rect 12805 17493 12817 17496
rect 12851 17524 12863 17527
rect 13170 17524 13176 17536
rect 12851 17496 13176 17524
rect 12851 17493 12863 17496
rect 12805 17487 12863 17493
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 13538 17484 13544 17536
rect 13596 17524 13602 17536
rect 13633 17527 13691 17533
rect 13633 17524 13645 17527
rect 13596 17496 13645 17524
rect 13596 17484 13602 17496
rect 13633 17493 13645 17496
rect 13679 17493 13691 17527
rect 13633 17487 13691 17493
rect 13722 17484 13728 17536
rect 13780 17524 13786 17536
rect 16500 17524 16528 17564
rect 13780 17496 16528 17524
rect 13780 17484 13786 17496
rect 16574 17484 16580 17536
rect 16632 17484 16638 17536
rect 16942 17484 16948 17536
rect 17000 17524 17006 17536
rect 17037 17527 17095 17533
rect 17037 17524 17049 17527
rect 17000 17496 17049 17524
rect 17000 17484 17006 17496
rect 17037 17493 17049 17496
rect 17083 17493 17095 17527
rect 17236 17524 17264 17564
rect 18138 17552 18144 17604
rect 18196 17592 18202 17604
rect 18877 17595 18935 17601
rect 18877 17592 18889 17595
rect 18196 17564 18889 17592
rect 18196 17552 18202 17564
rect 18877 17561 18889 17564
rect 18923 17561 18935 17595
rect 18877 17555 18935 17561
rect 20432 17595 20490 17601
rect 20432 17561 20444 17595
rect 20478 17592 20490 17595
rect 21082 17592 21088 17604
rect 20478 17564 21088 17592
rect 20478 17561 20490 17564
rect 20432 17555 20490 17561
rect 21082 17552 21088 17564
rect 21140 17552 21146 17604
rect 19521 17527 19579 17533
rect 19521 17524 19533 17527
rect 17236 17496 19533 17524
rect 17037 17487 17095 17493
rect 19521 17493 19533 17496
rect 19567 17524 19579 17527
rect 19794 17524 19800 17536
rect 19567 17496 19800 17524
rect 19567 17493 19579 17496
rect 19521 17487 19579 17493
rect 19794 17484 19800 17496
rect 19852 17484 19858 17536
rect 19999 17527 20057 17533
rect 19999 17493 20011 17527
rect 20045 17524 20057 17527
rect 20254 17524 20260 17536
rect 20045 17496 20260 17524
rect 20045 17493 20057 17496
rect 19999 17487 20057 17493
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 1104 17434 21988 17456
rect 1104 17382 4220 17434
rect 4272 17382 4284 17434
rect 4336 17382 4348 17434
rect 4400 17382 4412 17434
rect 4464 17382 4476 17434
rect 4528 17382 9441 17434
rect 9493 17382 9505 17434
rect 9557 17382 9569 17434
rect 9621 17382 9633 17434
rect 9685 17382 9697 17434
rect 9749 17382 14662 17434
rect 14714 17382 14726 17434
rect 14778 17382 14790 17434
rect 14842 17382 14854 17434
rect 14906 17382 14918 17434
rect 14970 17382 19883 17434
rect 19935 17382 19947 17434
rect 19999 17382 20011 17434
rect 20063 17382 20075 17434
rect 20127 17382 20139 17434
rect 20191 17382 21988 17434
rect 1104 17360 21988 17382
rect 1854 17280 1860 17332
rect 1912 17320 1918 17332
rect 2682 17320 2688 17332
rect 1912 17292 2688 17320
rect 1912 17280 1918 17292
rect 2682 17280 2688 17292
rect 2740 17320 2746 17332
rect 5187 17323 5245 17329
rect 2740 17292 3832 17320
rect 2740 17280 2746 17292
rect 2777 17255 2835 17261
rect 2777 17221 2789 17255
rect 2823 17252 2835 17255
rect 2866 17252 2872 17264
rect 2823 17224 2872 17252
rect 2823 17221 2835 17224
rect 2777 17215 2835 17221
rect 2866 17212 2872 17224
rect 2924 17212 2930 17264
rect 3050 17212 3056 17264
rect 3108 17212 3114 17264
rect 3804 17261 3832 17292
rect 5187 17289 5199 17323
rect 5233 17320 5245 17323
rect 6454 17320 6460 17332
rect 5233 17292 6460 17320
rect 5233 17289 5245 17292
rect 5187 17283 5245 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 7083 17323 7141 17329
rect 7083 17320 7095 17323
rect 6972 17292 7095 17320
rect 6972 17280 6978 17292
rect 7083 17289 7095 17292
rect 7129 17289 7141 17323
rect 8202 17320 8208 17332
rect 7083 17283 7141 17289
rect 7208 17292 8208 17320
rect 3789 17255 3847 17261
rect 3789 17221 3801 17255
rect 3835 17221 3847 17255
rect 3789 17215 3847 17221
rect 4709 17255 4767 17261
rect 4709 17221 4721 17255
rect 4755 17221 4767 17255
rect 4709 17215 4767 17221
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2593 17187 2651 17193
rect 2179 17156 2360 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 1946 17008 1952 17060
rect 2004 17008 2010 17060
rect 2332 17057 2360 17156
rect 2593 17153 2605 17187
rect 2639 17184 2651 17187
rect 3234 17184 3240 17196
rect 2639 17156 3240 17184
rect 2639 17153 2651 17156
rect 2593 17147 2651 17153
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 4724 17184 4752 17215
rect 4890 17212 4896 17264
rect 4948 17252 4954 17264
rect 5629 17255 5687 17261
rect 5629 17252 5641 17255
rect 4948 17224 5641 17252
rect 4948 17212 4954 17224
rect 5629 17221 5641 17224
rect 5675 17221 5687 17255
rect 5629 17215 5687 17221
rect 5994 17212 6000 17264
rect 6052 17252 6058 17264
rect 7208 17252 7236 17292
rect 8202 17280 8208 17292
rect 8260 17320 8266 17332
rect 11241 17323 11299 17329
rect 8260 17292 11100 17320
rect 8260 17280 8266 17292
rect 6052 17224 7236 17252
rect 7561 17255 7619 17261
rect 6052 17212 6058 17224
rect 7561 17221 7573 17255
rect 7607 17252 7619 17255
rect 7926 17252 7932 17264
rect 7607 17224 7932 17252
rect 7607 17221 7619 17224
rect 7561 17215 7619 17221
rect 7926 17212 7932 17224
rect 7984 17212 7990 17264
rect 8018 17212 8024 17264
rect 8076 17212 8082 17264
rect 10128 17255 10186 17261
rect 10128 17221 10140 17255
rect 10174 17252 10186 17255
rect 10502 17252 10508 17264
rect 10174 17224 10508 17252
rect 10174 17221 10186 17224
rect 10128 17215 10186 17221
rect 10502 17212 10508 17224
rect 10560 17212 10566 17264
rect 11072 17252 11100 17292
rect 11241 17289 11253 17323
rect 11287 17320 11299 17323
rect 11422 17320 11428 17332
rect 11287 17292 11428 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 11422 17280 11428 17292
rect 11480 17280 11486 17332
rect 11790 17280 11796 17332
rect 11848 17320 11854 17332
rect 13354 17320 13360 17332
rect 11848 17292 13360 17320
rect 11848 17280 11854 17292
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 13446 17280 13452 17332
rect 13504 17320 13510 17332
rect 14075 17323 14133 17329
rect 14075 17320 14087 17323
rect 13504 17292 14087 17320
rect 13504 17280 13510 17292
rect 14075 17289 14087 17292
rect 14121 17289 14133 17323
rect 14075 17283 14133 17289
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 16301 17323 16359 17329
rect 16301 17320 16313 17323
rect 15528 17292 16313 17320
rect 15528 17280 15534 17292
rect 16301 17289 16313 17292
rect 16347 17320 16359 17323
rect 17954 17320 17960 17332
rect 16347 17292 17960 17320
rect 16347 17289 16359 17292
rect 16301 17283 16359 17289
rect 17954 17280 17960 17292
rect 18012 17280 18018 17332
rect 18966 17280 18972 17332
rect 19024 17320 19030 17332
rect 19429 17323 19487 17329
rect 19429 17320 19441 17323
rect 19024 17292 19441 17320
rect 19024 17280 19030 17292
rect 19429 17289 19441 17292
rect 19475 17289 19487 17323
rect 19429 17283 19487 17289
rect 19702 17280 19708 17332
rect 19760 17320 19766 17332
rect 20162 17320 20168 17332
rect 19760 17292 20168 17320
rect 19760 17280 19766 17292
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 21545 17323 21603 17329
rect 21545 17320 21557 17323
rect 21324 17292 21557 17320
rect 21324 17280 21330 17292
rect 21545 17289 21557 17292
rect 21591 17289 21603 17323
rect 21545 17283 21603 17289
rect 11698 17252 11704 17264
rect 11072 17224 11704 17252
rect 11698 17212 11704 17224
rect 11756 17252 11762 17264
rect 12069 17255 12127 17261
rect 12069 17252 12081 17255
rect 11756 17224 12081 17252
rect 11756 17212 11762 17224
rect 12069 17221 12081 17224
rect 12115 17252 12127 17255
rect 12704 17255 12762 17261
rect 12115 17224 12434 17252
rect 12115 17221 12127 17224
rect 12069 17215 12127 17221
rect 4724 17156 4936 17184
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 4062 17116 4068 17128
rect 2915 17088 4068 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17116 4675 17119
rect 4706 17116 4712 17128
rect 4663 17088 4712 17116
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17085 4859 17119
rect 4908 17116 4936 17156
rect 5350 17144 5356 17196
rect 5408 17144 5414 17196
rect 5534 17144 5540 17196
rect 5592 17144 5598 17196
rect 5773 17187 5831 17193
rect 5773 17153 5785 17187
rect 5819 17184 5831 17187
rect 5902 17184 5908 17196
rect 5819 17156 5908 17184
rect 5819 17153 5831 17156
rect 5773 17147 5831 17153
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 6546 17144 6552 17196
rect 6604 17144 6610 17196
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 7834 17184 7840 17196
rect 6779 17156 7840 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 9582 17144 9588 17196
rect 9640 17184 9646 17196
rect 11790 17184 11796 17196
rect 9640 17156 11796 17184
rect 9640 17144 9646 17156
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 11882 17144 11888 17196
rect 11940 17144 11946 17196
rect 12406 17184 12434 17224
rect 12704 17221 12716 17255
rect 12750 17252 12762 17255
rect 12802 17252 12808 17264
rect 12750 17224 12808 17252
rect 12750 17221 12762 17224
rect 12704 17215 12762 17221
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 13722 17252 13728 17264
rect 13556 17224 13728 17252
rect 13556 17184 13584 17224
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 13814 17212 13820 17264
rect 13872 17252 13878 17264
rect 15194 17261 15200 17264
rect 14553 17255 14611 17261
rect 14553 17252 14565 17255
rect 13872 17224 14565 17252
rect 13872 17212 13878 17224
rect 14553 17221 14565 17224
rect 14599 17221 14611 17255
rect 15188 17252 15200 17261
rect 15155 17224 15200 17252
rect 14553 17215 14611 17221
rect 15188 17215 15200 17224
rect 15194 17212 15200 17215
rect 15252 17212 15258 17264
rect 17034 17212 17040 17264
rect 17092 17252 17098 17264
rect 17221 17255 17279 17261
rect 17221 17252 17233 17255
rect 17092 17224 17233 17252
rect 17092 17212 17098 17224
rect 17221 17221 17233 17224
rect 17267 17221 17279 17255
rect 17221 17215 17279 17221
rect 17402 17212 17408 17264
rect 17460 17252 17466 17264
rect 19058 17252 19064 17264
rect 17460 17224 19064 17252
rect 17460 17212 17466 17224
rect 12406 17156 13584 17184
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 14921 17187 14979 17193
rect 14921 17184 14933 17187
rect 13688 17156 14933 17184
rect 13688 17144 13694 17156
rect 14921 17153 14933 17156
rect 14967 17153 14979 17187
rect 17310 17184 17316 17196
rect 14921 17147 14979 17153
rect 15028 17156 17316 17184
rect 6822 17116 6828 17128
rect 4908 17088 6828 17116
rect 4801 17079 4859 17085
rect 2317 17051 2375 17057
rect 2317 17017 2329 17051
rect 2363 17017 2375 17051
rect 4816 17048 4844 17079
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 7558 17076 7564 17128
rect 7616 17076 7622 17128
rect 7653 17119 7711 17125
rect 7653 17085 7665 17119
rect 7699 17116 7711 17119
rect 8110 17116 8116 17128
rect 7699 17088 8116 17116
rect 7699 17085 7711 17088
rect 7653 17079 7711 17085
rect 8110 17076 8116 17088
rect 8168 17076 8174 17128
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17116 8907 17119
rect 9306 17116 9312 17128
rect 8895 17088 9312 17116
rect 8895 17085 8907 17088
rect 8849 17079 8907 17085
rect 9306 17076 9312 17088
rect 9364 17116 9370 17128
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 9364 17088 9873 17116
rect 9364 17076 9370 17088
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 9861 17079 9919 17085
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11606 17116 11612 17128
rect 11112 17088 11612 17116
rect 11112 17076 11118 17088
rect 11606 17076 11612 17088
rect 11664 17116 11670 17128
rect 12161 17119 12219 17125
rect 12161 17116 12173 17119
rect 11664 17088 12173 17116
rect 11664 17076 11670 17088
rect 12161 17085 12173 17088
rect 12207 17085 12219 17119
rect 12161 17079 12219 17085
rect 12434 17076 12440 17128
rect 12492 17076 12498 17128
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17085 14611 17119
rect 14553 17079 14611 17085
rect 6270 17048 6276 17060
rect 4816 17020 6276 17048
rect 2317 17011 2375 17017
rect 6270 17008 6276 17020
rect 6328 17008 6334 17060
rect 6546 17008 6552 17060
rect 6604 17048 6610 17060
rect 9582 17048 9588 17060
rect 6604 17020 9588 17048
rect 6604 17008 6610 17020
rect 9582 17008 9588 17020
rect 9640 17008 9646 17060
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 13817 17051 13875 17057
rect 13817 17048 13829 17051
rect 13596 17020 13829 17048
rect 13596 17008 13602 17020
rect 13817 17017 13829 17020
rect 13863 17017 13875 17051
rect 13817 17011 13875 17017
rect 14568 16992 14596 17079
rect 14642 17076 14648 17128
rect 14700 17116 14706 17128
rect 15028 17116 15056 17156
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 17865 17187 17923 17193
rect 17865 17153 17877 17187
rect 17911 17184 17923 17187
rect 17954 17184 17960 17196
rect 17911 17156 17960 17184
rect 17911 17153 17923 17156
rect 17865 17147 17923 17153
rect 17954 17144 17960 17156
rect 18012 17144 18018 17196
rect 18064 17193 18092 17224
rect 19058 17212 19064 17224
rect 19116 17212 19122 17264
rect 21450 17252 21456 17264
rect 19812 17224 21456 17252
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18316 17187 18374 17193
rect 18316 17153 18328 17187
rect 18362 17184 18374 17187
rect 18598 17184 18604 17196
rect 18362 17156 18604 17184
rect 18362 17153 18374 17156
rect 18316 17147 18374 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 19812 17193 19840 17224
rect 21450 17212 21456 17224
rect 21508 17212 21514 17264
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17153 19855 17187
rect 19797 17147 19855 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20254 17184 20260 17196
rect 20119 17156 20260 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 20254 17144 20260 17156
rect 20312 17144 20318 17196
rect 20438 17193 20444 17196
rect 20432 17184 20444 17193
rect 20399 17156 20444 17184
rect 20432 17147 20444 17156
rect 20438 17144 20444 17147
rect 20496 17144 20502 17196
rect 14700 17088 15056 17116
rect 14700 17076 14706 17088
rect 15930 17076 15936 17128
rect 15988 17116 15994 17128
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 15988 17088 17141 17116
rect 15988 17076 15994 17088
rect 17129 17085 17141 17088
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 19116 17088 20177 17116
rect 19116 17076 19122 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 5905 16983 5963 16989
rect 5905 16980 5917 16983
rect 5592 16952 5917 16980
rect 5592 16940 5598 16952
rect 5905 16949 5917 16952
rect 5951 16949 5963 16983
rect 5905 16943 5963 16949
rect 6365 16983 6423 16989
rect 6365 16949 6377 16983
rect 6411 16980 6423 16983
rect 6454 16980 6460 16992
rect 6411 16952 6460 16980
rect 6411 16949 6423 16952
rect 6365 16943 6423 16949
rect 6454 16940 6460 16952
rect 6512 16940 6518 16992
rect 6914 16940 6920 16992
rect 6972 16940 6978 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 11609 16983 11667 16989
rect 11609 16980 11621 16983
rect 9732 16952 11621 16980
rect 9732 16940 9738 16952
rect 11609 16949 11621 16952
rect 11655 16949 11667 16983
rect 11609 16943 11667 16949
rect 12250 16940 12256 16992
rect 12308 16980 12314 16992
rect 14458 16980 14464 16992
rect 12308 16952 14464 16980
rect 12308 16940 12314 16952
rect 14458 16940 14464 16952
rect 14516 16940 14522 16992
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 15654 16980 15660 16992
rect 14608 16952 15660 16980
rect 14608 16940 14614 16952
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 16758 16940 16764 16992
rect 16816 16940 16822 16992
rect 17678 16940 17684 16992
rect 17736 16940 17742 16992
rect 19610 16940 19616 16992
rect 19668 16940 19674 16992
rect 19702 16940 19708 16992
rect 19760 16980 19766 16992
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 19760 16952 19901 16980
rect 19760 16940 19766 16952
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 1104 16890 21988 16912
rect 1104 16838 3560 16890
rect 3612 16838 3624 16890
rect 3676 16838 3688 16890
rect 3740 16838 3752 16890
rect 3804 16838 3816 16890
rect 3868 16838 8781 16890
rect 8833 16838 8845 16890
rect 8897 16838 8909 16890
rect 8961 16838 8973 16890
rect 9025 16838 9037 16890
rect 9089 16838 14002 16890
rect 14054 16838 14066 16890
rect 14118 16838 14130 16890
rect 14182 16838 14194 16890
rect 14246 16838 14258 16890
rect 14310 16838 19223 16890
rect 19275 16838 19287 16890
rect 19339 16838 19351 16890
rect 19403 16838 19415 16890
rect 19467 16838 19479 16890
rect 19531 16838 21988 16890
rect 1104 16816 21988 16838
rect 5350 16736 5356 16788
rect 5408 16736 5414 16788
rect 6546 16776 6552 16788
rect 5828 16748 6552 16776
rect 5828 16708 5856 16748
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 9306 16776 9312 16788
rect 6840 16748 9312 16776
rect 4264 16680 5856 16708
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4264 16640 4292 16680
rect 4120 16612 4292 16640
rect 4120 16600 4126 16612
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16572 1455 16575
rect 2682 16572 2688 16584
rect 1443 16544 2688 16572
rect 1443 16541 1455 16544
rect 1397 16535 1455 16541
rect 2682 16532 2688 16544
rect 2740 16532 2746 16584
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3605 16575 3663 16581
rect 3191 16544 3556 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 1670 16513 1676 16516
rect 1664 16467 1676 16513
rect 1670 16464 1676 16467
rect 1728 16464 1734 16516
rect 2774 16396 2780 16448
rect 2832 16396 2838 16448
rect 2958 16396 2964 16448
rect 3016 16396 3022 16448
rect 3418 16396 3424 16448
rect 3476 16396 3482 16448
rect 3528 16436 3556 16544
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 3878 16572 3884 16584
rect 3651 16544 3884 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4264 16572 4292 16612
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 4614 16640 4620 16652
rect 4387 16612 4620 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 4706 16600 4712 16652
rect 4764 16640 4770 16652
rect 5626 16640 5632 16652
rect 4764 16612 5632 16640
rect 4764 16600 4770 16612
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 6730 16600 6736 16652
rect 6788 16640 6794 16652
rect 6840 16649 6868 16748
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 9582 16736 9588 16788
rect 9640 16776 9646 16788
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 9640 16748 10057 16776
rect 9640 16736 9646 16748
rect 10045 16745 10057 16748
rect 10091 16745 10103 16779
rect 11514 16776 11520 16788
rect 10045 16739 10103 16745
rect 10428 16748 11520 16776
rect 7926 16668 7932 16720
rect 7984 16708 7990 16720
rect 8205 16711 8263 16717
rect 8205 16708 8217 16711
rect 7984 16680 8217 16708
rect 7984 16668 7990 16680
rect 8205 16677 8217 16680
rect 8251 16677 8263 16711
rect 8205 16671 8263 16677
rect 8386 16668 8392 16720
rect 8444 16708 8450 16720
rect 9217 16711 9275 16717
rect 9217 16708 9229 16711
rect 8444 16680 9229 16708
rect 8444 16668 8450 16680
rect 9217 16677 9229 16680
rect 9263 16708 9275 16711
rect 10428 16708 10456 16748
rect 11514 16736 11520 16748
rect 11572 16736 11578 16788
rect 11793 16779 11851 16785
rect 11793 16745 11805 16779
rect 11839 16776 11851 16779
rect 11882 16776 11888 16788
rect 11839 16748 11888 16776
rect 11839 16745 11851 16748
rect 11793 16739 11851 16745
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 13814 16736 13820 16788
rect 13872 16736 13878 16788
rect 14108 16748 15884 16776
rect 9263 16680 10456 16708
rect 9263 16677 9275 16680
rect 9217 16671 9275 16677
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 6788 16612 6837 16640
rect 6788 16600 6794 16612
rect 6825 16609 6837 16612
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 9306 16600 9312 16652
rect 9364 16640 9370 16652
rect 14108 16649 14136 16748
rect 15473 16711 15531 16717
rect 15473 16677 15485 16711
rect 15519 16708 15531 16711
rect 15654 16708 15660 16720
rect 15519 16680 15660 16708
rect 15519 16677 15531 16680
rect 15473 16671 15531 16677
rect 15654 16668 15660 16680
rect 15712 16668 15718 16720
rect 15856 16649 15884 16748
rect 20530 16736 20536 16788
rect 20588 16776 20594 16788
rect 20625 16779 20683 16785
rect 20625 16776 20637 16779
rect 20588 16748 20637 16776
rect 20588 16736 20594 16748
rect 20625 16745 20637 16748
rect 20671 16745 20683 16779
rect 20625 16739 20683 16745
rect 10413 16643 10471 16649
rect 10413 16640 10425 16643
rect 9364 16612 10425 16640
rect 9364 16600 9370 16612
rect 10413 16609 10425 16612
rect 10459 16609 10471 16643
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 10413 16603 10471 16609
rect 13648 16612 14105 16640
rect 13648 16584 13676 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 15841 16643 15899 16649
rect 15841 16609 15853 16643
rect 15887 16609 15899 16643
rect 15841 16603 15899 16609
rect 17402 16600 17408 16652
rect 17460 16600 17466 16652
rect 19058 16600 19064 16652
rect 19116 16640 19122 16652
rect 19245 16643 19303 16649
rect 19245 16640 19257 16643
rect 19116 16612 19257 16640
rect 19116 16600 19122 16612
rect 19245 16609 19257 16612
rect 19291 16640 19303 16643
rect 20640 16640 20668 16739
rect 21450 16736 21456 16788
rect 21508 16736 21514 16788
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 19291 16612 19380 16640
rect 20640 16612 21005 16640
rect 19291 16609 19303 16612
rect 19245 16603 19303 16609
rect 19352 16584 19380 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 4433 16575 4491 16581
rect 4433 16572 4445 16575
rect 4264 16544 4445 16572
rect 4433 16541 4445 16544
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 6454 16532 6460 16584
rect 6512 16581 6518 16584
rect 6512 16572 6524 16581
rect 6512 16544 6557 16572
rect 6512 16535 6524 16544
rect 6512 16532 6518 16535
rect 6914 16532 6920 16584
rect 6972 16572 6978 16584
rect 7081 16575 7139 16581
rect 7081 16572 7093 16575
rect 6972 16544 7093 16572
rect 6972 16532 6978 16544
rect 7081 16541 7093 16544
rect 7127 16541 7139 16575
rect 7081 16535 7139 16541
rect 8478 16532 8484 16584
rect 8536 16532 8542 16584
rect 8662 16532 8668 16584
rect 8720 16572 8726 16584
rect 9033 16575 9091 16581
rect 9033 16572 9045 16575
rect 8720 16544 9045 16572
rect 8720 16532 8726 16544
rect 9033 16541 9045 16544
rect 9079 16541 9091 16575
rect 9033 16535 9091 16541
rect 9585 16575 9643 16581
rect 9585 16541 9597 16575
rect 9631 16572 9643 16575
rect 9674 16572 9680 16584
rect 9631 16544 9680 16572
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 10669 16575 10727 16581
rect 10669 16572 10681 16575
rect 9876 16544 10681 16572
rect 3863 16439 3921 16445
rect 3863 16436 3875 16439
rect 3528 16408 3875 16436
rect 3863 16405 3875 16408
rect 3909 16405 3921 16439
rect 3863 16399 3921 16405
rect 4341 16439 4399 16445
rect 4341 16405 4353 16439
rect 4387 16436 4399 16439
rect 4706 16436 4712 16448
rect 4387 16408 4712 16436
rect 4387 16405 4399 16408
rect 4341 16399 4399 16405
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 8665 16439 8723 16445
rect 8665 16405 8677 16439
rect 8711 16436 8723 16439
rect 8938 16436 8944 16448
rect 8711 16408 8944 16436
rect 8711 16405 8723 16408
rect 8665 16399 8723 16405
rect 8938 16396 8944 16408
rect 8996 16396 9002 16448
rect 9769 16439 9827 16445
rect 9769 16405 9781 16439
rect 9815 16436 9827 16439
rect 9876 16436 9904 16544
rect 10669 16541 10681 16544
rect 10715 16541 10727 16575
rect 10669 16535 10727 16541
rect 12158 16532 12164 16584
rect 12216 16532 12222 16584
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 13630 16572 13636 16584
rect 12492 16544 13636 16572
rect 12492 16532 12498 16544
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 14366 16581 14372 16584
rect 14360 16572 14372 16581
rect 14327 16544 14372 16572
rect 14360 16535 14372 16544
rect 14366 16532 14372 16535
rect 14424 16532 14430 16584
rect 16108 16575 16166 16581
rect 16108 16541 16120 16575
rect 16154 16572 16166 16575
rect 16574 16572 16580 16584
rect 16154 16544 16580 16572
rect 16154 16541 16166 16544
rect 16108 16535 16166 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 17678 16581 17684 16584
rect 17672 16572 17684 16581
rect 17639 16544 17684 16572
rect 17672 16535 17684 16544
rect 17678 16532 17684 16535
rect 17736 16532 17742 16584
rect 19334 16532 19340 16584
rect 19392 16532 19398 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 19444 16544 20913 16572
rect 9950 16464 9956 16516
rect 10008 16464 10014 16516
rect 12682 16507 12740 16513
rect 12682 16504 12694 16507
rect 12360 16476 12694 16504
rect 12360 16445 12388 16476
rect 12682 16473 12694 16476
rect 12728 16473 12740 16507
rect 12682 16467 12740 16473
rect 18874 16464 18880 16516
rect 18932 16504 18938 16516
rect 19444 16504 19472 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 18932 16476 19472 16504
rect 19512 16507 19570 16513
rect 18932 16464 18938 16476
rect 19512 16473 19524 16507
rect 19558 16504 19570 16507
rect 19610 16504 19616 16516
rect 19558 16476 19616 16504
rect 19558 16473 19570 16476
rect 19512 16467 19570 16473
rect 19610 16464 19616 16476
rect 19668 16464 19674 16516
rect 9815 16408 9904 16436
rect 12345 16439 12403 16445
rect 9815 16405 9827 16408
rect 9769 16399 9827 16405
rect 12345 16405 12357 16439
rect 12391 16405 12403 16439
rect 12345 16399 12403 16405
rect 16574 16396 16580 16448
rect 16632 16436 16638 16448
rect 17218 16436 17224 16448
rect 16632 16408 17224 16436
rect 16632 16396 16638 16408
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 18598 16396 18604 16448
rect 18656 16436 18662 16448
rect 18785 16439 18843 16445
rect 18785 16436 18797 16439
rect 18656 16408 18797 16436
rect 18656 16396 18662 16408
rect 18785 16405 18797 16408
rect 18831 16436 18843 16439
rect 20346 16436 20352 16448
rect 18831 16408 20352 16436
rect 18831 16405 18843 16408
rect 18785 16399 18843 16405
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 20993 16439 21051 16445
rect 20993 16436 21005 16439
rect 20956 16408 21005 16436
rect 20956 16396 20962 16408
rect 20993 16405 21005 16408
rect 21039 16405 21051 16439
rect 20993 16399 21051 16405
rect 1104 16346 21988 16368
rect 1104 16294 4220 16346
rect 4272 16294 4284 16346
rect 4336 16294 4348 16346
rect 4400 16294 4412 16346
rect 4464 16294 4476 16346
rect 4528 16294 9441 16346
rect 9493 16294 9505 16346
rect 9557 16294 9569 16346
rect 9621 16294 9633 16346
rect 9685 16294 9697 16346
rect 9749 16294 14662 16346
rect 14714 16294 14726 16346
rect 14778 16294 14790 16346
rect 14842 16294 14854 16346
rect 14906 16294 14918 16346
rect 14970 16294 19883 16346
rect 19935 16294 19947 16346
rect 19999 16294 20011 16346
rect 20063 16294 20075 16346
rect 20127 16294 20139 16346
rect 20191 16294 21988 16346
rect 1104 16272 21988 16294
rect 1670 16192 1676 16244
rect 1728 16192 1734 16244
rect 2501 16235 2559 16241
rect 2501 16201 2513 16235
rect 2547 16232 2559 16235
rect 2774 16232 2780 16244
rect 2547 16204 2780 16232
rect 2547 16201 2559 16204
rect 2501 16195 2559 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4246 16232 4252 16244
rect 4203 16204 4252 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4246 16192 4252 16204
rect 4304 16232 4310 16244
rect 4798 16232 4804 16244
rect 4304 16204 4804 16232
rect 4304 16192 4310 16204
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 7616 16204 7757 16232
rect 7616 16192 7622 16204
rect 7745 16201 7757 16204
rect 7791 16201 7803 16235
rect 7745 16195 7803 16201
rect 8478 16192 8484 16244
rect 8536 16232 8542 16244
rect 9858 16232 9864 16244
rect 8536 16204 9864 16232
rect 8536 16192 8542 16204
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 10321 16235 10379 16241
rect 10321 16201 10333 16235
rect 10367 16232 10379 16235
rect 10367 16204 11284 16232
rect 10367 16201 10379 16204
rect 10321 16195 10379 16201
rect 3044 16167 3102 16173
rect 3044 16133 3056 16167
rect 3090 16164 3102 16167
rect 3418 16164 3424 16176
rect 3090 16136 3424 16164
rect 3090 16133 3102 16136
rect 3044 16127 3102 16133
rect 3418 16124 3424 16136
rect 3476 16124 3482 16176
rect 5534 16124 5540 16176
rect 5592 16173 5598 16176
rect 5592 16164 5604 16173
rect 6730 16164 6736 16176
rect 5592 16136 5637 16164
rect 6380 16136 6736 16164
rect 5592 16127 5604 16136
rect 5592 16124 5598 16127
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 2317 16099 2375 16105
rect 1903 16068 2084 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 2056 15969 2084 16068
rect 2317 16065 2329 16099
rect 2363 16096 2375 16099
rect 2866 16096 2872 16108
rect 2363 16068 2872 16096
rect 2363 16065 2375 16068
rect 2317 16059 2375 16065
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5776 16068 5825 16096
rect 5776 16056 5782 16068
rect 5813 16065 5825 16068
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5902 16056 5908 16108
rect 5960 16056 5966 16108
rect 6380 16105 6408 16136
rect 6730 16124 6736 16136
rect 6788 16124 6794 16176
rect 7926 16124 7932 16176
rect 7984 16164 7990 16176
rect 8297 16167 8355 16173
rect 8297 16164 8309 16167
rect 7984 16136 8309 16164
rect 7984 16124 7990 16136
rect 8297 16133 8309 16136
rect 8343 16133 8355 16167
rect 9306 16164 9312 16176
rect 8297 16127 8355 16133
rect 8956 16136 9312 16164
rect 8956 16105 8984 16136
rect 9306 16124 9312 16136
rect 9364 16124 9370 16176
rect 11256 16173 11284 16204
rect 11882 16192 11888 16244
rect 11940 16232 11946 16244
rect 12069 16235 12127 16241
rect 12069 16232 12081 16235
rect 11940 16204 12081 16232
rect 11940 16192 11946 16204
rect 12069 16201 12081 16204
rect 12115 16201 12127 16235
rect 12069 16195 12127 16201
rect 12805 16235 12863 16241
rect 12805 16201 12817 16235
rect 12851 16232 12863 16235
rect 16758 16232 16764 16244
rect 12851 16204 13584 16232
rect 12851 16201 12863 16204
rect 12805 16195 12863 16201
rect 11241 16167 11299 16173
rect 11241 16133 11253 16167
rect 11287 16164 11299 16167
rect 12161 16167 12219 16173
rect 11287 16136 11928 16164
rect 11287 16133 11299 16136
rect 11241 16127 11299 16133
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16065 6423 16099
rect 6621 16099 6679 16105
rect 6621 16096 6633 16099
rect 6365 16059 6423 16065
rect 6472 16068 6633 16096
rect 2406 15988 2412 16040
rect 2464 16028 2470 16040
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 2464 16000 2605 16028
rect 2464 15988 2470 16000
rect 2593 15997 2605 16000
rect 2639 15997 2651 16031
rect 2593 15991 2651 15997
rect 2041 15963 2099 15969
rect 2041 15929 2053 15963
rect 2087 15929 2099 15963
rect 2041 15923 2099 15929
rect 2608 15892 2636 15991
rect 2682 15988 2688 16040
rect 2740 16028 2746 16040
rect 2777 16031 2835 16037
rect 2777 16028 2789 16031
rect 2740 16000 2789 16028
rect 2740 15988 2746 16000
rect 2777 15997 2789 16000
rect 2823 15997 2835 16031
rect 6472 16028 6500 16068
rect 6621 16065 6633 16068
rect 6667 16065 6679 16099
rect 6621 16059 6679 16065
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16065 8999 16099
rect 8941 16059 8999 16065
rect 9030 16056 9036 16108
rect 9088 16096 9094 16108
rect 11900 16105 11928 16136
rect 12161 16133 12173 16167
rect 12207 16164 12219 16167
rect 12250 16164 12256 16176
rect 12207 16136 12256 16164
rect 12207 16133 12219 16136
rect 12161 16127 12219 16133
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 13446 16124 13452 16176
rect 13504 16124 13510 16176
rect 13556 16164 13584 16204
rect 16132 16204 16764 16232
rect 13970 16167 14028 16173
rect 13970 16164 13982 16167
rect 13556 16136 13982 16164
rect 13970 16133 13982 16136
rect 14016 16133 14028 16167
rect 13970 16127 14028 16133
rect 15838 16124 15844 16176
rect 15896 16124 15902 16176
rect 16132 16173 16160 16204
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 20990 16232 20996 16244
rect 20855 16204 20996 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 15933 16167 15991 16173
rect 15933 16133 15945 16167
rect 15979 16133 15991 16167
rect 15933 16127 15991 16133
rect 16117 16167 16175 16173
rect 16117 16133 16129 16167
rect 16163 16133 16175 16167
rect 17218 16164 17224 16176
rect 16117 16127 16175 16133
rect 16684 16136 17224 16164
rect 9197 16099 9255 16105
rect 9197 16096 9209 16099
rect 9088 16068 9209 16096
rect 9088 16056 9094 16068
rect 9197 16065 9209 16068
rect 9243 16065 9255 16099
rect 9197 16059 9255 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16096 11943 16099
rect 12066 16096 12072 16108
rect 11931 16068 12072 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 12066 16056 12072 16068
rect 12124 16056 12130 16108
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 12667 16068 13032 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 2777 15991 2835 15997
rect 6104 16000 6500 16028
rect 8573 16031 8631 16037
rect 4798 15960 4804 15972
rect 4356 15932 4804 15960
rect 4356 15892 4384 15932
rect 4798 15920 4804 15932
rect 4856 15920 4862 15972
rect 6104 15969 6132 16000
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 8619 16000 8984 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 6089 15963 6147 15969
rect 6089 15929 6101 15963
rect 6135 15929 6147 15963
rect 6089 15923 6147 15929
rect 7834 15920 7840 15972
rect 7892 15960 7898 15972
rect 8021 15963 8079 15969
rect 8021 15960 8033 15963
rect 7892 15932 8033 15960
rect 7892 15920 7898 15932
rect 8021 15929 8033 15932
rect 8067 15929 8079 15963
rect 8021 15923 8079 15929
rect 2608 15864 4384 15892
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 4890 15892 4896 15904
rect 4479 15864 4896 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 8956 15892 8984 16000
rect 11330 15920 11336 15972
rect 11388 15960 11394 15972
rect 13004 15969 13032 16068
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 13136 16068 13553 16096
rect 13136 16056 13142 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 15470 16056 15476 16108
rect 15528 16056 15534 16108
rect 15948 16096 15976 16127
rect 16574 16096 16580 16108
rect 15948 16068 16580 16096
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 16684 16105 16712 16136
rect 17218 16124 17224 16136
rect 17276 16164 17282 16176
rect 17402 16164 17408 16176
rect 17276 16136 17408 16164
rect 17276 16124 17282 16136
rect 17402 16124 17408 16136
rect 17460 16124 17466 16176
rect 18598 16124 18604 16176
rect 18656 16124 18662 16176
rect 18785 16167 18843 16173
rect 18785 16133 18797 16167
rect 18831 16133 18843 16167
rect 19794 16164 19800 16176
rect 18785 16127 18843 16133
rect 19444 16136 19800 16164
rect 16942 16105 16948 16108
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 16936 16059 16948 16105
rect 17000 16096 17006 16108
rect 17000 16068 17036 16096
rect 16942 16056 16948 16059
rect 17000 16056 17006 16068
rect 18046 16056 18052 16108
rect 18104 16096 18110 16108
rect 18800 16096 18828 16127
rect 18104 16068 18828 16096
rect 18104 16056 18110 16068
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19444 16105 19472 16136
rect 19794 16124 19800 16136
rect 19852 16124 19858 16176
rect 21361 16167 21419 16173
rect 21361 16133 21373 16167
rect 21407 16164 21419 16167
rect 21542 16164 21548 16176
rect 21407 16136 21548 16164
rect 21407 16133 21419 16136
rect 21361 16127 21419 16133
rect 21542 16124 21548 16136
rect 21600 16124 21606 16176
rect 19429 16099 19487 16105
rect 19429 16096 19441 16099
rect 19392 16068 19441 16096
rect 19392 16056 19398 16068
rect 19429 16065 19441 16068
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 19696 16099 19754 16105
rect 19696 16096 19708 16099
rect 19576 16068 19708 16096
rect 19576 16056 19582 16068
rect 19696 16065 19708 16068
rect 19742 16065 19754 16099
rect 19696 16059 19754 16065
rect 21174 16056 21180 16108
rect 21232 16105 21238 16108
rect 21232 16099 21275 16105
rect 21263 16065 21275 16099
rect 21232 16059 21275 16065
rect 21232 16056 21238 16059
rect 21450 16056 21456 16108
rect 21508 16056 21514 16108
rect 21634 16056 21640 16108
rect 21692 16056 21698 16108
rect 13449 16031 13507 16037
rect 13449 15997 13461 16031
rect 13495 16028 13507 16031
rect 13495 16000 13584 16028
rect 13495 15997 13507 16000
rect 13449 15991 13507 15997
rect 11609 15963 11667 15969
rect 11609 15960 11621 15963
rect 11388 15932 11621 15960
rect 11388 15920 11394 15932
rect 11609 15929 11621 15932
rect 11655 15929 11667 15963
rect 11609 15923 11667 15929
rect 12989 15963 13047 15969
rect 12989 15929 13001 15963
rect 13035 15929 13047 15963
rect 12989 15923 13047 15929
rect 10870 15892 10876 15904
rect 8956 15864 10876 15892
rect 10870 15852 10876 15864
rect 10928 15892 10934 15904
rect 11054 15892 11060 15904
rect 10928 15864 11060 15892
rect 10928 15852 10934 15864
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 11698 15892 11704 15904
rect 11195 15864 11704 15892
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 13556 15892 13584 16000
rect 13630 15988 13636 16040
rect 13688 16028 13694 16040
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 13688 16000 13737 16028
rect 13688 15988 13694 16000
rect 13725 15997 13737 16000
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 18874 15988 18880 16040
rect 18932 15988 18938 16040
rect 15105 15963 15163 15969
rect 15105 15929 15117 15963
rect 15151 15960 15163 15963
rect 15930 15960 15936 15972
rect 15151 15932 15936 15960
rect 15151 15929 15163 15932
rect 15105 15923 15163 15929
rect 15930 15920 15936 15932
rect 15988 15920 15994 15972
rect 16393 15963 16451 15969
rect 16393 15929 16405 15963
rect 16439 15960 16451 15963
rect 16666 15960 16672 15972
rect 16439 15932 16672 15960
rect 16439 15929 16451 15932
rect 16393 15923 16451 15929
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 17954 15920 17960 15972
rect 18012 15960 18018 15972
rect 18325 15963 18383 15969
rect 18325 15960 18337 15963
rect 18012 15932 18337 15960
rect 18012 15920 18018 15932
rect 18325 15929 18337 15932
rect 18371 15929 18383 15963
rect 18325 15923 18383 15929
rect 21082 15920 21088 15972
rect 21140 15920 21146 15972
rect 14458 15892 14464 15904
rect 13556 15864 14464 15892
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 15654 15852 15660 15904
rect 15712 15852 15718 15904
rect 17034 15852 17040 15904
rect 17092 15892 17098 15904
rect 18049 15895 18107 15901
rect 18049 15892 18061 15895
rect 17092 15864 18061 15892
rect 17092 15852 17098 15864
rect 18049 15861 18061 15864
rect 18095 15861 18107 15895
rect 18049 15855 18107 15861
rect 1104 15802 21988 15824
rect 1104 15750 3560 15802
rect 3612 15750 3624 15802
rect 3676 15750 3688 15802
rect 3740 15750 3752 15802
rect 3804 15750 3816 15802
rect 3868 15750 8781 15802
rect 8833 15750 8845 15802
rect 8897 15750 8909 15802
rect 8961 15750 8973 15802
rect 9025 15750 9037 15802
rect 9089 15750 14002 15802
rect 14054 15750 14066 15802
rect 14118 15750 14130 15802
rect 14182 15750 14194 15802
rect 14246 15750 14258 15802
rect 14310 15750 19223 15802
rect 19275 15750 19287 15802
rect 19339 15750 19351 15802
rect 19403 15750 19415 15802
rect 19467 15750 19479 15802
rect 19531 15750 21988 15802
rect 1104 15728 21988 15750
rect 3878 15648 3884 15700
rect 3936 15648 3942 15700
rect 5902 15648 5908 15700
rect 5960 15688 5966 15700
rect 6089 15691 6147 15697
rect 6089 15688 6101 15691
rect 5960 15660 6101 15688
rect 5960 15648 5966 15660
rect 6089 15657 6101 15660
rect 6135 15657 6147 15691
rect 7285 15691 7343 15697
rect 7285 15688 7297 15691
rect 6089 15651 6147 15657
rect 7116 15660 7297 15688
rect 3513 15623 3571 15629
rect 3513 15589 3525 15623
rect 3559 15620 3571 15623
rect 4614 15620 4620 15632
rect 3559 15592 4620 15620
rect 3559 15589 3571 15592
rect 3513 15583 3571 15589
rect 4614 15580 4620 15592
rect 4672 15580 4678 15632
rect 4246 15512 4252 15564
rect 4304 15512 4310 15564
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4982 15552 4988 15564
rect 4479 15524 4988 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15552 5595 15555
rect 5626 15552 5632 15564
rect 5583 15524 5632 15552
rect 5583 15521 5595 15524
rect 5537 15515 5595 15521
rect 5626 15512 5632 15524
rect 5684 15512 5690 15564
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15484 2191 15487
rect 2682 15484 2688 15496
rect 2179 15456 2688 15484
rect 2179 15453 2191 15456
rect 2133 15447 2191 15453
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 5994 15484 6000 15496
rect 5859 15456 6000 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 2400 15419 2458 15425
rect 2400 15385 2412 15419
rect 2446 15416 2458 15419
rect 2958 15416 2964 15428
rect 2446 15388 2964 15416
rect 2446 15385 2458 15388
rect 2400 15379 2458 15385
rect 2958 15376 2964 15388
rect 3016 15376 3022 15428
rect 4341 15419 4399 15425
rect 4341 15385 4353 15419
rect 4387 15416 4399 15419
rect 4706 15416 4712 15428
rect 4387 15388 4712 15416
rect 4387 15385 4399 15388
rect 4341 15379 4399 15385
rect 4706 15376 4712 15388
rect 4764 15416 4770 15428
rect 5629 15419 5687 15425
rect 5629 15416 5641 15419
rect 4764 15388 5641 15416
rect 4764 15376 4770 15388
rect 5629 15385 5641 15388
rect 5675 15416 5687 15419
rect 7116 15416 7144 15660
rect 7285 15657 7297 15660
rect 7331 15688 7343 15691
rect 8478 15688 8484 15700
rect 7331 15660 8484 15688
rect 7331 15657 7343 15660
rect 7285 15651 7343 15657
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 10008 15660 10057 15688
rect 10008 15648 10014 15660
rect 10045 15657 10057 15660
rect 10091 15657 10103 15691
rect 10045 15651 10103 15657
rect 10229 15691 10287 15697
rect 10229 15657 10241 15691
rect 10275 15688 10287 15691
rect 10502 15688 10508 15700
rect 10275 15660 10508 15688
rect 10275 15657 10287 15660
rect 10229 15651 10287 15657
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 10652 15660 11069 15688
rect 10652 15648 10658 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11057 15651 11115 15657
rect 12158 15648 12164 15700
rect 12216 15688 12222 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 12216 15660 13185 15688
rect 12216 15648 12222 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 13173 15651 13231 15657
rect 15013 15691 15071 15697
rect 15013 15657 15025 15691
rect 15059 15688 15071 15691
rect 15102 15688 15108 15700
rect 15059 15660 15108 15688
rect 15059 15657 15071 15660
rect 15013 15651 15071 15657
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 16577 15691 16635 15697
rect 16577 15657 16589 15691
rect 16623 15688 16635 15691
rect 16850 15688 16856 15700
rect 16623 15660 16856 15688
rect 16623 15657 16635 15660
rect 16577 15651 16635 15657
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 9585 15623 9643 15629
rect 9585 15589 9597 15623
rect 9631 15620 9643 15623
rect 10962 15620 10968 15632
rect 9631 15592 10968 15620
rect 9631 15589 9643 15592
rect 9585 15583 9643 15589
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 7558 15484 7564 15496
rect 7515 15456 7564 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8720 15456 8953 15484
rect 8720 15444 8726 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9600 15416 9628 15583
rect 10962 15580 10968 15592
rect 11020 15620 11026 15632
rect 11020 15592 14504 15620
rect 11020 15580 11026 15592
rect 13633 15555 13691 15561
rect 13633 15521 13645 15555
rect 13679 15552 13691 15555
rect 13814 15552 13820 15564
rect 13679 15524 13820 15552
rect 13679 15521 13691 15524
rect 13633 15515 13691 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 14476 15561 14504 15592
rect 15654 15580 15660 15632
rect 15712 15620 15718 15632
rect 18874 15620 18880 15632
rect 15712 15592 18880 15620
rect 15712 15580 15718 15592
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 20254 15580 20260 15632
rect 20312 15620 20318 15632
rect 20717 15623 20775 15629
rect 20717 15620 20729 15623
rect 20312 15592 20729 15620
rect 20312 15580 20318 15592
rect 20717 15589 20729 15592
rect 20763 15589 20775 15623
rect 20717 15583 20775 15589
rect 14461 15555 14519 15561
rect 14461 15521 14473 15555
rect 14507 15521 14519 15555
rect 14461 15515 14519 15521
rect 14550 15512 14556 15564
rect 14608 15512 14614 15564
rect 17034 15512 17040 15564
rect 17092 15512 17098 15564
rect 17126 15512 17132 15564
rect 17184 15512 17190 15564
rect 21177 15555 21235 15561
rect 21177 15521 21189 15555
rect 21223 15552 21235 15555
rect 21542 15552 21548 15564
rect 21223 15524 21548 15552
rect 21223 15521 21235 15524
rect 21177 15515 21235 15521
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10244 15456 10701 15484
rect 5675 15388 7144 15416
rect 7392 15388 9628 15416
rect 9769 15419 9827 15425
rect 5675 15385 5687 15388
rect 5629 15379 5687 15385
rect 4982 15308 4988 15360
rect 5040 15348 5046 15360
rect 7392 15348 7420 15388
rect 9769 15385 9781 15419
rect 9815 15416 9827 15419
rect 10042 15416 10048 15428
rect 9815 15388 10048 15416
rect 9815 15385 9827 15388
rect 9769 15379 9827 15385
rect 10042 15376 10048 15388
rect 10100 15376 10106 15428
rect 10244 15360 10272 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 11296 15456 11345 15484
rect 11296 15444 11302 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 11606 15444 11612 15496
rect 11664 15444 11670 15496
rect 13354 15444 13360 15496
rect 13412 15484 13418 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13412 15456 13737 15484
rect 13412 15444 13418 15456
rect 13725 15453 13737 15456
rect 13771 15453 13783 15487
rect 15930 15484 15936 15496
rect 13725 15447 13783 15453
rect 14568 15456 15936 15484
rect 10594 15376 10600 15428
rect 10652 15376 10658 15428
rect 14568 15425 14596 15456
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15484 17923 15487
rect 18230 15484 18236 15496
rect 17911 15456 18236 15484
rect 17911 15453 17923 15456
rect 17865 15447 17923 15453
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 14553 15419 14611 15425
rect 14553 15385 14565 15419
rect 14599 15385 14611 15419
rect 18046 15416 18052 15428
rect 14553 15379 14611 15385
rect 17052 15388 18052 15416
rect 5040 15320 7420 15348
rect 5040 15308 5046 15320
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 10226 15357 10232 15360
rect 10220 15348 10232 15357
rect 10187 15320 10232 15348
rect 10220 15311 10232 15320
rect 10226 15308 10232 15311
rect 10284 15308 10290 15360
rect 10502 15308 10508 15360
rect 10560 15348 10566 15360
rect 11066 15351 11124 15357
rect 11066 15348 11078 15351
rect 10560 15320 11078 15348
rect 10560 15308 10566 15320
rect 11066 15317 11078 15320
rect 11112 15317 11124 15351
rect 11066 15311 11124 15317
rect 11422 15308 11428 15360
rect 11480 15308 11486 15360
rect 12802 15308 12808 15360
rect 12860 15348 12866 15360
rect 13446 15348 13452 15360
rect 12860 15320 13452 15348
rect 12860 15308 12866 15320
rect 13446 15308 13452 15320
rect 13504 15348 13510 15360
rect 17052 15357 17080 15388
rect 18046 15376 18052 15388
rect 18104 15376 18110 15428
rect 21269 15419 21327 15425
rect 21269 15385 21281 15419
rect 21315 15416 21327 15419
rect 21450 15416 21456 15428
rect 21315 15388 21456 15416
rect 21315 15385 21327 15388
rect 21269 15379 21327 15385
rect 21450 15376 21456 15388
rect 21508 15376 21514 15428
rect 13633 15351 13691 15357
rect 13633 15348 13645 15351
rect 13504 15320 13645 15348
rect 13504 15308 13510 15320
rect 13633 15317 13645 15320
rect 13679 15348 13691 15351
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 13679 15320 16129 15348
rect 13679 15317 13691 15320
rect 13633 15311 13691 15317
rect 16117 15317 16129 15320
rect 16163 15348 16175 15351
rect 17037 15351 17095 15357
rect 17037 15348 17049 15351
rect 16163 15320 17049 15348
rect 16163 15317 16175 15320
rect 16117 15311 16175 15317
rect 17037 15317 17049 15320
rect 17083 15317 17095 15351
rect 17037 15311 17095 15317
rect 17678 15308 17684 15360
rect 17736 15308 17742 15360
rect 21174 15308 21180 15360
rect 21232 15308 21238 15360
rect 1104 15258 21988 15280
rect 1104 15206 4220 15258
rect 4272 15206 4284 15258
rect 4336 15206 4348 15258
rect 4400 15206 4412 15258
rect 4464 15206 4476 15258
rect 4528 15206 9441 15258
rect 9493 15206 9505 15258
rect 9557 15206 9569 15258
rect 9621 15206 9633 15258
rect 9685 15206 9697 15258
rect 9749 15206 14662 15258
rect 14714 15206 14726 15258
rect 14778 15206 14790 15258
rect 14842 15206 14854 15258
rect 14906 15206 14918 15258
rect 14970 15206 19883 15258
rect 19935 15206 19947 15258
rect 19999 15206 20011 15258
rect 20063 15206 20075 15258
rect 20127 15206 20139 15258
rect 20191 15206 21988 15258
rect 1104 15184 21988 15206
rect 3697 15147 3755 15153
rect 3697 15113 3709 15147
rect 3743 15144 3755 15147
rect 4614 15144 4620 15156
rect 3743 15116 4620 15144
rect 3743 15113 3755 15116
rect 3697 15107 3755 15113
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 9306 15144 9312 15156
rect 8128 15116 9312 15144
rect 3513 15079 3571 15085
rect 3513 15045 3525 15079
rect 3559 15076 3571 15079
rect 4062 15076 4068 15088
rect 3559 15048 4068 15076
rect 3559 15045 3571 15048
rect 3513 15039 3571 15045
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 3418 15008 3424 15020
rect 3099 14980 3424 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 3418 14968 3424 14980
rect 3476 14968 3482 15020
rect 8128 15017 8156 15116
rect 9306 15104 9312 15116
rect 9364 15104 9370 15156
rect 10689 15147 10747 15153
rect 10689 15113 10701 15147
rect 10735 15144 10747 15147
rect 15470 15144 15476 15156
rect 10735 15116 15476 15144
rect 10735 15113 10747 15116
rect 10689 15107 10747 15113
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 20073 15147 20131 15153
rect 20073 15113 20085 15147
rect 20119 15113 20131 15147
rect 20073 15107 20131 15113
rect 9030 15036 9036 15088
rect 9088 15036 9094 15088
rect 10226 15036 10232 15088
rect 10284 15076 10290 15088
rect 10321 15079 10379 15085
rect 10321 15076 10333 15079
rect 10284 15048 10333 15076
rect 10284 15036 10290 15048
rect 10321 15045 10333 15048
rect 10367 15045 10379 15079
rect 10321 15039 10379 15045
rect 10502 15036 10508 15088
rect 10560 15036 10566 15088
rect 10870 15036 10876 15088
rect 10928 15036 10934 15088
rect 11238 15036 11244 15088
rect 11296 15036 11302 15088
rect 12066 15036 12072 15088
rect 12124 15036 12130 15088
rect 13449 15079 13507 15085
rect 13449 15076 13461 15079
rect 12912 15048 13461 15076
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 11974 15008 11980 15020
rect 11931 14980 11980 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 11974 14968 11980 14980
rect 12032 15008 12038 15020
rect 12912 15008 12940 15048
rect 13449 15045 13461 15048
rect 13495 15045 13507 15079
rect 13449 15039 13507 15045
rect 15838 15036 15844 15088
rect 15896 15076 15902 15088
rect 16301 15079 16359 15085
rect 16301 15076 16313 15079
rect 15896 15048 16313 15076
rect 15896 15036 15902 15048
rect 16301 15045 16313 15048
rect 16347 15045 16359 15079
rect 17954 15076 17960 15088
rect 16301 15039 16359 15045
rect 17144 15048 17960 15076
rect 12032 14980 12940 15008
rect 12032 14968 12038 14980
rect 13170 14968 13176 15020
rect 13228 14968 13234 15020
rect 15470 14968 15476 15020
rect 15528 14968 15534 15020
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 15008 16175 15011
rect 17144 15008 17172 15048
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 20088 15076 20116 15107
rect 20410 15079 20468 15085
rect 20410 15076 20422 15079
rect 20088 15048 20422 15076
rect 20410 15045 20422 15048
rect 20456 15045 20468 15079
rect 20410 15039 20468 15045
rect 16163 14980 17172 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 17218 14968 17224 15020
rect 17276 14968 17282 15020
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 17477 15011 17535 15017
rect 17477 15008 17489 15011
rect 17368 14980 17489 15008
rect 17368 14968 17374 14980
rect 17477 14977 17489 14980
rect 17523 14977 17535 15011
rect 17477 14971 17535 14977
rect 19613 15011 19671 15017
rect 19613 14977 19625 15011
rect 19659 15008 19671 15011
rect 19889 15011 19947 15017
rect 19659 14980 19748 15008
rect 19659 14977 19671 14980
rect 19613 14971 19671 14977
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 5074 14940 5080 14952
rect 3835 14912 5080 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 5074 14900 5080 14912
rect 5132 14940 5138 14952
rect 5350 14940 5356 14952
rect 5132 14912 5356 14940
rect 5132 14900 5138 14912
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 8389 14943 8447 14949
rect 8389 14940 8401 14943
rect 7800 14912 8401 14940
rect 7800 14900 7806 14912
rect 8389 14909 8401 14912
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12618 14940 12624 14952
rect 12207 14912 12624 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14940 13415 14943
rect 13538 14940 13544 14952
rect 13403 14912 13544 14940
rect 13403 14909 13415 14912
rect 13357 14903 13415 14909
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 16393 14943 16451 14949
rect 16393 14909 16405 14943
rect 16439 14940 16451 14943
rect 16574 14940 16580 14952
rect 16439 14912 16580 14940
rect 16439 14909 16451 14912
rect 16393 14903 16451 14909
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 2866 14832 2872 14884
rect 2924 14872 2930 14884
rect 3237 14875 3295 14881
rect 3237 14872 3249 14875
rect 2924 14844 3249 14872
rect 2924 14832 2930 14844
rect 3237 14841 3249 14844
rect 3283 14841 3295 14875
rect 10686 14872 10692 14884
rect 3237 14835 3295 14841
rect 9784 14844 10692 14872
rect 2958 14764 2964 14816
rect 3016 14764 3022 14816
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 9784 14804 9812 14844
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 11606 14832 11612 14884
rect 11664 14832 11670 14884
rect 14734 14832 14740 14884
rect 14792 14872 14798 14884
rect 15841 14875 15899 14881
rect 15841 14872 15853 14875
rect 14792 14844 15853 14872
rect 14792 14832 14798 14844
rect 15841 14841 15853 14844
rect 15887 14841 15899 14875
rect 19720 14872 19748 14980
rect 19889 14977 19901 15011
rect 19935 15008 19947 15011
rect 20254 15008 20260 15020
rect 19935 14980 20260 15008
rect 19935 14977 19947 14980
rect 19889 14971 19947 14977
rect 20254 14968 20260 14980
rect 20312 14968 20318 15020
rect 19794 14900 19800 14952
rect 19852 14940 19858 14952
rect 20165 14943 20223 14949
rect 20165 14940 20177 14943
rect 19852 14912 20177 14940
rect 19852 14900 19858 14912
rect 20165 14909 20177 14912
rect 20211 14909 20223 14943
rect 20165 14903 20223 14909
rect 19886 14872 19892 14884
rect 19720 14844 19892 14872
rect 15841 14835 15899 14841
rect 19886 14832 19892 14844
rect 19944 14832 19950 14884
rect 5868 14776 9812 14804
rect 9861 14807 9919 14813
rect 5868 14764 5874 14776
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 10410 14804 10416 14816
rect 9907 14776 10416 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 10505 14807 10563 14813
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 10594 14804 10600 14816
rect 10551 14776 10600 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 12986 14764 12992 14816
rect 13044 14764 13050 14816
rect 13446 14764 13452 14816
rect 13504 14764 13510 14816
rect 15286 14764 15292 14816
rect 15344 14764 15350 14816
rect 18598 14764 18604 14816
rect 18656 14764 18662 14816
rect 19429 14807 19487 14813
rect 19429 14773 19441 14807
rect 19475 14804 19487 14807
rect 19610 14804 19616 14816
rect 19475 14776 19616 14804
rect 19475 14773 19487 14776
rect 19429 14767 19487 14773
rect 19610 14764 19616 14776
rect 19668 14764 19674 14816
rect 21542 14764 21548 14816
rect 21600 14764 21606 14816
rect 1104 14714 21988 14736
rect 1104 14662 3560 14714
rect 3612 14662 3624 14714
rect 3676 14662 3688 14714
rect 3740 14662 3752 14714
rect 3804 14662 3816 14714
rect 3868 14662 8781 14714
rect 8833 14662 8845 14714
rect 8897 14662 8909 14714
rect 8961 14662 8973 14714
rect 9025 14662 9037 14714
rect 9089 14662 14002 14714
rect 14054 14662 14066 14714
rect 14118 14662 14130 14714
rect 14182 14662 14194 14714
rect 14246 14662 14258 14714
rect 14310 14662 19223 14714
rect 19275 14662 19287 14714
rect 19339 14662 19351 14714
rect 19403 14662 19415 14714
rect 19467 14662 19479 14714
rect 19531 14662 21988 14714
rect 1104 14640 21988 14662
rect 5810 14560 5816 14612
rect 5868 14560 5874 14612
rect 7650 14600 7656 14612
rect 7300 14572 7656 14600
rect 5074 14532 5080 14544
rect 4540 14504 5080 14532
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 2590 14464 2596 14476
rect 1627 14436 2596 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 3326 14424 3332 14476
rect 3384 14464 3390 14476
rect 4540 14464 4568 14504
rect 5074 14492 5080 14504
rect 5132 14492 5138 14544
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 7300 14532 7328 14572
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 10318 14600 10324 14612
rect 10091 14572 10324 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10318 14560 10324 14572
rect 10376 14600 10382 14612
rect 10594 14600 10600 14612
rect 10376 14572 10600 14600
rect 10376 14560 10382 14572
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 11974 14560 11980 14612
rect 12032 14560 12038 14612
rect 12894 14560 12900 14612
rect 12952 14600 12958 14612
rect 16022 14600 16028 14612
rect 12952 14572 16028 14600
rect 12952 14560 12958 14572
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 16632 14572 17540 14600
rect 16632 14560 16638 14572
rect 9033 14535 9091 14541
rect 9033 14532 9045 14535
rect 5684 14504 7328 14532
rect 7392 14504 9045 14532
rect 5684 14492 5690 14504
rect 3384 14436 4568 14464
rect 3384 14424 3390 14436
rect 2958 14356 2964 14408
rect 3016 14356 3022 14408
rect 3970 14356 3976 14408
rect 4028 14356 4034 14408
rect 4540 14405 4568 14436
rect 4982 14424 4988 14476
rect 5040 14464 5046 14476
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 5040 14436 5365 14464
rect 5040 14424 5046 14436
rect 5353 14433 5365 14436
rect 5399 14464 5411 14467
rect 5399 14436 6684 14464
rect 5399 14433 5411 14436
rect 5353 14427 5411 14433
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4433 14399 4491 14405
rect 4203 14368 4384 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 1578 14288 1584 14340
rect 1636 14328 1642 14340
rect 1857 14331 1915 14337
rect 1857 14328 1869 14331
rect 1636 14300 1869 14328
rect 1636 14288 1642 14300
rect 1857 14297 1869 14300
rect 1903 14297 1915 14331
rect 1857 14291 1915 14297
rect 3234 14288 3240 14340
rect 3292 14328 3298 14340
rect 3789 14331 3847 14337
rect 3789 14328 3801 14331
rect 3292 14300 3801 14328
rect 3292 14288 3298 14300
rect 3789 14297 3801 14300
rect 3835 14297 3847 14331
rect 3789 14291 3847 14297
rect 2866 14220 2872 14272
rect 2924 14260 2930 14272
rect 3326 14260 3332 14272
rect 2924 14232 3332 14260
rect 2924 14220 2930 14232
rect 3326 14220 3332 14232
rect 3384 14220 3390 14272
rect 4356 14260 4384 14368
rect 4433 14365 4445 14399
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4448 14328 4476 14359
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 4893 14399 4951 14405
rect 4893 14396 4905 14399
rect 4672 14368 4905 14396
rect 4672 14356 4678 14368
rect 4893 14365 4905 14368
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5166 14396 5172 14408
rect 5123 14368 5172 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5166 14356 5172 14368
rect 5224 14396 5230 14408
rect 5534 14396 5540 14408
rect 5224 14368 5540 14396
rect 5224 14356 5230 14368
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5626 14356 5632 14408
rect 5684 14356 5690 14408
rect 6656 14405 6684 14436
rect 7392 14405 7420 14504
rect 9033 14501 9045 14504
rect 9079 14501 9091 14535
rect 10410 14532 10416 14544
rect 9033 14495 9091 14501
rect 9232 14504 10416 14532
rect 7742 14424 7748 14476
rect 7800 14424 7806 14476
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14464 8539 14467
rect 9232 14464 9260 14504
rect 10410 14492 10416 14504
rect 10468 14492 10474 14544
rect 17512 14532 17540 14572
rect 17954 14560 17960 14612
rect 18012 14560 18018 14612
rect 18230 14560 18236 14612
rect 18288 14560 18294 14612
rect 19518 14600 19524 14612
rect 18892 14572 19524 14600
rect 18892 14532 18920 14572
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19886 14560 19892 14612
rect 19944 14600 19950 14612
rect 20901 14603 20959 14609
rect 20901 14600 20913 14603
rect 19944 14572 20913 14600
rect 19944 14560 19950 14572
rect 20901 14569 20913 14572
rect 20947 14569 20959 14603
rect 20901 14563 20959 14569
rect 17512 14504 18920 14532
rect 8527 14436 9260 14464
rect 8527 14433 8539 14436
rect 8481 14427 8539 14433
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 9364 14436 10609 14464
rect 9364 14424 9370 14436
rect 10597 14433 10609 14436
rect 10643 14433 10655 14467
rect 10597 14427 10655 14433
rect 13630 14424 13636 14476
rect 13688 14464 13694 14476
rect 14366 14464 14372 14476
rect 13688 14436 14372 14464
rect 13688 14424 13694 14436
rect 14366 14424 14372 14436
rect 14424 14464 14430 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14424 14436 15025 14464
rect 14424 14424 14430 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15013 14427 15071 14433
rect 18785 14467 18843 14473
rect 18785 14433 18797 14467
rect 18831 14464 18843 14467
rect 18892 14464 18920 14504
rect 20625 14535 20683 14541
rect 20625 14501 20637 14535
rect 20671 14501 20683 14535
rect 20625 14495 20683 14501
rect 18831 14436 18920 14464
rect 20640 14464 20668 14495
rect 21358 14464 21364 14476
rect 20640 14436 21364 14464
rect 18831 14433 18843 14436
rect 18785 14427 18843 14433
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 21450 14424 21456 14476
rect 21508 14424 21514 14476
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14396 6699 14399
rect 7377 14399 7435 14405
rect 6687 14368 6960 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 4706 14328 4712 14340
rect 4448 14300 4712 14328
rect 4706 14288 4712 14300
rect 4764 14288 4770 14340
rect 4801 14331 4859 14337
rect 4801 14297 4813 14331
rect 4847 14328 4859 14331
rect 5258 14328 5264 14340
rect 4847 14300 5264 14328
rect 4847 14297 4859 14300
rect 4801 14291 4859 14297
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 6472 14328 6500 14359
rect 6822 14328 6828 14340
rect 6472 14300 6828 14328
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 6932 14328 6960 14368
rect 7377 14365 7389 14399
rect 7423 14365 7435 14399
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 7377 14359 7435 14365
rect 8588 14328 8616 14382
rect 8772 14368 9781 14396
rect 8772 14328 8800 14368
rect 9769 14365 9781 14368
rect 9815 14365 9827 14399
rect 9769 14359 9827 14365
rect 10864 14399 10922 14405
rect 10864 14365 10876 14399
rect 10910 14396 10922 14399
rect 11422 14396 11428 14408
rect 10910 14368 11428 14396
rect 10910 14365 10922 14368
rect 10864 14359 10922 14365
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12250 14396 12256 14408
rect 12207 14368 12256 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12250 14356 12256 14368
rect 12308 14396 12314 14408
rect 13648 14396 13676 14424
rect 12308 14368 13676 14396
rect 12308 14356 12314 14368
rect 13722 14356 13728 14408
rect 13780 14356 13786 14408
rect 14734 14356 14740 14408
rect 14792 14356 14798 14408
rect 15286 14405 15292 14408
rect 15280 14396 15292 14405
rect 15247 14368 15292 14396
rect 15280 14359 15292 14368
rect 15286 14356 15292 14359
rect 15344 14356 15350 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 17218 14396 17224 14408
rect 16623 14368 17224 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14396 18567 14399
rect 18690 14396 18696 14408
rect 18555 14368 18696 14396
rect 18555 14365 18567 14368
rect 18509 14359 18567 14365
rect 18690 14356 18696 14368
rect 18748 14396 18754 14408
rect 19245 14399 19303 14405
rect 18748 14368 19196 14396
rect 18748 14356 18754 14368
rect 6932 14300 7972 14328
rect 8588 14300 8800 14328
rect 4890 14260 4896 14272
rect 4356 14232 4896 14260
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 6273 14263 6331 14269
rect 6273 14260 6285 14263
rect 6052 14232 6285 14260
rect 6052 14220 6058 14232
rect 6273 14229 6285 14232
rect 6319 14229 6331 14263
rect 6273 14223 6331 14229
rect 6733 14263 6791 14269
rect 6733 14229 6745 14263
rect 6779 14260 6791 14263
rect 7006 14260 7012 14272
rect 6779 14232 7012 14260
rect 6779 14229 6791 14232
rect 6733 14223 6791 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 7834 14260 7840 14272
rect 7607 14232 7840 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 7944 14260 7972 14300
rect 9214 14288 9220 14340
rect 9272 14328 9278 14340
rect 9309 14331 9367 14337
rect 9309 14328 9321 14331
rect 9272 14300 9321 14328
rect 9272 14288 9278 14300
rect 9309 14297 9321 14300
rect 9355 14297 9367 14331
rect 9309 14291 9367 14297
rect 9585 14331 9643 14337
rect 9585 14297 9597 14331
rect 9631 14328 9643 14331
rect 10045 14331 10103 14337
rect 10045 14328 10057 14331
rect 9631 14300 10057 14328
rect 9631 14297 9643 14300
rect 9585 14291 9643 14297
rect 9784 14272 9812 14300
rect 10045 14297 10057 14300
rect 10091 14297 10103 14331
rect 10045 14291 10103 14297
rect 10226 14288 10232 14340
rect 10284 14288 10290 14340
rect 12434 14337 12440 14340
rect 12428 14291 12440 14337
rect 12434 14288 12440 14291
rect 12492 14288 12498 14340
rect 16822 14331 16880 14337
rect 16822 14328 16834 14331
rect 14936 14300 16834 14328
rect 8662 14260 8668 14272
rect 7944 14232 8668 14260
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 9493 14263 9551 14269
rect 9493 14260 9505 14263
rect 9180 14232 9505 14260
rect 9180 14220 9186 14232
rect 9493 14229 9505 14232
rect 9539 14229 9551 14263
rect 9493 14223 9551 14229
rect 9766 14220 9772 14272
rect 9824 14220 9830 14272
rect 13538 14220 13544 14272
rect 13596 14220 13602 14272
rect 13906 14220 13912 14272
rect 13964 14220 13970 14272
rect 14936 14269 14964 14300
rect 16822 14297 16834 14300
rect 16868 14297 16880 14331
rect 19168 14328 19196 14368
rect 19245 14365 19257 14399
rect 19291 14396 19303 14399
rect 19334 14396 19340 14408
rect 19291 14368 19340 14396
rect 19291 14365 19303 14368
rect 19245 14359 19303 14365
rect 19334 14356 19340 14368
rect 19392 14396 19398 14408
rect 19794 14396 19800 14408
rect 19392 14368 19800 14396
rect 19392 14356 19398 14368
rect 19794 14356 19800 14368
rect 19852 14356 19858 14408
rect 19512 14331 19570 14337
rect 19168 14300 19472 14328
rect 16822 14291 16880 14297
rect 14921 14263 14979 14269
rect 14921 14229 14933 14263
rect 14967 14229 14979 14263
rect 14921 14223 14979 14229
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15896 14232 16405 14260
rect 15896 14220 15902 14232
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 18230 14220 18236 14272
rect 18288 14260 18294 14272
rect 18598 14260 18604 14272
rect 18288 14232 18604 14260
rect 18288 14220 18294 14232
rect 18598 14220 18604 14232
rect 18656 14260 18662 14272
rect 18693 14263 18751 14269
rect 18693 14260 18705 14263
rect 18656 14232 18705 14260
rect 18656 14220 18662 14232
rect 18693 14229 18705 14232
rect 18739 14229 18751 14263
rect 19444 14260 19472 14300
rect 19512 14297 19524 14331
rect 19558 14328 19570 14331
rect 19610 14328 19616 14340
rect 19558 14300 19616 14328
rect 19558 14297 19570 14300
rect 19512 14291 19570 14297
rect 19610 14288 19616 14300
rect 19668 14288 19674 14340
rect 20714 14260 20720 14272
rect 19444 14232 20720 14260
rect 18693 14223 18751 14229
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 20806 14220 20812 14272
rect 20864 14260 20870 14272
rect 21361 14263 21419 14269
rect 21361 14260 21373 14263
rect 20864 14232 21373 14260
rect 20864 14220 20870 14232
rect 21361 14229 21373 14232
rect 21407 14229 21419 14263
rect 21361 14223 21419 14229
rect 1104 14170 21988 14192
rect 1104 14118 4220 14170
rect 4272 14118 4284 14170
rect 4336 14118 4348 14170
rect 4400 14118 4412 14170
rect 4464 14118 4476 14170
rect 4528 14118 9441 14170
rect 9493 14118 9505 14170
rect 9557 14118 9569 14170
rect 9621 14118 9633 14170
rect 9685 14118 9697 14170
rect 9749 14118 14662 14170
rect 14714 14118 14726 14170
rect 14778 14118 14790 14170
rect 14842 14118 14854 14170
rect 14906 14118 14918 14170
rect 14970 14118 19883 14170
rect 19935 14118 19947 14170
rect 19999 14118 20011 14170
rect 20063 14118 20075 14170
rect 20127 14118 20139 14170
rect 20191 14118 21988 14170
rect 1104 14096 21988 14118
rect 1578 14016 1584 14068
rect 1636 14016 1642 14068
rect 2682 14016 2688 14068
rect 2740 14056 2746 14068
rect 5718 14056 5724 14068
rect 2740 14028 5724 14056
rect 2740 14016 2746 14028
rect 2038 13948 2044 14000
rect 2096 13948 2102 14000
rect 2866 13988 2872 14000
rect 2148 13960 2872 13988
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 2148 13920 2176 13960
rect 2866 13948 2872 13960
rect 2924 13948 2930 14000
rect 3068 13988 3096 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 5810 14016 5816 14068
rect 5868 14016 5874 14068
rect 6546 14016 6552 14068
rect 6604 14016 6610 14068
rect 9306 14056 9312 14068
rect 7576 14028 9312 14056
rect 2976 13960 3096 13988
rect 1719 13906 2176 13920
rect 1719 13892 2162 13906
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 2774 13880 2780 13932
rect 2832 13880 2838 13932
rect 2976 13929 3004 13960
rect 3234 13948 3240 14000
rect 3292 13948 3298 14000
rect 4522 13988 4528 14000
rect 4462 13960 4528 13988
rect 4522 13948 4528 13960
rect 4580 13948 4586 14000
rect 4614 13948 4620 14000
rect 4672 13988 4678 14000
rect 5353 13991 5411 13997
rect 5353 13988 5365 13991
rect 4672 13960 5365 13988
rect 4672 13948 4678 13960
rect 5353 13957 5365 13960
rect 5399 13957 5411 13991
rect 5353 13951 5411 13957
rect 5626 13948 5632 14000
rect 5684 13948 5690 14000
rect 6730 13988 6736 14000
rect 6564 13960 6736 13988
rect 6564 13929 6592 13960
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 2961 13883 3019 13889
rect 4724 13892 5181 13920
rect 4724 13864 4752 13892
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 6181 13923 6239 13929
rect 6181 13889 6193 13923
rect 6227 13920 6239 13923
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6227 13892 6561 13920
rect 6227 13889 6239 13892
rect 6181 13883 6239 13889
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 6549 13883 6607 13889
rect 6656 13892 7113 13920
rect 4706 13812 4712 13864
rect 4764 13812 4770 13864
rect 4893 13855 4951 13861
rect 4893 13821 4905 13855
rect 4939 13821 4951 13855
rect 4893 13815 4951 13821
rect 4908 13784 4936 13815
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 5132 13824 5273 13852
rect 5132 13812 5138 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5261 13815 5319 13821
rect 5460 13824 6101 13852
rect 5166 13784 5172 13796
rect 4908 13756 5172 13784
rect 5166 13744 5172 13756
rect 5224 13784 5230 13796
rect 5460 13784 5488 13824
rect 6089 13821 6101 13824
rect 6135 13821 6147 13855
rect 6089 13815 6147 13821
rect 6365 13855 6423 13861
rect 6365 13821 6377 13855
rect 6411 13821 6423 13855
rect 6656 13852 6684 13892
rect 7101 13889 7113 13892
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7374 13880 7380 13932
rect 7432 13880 7438 13932
rect 7576 13929 7604 14028
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 11793 14059 11851 14065
rect 11793 14025 11805 14059
rect 11839 14056 11851 14059
rect 12342 14056 12348 14068
rect 11839 14028 12348 14056
rect 11839 14025 11851 14028
rect 11793 14019 11851 14025
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12894 14056 12900 14068
rect 12544 14028 12900 14056
rect 7834 13948 7840 14000
rect 7892 13948 7898 14000
rect 8570 13948 8576 14000
rect 8628 13948 8634 14000
rect 10413 13991 10471 13997
rect 10413 13957 10425 13991
rect 10459 13988 10471 13991
rect 10502 13988 10508 14000
rect 10459 13960 10508 13988
rect 10459 13957 10471 13960
rect 10413 13951 10471 13957
rect 10502 13948 10508 13960
rect 10560 13988 10566 14000
rect 10560 13960 10824 13988
rect 10560 13948 10566 13960
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13889 7619 13923
rect 9766 13920 9772 13932
rect 7561 13883 7619 13889
rect 9324 13892 9772 13920
rect 6365 13815 6423 13821
rect 6472 13824 6684 13852
rect 5224 13756 5488 13784
rect 5224 13744 5230 13756
rect 5626 13744 5632 13796
rect 5684 13784 5690 13796
rect 6380 13784 6408 13815
rect 5684 13756 6408 13784
rect 5684 13744 5690 13756
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 5997 13719 6055 13725
rect 5997 13716 6009 13719
rect 5316 13688 6009 13716
rect 5316 13676 5322 13688
rect 5997 13685 6009 13688
rect 6043 13716 6055 13719
rect 6472 13716 6500 13824
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 7466 13812 7472 13864
rect 7524 13812 7530 13864
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 9324 13861 9352 13892
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 10134 13920 10140 13932
rect 9999 13892 10140 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 9309 13855 9367 13861
rect 8352 13824 8892 13852
rect 8352 13812 8358 13824
rect 8864 13784 8892 13824
rect 9309 13821 9321 13855
rect 9355 13821 9367 13855
rect 10336 13852 10364 13883
rect 10686 13880 10692 13932
rect 10744 13880 10750 13932
rect 10796 13929 10824 13960
rect 10870 13948 10876 14000
rect 10928 13988 10934 14000
rect 12437 13991 12495 13997
rect 10928 13960 11284 13988
rect 10928 13948 10934 13960
rect 11256 13929 11284 13960
rect 12437 13957 12449 13991
rect 12483 13988 12495 13991
rect 12544 13988 12572 14028
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 13538 14016 13544 14068
rect 13596 14056 13602 14068
rect 17221 14059 17279 14065
rect 13596 14028 14688 14056
rect 13596 14016 13602 14028
rect 12483 13960 12572 13988
rect 12483 13957 12495 13960
rect 12437 13951 12495 13957
rect 12618 13948 12624 14000
rect 12676 13988 12682 14000
rect 13170 13988 13176 14000
rect 12676 13960 13176 13988
rect 12676 13948 12682 13960
rect 13170 13948 13176 13960
rect 13228 13988 13234 14000
rect 13228 13960 13584 13988
rect 13228 13948 13234 13960
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11241 13923 11299 13929
rect 11241 13889 11253 13923
rect 11287 13889 11299 13923
rect 11241 13883 11299 13889
rect 11609 13923 11667 13929
rect 11609 13889 11621 13923
rect 11655 13920 11667 13923
rect 11959 13923 12017 13929
rect 11959 13920 11971 13923
rect 11655 13892 11971 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 11959 13889 11971 13892
rect 12005 13889 12017 13923
rect 11959 13883 12017 13889
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 13446 13920 13452 13932
rect 12299 13892 13452 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 10410 13852 10416 13864
rect 10336 13824 10416 13852
rect 9309 13815 9367 13821
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 11072 13852 11100 13883
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 13556 13920 13584 13960
rect 13906 13948 13912 14000
rect 13964 13997 13970 14000
rect 14660 13997 14688 14028
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 17310 14056 17316 14068
rect 17267 14028 17316 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 18690 14016 18696 14068
rect 18748 14016 18754 14068
rect 18782 14016 18788 14068
rect 18840 14056 18846 14068
rect 18840 14028 19472 14056
rect 18840 14016 18846 14028
rect 13964 13988 13976 13997
rect 14645 13991 14703 13997
rect 13964 13960 14009 13988
rect 13964 13951 13976 13960
rect 14645 13957 14657 13991
rect 14691 13957 14703 13991
rect 14645 13951 14703 13957
rect 13964 13948 13970 13951
rect 14826 13948 14832 14000
rect 14884 13948 14890 14000
rect 15838 13948 15844 14000
rect 15896 13948 15902 14000
rect 16022 13948 16028 14000
rect 16080 13948 16086 14000
rect 17580 13991 17638 13997
rect 17580 13957 17592 13991
rect 17626 13988 17638 13991
rect 17678 13988 17684 14000
rect 17626 13960 17684 13988
rect 17626 13957 17638 13960
rect 17580 13951 17638 13957
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 19334 13988 19340 14000
rect 18892 13960 19340 13988
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 13556 13892 14933 13920
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 16040 13920 16068 13948
rect 15712 13892 16068 13920
rect 15712 13880 15718 13892
rect 17034 13880 17040 13932
rect 17092 13880 17098 13932
rect 17218 13880 17224 13932
rect 17276 13920 17282 13932
rect 18892 13929 18920 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 17313 13923 17371 13929
rect 17313 13920 17325 13923
rect 17276 13892 17325 13920
rect 17276 13880 17282 13892
rect 17313 13889 17325 13892
rect 17359 13889 17371 13923
rect 17313 13883 17371 13889
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 18966 13880 18972 13932
rect 19024 13920 19030 13932
rect 19133 13923 19191 13929
rect 19133 13920 19145 13923
rect 19024 13892 19145 13920
rect 19024 13880 19030 13892
rect 19133 13889 19145 13892
rect 19179 13889 19191 13923
rect 19444 13920 19472 14028
rect 20254 14016 20260 14068
rect 20312 14056 20318 14068
rect 21269 14059 21327 14065
rect 21269 14056 21281 14059
rect 20312 14028 21281 14056
rect 20312 14016 20318 14028
rect 21269 14025 21281 14028
rect 21315 14025 21327 14059
rect 21269 14019 21327 14025
rect 20622 13948 20628 14000
rect 20680 13948 20686 14000
rect 20806 13948 20812 14000
rect 20864 13948 20870 14000
rect 19444 13892 20668 13920
rect 19133 13883 19191 13889
rect 12529 13855 12587 13861
rect 12529 13852 12541 13855
rect 11072 13824 12541 13852
rect 12529 13821 12541 13824
rect 12575 13852 12587 13855
rect 12618 13852 12624 13864
rect 12575 13824 12624 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 12618 13812 12624 13824
rect 12676 13812 12682 13864
rect 14185 13855 14243 13861
rect 14185 13821 14197 13855
rect 14231 13852 14243 13855
rect 14366 13852 14372 13864
rect 14231 13824 14372 13852
rect 14231 13821 14243 13824
rect 14185 13815 14243 13821
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 15528 13824 15608 13852
rect 15528 13812 15534 13824
rect 11790 13784 11796 13796
rect 8864 13756 11796 13784
rect 11790 13744 11796 13756
rect 11848 13744 11854 13796
rect 15580 13793 15608 13824
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15988 13824 16129 13852
rect 15988 13812 15994 13824
rect 16117 13821 16129 13824
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 20530 13812 20536 13864
rect 20588 13812 20594 13864
rect 20640 13852 20668 13892
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 21453 13923 21511 13929
rect 21453 13920 21465 13923
rect 20772 13892 21465 13920
rect 20772 13880 20778 13892
rect 21453 13889 21465 13892
rect 21499 13889 21511 13923
rect 21453 13883 21511 13889
rect 20898 13852 20904 13864
rect 20640 13824 20904 13852
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 15565 13787 15623 13793
rect 15565 13753 15577 13787
rect 15611 13753 15623 13787
rect 15565 13747 15623 13753
rect 19886 13744 19892 13796
rect 19944 13784 19950 13796
rect 21085 13787 21143 13793
rect 21085 13784 21097 13787
rect 19944 13756 21097 13784
rect 19944 13744 19950 13756
rect 21085 13753 21097 13756
rect 21131 13753 21143 13787
rect 21085 13747 21143 13753
rect 6043 13688 6500 13716
rect 6043 13685 6055 13688
rect 5997 13679 6055 13685
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 9214 13716 9220 13728
rect 8536 13688 9220 13716
rect 8536 13676 8542 13688
rect 9214 13676 9220 13688
rect 9272 13716 9278 13728
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 9272 13688 9597 13716
rect 9272 13676 9278 13688
rect 9585 13685 9597 13688
rect 9631 13716 9643 13719
rect 10226 13716 10232 13728
rect 9631 13688 10232 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 12805 13719 12863 13725
rect 12805 13685 12817 13719
rect 12851 13716 12863 13719
rect 13262 13716 13268 13728
rect 12851 13688 13268 13716
rect 12851 13685 12863 13688
rect 12805 13679 12863 13685
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 14369 13719 14427 13725
rect 14369 13716 14381 13719
rect 13872 13688 14381 13716
rect 13872 13676 13878 13688
rect 14369 13685 14381 13688
rect 14415 13685 14427 13719
rect 14369 13679 14427 13685
rect 20257 13719 20315 13725
rect 20257 13685 20269 13719
rect 20303 13716 20315 13719
rect 20806 13716 20812 13728
rect 20303 13688 20812 13716
rect 20303 13685 20315 13688
rect 20257 13679 20315 13685
rect 20806 13676 20812 13688
rect 20864 13676 20870 13728
rect 1104 13626 21988 13648
rect 1104 13574 3560 13626
rect 3612 13574 3624 13626
rect 3676 13574 3688 13626
rect 3740 13574 3752 13626
rect 3804 13574 3816 13626
rect 3868 13574 8781 13626
rect 8833 13574 8845 13626
rect 8897 13574 8909 13626
rect 8961 13574 8973 13626
rect 9025 13574 9037 13626
rect 9089 13574 14002 13626
rect 14054 13574 14066 13626
rect 14118 13574 14130 13626
rect 14182 13574 14194 13626
rect 14246 13574 14258 13626
rect 14310 13574 19223 13626
rect 19275 13574 19287 13626
rect 19339 13574 19351 13626
rect 19403 13574 19415 13626
rect 19467 13574 19479 13626
rect 19531 13574 21988 13626
rect 1104 13552 21988 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3513 13515 3571 13521
rect 3513 13512 3525 13515
rect 2832 13484 3525 13512
rect 2832 13472 2838 13484
rect 3513 13481 3525 13484
rect 3559 13481 3571 13515
rect 3513 13475 3571 13481
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13376 1823 13379
rect 2682 13376 2688 13388
rect 1811 13348 2688 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 3528 13376 3556 13475
rect 4522 13472 4528 13524
rect 4580 13472 4586 13524
rect 4798 13472 4804 13524
rect 4856 13512 4862 13524
rect 4893 13515 4951 13521
rect 4893 13512 4905 13515
rect 4856 13484 4905 13512
rect 4856 13472 4862 13484
rect 4893 13481 4905 13484
rect 4939 13481 4951 13515
rect 4893 13475 4951 13481
rect 5166 13472 5172 13524
rect 5224 13472 5230 13524
rect 5258 13472 5264 13524
rect 5316 13472 5322 13524
rect 7098 13512 7104 13524
rect 5368 13484 7104 13512
rect 4341 13379 4399 13385
rect 3528 13348 4016 13376
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 3786 13308 3792 13320
rect 3384 13280 3792 13308
rect 3384 13268 3390 13280
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 3988 13317 4016 13348
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 4706 13376 4712 13388
rect 4387 13348 4712 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 5368 13385 5396 13484
rect 7098 13472 7104 13484
rect 7156 13472 7162 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 7432 13484 7757 13512
rect 7432 13472 7438 13484
rect 7745 13481 7757 13484
rect 7791 13481 7803 13515
rect 8294 13512 8300 13524
rect 7745 13475 7803 13481
rect 7852 13484 8300 13512
rect 7852 13444 7880 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8570 13472 8576 13524
rect 8628 13472 8634 13524
rect 9122 13472 9128 13524
rect 9180 13472 9186 13524
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10100 13484 10793 13512
rect 10100 13472 10106 13484
rect 10781 13481 10793 13484
rect 10827 13481 10839 13515
rect 10781 13475 10839 13481
rect 12161 13515 12219 13521
rect 12161 13481 12173 13515
rect 12207 13512 12219 13515
rect 12434 13512 12440 13524
rect 12207 13484 12440 13512
rect 12207 13481 12219 13484
rect 12161 13475 12219 13481
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13504 13484 13645 13512
rect 13504 13472 13510 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 17034 13472 17040 13524
rect 17092 13512 17098 13524
rect 17773 13515 17831 13521
rect 17773 13512 17785 13515
rect 17092 13484 17785 13512
rect 17092 13472 17098 13484
rect 17773 13481 17785 13484
rect 17819 13481 17831 13515
rect 17773 13475 17831 13481
rect 18966 13472 18972 13524
rect 19024 13512 19030 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 19024 13484 19257 13512
rect 19024 13472 19030 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 21174 13472 21180 13524
rect 21232 13512 21238 13524
rect 21361 13515 21419 13521
rect 21361 13512 21373 13515
rect 21232 13484 21373 13512
rect 21232 13472 21238 13484
rect 21361 13481 21373 13484
rect 21407 13481 21419 13515
rect 21361 13475 21419 13481
rect 10134 13444 10140 13456
rect 7024 13416 7880 13444
rect 7944 13416 10140 13444
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 5626 13336 5632 13388
rect 5684 13336 5690 13388
rect 5718 13336 5724 13388
rect 5776 13336 5782 13388
rect 5994 13336 6000 13388
rect 6052 13336 6058 13388
rect 6086 13336 6092 13388
rect 6144 13376 6150 13388
rect 7024 13376 7052 13416
rect 6144 13348 7052 13376
rect 6144 13336 6150 13348
rect 7374 13336 7380 13388
rect 7432 13376 7438 13388
rect 7944 13385 7972 13416
rect 10134 13404 10140 13416
rect 10192 13404 10198 13456
rect 16761 13447 16819 13453
rect 16761 13413 16773 13447
rect 16807 13444 16819 13447
rect 16850 13444 16856 13456
rect 16807 13416 16856 13444
rect 16807 13413 16819 13416
rect 16761 13407 16819 13413
rect 16850 13404 16856 13416
rect 16908 13404 16914 13456
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7432 13348 7481 13376
rect 7432 13336 7438 13348
rect 7469 13345 7481 13348
rect 7515 13376 7527 13379
rect 7929 13379 7987 13385
rect 7929 13376 7941 13379
rect 7515 13348 7941 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 7929 13345 7941 13348
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 8113 13379 8171 13385
rect 8113 13345 8125 13379
rect 8159 13376 8171 13379
rect 8570 13376 8576 13388
rect 8159 13348 8576 13376
rect 8159 13345 8171 13348
rect 8113 13339 8171 13345
rect 8570 13336 8576 13348
rect 8628 13336 8634 13388
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13376 9735 13379
rect 9861 13379 9919 13385
rect 9861 13376 9873 13379
rect 9723 13348 9873 13376
rect 9723 13345 9735 13348
rect 9677 13339 9735 13345
rect 9861 13345 9873 13348
rect 9907 13345 9919 13379
rect 9861 13339 9919 13345
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 10008 13348 10425 13376
rect 10008 13336 10014 13348
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 10413 13339 10471 13345
rect 12250 13336 12256 13388
rect 12308 13336 12314 13388
rect 15930 13336 15936 13388
rect 15988 13376 15994 13388
rect 15988 13348 18184 13376
rect 15988 13336 15994 13348
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4522 13308 4528 13320
rect 4019 13280 4528 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 4982 13308 4988 13320
rect 4663 13280 4988 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 2038 13200 2044 13252
rect 2096 13200 2102 13252
rect 3050 13200 3056 13252
rect 3108 13200 3114 13252
rect 3418 13200 3424 13252
rect 3476 13240 3482 13252
rect 4632 13240 4660 13271
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 3476 13212 4660 13240
rect 3476 13200 3482 13212
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 6086 13240 6092 13252
rect 5408 13212 6092 13240
rect 5408 13200 5414 13212
rect 6086 13200 6092 13212
rect 6144 13200 6150 13252
rect 7006 13200 7012 13252
rect 7064 13200 7070 13252
rect 3970 13132 3976 13184
rect 4028 13132 4034 13184
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 6730 13172 6736 13184
rect 5583 13144 6736 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 8220 13172 8248 13271
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 8481 13311 8539 13317
rect 8481 13308 8493 13311
rect 8352 13280 8493 13308
rect 8352 13268 8358 13280
rect 8481 13277 8493 13280
rect 8527 13308 8539 13311
rect 8662 13308 8668 13320
rect 8527 13280 8668 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9585 13311 9643 13317
rect 9272 13280 9317 13308
rect 9272 13268 9278 13280
rect 9585 13277 9597 13311
rect 9631 13277 9643 13311
rect 9585 13271 9643 13277
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 10042 13308 10048 13320
rect 9815 13280 10048 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 9600 13240 9628 13271
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13308 10195 13311
rect 10226 13308 10232 13320
rect 10183 13280 10232 13308
rect 10183 13277 10195 13280
rect 10137 13271 10195 13277
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10318 13268 10324 13320
rect 10376 13268 10382 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 10686 13308 10692 13320
rect 10643 13280 10692 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 11977 13311 12035 13317
rect 11977 13277 11989 13311
rect 12023 13308 12035 13311
rect 13814 13308 13820 13320
rect 12023 13280 13820 13308
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 15703 13280 16344 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 16316 13252 16344 13280
rect 18156 13252 18184 13348
rect 18230 13336 18236 13388
rect 18288 13336 18294 13388
rect 19794 13336 19800 13388
rect 19852 13376 19858 13388
rect 19981 13379 20039 13385
rect 19981 13376 19993 13379
rect 19852 13348 19993 13376
rect 19852 13336 19858 13348
rect 19981 13345 19993 13348
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 19886 13308 19892 13320
rect 19475 13280 19892 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 20254 13317 20260 13320
rect 20248 13308 20260 13317
rect 20215 13280 20260 13308
rect 20248 13271 20260 13280
rect 20254 13268 20260 13271
rect 20312 13268 20318 13320
rect 10870 13240 10876 13252
rect 9600 13212 10876 13240
rect 10870 13200 10876 13212
rect 10928 13200 10934 13252
rect 12342 13200 12348 13252
rect 12400 13240 12406 13252
rect 12498 13243 12556 13249
rect 12498 13240 12510 13243
rect 12400 13212 12510 13240
rect 12400 13200 12406 13212
rect 12498 13209 12510 13212
rect 12544 13209 12556 13243
rect 12498 13203 12556 13209
rect 14458 13200 14464 13252
rect 14516 13240 14522 13252
rect 15841 13243 15899 13249
rect 15841 13240 15853 13243
rect 14516 13212 15853 13240
rect 14516 13200 14522 13212
rect 15841 13209 15853 13212
rect 15887 13209 15899 13243
rect 15841 13203 15899 13209
rect 16209 13243 16267 13249
rect 16209 13209 16221 13243
rect 16255 13209 16267 13243
rect 16209 13203 16267 13209
rect 9858 13172 9864 13184
rect 8220 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13172 9922 13184
rect 10410 13172 10416 13184
rect 9916 13144 10416 13172
rect 9916 13132 9922 13144
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 15363 13175 15421 13181
rect 15363 13172 15375 13175
rect 14608 13144 15375 13172
rect 14608 13132 14614 13144
rect 15363 13141 15375 13144
rect 15409 13141 15421 13175
rect 16224 13172 16252 13203
rect 16298 13200 16304 13252
rect 16356 13200 16362 13252
rect 16482 13200 16488 13252
rect 16540 13200 16546 13252
rect 18138 13200 18144 13252
rect 18196 13240 18202 13252
rect 18325 13243 18383 13249
rect 18325 13240 18337 13243
rect 18196 13212 18337 13240
rect 18196 13200 18202 13212
rect 18325 13209 18337 13212
rect 18371 13240 18383 13243
rect 20530 13240 20536 13252
rect 18371 13212 20536 13240
rect 18371 13209 18383 13212
rect 18325 13203 18383 13209
rect 20530 13200 20536 13212
rect 20588 13200 20594 13252
rect 16574 13172 16580 13184
rect 16224 13144 16580 13172
rect 15363 13135 15421 13141
rect 16574 13132 16580 13144
rect 16632 13172 16638 13184
rect 17310 13172 17316 13184
rect 16632 13144 17316 13172
rect 16632 13132 16638 13144
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 18230 13132 18236 13184
rect 18288 13172 18294 13184
rect 18414 13172 18420 13184
rect 18288 13144 18420 13172
rect 18288 13132 18294 13144
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 1104 13082 21988 13104
rect 1104 13030 4220 13082
rect 4272 13030 4284 13082
rect 4336 13030 4348 13082
rect 4400 13030 4412 13082
rect 4464 13030 4476 13082
rect 4528 13030 9441 13082
rect 9493 13030 9505 13082
rect 9557 13030 9569 13082
rect 9621 13030 9633 13082
rect 9685 13030 9697 13082
rect 9749 13030 14662 13082
rect 14714 13030 14726 13082
rect 14778 13030 14790 13082
rect 14842 13030 14854 13082
rect 14906 13030 14918 13082
rect 14970 13030 19883 13082
rect 19935 13030 19947 13082
rect 19999 13030 20011 13082
rect 20063 13030 20075 13082
rect 20127 13030 20139 13082
rect 20191 13030 21988 13082
rect 1104 13008 21988 13030
rect 3050 12928 3056 12980
rect 3108 12928 3114 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12937 4215 12971
rect 4157 12931 4215 12937
rect 4341 12971 4399 12977
rect 4341 12937 4353 12971
rect 4387 12968 4399 12971
rect 4706 12968 4712 12980
rect 4387 12940 4712 12968
rect 4387 12937 4399 12940
rect 4341 12931 4399 12937
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12832 3203 12835
rect 3418 12832 3424 12844
rect 3191 12804 3424 12832
rect 3191 12801 3203 12804
rect 3145 12795 3203 12801
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 4172 12764 4200 12931
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5445 12971 5503 12977
rect 5445 12937 5457 12971
rect 5491 12968 5503 12971
rect 5626 12968 5632 12980
rect 5491 12940 5632 12968
rect 5491 12937 5503 12940
rect 5445 12931 5503 12937
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 6454 12928 6460 12980
rect 6512 12928 6518 12980
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7098 12968 7104 12980
rect 6972 12940 7104 12968
rect 6972 12928 6978 12940
rect 7098 12928 7104 12940
rect 7156 12968 7162 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 7156 12940 11897 12968
rect 7156 12928 7162 12940
rect 11885 12937 11897 12940
rect 11931 12937 11943 12971
rect 14737 12971 14795 12977
rect 11885 12931 11943 12937
rect 12406 12940 13308 12968
rect 4525 12903 4583 12909
rect 4525 12869 4537 12903
rect 4571 12900 4583 12903
rect 4614 12900 4620 12912
rect 4571 12872 4620 12900
rect 4571 12869 4583 12872
rect 4525 12863 4583 12869
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 5810 12900 5816 12912
rect 5092 12872 5816 12900
rect 5092 12841 5120 12872
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 6181 12903 6239 12909
rect 6181 12869 6193 12903
rect 6227 12900 6239 12903
rect 6546 12900 6552 12912
rect 6227 12872 6552 12900
rect 6227 12869 6239 12872
rect 6181 12863 6239 12869
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 7282 12860 7288 12912
rect 7340 12860 7346 12912
rect 7377 12903 7435 12909
rect 7377 12869 7389 12903
rect 7423 12900 7435 12903
rect 7466 12900 7472 12912
rect 7423 12872 7472 12900
rect 7423 12869 7435 12872
rect 7377 12863 7435 12869
rect 7466 12860 7472 12872
rect 7524 12900 7530 12912
rect 9306 12900 9312 12912
rect 7524 12872 9312 12900
rect 7524 12860 7530 12872
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5350 12792 5356 12844
rect 5408 12792 5414 12844
rect 5902 12792 5908 12844
rect 5960 12792 5966 12844
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12801 6147 12835
rect 6089 12795 6147 12801
rect 4890 12764 4896 12776
rect 4172 12736 4896 12764
rect 4890 12724 4896 12736
rect 4948 12764 4954 12776
rect 6104 12764 6132 12795
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6638 12832 6644 12844
rect 6328 12804 6644 12832
rect 6328 12792 6334 12804
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 6788 12804 7512 12832
rect 6788 12792 6794 12804
rect 7006 12764 7012 12776
rect 4948 12736 7012 12764
rect 4948 12724 4954 12736
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12764 7343 12767
rect 7374 12764 7380 12776
rect 7331 12736 7380 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 7484 12764 7512 12804
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 8128 12841 8156 12872
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7708 12804 7757 12832
rect 7708 12792 7714 12804
rect 7745 12801 7757 12804
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12832 8447 12835
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 8435 12804 8585 12832
rect 8435 12801 8447 12804
rect 8389 12795 8447 12801
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 8662 12792 8668 12844
rect 8720 12832 8726 12844
rect 9140 12841 9168 12872
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 10134 12900 10140 12912
rect 9876 12872 10140 12900
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8720 12804 8953 12832
rect 8720 12792 8726 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12801 9183 12835
rect 9876 12832 9904 12872
rect 10060 12841 10088 12872
rect 10134 12860 10140 12872
rect 10192 12860 10198 12912
rect 10321 12903 10379 12909
rect 10321 12869 10333 12903
rect 10367 12900 10379 12903
rect 10870 12900 10876 12912
rect 10367 12872 10876 12900
rect 10367 12869 10379 12872
rect 10321 12863 10379 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 12406 12900 12434 12940
rect 10980 12872 12434 12900
rect 9125 12795 9183 12801
rect 9232 12804 9904 12832
rect 10045 12835 10103 12841
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7484 12736 7941 12764
rect 7929 12733 7941 12736
rect 7975 12764 7987 12767
rect 8481 12767 8539 12773
rect 7975 12736 8156 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 6546 12656 6552 12708
rect 6604 12696 6610 12708
rect 7653 12699 7711 12705
rect 7653 12696 7665 12699
rect 6604 12668 7665 12696
rect 6604 12656 6610 12668
rect 7653 12665 7665 12668
rect 7699 12665 7711 12699
rect 7653 12659 7711 12665
rect 3786 12588 3792 12640
rect 3844 12628 3850 12640
rect 4341 12631 4399 12637
rect 4341 12628 4353 12631
rect 3844 12600 4353 12628
rect 3844 12588 3850 12600
rect 4341 12597 4353 12600
rect 4387 12597 4399 12631
rect 4341 12591 4399 12597
rect 4890 12588 4896 12640
rect 4948 12588 4954 12640
rect 5718 12588 5724 12640
rect 5776 12588 5782 12640
rect 6822 12588 6828 12640
rect 6880 12588 6886 12640
rect 8128 12628 8156 12736
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 8680 12764 8708 12792
rect 8527 12736 8708 12764
rect 8956 12764 8984 12795
rect 9232 12764 9260 12804
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10505 12795 10563 12801
rect 10612 12804 10701 12832
rect 8956 12736 9260 12764
rect 9769 12767 9827 12773
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 9769 12733 9781 12767
rect 9815 12733 9827 12767
rect 9769 12727 9827 12733
rect 8570 12656 8576 12708
rect 8628 12696 8634 12708
rect 8665 12699 8723 12705
rect 8665 12696 8677 12699
rect 8628 12668 8677 12696
rect 8628 12656 8634 12668
rect 8665 12665 8677 12668
rect 8711 12665 8723 12699
rect 9784 12696 9812 12727
rect 9858 12724 9864 12776
rect 9916 12724 9922 12776
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12764 10011 12767
rect 10226 12764 10232 12776
rect 9999 12736 10232 12764
rect 9999 12733 10011 12736
rect 9953 12727 10011 12733
rect 10226 12724 10232 12736
rect 10284 12764 10290 12776
rect 10520 12764 10548 12795
rect 10284 12736 10548 12764
rect 10284 12724 10290 12736
rect 10612 12708 10640 12804
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 10980 12832 11008 12872
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 13170 12900 13176 12912
rect 12768 12872 13176 12900
rect 12768 12860 12774 12872
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 13280 12909 13308 12940
rect 14737 12937 14749 12971
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 16209 12971 16267 12977
rect 16209 12937 16221 12971
rect 16255 12968 16267 12971
rect 16298 12968 16304 12980
rect 16255 12940 16304 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 13265 12903 13323 12909
rect 13265 12869 13277 12903
rect 13311 12900 13323 12903
rect 14752 12900 14780 12931
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 18046 12928 18052 12980
rect 18104 12928 18110 12980
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 20346 12968 20352 12980
rect 20303 12940 20352 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 20346 12928 20352 12940
rect 20404 12928 20410 12980
rect 15074 12903 15132 12909
rect 15074 12900 15086 12903
rect 13311 12872 14688 12900
rect 14752 12872 15086 12900
rect 13311 12869 13323 12872
rect 13265 12863 13323 12869
rect 10836 12804 11008 12832
rect 10836 12792 10842 12804
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 11848 12804 12173 12832
rect 11848 12792 11854 12804
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 12526 12792 12532 12844
rect 12584 12792 12590 12844
rect 14550 12792 14556 12844
rect 14608 12792 14614 12844
rect 14660 12832 14688 12872
rect 15074 12869 15086 12872
rect 15120 12869 15132 12903
rect 15074 12863 15132 12869
rect 18138 12860 18144 12912
rect 18196 12860 18202 12912
rect 18506 12900 18512 12912
rect 18432 12872 18512 12900
rect 14660 12804 15884 12832
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12764 12403 12767
rect 12986 12764 12992 12776
rect 12391 12736 12992 12764
rect 12391 12733 12403 12736
rect 12345 12727 12403 12733
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 13262 12724 13268 12776
rect 13320 12724 13326 12776
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 14829 12767 14887 12773
rect 14829 12764 14841 12767
rect 14424 12736 14841 12764
rect 14424 12724 14430 12736
rect 14829 12733 14841 12736
rect 14875 12733 14887 12767
rect 14829 12727 14887 12733
rect 10042 12696 10048 12708
rect 9784 12668 10048 12696
rect 8665 12659 8723 12665
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 10134 12656 10140 12708
rect 10192 12696 10198 12708
rect 10318 12696 10324 12708
rect 10192 12668 10324 12696
rect 10192 12656 10198 12668
rect 10318 12656 10324 12668
rect 10376 12696 10382 12708
rect 10594 12696 10600 12708
rect 10376 12668 10600 12696
rect 10376 12656 10382 12668
rect 10594 12656 10600 12668
rect 10652 12656 10658 12708
rect 12253 12699 12311 12705
rect 12253 12665 12265 12699
rect 12299 12696 12311 12699
rect 13630 12696 13636 12708
rect 12299 12668 13636 12696
rect 12299 12665 12311 12668
rect 12253 12659 12311 12665
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 13722 12656 13728 12708
rect 13780 12656 13786 12708
rect 15856 12696 15884 12804
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 18432 12832 18460 12872
rect 18506 12860 18512 12872
rect 18564 12900 18570 12912
rect 18877 12903 18935 12909
rect 18877 12900 18889 12903
rect 18564 12872 18889 12900
rect 18564 12860 18570 12872
rect 18877 12869 18889 12872
rect 18923 12869 18935 12903
rect 18877 12863 18935 12869
rect 20441 12903 20499 12909
rect 20441 12869 20453 12903
rect 20487 12900 20499 12903
rect 21174 12900 21180 12912
rect 20487 12872 21180 12900
rect 20487 12869 20499 12872
rect 20441 12863 20499 12869
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 18064 12804 18460 12832
rect 18064 12773 18092 12804
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 18656 12804 18705 12832
rect 18656 12792 18662 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12832 20223 12835
rect 20346 12832 20352 12844
rect 20211 12804 20352 12832
rect 20211 12801 20223 12804
rect 20165 12795 20223 12801
rect 20346 12792 20352 12804
rect 20404 12832 20410 12844
rect 20530 12832 20536 12844
rect 20404 12804 20536 12832
rect 20404 12792 20410 12804
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 18966 12724 18972 12776
rect 19024 12724 19030 12776
rect 18230 12696 18236 12708
rect 15856 12668 18236 12696
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 20714 12656 20720 12708
rect 20772 12656 20778 12708
rect 9214 12628 9220 12640
rect 8128 12600 9220 12628
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 10226 12588 10232 12640
rect 10284 12588 10290 12640
rect 12434 12588 12440 12640
rect 12492 12588 12498 12640
rect 16666 12588 16672 12640
rect 16724 12588 16730 12640
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17589 12631 17647 12637
rect 17589 12628 17601 12631
rect 16908 12600 17601 12628
rect 16908 12588 16914 12600
rect 17589 12597 17601 12600
rect 17635 12597 17647 12631
rect 17589 12591 17647 12597
rect 18414 12588 18420 12640
rect 18472 12588 18478 12640
rect 1104 12538 21988 12560
rect 1104 12486 3560 12538
rect 3612 12486 3624 12538
rect 3676 12486 3688 12538
rect 3740 12486 3752 12538
rect 3804 12486 3816 12538
rect 3868 12486 8781 12538
rect 8833 12486 8845 12538
rect 8897 12486 8909 12538
rect 8961 12486 8973 12538
rect 9025 12486 9037 12538
rect 9089 12486 14002 12538
rect 14054 12486 14066 12538
rect 14118 12486 14130 12538
rect 14182 12486 14194 12538
rect 14246 12486 14258 12538
rect 14310 12486 19223 12538
rect 19275 12486 19287 12538
rect 19339 12486 19351 12538
rect 19403 12486 19415 12538
rect 19467 12486 19479 12538
rect 19531 12486 21988 12538
rect 1104 12464 21988 12486
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 6733 12427 6791 12433
rect 6733 12424 6745 12427
rect 6696 12396 6745 12424
rect 6696 12384 6702 12396
rect 6733 12393 6745 12396
rect 6779 12393 6791 12427
rect 6733 12387 6791 12393
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 9180 12396 10548 12424
rect 9180 12384 9186 12396
rect 2409 12359 2467 12365
rect 2409 12325 2421 12359
rect 2455 12325 2467 12359
rect 9033 12359 9091 12365
rect 9033 12356 9045 12359
rect 2409 12319 2467 12325
rect 8588 12328 9045 12356
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2424 12220 2452 12319
rect 2866 12248 2872 12300
rect 2924 12248 2930 12300
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 4985 12291 5043 12297
rect 4985 12288 4997 12291
rect 4672 12260 4997 12288
rect 4672 12248 4678 12260
rect 4985 12257 4997 12260
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 5718 12288 5724 12300
rect 5307 12260 5724 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 7432 12260 7941 12288
rect 7432 12248 7438 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 2179 12192 2452 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 2832 12192 4353 12220
rect 2832 12180 2838 12192
rect 4341 12189 4353 12192
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7248 12192 7665 12220
rect 7248 12180 7254 12192
rect 7653 12189 7665 12192
rect 7699 12220 7711 12223
rect 8202 12220 8208 12232
rect 7699 12192 8208 12220
rect 7699 12189 7711 12192
rect 7653 12183 7711 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8478 12180 8484 12232
rect 8536 12180 8542 12232
rect 8588 12229 8616 12328
rect 9033 12325 9045 12328
rect 9079 12356 9091 12359
rect 9858 12356 9864 12368
rect 9079 12328 9864 12356
rect 9079 12325 9091 12328
rect 9033 12319 9091 12325
rect 9858 12316 9864 12328
rect 9916 12356 9922 12368
rect 10410 12356 10416 12368
rect 9916 12328 10416 12356
rect 9916 12316 9922 12328
rect 10410 12316 10416 12328
rect 10468 12316 10474 12368
rect 10520 12356 10548 12396
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 11149 12427 11207 12433
rect 11149 12424 11161 12427
rect 10652 12396 11161 12424
rect 10652 12384 10658 12396
rect 11149 12393 11161 12396
rect 11195 12393 11207 12427
rect 11149 12387 11207 12393
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12986 12424 12992 12436
rect 12492 12396 12992 12424
rect 12492 12384 12498 12396
rect 12986 12384 12992 12396
rect 13044 12424 13050 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13044 12396 13737 12424
rect 13044 12384 13050 12396
rect 13725 12393 13737 12396
rect 13771 12393 13783 12427
rect 13725 12387 13783 12393
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16482 12424 16488 12436
rect 16347 12396 16488 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 18414 12424 18420 12436
rect 16592 12396 18420 12424
rect 10781 12359 10839 12365
rect 10781 12356 10793 12359
rect 10520 12328 10793 12356
rect 10781 12325 10793 12328
rect 10827 12325 10839 12359
rect 10781 12319 10839 12325
rect 10597 12291 10655 12297
rect 10597 12288 10609 12291
rect 9416 12260 10609 12288
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12189 8631 12223
rect 8573 12183 8631 12189
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 9416 12229 9444 12260
rect 10597 12257 10609 12260
rect 10643 12288 10655 12291
rect 10643 12260 11008 12288
rect 10643 12257 10655 12260
rect 10597 12251 10655 12257
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 9364 12192 9413 12220
rect 9364 12180 9370 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10100 12192 10149 12220
rect 10100 12180 10106 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10410 12180 10416 12232
rect 10468 12180 10474 12232
rect 10980 12229 11008 12260
rect 13262 12248 13268 12300
rect 13320 12248 13326 12300
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 11112 12192 11437 12220
rect 11112 12180 11118 12192
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 11514 12180 11520 12232
rect 11572 12180 11578 12232
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 13817 12223 13875 12229
rect 13817 12220 13829 12223
rect 13780 12192 13829 12220
rect 13780 12180 13786 12192
rect 13817 12189 13829 12192
rect 13863 12189 13875 12223
rect 13817 12183 13875 12189
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12220 14979 12223
rect 15010 12220 15016 12232
rect 14967 12192 15016 12220
rect 14967 12189 14979 12192
rect 14921 12183 14979 12189
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 16592 12229 16620 12396
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 18509 12359 18567 12365
rect 18509 12325 18521 12359
rect 18555 12356 18567 12359
rect 18598 12356 18604 12368
rect 18555 12328 18604 12356
rect 18555 12325 18567 12328
rect 18509 12319 18567 12325
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 18966 12316 18972 12368
rect 19024 12356 19030 12368
rect 21177 12359 21235 12365
rect 19024 12328 19334 12356
rect 19024 12316 19030 12328
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 16850 12180 16856 12232
rect 16908 12180 16914 12232
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 19306 12220 19334 12328
rect 21177 12325 21189 12359
rect 21223 12356 21235 12359
rect 21266 12356 21272 12368
rect 21223 12328 21272 12356
rect 21223 12325 21235 12328
rect 21177 12319 21235 12325
rect 21266 12316 21272 12328
rect 21324 12316 21330 12368
rect 19702 12248 19708 12300
rect 19760 12288 19766 12300
rect 20257 12291 20315 12297
rect 20257 12288 20269 12291
rect 19760 12260 20269 12288
rect 19760 12248 19766 12260
rect 20257 12257 20269 12260
rect 20303 12288 20315 12291
rect 20438 12288 20444 12300
rect 20303 12260 20444 12288
rect 20303 12257 20315 12260
rect 20257 12251 20315 12257
rect 20438 12248 20444 12260
rect 20496 12248 20502 12300
rect 20530 12220 20536 12232
rect 19306 12192 20536 12220
rect 20530 12180 20536 12192
rect 20588 12220 20594 12232
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 20588 12192 20637 12220
rect 20588 12180 20594 12192
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 2961 12155 3019 12161
rect 2961 12121 2973 12155
rect 3007 12152 3019 12155
rect 3050 12152 3056 12164
rect 3007 12124 3056 12152
rect 3007 12121 3019 12124
rect 2961 12115 3019 12121
rect 3050 12112 3056 12124
rect 3108 12152 3114 12164
rect 4617 12155 4675 12161
rect 4617 12152 4629 12155
rect 3108 12124 4629 12152
rect 3108 12112 3114 12124
rect 4617 12121 4629 12124
rect 4663 12152 4675 12155
rect 4890 12152 4896 12164
rect 4663 12124 4896 12152
rect 4663 12121 4675 12124
rect 4617 12115 4675 12121
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 6546 12152 6552 12164
rect 6486 12124 6552 12152
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 9784 12152 9812 12180
rect 10318 12152 10324 12164
rect 9784 12124 10324 12152
rect 10318 12112 10324 12124
rect 10376 12152 10382 12164
rect 10505 12155 10563 12161
rect 10505 12152 10517 12155
rect 10376 12124 10517 12152
rect 10376 12112 10382 12124
rect 10505 12121 10517 12124
rect 10551 12121 10563 12155
rect 10505 12115 10563 12121
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 13170 12152 13176 12164
rect 12676 12124 13176 12152
rect 12676 12112 12682 12124
rect 13170 12112 13176 12124
rect 13228 12112 13234 12164
rect 15188 12155 15246 12161
rect 15188 12121 15200 12155
rect 15234 12152 15246 12155
rect 16666 12152 16672 12164
rect 15234 12124 16672 12152
rect 15234 12121 15246 12124
rect 15188 12115 15246 12121
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 17374 12155 17432 12161
rect 17374 12152 17386 12155
rect 16776 12124 17386 12152
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 1949 12087 2007 12093
rect 1949 12084 1961 12087
rect 1912 12056 1961 12084
rect 1912 12044 1918 12056
rect 1949 12053 1961 12056
rect 1995 12053 2007 12087
rect 1949 12047 2007 12053
rect 2866 12044 2872 12096
rect 2924 12044 2930 12096
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 4047 12087 4105 12093
rect 4047 12084 4059 12087
rect 3384 12056 4059 12084
rect 3384 12044 3390 12056
rect 4047 12053 4059 12056
rect 4093 12053 4105 12087
rect 4047 12047 4105 12053
rect 4525 12087 4583 12093
rect 4525 12053 4537 12087
rect 4571 12084 4583 12087
rect 4982 12084 4988 12096
rect 4571 12056 4988 12084
rect 4571 12053 4583 12056
rect 4525 12047 4583 12053
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 7742 12044 7748 12096
rect 7800 12044 7806 12096
rect 8110 12044 8116 12096
rect 8168 12044 8174 12096
rect 9950 12044 9956 12096
rect 10008 12044 10014 12096
rect 11238 12044 11244 12096
rect 11296 12044 11302 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 12434 12084 12440 12096
rect 11388 12056 12440 12084
rect 11388 12044 11394 12056
rect 12434 12044 12440 12056
rect 12492 12084 12498 12096
rect 12710 12084 12716 12096
rect 12492 12056 12716 12084
rect 12492 12044 12498 12056
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 16776 12093 16804 12124
rect 17374 12121 17386 12124
rect 17420 12121 17432 12155
rect 17374 12115 17432 12121
rect 20349 12155 20407 12161
rect 20349 12121 20361 12155
rect 20395 12152 20407 12155
rect 20806 12152 20812 12164
rect 20395 12124 20812 12152
rect 20395 12121 20407 12124
rect 20349 12115 20407 12121
rect 20806 12112 20812 12124
rect 20864 12112 20870 12164
rect 20901 12155 20959 12161
rect 20901 12121 20913 12155
rect 20947 12152 20959 12155
rect 21358 12152 21364 12164
rect 20947 12124 21364 12152
rect 20947 12121 20959 12124
rect 20901 12115 20959 12121
rect 21358 12112 21364 12124
rect 21416 12112 21422 12164
rect 13541 12087 13599 12093
rect 13541 12084 13553 12087
rect 13504 12056 13553 12084
rect 13504 12044 13510 12056
rect 13541 12053 13553 12056
rect 13587 12053 13599 12087
rect 13541 12047 13599 12053
rect 16761 12087 16819 12093
rect 16761 12053 16773 12087
rect 16807 12053 16819 12087
rect 16761 12047 16819 12053
rect 17034 12044 17040 12096
rect 17092 12044 17098 12096
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19779 12087 19837 12093
rect 19779 12084 19791 12087
rect 19300 12056 19791 12084
rect 19300 12044 19306 12056
rect 19779 12053 19791 12056
rect 19825 12053 19837 12087
rect 19779 12047 19837 12053
rect 20257 12087 20315 12093
rect 20257 12053 20269 12087
rect 20303 12084 20315 12087
rect 20714 12084 20720 12096
rect 20303 12056 20720 12084
rect 20303 12053 20315 12056
rect 20257 12047 20315 12053
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 1104 11994 21988 12016
rect 1104 11942 4220 11994
rect 4272 11942 4284 11994
rect 4336 11942 4348 11994
rect 4400 11942 4412 11994
rect 4464 11942 4476 11994
rect 4528 11942 9441 11994
rect 9493 11942 9505 11994
rect 9557 11942 9569 11994
rect 9621 11942 9633 11994
rect 9685 11942 9697 11994
rect 9749 11942 14662 11994
rect 14714 11942 14726 11994
rect 14778 11942 14790 11994
rect 14842 11942 14854 11994
rect 14906 11942 14918 11994
rect 14970 11942 19883 11994
rect 19935 11942 19947 11994
rect 19999 11942 20011 11994
rect 20063 11942 20075 11994
rect 20127 11942 20139 11994
rect 20191 11942 21988 11994
rect 1104 11920 21988 11942
rect 3513 11883 3571 11889
rect 3513 11849 3525 11883
rect 3559 11849 3571 11883
rect 3513 11843 3571 11849
rect 3528 11812 3556 11843
rect 9306 11840 9312 11892
rect 9364 11840 9370 11892
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10137 11883 10195 11889
rect 10137 11880 10149 11883
rect 10100 11852 10149 11880
rect 10100 11840 10106 11852
rect 10137 11849 10149 11852
rect 10183 11849 10195 11883
rect 10137 11843 10195 11849
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 11701 11883 11759 11889
rect 11701 11880 11713 11883
rect 10652 11852 11713 11880
rect 10652 11840 10658 11852
rect 11701 11849 11713 11852
rect 11747 11849 11759 11883
rect 13262 11880 13268 11892
rect 11701 11843 11759 11849
rect 11900 11852 13268 11880
rect 3850 11815 3908 11821
rect 3850 11812 3862 11815
rect 1596 11784 2774 11812
rect 3528 11784 3862 11812
rect 1596 11753 1624 11784
rect 1854 11753 1860 11756
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1848 11744 1860 11753
rect 1815 11716 1860 11744
rect 1581 11707 1639 11713
rect 1848 11707 1860 11716
rect 1854 11704 1860 11707
rect 1912 11704 1918 11756
rect 2746 11676 2774 11784
rect 3850 11781 3862 11784
rect 3896 11781 3908 11815
rect 3850 11775 3908 11781
rect 7742 11772 7748 11824
rect 7800 11812 7806 11824
rect 7800 11784 8326 11812
rect 7800 11772 7806 11784
rect 3326 11704 3332 11756
rect 3384 11704 3390 11756
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 5353 11747 5411 11753
rect 5353 11744 5365 11747
rect 5132 11716 5365 11744
rect 5132 11704 5138 11716
rect 5353 11713 5365 11716
rect 5399 11713 5411 11747
rect 9324 11744 9352 11840
rect 10229 11815 10287 11821
rect 10229 11781 10241 11815
rect 10275 11812 10287 11815
rect 10318 11812 10324 11824
rect 10275 11784 10324 11812
rect 10275 11781 10287 11784
rect 10229 11775 10287 11781
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 11146 11772 11152 11824
rect 11204 11772 11210 11824
rect 11241 11815 11299 11821
rect 11241 11781 11253 11815
rect 11287 11812 11299 11815
rect 11330 11812 11336 11824
rect 11287 11784 11336 11812
rect 11287 11781 11299 11784
rect 11241 11775 11299 11781
rect 11330 11772 11336 11784
rect 11388 11772 11394 11824
rect 11900 11753 11928 11852
rect 13262 11840 13268 11852
rect 13320 11880 13326 11892
rect 13722 11880 13728 11892
rect 13320 11852 13728 11880
rect 13320 11840 13326 11852
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 15289 11883 15347 11889
rect 15289 11849 15301 11883
rect 15335 11880 15347 11883
rect 15930 11880 15936 11892
rect 15335 11852 15936 11880
rect 15335 11849 15347 11852
rect 15289 11843 15347 11849
rect 15930 11840 15936 11852
rect 15988 11840 15994 11892
rect 18506 11840 18512 11892
rect 18564 11840 18570 11892
rect 19429 11883 19487 11889
rect 19429 11849 19441 11883
rect 19475 11849 19487 11883
rect 19429 11843 19487 11849
rect 11992 11784 15148 11812
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 9324 11716 10057 11744
rect 5353 11707 5411 11713
rect 10045 11713 10057 11716
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 3605 11679 3663 11685
rect 3605 11676 3617 11679
rect 2746 11648 3617 11676
rect 3605 11645 3617 11648
rect 3651 11645 3663 11679
rect 3605 11639 3663 11645
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11676 7895 11679
rect 8570 11676 8576 11688
rect 7883 11648 8576 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 2958 11500 2964 11552
rect 3016 11500 3022 11552
rect 3620 11540 3648 11639
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 6086 11608 6092 11620
rect 5040 11580 6092 11608
rect 5040 11568 5046 11580
rect 6086 11568 6092 11580
rect 6144 11568 6150 11620
rect 4614 11540 4620 11552
rect 3620 11512 4620 11540
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 5166 11500 5172 11552
rect 5224 11500 5230 11552
rect 7576 11540 7604 11639
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9582 11676 9588 11688
rect 9539 11648 9588 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 9858 11676 9864 11688
rect 9723 11648 9864 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11676 11207 11679
rect 11195 11648 11468 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 11054 11608 11060 11620
rect 10735 11580 11060 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 11054 11568 11060 11580
rect 11112 11568 11118 11620
rect 10502 11540 10508 11552
rect 7576 11512 10508 11540
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 11440 11540 11468 11648
rect 11532 11608 11560 11707
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 11992 11676 12020 11784
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11744 12219 11747
rect 12207 11716 12572 11744
rect 12207 11713 12219 11716
rect 12161 11707 12219 11713
rect 12544 11688 12572 11716
rect 13446 11704 13452 11756
rect 13504 11753 13510 11756
rect 13504 11744 13516 11753
rect 13504 11716 13549 11744
rect 13504 11707 13516 11716
rect 13504 11704 13510 11707
rect 13814 11704 13820 11756
rect 13872 11704 13878 11756
rect 15120 11753 15148 11784
rect 16022 11772 16028 11824
rect 16080 11772 16086 11824
rect 17034 11772 17040 11824
rect 17092 11812 17098 11824
rect 17374 11815 17432 11821
rect 17374 11812 17386 11815
rect 17092 11784 17386 11812
rect 17092 11772 17098 11784
rect 17374 11781 17386 11784
rect 17420 11781 17432 11815
rect 19444 11812 19472 11843
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 20772 11852 20913 11880
rect 20772 11840 20778 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 20901 11843 20959 11849
rect 19766 11815 19824 11821
rect 19766 11812 19778 11815
rect 19444 11784 19778 11812
rect 17374 11775 17432 11781
rect 19766 11781 19778 11784
rect 19812 11781 19824 11815
rect 19766 11775 19824 11781
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11713 15163 11747
rect 15105 11707 15163 11713
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 15712 11716 15853 11744
rect 15712 11704 15718 11716
rect 15841 11713 15853 11716
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 16482 11704 16488 11756
rect 16540 11704 16546 11756
rect 17126 11704 17132 11756
rect 17184 11704 17190 11756
rect 19242 11704 19248 11756
rect 19300 11704 19306 11756
rect 21266 11704 21272 11756
rect 21324 11704 21330 11756
rect 11664 11648 12020 11676
rect 11664 11636 11670 11648
rect 12526 11636 12532 11688
rect 12584 11636 12590 11688
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 13771 11648 15148 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 15120 11620 15148 11648
rect 16114 11636 16120 11688
rect 16172 11636 16178 11688
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19521 11679 19579 11685
rect 19521 11676 19533 11679
rect 19116 11648 19533 11676
rect 19116 11636 19122 11648
rect 19521 11645 19533 11648
rect 19567 11645 19579 11679
rect 19521 11639 19579 11645
rect 12345 11611 12403 11617
rect 12345 11608 12357 11611
rect 11532 11580 12357 11608
rect 12345 11577 12357 11580
rect 12391 11577 12403 11611
rect 12345 11571 12403 11577
rect 11882 11540 11888 11552
rect 11440 11512 11888 11540
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 12360 11540 12388 11571
rect 15102 11568 15108 11620
rect 15160 11568 15166 11620
rect 12618 11540 12624 11552
rect 12360 11512 12624 11540
rect 12618 11500 12624 11512
rect 12676 11540 12682 11552
rect 13078 11540 13084 11552
rect 12676 11512 13084 11540
rect 12676 11500 12682 11512
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 14001 11543 14059 11549
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 14366 11540 14372 11552
rect 14047 11512 14372 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 15562 11500 15568 11552
rect 15620 11500 15626 11552
rect 16298 11500 16304 11552
rect 16356 11500 16362 11552
rect 21082 11500 21088 11552
rect 21140 11500 21146 11552
rect 1104 11450 21988 11472
rect 1104 11398 3560 11450
rect 3612 11398 3624 11450
rect 3676 11398 3688 11450
rect 3740 11398 3752 11450
rect 3804 11398 3816 11450
rect 3868 11398 8781 11450
rect 8833 11398 8845 11450
rect 8897 11398 8909 11450
rect 8961 11398 8973 11450
rect 9025 11398 9037 11450
rect 9089 11398 14002 11450
rect 14054 11398 14066 11450
rect 14118 11398 14130 11450
rect 14182 11398 14194 11450
rect 14246 11398 14258 11450
rect 14310 11398 19223 11450
rect 19275 11398 19287 11450
rect 19339 11398 19351 11450
rect 19403 11398 19415 11450
rect 19467 11398 19479 11450
rect 19531 11398 21988 11450
rect 1104 11376 21988 11398
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11336 4399 11339
rect 4798 11336 4804 11348
rect 4387 11308 4804 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 7098 11336 7104 11348
rect 4948 11308 7104 11336
rect 4948 11296 4954 11308
rect 7098 11296 7104 11308
rect 7156 11336 7162 11348
rect 8294 11336 8300 11348
rect 7156 11308 8300 11336
rect 7156 11296 7162 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 9769 11339 9827 11345
rect 9769 11305 9781 11339
rect 9815 11305 9827 11339
rect 9769 11299 9827 11305
rect 10597 11339 10655 11345
rect 10597 11305 10609 11339
rect 10643 11336 10655 11339
rect 11606 11336 11612 11348
rect 10643 11308 11612 11336
rect 10643 11305 10655 11308
rect 10597 11299 10655 11305
rect 1673 11271 1731 11277
rect 1673 11237 1685 11271
rect 1719 11237 1731 11271
rect 1673 11231 1731 11237
rect 1688 11200 1716 11231
rect 6638 11228 6644 11280
rect 6696 11228 6702 11280
rect 7282 11228 7288 11280
rect 7340 11228 7346 11280
rect 9214 11228 9220 11280
rect 9272 11228 9278 11280
rect 9784 11268 9812 11299
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 12345 11339 12403 11345
rect 12345 11336 12357 11339
rect 11940 11308 12357 11336
rect 11940 11296 11946 11308
rect 12345 11305 12357 11308
rect 12391 11305 12403 11339
rect 12345 11299 12403 11305
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13354 11336 13360 11348
rect 13311 11308 13360 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 9784 11240 10640 11268
rect 6914 11200 6920 11212
rect 1688 11172 1900 11200
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11101 1547 11135
rect 1489 11095 1547 11101
rect 1504 11064 1532 11095
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 1765 11135 1823 11141
rect 1765 11132 1777 11135
rect 1728 11104 1777 11132
rect 1728 11092 1734 11104
rect 1765 11101 1777 11104
rect 1811 11101 1823 11135
rect 1872 11132 1900 11172
rect 3988 11172 4476 11200
rect 2021 11135 2079 11141
rect 2021 11132 2033 11135
rect 1872 11104 2033 11132
rect 1765 11095 1823 11101
rect 2021 11101 2033 11104
rect 2067 11101 2079 11135
rect 2021 11095 2079 11101
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 3988 11141 4016 11172
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3016 11104 3801 11132
rect 3016 11092 3022 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4209 11135 4267 11141
rect 4209 11101 4221 11135
rect 4255 11132 4267 11135
rect 4255 11104 4384 11132
rect 4255 11101 4267 11104
rect 4209 11095 4267 11101
rect 3326 11064 3332 11076
rect 1504 11036 3332 11064
rect 3326 11024 3332 11036
rect 3384 11024 3390 11076
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11033 4123 11067
rect 4065 11027 4123 11033
rect 3145 10999 3203 11005
rect 3145 10965 3157 10999
rect 3191 10996 3203 10999
rect 3786 10996 3792 11008
rect 3191 10968 3792 10996
rect 3191 10965 3203 10968
rect 3145 10959 3203 10965
rect 3786 10956 3792 10968
rect 3844 10996 3850 11008
rect 4080 10996 4108 11027
rect 3844 10968 4108 10996
rect 4356 10996 4384 11104
rect 4448 11064 4476 11172
rect 6288 11172 6920 11200
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 4614 11132 4620 11144
rect 4571 11104 4620 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 4792 11135 4850 11141
rect 4792 11101 4804 11135
rect 4838 11132 4850 11135
rect 5166 11132 5172 11144
rect 4838 11104 5172 11132
rect 4838 11101 4850 11104
rect 4792 11095 4850 11101
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 5350 11064 5356 11076
rect 4448 11036 5356 11064
rect 5350 11024 5356 11036
rect 5408 11064 5414 11076
rect 6288 11073 6316 11172
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 9122 11200 9128 11212
rect 8588 11172 9128 11200
rect 6509 11135 6567 11141
rect 6509 11101 6521 11135
rect 6555 11132 6567 11135
rect 7024 11132 7236 11134
rect 8588 11132 8616 11172
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 9232 11200 9260 11228
rect 10612 11212 10640 11240
rect 9375 11203 9433 11209
rect 9375 11200 9387 11203
rect 9232 11172 9387 11200
rect 9375 11169 9387 11172
rect 9421 11169 9433 11203
rect 9950 11200 9956 11212
rect 9375 11163 9433 11169
rect 9508 11172 9956 11200
rect 6555 11106 8616 11132
rect 6555 11104 7052 11106
rect 7208 11104 8616 11106
rect 8665 11135 8723 11141
rect 6555 11101 6567 11104
rect 6509 11095 6567 11101
rect 8665 11101 8677 11135
rect 8711 11132 8723 11135
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 8711 11104 9229 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 9217 11101 9229 11104
rect 9263 11132 9275 11135
rect 9508 11132 9536 11172
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 10226 11160 10232 11212
rect 10284 11160 10290 11212
rect 10594 11160 10600 11212
rect 10652 11160 10658 11212
rect 9263 11104 9536 11132
rect 9585 11135 9643 11141
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 9585 11101 9597 11135
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11132 10103 11135
rect 10244 11132 10272 11160
rect 10091 11104 10272 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 6273 11067 6331 11073
rect 6273 11064 6285 11067
rect 5408 11036 6285 11064
rect 5408 11024 5414 11036
rect 6273 11033 6285 11036
rect 6319 11033 6331 11067
rect 6273 11027 6331 11033
rect 6365 11067 6423 11073
rect 6365 11033 6377 11067
rect 6411 11064 6423 11067
rect 6411 11036 6500 11064
rect 6411 11033 6423 11036
rect 6365 11027 6423 11033
rect 4890 10996 4896 11008
rect 4356 10968 4896 10996
rect 3844 10956 3850 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 5905 10999 5963 11005
rect 5905 10996 5917 10999
rect 5592 10968 5917 10996
rect 5592 10956 5598 10968
rect 5905 10965 5917 10968
rect 5951 10996 5963 10999
rect 6472 10996 6500 11036
rect 6914 11024 6920 11076
rect 6972 11024 6978 11076
rect 7098 11024 7104 11076
rect 7156 11024 7162 11076
rect 8113 11067 8171 11073
rect 8113 11033 8125 11067
rect 8159 11064 8171 11067
rect 9600 11064 9628 11095
rect 10318 11092 10324 11144
rect 10376 11132 10382 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 10376 11104 10425 11132
rect 10376 11092 10382 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10502 11092 10508 11144
rect 10560 11132 10566 11144
rect 11238 11141 11244 11144
rect 10965 11135 11023 11141
rect 10965 11132 10977 11135
rect 10560 11104 10977 11132
rect 10560 11092 10566 11104
rect 10965 11101 10977 11104
rect 11011 11101 11023 11135
rect 11232 11132 11244 11141
rect 11199 11104 11244 11132
rect 10965 11095 11023 11101
rect 11232 11095 11244 11104
rect 11238 11092 11244 11095
rect 11296 11092 11302 11144
rect 12360 11132 12388 11299
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 12802 11228 12808 11280
rect 12860 11268 12866 11280
rect 13630 11268 13636 11280
rect 12860 11240 13636 11268
rect 12860 11228 12866 11240
rect 13630 11228 13636 11240
rect 13688 11268 13694 11280
rect 13740 11268 13768 11299
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14185 11339 14243 11345
rect 14185 11336 14197 11339
rect 13872 11308 14197 11336
rect 13872 11296 13878 11308
rect 14185 11305 14197 11308
rect 14231 11305 14243 11339
rect 14185 11299 14243 11305
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 16540 11308 16773 11336
rect 16540 11296 16546 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 20714 11336 20720 11348
rect 16761 11299 16819 11305
rect 16868 11308 20720 11336
rect 13688 11240 13768 11268
rect 13688 11228 13694 11240
rect 16114 11228 16120 11280
rect 16172 11268 16178 11280
rect 16868 11268 16896 11308
rect 16172 11240 16896 11268
rect 16172 11228 16178 11240
rect 17586 11228 17592 11280
rect 17644 11268 17650 11280
rect 17681 11271 17739 11277
rect 17681 11268 17693 11271
rect 17644 11240 17693 11268
rect 17644 11228 17650 11240
rect 17681 11237 17693 11240
rect 17727 11237 17739 11271
rect 17681 11231 17739 11237
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 13320 11172 14565 11200
rect 13320 11160 13326 11172
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 17218 11200 17224 11212
rect 16632 11172 17224 11200
rect 16632 11160 16638 11172
rect 17218 11160 17224 11172
rect 17276 11160 17282 11212
rect 18248 11209 18276 11308
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 21358 11296 21364 11348
rect 21416 11296 21422 11348
rect 18233 11203 18291 11209
rect 18233 11169 18245 11203
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 19058 11160 19064 11212
rect 19116 11200 19122 11212
rect 19981 11203 20039 11209
rect 19981 11200 19993 11203
rect 19116 11172 19993 11200
rect 19116 11160 19122 11172
rect 19981 11169 19993 11172
rect 20027 11169 20039 11203
rect 19981 11163 20039 11169
rect 13633 11135 13691 11141
rect 13633 11132 13645 11135
rect 12360 11104 13645 11132
rect 13633 11101 13645 11104
rect 13679 11101 13691 11135
rect 13633 11095 13691 11101
rect 15102 11092 15108 11144
rect 15160 11092 15166 11144
rect 15372 11135 15430 11141
rect 15372 11101 15384 11135
rect 15418 11132 15430 11135
rect 16298 11132 16304 11144
rect 15418 11104 16304 11132
rect 15418 11101 15430 11104
rect 15372 11095 15430 11101
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 19705 11135 19763 11141
rect 16408 11104 17172 11132
rect 10778 11064 10784 11076
rect 8159 11036 8616 11064
rect 9600 11036 10784 11064
rect 8159 11033 8171 11036
rect 8113 11027 8171 11033
rect 5951 10968 6500 10996
rect 6932 10996 6960 11024
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 6932 10968 7849 10996
rect 5951 10965 5963 10968
rect 5905 10959 5963 10965
rect 7837 10965 7849 10968
rect 7883 10996 7895 10999
rect 8202 10996 8208 11008
rect 7883 10968 8208 10996
rect 7883 10965 7895 10968
rect 7837 10959 7895 10965
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8389 10999 8447 11005
rect 8389 10965 8401 10999
rect 8435 10996 8447 10999
rect 8478 10996 8484 11008
rect 8435 10968 8484 10996
rect 8435 10965 8447 10968
rect 8389 10959 8447 10965
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 8588 10996 8616 11036
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 12713 11067 12771 11073
rect 12713 11064 12725 11067
rect 12492 11036 12725 11064
rect 12492 11024 12498 11036
rect 12713 11033 12725 11036
rect 12759 11064 12771 11067
rect 12989 11067 13047 11073
rect 12759 11036 12940 11064
rect 12759 11033 12771 11036
rect 12713 11027 12771 11033
rect 9122 10996 9128 11008
rect 8588 10968 9128 10996
rect 9122 10956 9128 10968
rect 9180 10996 9186 11008
rect 9861 10999 9919 11005
rect 9861 10996 9873 10999
rect 9180 10968 9873 10996
rect 9180 10956 9186 10968
rect 9861 10965 9873 10968
rect 9907 10965 9919 10999
rect 9861 10959 9919 10965
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 12805 10999 12863 11005
rect 12805 10996 12817 10999
rect 12676 10968 12817 10996
rect 12676 10956 12682 10968
rect 12805 10965 12817 10968
rect 12851 10965 12863 10999
rect 12912 10996 12940 11036
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 13078 11064 13084 11076
rect 13035 11036 13084 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 13446 11024 13452 11076
rect 13504 11024 13510 11076
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 13556 11036 14749 11064
rect 13556 10996 13584 11036
rect 14737 11033 14749 11036
rect 14783 11033 14795 11067
rect 14737 11027 14795 11033
rect 16022 11024 16028 11076
rect 16080 11064 16086 11076
rect 16408 11064 16436 11104
rect 16574 11064 16580 11076
rect 16080 11036 16436 11064
rect 16500 11036 16580 11064
rect 16080 11024 16086 11036
rect 12912 10968 13584 10996
rect 12805 10959 12863 10965
rect 14458 10956 14464 11008
rect 14516 10996 14522 11008
rect 14645 10999 14703 11005
rect 14645 10996 14657 10999
rect 14516 10968 14657 10996
rect 14516 10956 14522 10968
rect 14645 10965 14657 10968
rect 14691 10996 14703 10999
rect 15010 10996 15016 11008
rect 14691 10968 15016 10996
rect 14691 10965 14703 10968
rect 14645 10959 14703 10965
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 16500 11005 16528 11036
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 16485 10999 16543 11005
rect 16485 10965 16497 10999
rect 16531 10965 16543 10999
rect 17144 10996 17172 11104
rect 19705 11101 19717 11135
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 20248 11135 20306 11141
rect 20248 11101 20260 11135
rect 20294 11132 20306 11135
rect 21082 11132 21088 11144
rect 20294 11104 21088 11132
rect 20294 11101 20306 11104
rect 20248 11095 20306 11101
rect 17310 11024 17316 11076
rect 17368 11024 17374 11076
rect 17954 11024 17960 11076
rect 18012 11024 18018 11076
rect 19720 11064 19748 11095
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 20898 11064 20904 11076
rect 19720 11036 20904 11064
rect 20898 11024 20904 11036
rect 20956 11024 20962 11076
rect 17221 10999 17279 11005
rect 17221 10996 17233 10999
rect 17144 10968 17233 10996
rect 16485 10959 16543 10965
rect 17221 10965 17233 10968
rect 17267 10965 17279 10999
rect 17221 10959 17279 10965
rect 18138 10956 18144 11008
rect 18196 10956 18202 11008
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 19889 10999 19947 11005
rect 19889 10996 19901 10999
rect 19852 10968 19901 10996
rect 19852 10956 19858 10968
rect 19889 10965 19901 10968
rect 19935 10965 19947 10999
rect 19889 10959 19947 10965
rect 1104 10906 21988 10928
rect 1104 10854 4220 10906
rect 4272 10854 4284 10906
rect 4336 10854 4348 10906
rect 4400 10854 4412 10906
rect 4464 10854 4476 10906
rect 4528 10854 9441 10906
rect 9493 10854 9505 10906
rect 9557 10854 9569 10906
rect 9621 10854 9633 10906
rect 9685 10854 9697 10906
rect 9749 10854 14662 10906
rect 14714 10854 14726 10906
rect 14778 10854 14790 10906
rect 14842 10854 14854 10906
rect 14906 10854 14918 10906
rect 14970 10854 19883 10906
rect 19935 10854 19947 10906
rect 19999 10854 20011 10906
rect 20063 10854 20075 10906
rect 20127 10854 20139 10906
rect 20191 10854 21988 10906
rect 1104 10832 21988 10854
rect 3786 10752 3792 10804
rect 3844 10752 3850 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 5258 10792 5264 10804
rect 4212 10764 5264 10792
rect 4212 10752 4218 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5534 10752 5540 10804
rect 5592 10752 5598 10804
rect 11790 10792 11796 10804
rect 11164 10764 11796 10792
rect 3234 10684 3240 10736
rect 3292 10724 3298 10736
rect 3605 10727 3663 10733
rect 3605 10724 3617 10727
rect 3292 10696 3617 10724
rect 3292 10684 3298 10696
rect 3605 10693 3617 10696
rect 3651 10693 3663 10727
rect 3605 10687 3663 10693
rect 4341 10727 4399 10733
rect 4341 10693 4353 10727
rect 4387 10724 4399 10727
rect 4706 10724 4712 10736
rect 4387 10696 4712 10724
rect 4387 10693 4399 10696
rect 4341 10687 4399 10693
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 5353 10727 5411 10733
rect 5353 10693 5365 10727
rect 5399 10724 5411 10727
rect 5442 10724 5448 10736
rect 5399 10696 5448 10724
rect 5399 10693 5411 10696
rect 5353 10687 5411 10693
rect 5442 10684 5448 10696
rect 5500 10684 5506 10736
rect 7469 10727 7527 10733
rect 7469 10693 7481 10727
rect 7515 10724 7527 10727
rect 10137 10727 10195 10733
rect 7515 10696 8156 10724
rect 7515 10693 7527 10696
rect 7469 10687 7527 10693
rect 8128 10668 8156 10696
rect 10137 10693 10149 10727
rect 10183 10724 10195 10727
rect 11164 10724 11192 10764
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12584 10764 12909 10792
rect 12584 10752 12590 10764
rect 12897 10761 12909 10764
rect 12943 10792 12955 10795
rect 13446 10792 13452 10804
rect 12943 10764 13452 10792
rect 12943 10761 12955 10764
rect 12897 10755 12955 10761
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16393 10795 16451 10801
rect 16393 10792 16405 10795
rect 16080 10764 16405 10792
rect 16080 10752 16086 10764
rect 16393 10761 16405 10764
rect 16439 10761 16451 10795
rect 16393 10755 16451 10761
rect 19153 10795 19211 10801
rect 19153 10761 19165 10795
rect 19199 10761 19211 10795
rect 19153 10755 19211 10761
rect 20625 10795 20683 10801
rect 20625 10761 20637 10795
rect 20671 10761 20683 10795
rect 20625 10755 20683 10761
rect 10183 10696 11192 10724
rect 10183 10693 10195 10696
rect 10137 10687 10195 10693
rect 1946 10665 1952 10668
rect 1940 10619 1952 10665
rect 1946 10616 1952 10619
rect 2004 10616 2010 10668
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 5902 10656 5908 10668
rect 4663 10628 5908 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 5902 10616 5908 10628
rect 5960 10656 5966 10668
rect 6822 10656 6828 10668
rect 5960 10628 6828 10656
rect 5960 10616 5966 10628
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7064 10628 7665 10656
rect 7064 10616 7070 10628
rect 7653 10625 7665 10628
rect 7699 10656 7711 10659
rect 7926 10656 7932 10668
rect 7699 10628 7932 10656
rect 7699 10625 7711 10628
rect 7653 10619 7711 10625
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8110 10616 8116 10668
rect 8168 10616 8174 10668
rect 8478 10616 8484 10668
rect 8536 10616 8542 10668
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9214 10616 9220 10668
rect 9272 10656 9278 10668
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 9272 10628 9321 10656
rect 9272 10616 9278 10628
rect 9309 10625 9321 10628
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 9858 10616 9864 10668
rect 9916 10616 9922 10668
rect 10594 10616 10600 10668
rect 10652 10616 10658 10668
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 11164 10665 11192 10696
rect 14366 10684 14372 10736
rect 14424 10733 14430 10736
rect 14424 10724 14436 10733
rect 16114 10724 16120 10736
rect 14424 10696 14469 10724
rect 14568 10696 16120 10724
rect 14424 10687 14436 10696
rect 14424 10684 14430 10687
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 1670 10548 1676 10600
rect 1728 10548 1734 10600
rect 3881 10591 3939 10597
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 4154 10588 4160 10600
rect 3927 10560 4160 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10588 4583 10591
rect 4798 10588 4804 10600
rect 4571 10560 4804 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5442 10588 5448 10600
rect 4908 10560 5448 10588
rect 3326 10480 3332 10532
rect 3384 10480 3390 10532
rect 4908 10520 4936 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 4632 10492 4936 10520
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 4632 10461 4660 10492
rect 5074 10480 5080 10532
rect 5132 10480 5138 10532
rect 5258 10480 5264 10532
rect 5316 10520 5322 10532
rect 5644 10520 5672 10551
rect 10410 10548 10416 10600
rect 10468 10548 10474 10600
rect 5316 10492 5672 10520
rect 5316 10480 5322 10492
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 10686 10520 10692 10532
rect 10376 10492 10692 10520
rect 10376 10480 10382 10492
rect 10686 10480 10692 10492
rect 10744 10520 10750 10532
rect 10980 10520 11008 10619
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11773 10659 11831 10665
rect 11773 10656 11785 10659
rect 11296 10628 11785 10656
rect 11296 10616 11302 10628
rect 11773 10625 11785 10628
rect 11819 10625 11831 10659
rect 11773 10619 11831 10625
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 14568 10656 14596 10696
rect 16114 10684 16120 10696
rect 16172 10684 16178 10736
rect 17126 10684 17132 10736
rect 17184 10724 17190 10736
rect 19168 10724 19196 10755
rect 19490 10727 19548 10733
rect 19490 10724 19502 10727
rect 17184 10696 18644 10724
rect 19168 10696 19502 10724
rect 17184 10684 17190 10696
rect 12124 10628 14596 10656
rect 14645 10659 14703 10665
rect 12124 10616 12130 10628
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14691 10628 15025 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 15013 10625 15025 10628
rect 15059 10656 15071 10659
rect 15102 10656 15108 10668
rect 15059 10628 15108 10656
rect 15059 10625 15071 10628
rect 15013 10619 15071 10625
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 15286 10665 15292 10668
rect 15280 10619 15292 10665
rect 15286 10616 15292 10619
rect 15344 10616 15350 10668
rect 18616 10665 18644 10696
rect 19490 10693 19502 10696
rect 19536 10693 19548 10727
rect 20640 10724 20668 10755
rect 20993 10727 21051 10733
rect 20993 10724 21005 10727
rect 20640 10696 21005 10724
rect 19490 10687 19548 10693
rect 20993 10693 21005 10696
rect 21039 10724 21051 10727
rect 21358 10724 21364 10736
rect 21039 10696 21364 10724
rect 21039 10693 21051 10696
rect 20993 10687 21051 10693
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 18345 10659 18403 10665
rect 18345 10625 18357 10659
rect 18391 10656 18403 10659
rect 18601 10659 18659 10665
rect 18391 10628 18552 10656
rect 18391 10625 18403 10628
rect 18345 10619 18403 10625
rect 11514 10548 11520 10600
rect 11572 10548 11578 10600
rect 18524 10588 18552 10628
rect 18601 10625 18613 10659
rect 18647 10656 18659 10659
rect 18647 10628 18828 10656
rect 18647 10625 18659 10628
rect 18601 10619 18659 10625
rect 18800 10588 18828 10628
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10656 19027 10659
rect 19015 10628 21496 10656
rect 19015 10625 19027 10628
rect 18969 10619 19027 10625
rect 19058 10588 19064 10600
rect 18524 10560 18644 10588
rect 18800 10560 19064 10588
rect 10744 10492 11008 10520
rect 10744 10480 10750 10492
rect 13262 10480 13268 10532
rect 13320 10480 13326 10532
rect 18616 10520 18644 10560
rect 19058 10548 19064 10560
rect 19116 10588 19122 10600
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 19116 10560 19257 10588
rect 19116 10548 19122 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 20806 10548 20812 10600
rect 20864 10588 20870 10600
rect 20901 10591 20959 10597
rect 20901 10588 20913 10591
rect 20864 10560 20913 10588
rect 20864 10548 20870 10560
rect 20901 10557 20913 10560
rect 20947 10557 20959 10591
rect 20901 10551 20959 10557
rect 20990 10548 20996 10600
rect 21048 10548 21054 10600
rect 21468 10529 21496 10628
rect 18693 10523 18751 10529
rect 18693 10520 18705 10523
rect 18616 10492 18705 10520
rect 18693 10489 18705 10492
rect 18739 10489 18751 10523
rect 18693 10483 18751 10489
rect 21453 10523 21511 10529
rect 21453 10489 21465 10523
rect 21499 10489 21511 10523
rect 21453 10483 21511 10489
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2924 10424 3065 10452
rect 2924 10412 2930 10424
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 3053 10415 3111 10421
rect 4617 10455 4675 10461
rect 4617 10421 4629 10455
rect 4663 10421 4675 10455
rect 4617 10415 4675 10421
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5810 10452 5816 10464
rect 4847 10424 5816 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 7374 10452 7380 10464
rect 6052 10424 7380 10452
rect 6052 10412 6058 10424
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7742 10412 7748 10464
rect 7800 10412 7806 10464
rect 11057 10455 11115 10461
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 14366 10452 14372 10464
rect 11103 10424 14372 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 17221 10455 17279 10461
rect 17221 10421 17233 10455
rect 17267 10452 17279 10455
rect 17954 10452 17960 10464
rect 17267 10424 17960 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 1104 10362 21988 10384
rect 1104 10310 3560 10362
rect 3612 10310 3624 10362
rect 3676 10310 3688 10362
rect 3740 10310 3752 10362
rect 3804 10310 3816 10362
rect 3868 10310 8781 10362
rect 8833 10310 8845 10362
rect 8897 10310 8909 10362
rect 8961 10310 8973 10362
rect 9025 10310 9037 10362
rect 9089 10310 14002 10362
rect 14054 10310 14066 10362
rect 14118 10310 14130 10362
rect 14182 10310 14194 10362
rect 14246 10310 14258 10362
rect 14310 10310 19223 10362
rect 19275 10310 19287 10362
rect 19339 10310 19351 10362
rect 19403 10310 19415 10362
rect 19467 10310 19479 10362
rect 19531 10310 21988 10362
rect 1104 10288 21988 10310
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 2041 10251 2099 10257
rect 2041 10248 2053 10251
rect 2004 10220 2053 10248
rect 2004 10208 2010 10220
rect 2041 10217 2053 10220
rect 2087 10217 2099 10251
rect 2041 10211 2099 10217
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 6086 10248 6092 10260
rect 3200 10220 6092 10248
rect 3200 10208 3206 10220
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 6288 10220 6561 10248
rect 2409 10183 2467 10189
rect 2409 10149 2421 10183
rect 2455 10149 2467 10183
rect 2409 10143 2467 10149
rect 3513 10183 3571 10189
rect 3513 10149 3525 10183
rect 3559 10180 3571 10183
rect 4154 10180 4160 10192
rect 3559 10152 4160 10180
rect 3559 10149 3571 10152
rect 3513 10143 3571 10149
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2424 10044 2452 10143
rect 4154 10140 4160 10152
rect 4212 10140 4218 10192
rect 5442 10140 5448 10192
rect 5500 10180 5506 10192
rect 6288 10180 6316 10220
rect 6549 10217 6561 10220
rect 6595 10248 6607 10251
rect 7742 10248 7748 10260
rect 6595 10220 7748 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8113 10251 8171 10257
rect 8113 10217 8125 10251
rect 8159 10248 8171 10251
rect 8478 10248 8484 10260
rect 8159 10220 8484 10248
rect 8159 10217 8171 10220
rect 8113 10211 8171 10217
rect 5500 10152 6316 10180
rect 6365 10183 6423 10189
rect 5500 10140 5506 10152
rect 6365 10149 6377 10183
rect 6411 10149 6423 10183
rect 6365 10143 6423 10149
rect 5276 10084 5948 10112
rect 2271 10016 2452 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 3050 10004 3056 10056
rect 3108 10044 3114 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 3108 10016 3249 10044
rect 3108 10004 3114 10016
rect 3237 10013 3249 10016
rect 3283 10044 3295 10047
rect 3326 10044 3332 10056
rect 3283 10016 3332 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4154 10044 4160 10056
rect 4019 10016 4160 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 4295 10016 4660 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4632 9988 4660 10016
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5276 10044 5304 10084
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5132 10016 5304 10044
rect 5644 10016 5825 10044
rect 5132 10004 5138 10016
rect 1302 9936 1308 9988
rect 1360 9976 1366 9988
rect 2685 9979 2743 9985
rect 2685 9976 2697 9979
rect 1360 9948 2697 9976
rect 1360 9936 1366 9948
rect 2685 9945 2697 9948
rect 2731 9945 2743 9979
rect 2685 9939 2743 9945
rect 2958 9936 2964 9988
rect 3016 9936 3022 9988
rect 4494 9979 4552 9985
rect 4494 9976 4506 9979
rect 4172 9948 4506 9976
rect 2866 9868 2872 9920
rect 2924 9868 2930 9920
rect 4172 9917 4200 9948
rect 4494 9945 4506 9948
rect 4540 9945 4552 9979
rect 4494 9939 4552 9945
rect 4614 9936 4620 9988
rect 4672 9936 4678 9988
rect 5644 9920 5672 10016
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 5920 9976 5948 10084
rect 5994 10004 6000 10056
rect 6052 10004 6058 10056
rect 6086 10004 6092 10056
rect 6144 10004 6150 10056
rect 6233 10047 6291 10053
rect 6233 10013 6245 10047
rect 6279 10044 6291 10047
rect 6380 10044 6408 10143
rect 7374 10140 7380 10192
rect 7432 10180 7438 10192
rect 8021 10183 8079 10189
rect 8021 10180 8033 10183
rect 7432 10152 8033 10180
rect 7432 10140 7438 10152
rect 8021 10149 8033 10152
rect 8067 10149 8079 10183
rect 8021 10143 8079 10149
rect 6638 10072 6644 10124
rect 6696 10072 6702 10124
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6279 10013 6316 10044
rect 6380 10016 6561 10044
rect 6233 10007 6316 10013
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 6288 9976 6316 10007
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 7926 10004 7932 10056
rect 7984 10004 7990 10056
rect 8128 9976 8156 10211
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11238 10248 11244 10260
rect 10919 10220 11244 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 12066 10248 12072 10260
rect 11440 10220 12072 10248
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 11440 10180 11468 10220
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12986 10208 12992 10260
rect 13044 10208 13050 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15381 10251 15439 10257
rect 15381 10248 15393 10251
rect 15344 10220 15393 10248
rect 15344 10208 15350 10220
rect 15381 10217 15393 10220
rect 15427 10217 15439 10251
rect 15381 10211 15439 10217
rect 15746 10208 15752 10260
rect 15804 10208 15810 10260
rect 16945 10251 17003 10257
rect 16945 10217 16957 10251
rect 16991 10248 17003 10251
rect 17310 10248 17316 10260
rect 16991 10220 17316 10248
rect 16991 10217 17003 10220
rect 16945 10211 17003 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 18509 10251 18567 10257
rect 18509 10248 18521 10251
rect 18196 10220 18521 10248
rect 18196 10208 18202 10220
rect 18509 10217 18521 10220
rect 18555 10217 18567 10251
rect 18509 10211 18567 10217
rect 10244 10152 11468 10180
rect 11517 10183 11575 10189
rect 10244 10121 10272 10152
rect 11517 10149 11529 10183
rect 11563 10149 11575 10183
rect 11517 10143 11575 10149
rect 10229 10115 10287 10121
rect 8956 10084 10088 10112
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8956 10053 8984 10084
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8352 10016 8953 10044
rect 8352 10004 8358 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 10060 10053 10088 10084
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 9272 10016 9321 10044
rect 9272 10004 9278 10016
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 11532 10044 11560 10143
rect 11977 10115 12035 10121
rect 11977 10081 11989 10115
rect 12023 10112 12035 10115
rect 12526 10112 12532 10124
rect 12023 10084 12532 10112
rect 12023 10081 12035 10084
rect 11977 10075 12035 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 12894 10072 12900 10124
rect 12952 10072 12958 10124
rect 17126 10072 17132 10124
rect 17184 10072 17190 10124
rect 10735 10016 11560 10044
rect 12069 10047 12127 10053
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 12069 10013 12081 10047
rect 12115 10044 12127 10047
rect 12342 10044 12348 10056
rect 12115 10016 12348 10044
rect 12115 10013 12127 10016
rect 12069 10007 12127 10013
rect 5920 9948 8156 9976
rect 9968 9976 9996 10007
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 12912 10044 12940 10072
rect 12728 10016 12940 10044
rect 10318 9976 10324 9988
rect 9968 9948 10324 9976
rect 10318 9936 10324 9948
rect 10376 9936 10382 9988
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 12728 9976 12756 10016
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13280 10016 14289 10044
rect 10836 9948 12756 9976
rect 10836 9936 10842 9948
rect 12802 9936 12808 9988
rect 12860 9936 12866 9988
rect 4157 9911 4215 9917
rect 4157 9877 4169 9911
rect 4203 9877 4215 9911
rect 4157 9871 4215 9877
rect 4246 9868 4252 9920
rect 4304 9908 4310 9920
rect 4798 9908 4804 9920
rect 4304 9880 4804 9908
rect 4304 9868 4310 9880
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 5626 9868 5632 9920
rect 5684 9868 5690 9920
rect 7006 9868 7012 9920
rect 7064 9868 7070 9920
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 7432 9880 7665 9908
rect 7432 9868 7438 9880
rect 7653 9877 7665 9880
rect 7699 9908 7711 9911
rect 7926 9908 7932 9920
rect 7699 9880 7932 9908
rect 7699 9877 7711 9880
rect 7653 9871 7711 9877
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 11977 9911 12035 9917
rect 11977 9877 11989 9911
rect 12023 9908 12035 9911
rect 12434 9908 12440 9920
rect 12023 9880 12440 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 12434 9868 12440 9880
rect 12492 9908 12498 9920
rect 13170 9908 13176 9920
rect 12492 9880 13176 9908
rect 12492 9868 12498 9880
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 13280 9917 13308 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14366 10004 14372 10056
rect 14424 10044 14430 10056
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 14424 10016 14473 10044
rect 14424 10004 14430 10016
rect 14461 10013 14473 10016
rect 14507 10044 14519 10047
rect 15378 10044 15384 10056
rect 14507 10016 15384 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 15562 10004 15568 10056
rect 15620 10004 15626 10056
rect 19058 10004 19064 10056
rect 19116 10044 19122 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19116 10016 19809 10044
rect 19116 10004 19122 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 20053 10047 20111 10053
rect 20053 10044 20065 10047
rect 19944 10016 20065 10044
rect 19944 10004 19950 10016
rect 20053 10013 20065 10016
rect 20099 10013 20111 10047
rect 20053 10007 20111 10013
rect 20622 10004 20628 10056
rect 20680 10044 20686 10056
rect 21545 10047 21603 10053
rect 21545 10044 21557 10047
rect 20680 10016 21557 10044
rect 20680 10004 20686 10016
rect 21545 10013 21557 10016
rect 21591 10013 21603 10047
rect 21545 10007 21603 10013
rect 14645 9979 14703 9985
rect 14645 9945 14657 9979
rect 14691 9976 14703 9979
rect 16025 9979 16083 9985
rect 16025 9976 16037 9979
rect 14691 9948 16037 9976
rect 14691 9945 14703 9948
rect 14645 9939 14703 9945
rect 16025 9945 16037 9948
rect 16071 9976 16083 9979
rect 16206 9976 16212 9988
rect 16071 9948 16212 9976
rect 16071 9945 16083 9948
rect 16025 9939 16083 9945
rect 16206 9936 16212 9948
rect 16264 9976 16270 9988
rect 17402 9985 17408 9988
rect 16669 9979 16727 9985
rect 16669 9976 16681 9979
rect 16264 9948 16681 9976
rect 16264 9936 16270 9948
rect 16669 9945 16681 9948
rect 16715 9945 16727 9979
rect 16669 9939 16727 9945
rect 17396 9939 17408 9985
rect 17402 9936 17408 9939
rect 17460 9936 17466 9988
rect 20254 9936 20260 9988
rect 20312 9976 20318 9988
rect 20312 9948 21404 9976
rect 20312 9936 20318 9948
rect 13265 9911 13323 9917
rect 13265 9877 13277 9911
rect 13311 9877 13323 9911
rect 13265 9871 13323 9877
rect 21177 9911 21235 9917
rect 21177 9877 21189 9911
rect 21223 9908 21235 9911
rect 21266 9908 21272 9920
rect 21223 9880 21272 9908
rect 21223 9877 21235 9880
rect 21177 9871 21235 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 21376 9917 21404 9948
rect 21361 9911 21419 9917
rect 21361 9877 21373 9911
rect 21407 9877 21419 9911
rect 21361 9871 21419 9877
rect 1104 9818 21988 9840
rect 1104 9766 4220 9818
rect 4272 9766 4284 9818
rect 4336 9766 4348 9818
rect 4400 9766 4412 9818
rect 4464 9766 4476 9818
rect 4528 9766 9441 9818
rect 9493 9766 9505 9818
rect 9557 9766 9569 9818
rect 9621 9766 9633 9818
rect 9685 9766 9697 9818
rect 9749 9766 14662 9818
rect 14714 9766 14726 9818
rect 14778 9766 14790 9818
rect 14842 9766 14854 9818
rect 14906 9766 14918 9818
rect 14970 9766 19883 9818
rect 19935 9766 19947 9818
rect 19999 9766 20011 9818
rect 20063 9766 20075 9818
rect 20127 9766 20139 9818
rect 20191 9766 21988 9818
rect 1104 9744 21988 9766
rect 5997 9707 6055 9713
rect 5997 9673 6009 9707
rect 6043 9673 6055 9707
rect 5997 9667 6055 9673
rect 8297 9707 8355 9713
rect 8297 9673 8309 9707
rect 8343 9673 8355 9707
rect 8297 9667 8355 9673
rect 8941 9707 8999 9713
rect 8941 9673 8953 9707
rect 8987 9704 8999 9707
rect 9674 9704 9680 9716
rect 8987 9676 9680 9704
rect 8987 9673 8999 9676
rect 8941 9667 8999 9673
rect 1302 9596 1308 9648
rect 1360 9636 1366 9648
rect 2593 9639 2651 9645
rect 2593 9636 2605 9639
rect 1360 9608 2605 9636
rect 1360 9596 1366 9608
rect 2593 9605 2605 9608
rect 2639 9605 2651 9639
rect 2593 9599 2651 9605
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9605 2835 9639
rect 2777 9599 2835 9605
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9568 2191 9571
rect 2792 9568 2820 9599
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 2924 9608 3832 9636
rect 2924 9596 2930 9608
rect 3050 9568 3056 9580
rect 2179 9540 2360 9568
rect 2792 9540 3056 9568
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 2332 9441 2360 9540
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 3804 9577 3832 9608
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 5077 9639 5135 9645
rect 5077 9636 5089 9639
rect 3936 9608 5089 9636
rect 3936 9596 3942 9608
rect 5077 9605 5089 9608
rect 5123 9605 5135 9639
rect 5077 9599 5135 9605
rect 5261 9639 5319 9645
rect 5261 9605 5273 9639
rect 5307 9636 5319 9639
rect 5626 9636 5632 9648
rect 5307 9608 5632 9636
rect 5307 9605 5319 9608
rect 5261 9599 5319 9605
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 5810 9596 5816 9648
rect 5868 9596 5874 9648
rect 6012 9636 6040 9667
rect 6546 9636 6552 9648
rect 6012 9608 6552 9636
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 8312 9636 8340 9667
rect 9674 9664 9680 9676
rect 9732 9704 9738 9716
rect 10410 9704 10416 9716
rect 9732 9676 10416 9704
rect 9732 9664 9738 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 17402 9664 17408 9716
rect 17460 9664 17466 9716
rect 17957 9707 18015 9713
rect 17957 9673 17969 9707
rect 18003 9704 18015 9707
rect 18138 9704 18144 9716
rect 18003 9676 18144 9704
rect 18003 9673 18015 9676
rect 17957 9667 18015 9673
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 21358 9664 21364 9716
rect 21416 9664 21422 9716
rect 8478 9636 8484 9648
rect 6656 9608 7696 9636
rect 8312 9608 8484 9636
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 3970 9528 3976 9580
rect 4028 9528 4034 9580
rect 4062 9528 4068 9580
rect 4120 9528 4126 9580
rect 4209 9571 4267 9577
rect 4209 9537 4221 9571
rect 4255 9568 4267 9571
rect 4982 9568 4988 9580
rect 4255 9540 4988 9568
rect 4255 9537 4267 9540
rect 4209 9531 4267 9537
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5951 9571 6009 9577
rect 5951 9537 5963 9571
rect 5997 9568 6009 9571
rect 6086 9568 6092 9580
rect 5997 9540 6092 9568
rect 5997 9537 6009 9540
rect 5951 9531 6009 9537
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6656 9577 6684 9608
rect 7668 9580 7696 9608
rect 8478 9596 8484 9608
rect 8536 9636 8542 9648
rect 10045 9639 10103 9645
rect 8536 9608 9444 9636
rect 8536 9596 8542 9608
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 6457 9571 6515 9577
rect 6457 9568 6469 9571
rect 6227 9540 6469 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6457 9537 6469 9540
rect 6503 9537 6515 9571
rect 6457 9531 6515 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 6788 9540 6929 9568
rect 6788 9528 6794 9540
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 7184 9571 7242 9577
rect 7184 9537 7196 9571
rect 7230 9568 7242 9571
rect 7558 9568 7564 9580
rect 7230 9540 7564 9568
rect 7230 9537 7242 9540
rect 7184 9531 7242 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 7708 9540 8769 9568
rect 7708 9528 7714 9540
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9122 9568 9128 9580
rect 9079 9540 9128 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 2869 9503 2927 9509
rect 2869 9469 2881 9503
rect 2915 9500 2927 9503
rect 2958 9500 2964 9512
rect 2915 9472 2964 9500
rect 2915 9469 2927 9472
rect 2869 9463 2927 9469
rect 2958 9460 2964 9472
rect 3016 9500 3022 9512
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3016 9472 3617 9500
rect 3016 9460 3022 9472
rect 3605 9469 3617 9472
rect 3651 9500 3663 9503
rect 5353 9503 5411 9509
rect 5353 9500 5365 9503
rect 3651 9472 5365 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 5353 9469 5365 9472
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6871 9472 6960 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 2317 9435 2375 9441
rect 2317 9401 2329 9435
rect 2363 9401 2375 9435
rect 2317 9395 2375 9401
rect 4341 9435 4399 9441
rect 4341 9401 4353 9435
rect 4387 9432 4399 9435
rect 4706 9432 4712 9444
rect 4387 9404 4712 9432
rect 4387 9401 4399 9404
rect 4341 9395 4399 9401
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 4798 9392 4804 9444
rect 4856 9392 4862 9444
rect 5626 9392 5632 9444
rect 5684 9392 5690 9444
rect 1946 9324 1952 9376
rect 2004 9324 2010 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 5994 9364 6000 9376
rect 4028 9336 6000 9364
rect 4028 9324 4034 9336
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 6932 9364 6960 9472
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 9048 9500 9076 9531
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 9416 9577 9444 9608
rect 10045 9605 10057 9639
rect 10091 9636 10103 9639
rect 10594 9636 10600 9648
rect 10091 9608 10600 9636
rect 10091 9605 10103 9608
rect 10045 9599 10103 9605
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 12618 9596 12624 9648
rect 12676 9636 12682 9648
rect 13173 9639 13231 9645
rect 13173 9636 13185 9639
rect 12676 9608 13185 9636
rect 12676 9596 12682 9608
rect 13173 9605 13185 9608
rect 13219 9605 13231 9639
rect 13173 9599 13231 9605
rect 13265 9639 13323 9645
rect 13265 9605 13277 9639
rect 13311 9636 13323 9639
rect 13311 9608 14320 9636
rect 13311 9605 13323 9608
rect 13265 9599 13323 9605
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 10778 9568 10784 9580
rect 9907 9540 10784 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 13541 9571 13599 9577
rect 12575 9540 12756 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 7984 9472 9076 9500
rect 9585 9503 9643 9509
rect 7984 9460 7990 9472
rect 9585 9469 9597 9503
rect 9631 9469 9643 9503
rect 9585 9463 9643 9469
rect 8018 9392 8024 9444
rect 8076 9432 8082 9444
rect 8573 9435 8631 9441
rect 8573 9432 8585 9435
rect 8076 9404 8585 9432
rect 8076 9392 8082 9404
rect 8573 9401 8585 9404
rect 8619 9401 8631 9435
rect 8573 9395 8631 9401
rect 8662 9392 8668 9444
rect 8720 9432 8726 9444
rect 9600 9432 9628 9463
rect 12728 9441 12756 9540
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 14292 9568 14320 9608
rect 14366 9596 14372 9648
rect 14424 9596 14430 9648
rect 14461 9639 14519 9645
rect 14461 9605 14473 9639
rect 14507 9636 14519 9639
rect 15746 9636 15752 9648
rect 14507 9608 15752 9636
rect 14507 9605 14519 9608
rect 14461 9599 14519 9605
rect 14476 9568 14504 9599
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 16301 9639 16359 9645
rect 16301 9605 16313 9639
rect 16347 9636 16359 9639
rect 17034 9636 17040 9648
rect 16347 9608 17040 9636
rect 16347 9605 16359 9608
rect 16301 9599 16359 9605
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 19058 9596 19064 9648
rect 19116 9636 19122 9648
rect 19705 9639 19763 9645
rect 19705 9636 19717 9639
rect 19116 9608 19717 9636
rect 19116 9596 19122 9608
rect 19705 9605 19717 9608
rect 19751 9605 19763 9639
rect 19705 9599 19763 9605
rect 20165 9639 20223 9645
rect 20165 9605 20177 9639
rect 20211 9636 20223 9639
rect 20438 9636 20444 9648
rect 20211 9608 20444 9636
rect 20211 9605 20223 9608
rect 20165 9599 20223 9605
rect 20438 9596 20444 9608
rect 20496 9596 20502 9648
rect 20530 9596 20536 9648
rect 20588 9636 20594 9648
rect 21453 9639 21511 9645
rect 21453 9636 21465 9639
rect 20588 9608 21465 9636
rect 20588 9596 20594 9608
rect 21453 9605 21465 9608
rect 21499 9605 21511 9639
rect 21453 9599 21511 9605
rect 13587 9540 13952 9568
rect 14292 9540 14504 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9500 13231 9503
rect 13814 9500 13820 9512
rect 13219 9472 13820 9500
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 13924 9441 13952 9540
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 15436 9540 15608 9568
rect 15436 9528 15442 9540
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 15470 9500 15476 9512
rect 14415 9472 15476 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 15580 9500 15608 9540
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 15712 9540 16129 9568
rect 15712 9528 15718 9540
rect 16117 9537 16129 9540
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 17586 9528 17592 9580
rect 17644 9528 17650 9580
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 18969 9571 19027 9577
rect 18969 9568 18981 9571
rect 18196 9540 18981 9568
rect 18196 9528 18202 9540
rect 18969 9537 18981 9540
rect 19015 9537 19027 9571
rect 18969 9531 19027 9537
rect 20349 9571 20407 9577
rect 20349 9537 20361 9571
rect 20395 9568 20407 9571
rect 21174 9568 21180 9580
rect 20395 9540 21180 9568
rect 20395 9537 20407 9540
rect 20349 9531 20407 9537
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 15838 9500 15844 9512
rect 15580 9472 15844 9500
rect 15838 9460 15844 9472
rect 15896 9500 15902 9512
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 15896 9472 16405 9500
rect 15896 9460 15902 9472
rect 16393 9469 16405 9472
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 17310 9460 17316 9512
rect 17368 9500 17374 9512
rect 17865 9503 17923 9509
rect 17865 9500 17877 9503
rect 17368 9472 17877 9500
rect 17368 9460 17374 9472
rect 17865 9469 17877 9472
rect 17911 9469 17923 9503
rect 17865 9463 17923 9469
rect 8720 9404 9628 9432
rect 12713 9435 12771 9441
rect 8720 9392 8726 9404
rect 12713 9401 12725 9435
rect 12759 9401 12771 9435
rect 12713 9395 12771 9401
rect 13909 9435 13967 9441
rect 13909 9401 13921 9435
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 8294 9364 8300 9376
rect 6932 9336 8300 9364
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 9217 9367 9275 9373
rect 9217 9364 9229 9367
rect 8444 9336 9229 9364
rect 8444 9324 8450 9336
rect 9217 9333 9229 9336
rect 9263 9333 9275 9367
rect 9217 9327 9275 9333
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 10042 9364 10048 9376
rect 9815 9336 10048 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 12158 9324 12164 9376
rect 12216 9364 12222 9376
rect 12345 9367 12403 9373
rect 12345 9364 12357 9367
rect 12216 9336 12357 9364
rect 12216 9324 12222 9336
rect 12345 9333 12357 9336
rect 12391 9333 12403 9367
rect 12345 9327 12403 9333
rect 13722 9324 13728 9376
rect 13780 9324 13786 9376
rect 15841 9367 15899 9373
rect 15841 9333 15853 9367
rect 15887 9364 15899 9367
rect 16298 9364 16304 9376
rect 15887 9336 16304 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 17880 9364 17908 9463
rect 18046 9460 18052 9512
rect 18104 9460 18110 9512
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 18417 9435 18475 9441
rect 18417 9401 18429 9435
rect 18463 9432 18475 9435
rect 18874 9432 18880 9444
rect 18463 9404 18880 9432
rect 18463 9401 18475 9404
rect 18417 9395 18475 9401
rect 18874 9392 18880 9404
rect 18932 9392 18938 9444
rect 19886 9392 19892 9444
rect 19944 9432 19950 9444
rect 20088 9432 20116 9463
rect 21358 9460 21364 9512
rect 21416 9460 21422 9512
rect 20346 9432 20352 9444
rect 19944 9404 20352 9432
rect 19944 9392 19950 9404
rect 20346 9392 20352 9404
rect 20404 9392 20410 9444
rect 20622 9392 20628 9444
rect 20680 9392 20686 9444
rect 20898 9392 20904 9444
rect 20956 9392 20962 9444
rect 20530 9364 20536 9376
rect 17880 9336 20536 9364
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 1104 9274 21988 9296
rect 1104 9222 3560 9274
rect 3612 9222 3624 9274
rect 3676 9222 3688 9274
rect 3740 9222 3752 9274
rect 3804 9222 3816 9274
rect 3868 9222 8781 9274
rect 8833 9222 8845 9274
rect 8897 9222 8909 9274
rect 8961 9222 8973 9274
rect 9025 9222 9037 9274
rect 9089 9222 14002 9274
rect 14054 9222 14066 9274
rect 14118 9222 14130 9274
rect 14182 9222 14194 9274
rect 14246 9222 14258 9274
rect 14310 9222 19223 9274
rect 19275 9222 19287 9274
rect 19339 9222 19351 9274
rect 19403 9222 19415 9274
rect 19467 9222 19479 9274
rect 19531 9222 21988 9274
rect 1104 9200 21988 9222
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 7650 9160 7656 9172
rect 7423 9132 7656 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 17034 9120 17040 9172
rect 17092 9120 17098 9172
rect 18230 9120 18236 9172
rect 18288 9160 18294 9172
rect 18601 9163 18659 9169
rect 18601 9160 18613 9163
rect 18288 9132 18613 9160
rect 18288 9120 18294 9132
rect 18601 9129 18613 9132
rect 18647 9160 18659 9163
rect 20806 9160 20812 9172
rect 18647 9132 20812 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 20806 9120 20812 9132
rect 20864 9120 20870 9172
rect 4890 9052 4896 9104
rect 4948 9092 4954 9104
rect 4948 9064 5212 9092
rect 4948 9052 4954 9064
rect 1670 8916 1676 8968
rect 1728 8916 1734 8968
rect 1946 8965 1952 8968
rect 1940 8956 1952 8965
rect 1907 8928 1952 8956
rect 1940 8919 1952 8928
rect 1946 8916 1952 8919
rect 2004 8916 2010 8968
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 4706 8956 4712 8968
rect 3467 8928 4712 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 4890 8916 4896 8968
rect 4948 8916 4954 8968
rect 5184 8956 5212 9064
rect 7558 9052 7564 9104
rect 7616 9052 7622 9104
rect 7834 9052 7840 9104
rect 7892 9092 7898 9104
rect 8297 9095 8355 9101
rect 8297 9092 8309 9095
rect 7892 9064 8309 9092
rect 7892 9052 7898 9064
rect 8297 9061 8309 9064
rect 8343 9061 8355 9095
rect 8297 9055 8355 9061
rect 10965 9095 11023 9101
rect 10965 9061 10977 9095
rect 11011 9092 11023 9095
rect 11698 9092 11704 9104
rect 11011 9064 11704 9092
rect 11011 9061 11023 9064
rect 10965 9055 11023 9061
rect 11698 9052 11704 9064
rect 11756 9052 11762 9104
rect 13265 9095 13323 9101
rect 13265 9061 13277 9095
rect 13311 9092 13323 9095
rect 13906 9092 13912 9104
rect 13311 9064 13912 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 7340 8996 8708 9024
rect 7340 8984 7346 8996
rect 5313 8959 5371 8965
rect 5313 8956 5325 8959
rect 5184 8928 5325 8956
rect 5313 8925 5325 8928
rect 5359 8956 5371 8959
rect 5534 8956 5540 8968
rect 5359 8928 5540 8956
rect 5359 8925 5371 8928
rect 5313 8919 5371 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6730 8956 6736 8968
rect 6043 8928 6736 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7064 8928 7757 8956
rect 7064 8916 7070 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7883 8959 7941 8965
rect 7883 8925 7895 8959
rect 7929 8956 7941 8959
rect 8018 8956 8024 8968
rect 7929 8928 8024 8956
rect 7929 8925 7941 8928
rect 7883 8919 7941 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 8478 8916 8484 8968
rect 8536 8916 8542 8968
rect 3789 8891 3847 8897
rect 3789 8857 3801 8891
rect 3835 8888 3847 8891
rect 3878 8888 3884 8900
rect 3835 8860 3884 8888
rect 3835 8857 3847 8860
rect 3789 8851 3847 8857
rect 3878 8848 3884 8860
rect 3936 8848 3942 8900
rect 4614 8848 4620 8900
rect 4672 8848 4678 8900
rect 4798 8848 4804 8900
rect 4856 8888 4862 8900
rect 5074 8888 5080 8900
rect 4856 8860 5080 8888
rect 4856 8848 4862 8860
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 5166 8848 5172 8900
rect 5224 8848 5230 8900
rect 5626 8848 5632 8900
rect 5684 8888 5690 8900
rect 6242 8891 6300 8897
rect 6242 8888 6254 8891
rect 5684 8860 6254 8888
rect 5684 8848 5690 8860
rect 6242 8857 6254 8860
rect 6288 8857 6300 8891
rect 6242 8851 6300 8857
rect 8113 8891 8171 8897
rect 8113 8857 8125 8891
rect 8159 8888 8171 8891
rect 8386 8888 8392 8900
rect 8159 8860 8392 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 8386 8848 8392 8860
rect 8444 8848 8450 8900
rect 8680 8897 8708 8996
rect 10502 8984 10508 9036
rect 10560 8984 10566 9036
rect 11514 8984 11520 9036
rect 11572 9024 11578 9036
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 11572 8996 11897 9024
rect 11572 8984 11578 8996
rect 11885 8993 11897 8996
rect 11931 8993 11943 9027
rect 14090 9024 14096 9036
rect 11885 8987 11943 8993
rect 13556 8996 14096 9024
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9122 8956 9128 8968
rect 8803 8928 9128 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 11606 8956 11612 8968
rect 10827 8928 11612 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 11900 8956 11928 8987
rect 13556 8956 13584 8996
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 17126 8984 17132 9036
rect 17184 9024 17190 9036
rect 17221 9027 17279 9033
rect 17221 9024 17233 9027
rect 17184 8996 17233 9024
rect 17184 8984 17190 8996
rect 17221 8993 17233 8996
rect 17267 8993 17279 9027
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 17221 8987 17279 8993
rect 18340 8996 20177 9024
rect 11900 8928 13584 8956
rect 13633 8959 13691 8965
rect 12360 8900 12388 8928
rect 13633 8925 13645 8959
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 8665 8891 8723 8897
rect 8665 8857 8677 8891
rect 8711 8888 8723 8891
rect 9674 8888 9680 8900
rect 8711 8860 9680 8888
rect 8711 8857 8723 8860
rect 8665 8851 8723 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 10238 8891 10296 8897
rect 10238 8888 10250 8891
rect 10192 8860 10250 8888
rect 10192 8848 10198 8860
rect 10238 8857 10250 8860
rect 10284 8857 10296 8891
rect 10238 8851 10296 8857
rect 11238 8848 11244 8900
rect 11296 8848 11302 8900
rect 12158 8897 12164 8900
rect 11517 8891 11575 8897
rect 11517 8857 11529 8891
rect 11563 8857 11575 8891
rect 12152 8888 12164 8897
rect 12119 8860 12164 8888
rect 11517 8851 11575 8857
rect 12152 8851 12164 8860
rect 3050 8780 3056 8832
rect 3108 8780 3114 8832
rect 3605 8823 3663 8829
rect 3605 8789 3617 8823
rect 3651 8820 3663 8823
rect 4062 8820 4068 8832
rect 3651 8792 4068 8820
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 5462 8823 5520 8829
rect 5462 8789 5474 8823
rect 5508 8820 5520 8823
rect 5810 8820 5816 8832
rect 5508 8792 5816 8820
rect 5508 8789 5520 8792
rect 5462 8783 5520 8789
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 6822 8820 6828 8832
rect 6604 8792 6828 8820
rect 6604 8780 6610 8792
rect 6822 8780 6828 8792
rect 6880 8820 6886 8832
rect 7926 8820 7932 8832
rect 6880 8792 7932 8820
rect 6880 8780 6886 8792
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8820 9183 8823
rect 9306 8820 9312 8832
rect 9171 8792 9312 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 10594 8780 10600 8832
rect 10652 8780 10658 8832
rect 11422 8780 11428 8832
rect 11480 8780 11486 8832
rect 11532 8820 11560 8851
rect 12158 8848 12164 8851
rect 12216 8848 12222 8900
rect 12342 8848 12348 8900
rect 12400 8848 12406 8900
rect 13648 8888 13676 8919
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 14349 8959 14407 8965
rect 14349 8956 14361 8959
rect 13780 8928 14361 8956
rect 13780 8916 13786 8928
rect 14349 8925 14361 8928
rect 14395 8925 14407 8959
rect 14349 8919 14407 8925
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 15160 8928 15669 8956
rect 15160 8916 15166 8928
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 17236 8956 17264 8987
rect 18340 8968 18368 8996
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 18322 8956 18328 8968
rect 17236 8928 18328 8956
rect 15657 8919 15715 8925
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 18969 8959 19027 8965
rect 18969 8925 18981 8959
rect 19015 8956 19027 8959
rect 19319 8959 19377 8965
rect 19319 8956 19331 8959
rect 19015 8928 19331 8956
rect 19015 8925 19027 8928
rect 18969 8919 19027 8925
rect 19319 8925 19331 8928
rect 19365 8925 19377 8959
rect 19319 8919 19377 8925
rect 19886 8916 19892 8968
rect 19944 8916 19950 8968
rect 13814 8888 13820 8900
rect 13648 8860 13820 8888
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 15924 8891 15982 8897
rect 15924 8857 15936 8891
rect 15970 8888 15982 8891
rect 16114 8888 16120 8900
rect 15970 8860 16120 8888
rect 15970 8857 15982 8860
rect 15924 8851 15982 8857
rect 16114 8848 16120 8860
rect 16172 8848 16178 8900
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 17466 8891 17524 8897
rect 17466 8888 17478 8891
rect 16908 8860 17478 8888
rect 16908 8848 16914 8860
rect 17466 8857 17478 8860
rect 17512 8857 17524 8891
rect 17466 8851 17524 8857
rect 19613 8891 19671 8897
rect 19613 8857 19625 8891
rect 19659 8888 19671 8891
rect 19702 8888 19708 8900
rect 19659 8860 19708 8888
rect 19659 8857 19671 8860
rect 19613 8851 19671 8857
rect 19702 8848 19708 8860
rect 19760 8848 19766 8900
rect 20432 8891 20490 8897
rect 20432 8857 20444 8891
rect 20478 8888 20490 8891
rect 20990 8888 20996 8900
rect 20478 8860 20996 8888
rect 20478 8857 20490 8860
rect 20432 8851 20490 8857
rect 20990 8848 20996 8860
rect 21048 8848 21054 8900
rect 13170 8820 13176 8832
rect 11532 8792 13176 8820
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 18414 8820 18420 8832
rect 15528 8792 18420 8820
rect 15528 8780 15534 8792
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 18785 8823 18843 8829
rect 18785 8789 18797 8823
rect 18831 8820 18843 8823
rect 18874 8820 18880 8832
rect 18831 8792 18880 8820
rect 18831 8789 18843 8792
rect 18785 8783 18843 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19797 8823 19855 8829
rect 19797 8789 19809 8823
rect 19843 8820 19855 8823
rect 20530 8820 20536 8832
rect 19843 8792 20536 8820
rect 19843 8789 19855 8792
rect 19797 8783 19855 8789
rect 20530 8780 20536 8792
rect 20588 8820 20594 8832
rect 20898 8820 20904 8832
rect 20588 8792 20904 8820
rect 20588 8780 20594 8792
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 21358 8780 21364 8832
rect 21416 8820 21422 8832
rect 21545 8823 21603 8829
rect 21545 8820 21557 8823
rect 21416 8792 21557 8820
rect 21416 8780 21422 8792
rect 21545 8789 21557 8792
rect 21591 8789 21603 8823
rect 21545 8783 21603 8789
rect 1104 8730 21988 8752
rect 1104 8678 4220 8730
rect 4272 8678 4284 8730
rect 4336 8678 4348 8730
rect 4400 8678 4412 8730
rect 4464 8678 4476 8730
rect 4528 8678 9441 8730
rect 9493 8678 9505 8730
rect 9557 8678 9569 8730
rect 9621 8678 9633 8730
rect 9685 8678 9697 8730
rect 9749 8678 14662 8730
rect 14714 8678 14726 8730
rect 14778 8678 14790 8730
rect 14842 8678 14854 8730
rect 14906 8678 14918 8730
rect 14970 8678 19883 8730
rect 19935 8678 19947 8730
rect 19999 8678 20011 8730
rect 20063 8678 20075 8730
rect 20127 8678 20139 8730
rect 20191 8678 21988 8730
rect 1104 8656 21988 8678
rect 5166 8576 5172 8628
rect 5224 8616 5230 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5224 8588 5457 8616
rect 5224 8576 5230 8588
rect 5445 8585 5457 8588
rect 5491 8585 5503 8619
rect 5445 8579 5503 8585
rect 7282 8576 7288 8628
rect 7340 8576 7346 8628
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 7926 8576 7932 8628
rect 7984 8576 7990 8628
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 14366 8616 14372 8628
rect 14323 8588 14372 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 17092 8588 18061 8616
rect 17092 8576 17098 8588
rect 18049 8585 18061 8588
rect 18095 8585 18107 8619
rect 19610 8616 19616 8628
rect 18049 8579 18107 8585
rect 18156 8588 19616 8616
rect 1670 8508 1676 8560
rect 1728 8548 1734 8560
rect 4614 8548 4620 8560
rect 1728 8520 4620 8548
rect 1728 8508 1734 8520
rect 1762 8440 1768 8492
rect 1820 8440 1826 8492
rect 2056 8489 2084 8520
rect 4080 8489 4108 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 6086 8508 6092 8560
rect 6144 8548 6150 8560
rect 6917 8551 6975 8557
rect 6917 8548 6929 8551
rect 6144 8520 6929 8548
rect 6144 8508 6150 8520
rect 6917 8517 6929 8520
rect 6963 8517 6975 8551
rect 6917 8511 6975 8517
rect 7374 8508 7380 8560
rect 7432 8508 7438 8560
rect 7561 8551 7619 8557
rect 7561 8517 7573 8551
rect 7607 8548 7619 8551
rect 8450 8551 8508 8557
rect 8450 8548 8462 8551
rect 7607 8520 8462 8548
rect 7607 8517 7619 8520
rect 7561 8511 7619 8517
rect 8450 8517 8462 8520
rect 8496 8517 8508 8551
rect 10226 8548 10232 8560
rect 8450 8511 8508 8517
rect 9876 8520 10232 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 2297 8483 2355 8489
rect 2297 8480 2309 8483
rect 2041 8443 2099 8449
rect 2148 8452 2309 8480
rect 2148 8412 2176 8452
rect 2297 8449 2309 8452
rect 2343 8449 2355 8483
rect 2297 8443 2355 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4321 8483 4379 8489
rect 4321 8480 4333 8483
rect 4212 8452 4333 8480
rect 4212 8440 4218 8452
rect 4321 8449 4333 8452
rect 4367 8449 4379 8483
rect 4321 8443 4379 8449
rect 5626 8440 5632 8492
rect 5684 8440 5690 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 7098 8440 7104 8492
rect 7156 8440 7162 8492
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8294 8480 8300 8492
rect 8159 8452 8300 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 9876 8489 9904 8520
rect 10226 8508 10232 8520
rect 10284 8548 10290 8560
rect 10502 8548 10508 8560
rect 10284 8520 10508 8548
rect 10284 8508 10290 8520
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 12618 8508 12624 8560
rect 12676 8508 12682 8560
rect 13164 8551 13222 8557
rect 13164 8517 13176 8551
rect 13210 8548 13222 8551
rect 13446 8548 13452 8560
rect 13210 8520 13452 8548
rect 13210 8517 13222 8520
rect 13164 8511 13222 8517
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 14090 8508 14096 8560
rect 14148 8548 14154 8560
rect 14550 8548 14556 8560
rect 14148 8520 14556 8548
rect 14148 8508 14154 8520
rect 14550 8508 14556 8520
rect 14608 8548 14614 8560
rect 15102 8548 15108 8560
rect 14608 8520 15108 8548
rect 14608 8508 14614 8520
rect 15102 8508 15108 8520
rect 15160 8548 15166 8560
rect 15197 8551 15255 8557
rect 15197 8548 15209 8551
rect 15160 8520 15209 8548
rect 15160 8508 15166 8520
rect 15197 8517 15209 8520
rect 15243 8517 15255 8551
rect 15197 8511 15255 8517
rect 15838 8508 15844 8560
rect 15896 8508 15902 8560
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 16942 8548 16948 8560
rect 15979 8520 16948 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17218 8508 17224 8560
rect 17276 8508 17282 8560
rect 18156 8557 18184 8588
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 21174 8576 21180 8628
rect 21232 8616 21238 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 21232 8588 21373 8616
rect 21232 8576 21238 8588
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 20254 8557 20260 8560
rect 18141 8551 18199 8557
rect 18141 8517 18153 8551
rect 18187 8517 18199 8551
rect 20248 8548 20260 8557
rect 18141 8511 18199 8517
rect 18340 8520 20024 8548
rect 20215 8520 20260 8548
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10128 8483 10186 8489
rect 10128 8449 10140 8483
rect 10174 8480 10186 8483
rect 10594 8480 10600 8492
rect 10174 8452 10600 8480
rect 10174 8449 10186 8452
rect 10128 8443 10186 8449
rect 1964 8384 2176 8412
rect 1964 8353 1992 8384
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 6788 8384 8217 8412
rect 6788 8372 6794 8384
rect 8205 8381 8217 8384
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 1949 8347 2007 8353
rect 1949 8313 1961 8347
rect 1995 8313 2007 8347
rect 1949 8307 2007 8313
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 3421 8279 3479 8285
rect 3421 8276 3433 8279
rect 3200 8248 3433 8276
rect 3200 8236 3206 8248
rect 3421 8245 3433 8248
rect 3467 8245 3479 8279
rect 3421 8239 3479 8245
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 5442 8276 5448 8288
rect 5040 8248 5448 8276
rect 5040 8236 5046 8248
rect 5442 8236 5448 8248
rect 5500 8276 5506 8288
rect 5629 8279 5687 8285
rect 5629 8276 5641 8279
rect 5500 8248 5641 8276
rect 5500 8236 5506 8248
rect 5629 8245 5641 8248
rect 5675 8245 5687 8279
rect 5629 8239 5687 8245
rect 6086 8236 6092 8288
rect 6144 8236 6150 8288
rect 8220 8276 8248 8375
rect 9876 8344 9904 8443
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8480 11851 8483
rect 11839 8452 12204 8480
rect 11839 8449 11851 8452
rect 11793 8443 11851 8449
rect 9508 8316 9904 8344
rect 11241 8347 11299 8353
rect 9122 8276 9128 8288
rect 8220 8248 9128 8276
rect 9122 8236 9128 8248
rect 9180 8276 9186 8288
rect 9508 8276 9536 8316
rect 11241 8313 11253 8347
rect 11287 8344 11299 8347
rect 11422 8344 11428 8356
rect 11287 8316 11428 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 11422 8304 11428 8316
rect 11480 8344 11486 8356
rect 11882 8344 11888 8356
rect 11480 8316 11888 8344
rect 11480 8304 11486 8316
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 12176 8353 12204 8452
rect 12342 8440 12348 8492
rect 12400 8480 12406 8492
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12400 8452 12909 8480
rect 12400 8440 12406 8452
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13004 8452 14412 8480
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 12621 8415 12679 8421
rect 12621 8412 12633 8415
rect 12584 8384 12633 8412
rect 12584 8372 12590 8384
rect 12621 8381 12633 8384
rect 12667 8381 12679 8415
rect 12621 8375 12679 8381
rect 12161 8347 12219 8353
rect 12161 8313 12173 8347
rect 12207 8313 12219 8347
rect 12636 8344 12664 8375
rect 12710 8372 12716 8424
rect 12768 8372 12774 8424
rect 13004 8412 13032 8452
rect 12820 8384 13032 8412
rect 14384 8412 14412 8452
rect 14458 8440 14464 8492
rect 14516 8440 14522 8492
rect 15856 8480 15884 8508
rect 18340 8492 18368 8520
rect 17954 8480 17960 8492
rect 15856 8452 17960 8480
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18230 8480 18236 8492
rect 18064 8452 18236 8480
rect 15102 8412 15108 8424
rect 14384 8384 15108 8412
rect 12820 8344 12848 8384
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 15746 8372 15752 8424
rect 15804 8412 15810 8424
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15804 8384 15945 8412
rect 15804 8372 15810 8384
rect 15933 8381 15945 8384
rect 15979 8381 15991 8415
rect 15933 8375 15991 8381
rect 17126 8372 17132 8424
rect 17184 8372 17190 8424
rect 17310 8372 17316 8424
rect 17368 8372 17374 8424
rect 18064 8421 18092 8452
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 18322 8440 18328 8492
rect 18380 8440 18386 8492
rect 18592 8483 18650 8489
rect 18592 8449 18604 8483
rect 18638 8480 18650 8483
rect 18874 8480 18880 8492
rect 18638 8452 18880 8480
rect 18638 8449 18650 8452
rect 18592 8443 18650 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 19996 8489 20024 8520
rect 20248 8511 20260 8520
rect 20254 8508 20260 8511
rect 20312 8508 20318 8560
rect 19981 8483 20039 8489
rect 19981 8449 19993 8483
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 12636 8316 12848 8344
rect 12161 8307 12219 8313
rect 13906 8304 13912 8356
rect 13964 8344 13970 8356
rect 14458 8344 14464 8356
rect 13964 8316 14464 8344
rect 13964 8304 13970 8316
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 16393 8347 16451 8353
rect 16393 8313 16405 8347
rect 16439 8344 16451 8347
rect 18230 8344 18236 8356
rect 16439 8316 18236 8344
rect 16439 8313 16451 8316
rect 16393 8307 16451 8313
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 9180 8248 9536 8276
rect 9180 8236 9186 8248
rect 9582 8236 9588 8288
rect 9640 8236 9646 8288
rect 11514 8236 11520 8288
rect 11572 8236 11578 8288
rect 11977 8279 12035 8285
rect 11977 8245 11989 8279
rect 12023 8276 12035 8279
rect 12066 8276 12072 8288
rect 12023 8248 12072 8276
rect 12023 8245 12035 8248
rect 11977 8239 12035 8245
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 16758 8236 16764 8288
rect 16816 8236 16822 8288
rect 17586 8236 17592 8288
rect 17644 8236 17650 8288
rect 19702 8236 19708 8288
rect 19760 8236 19766 8288
rect 1104 8186 21988 8208
rect 1104 8134 3560 8186
rect 3612 8134 3624 8186
rect 3676 8134 3688 8186
rect 3740 8134 3752 8186
rect 3804 8134 3816 8186
rect 3868 8134 8781 8186
rect 8833 8134 8845 8186
rect 8897 8134 8909 8186
rect 8961 8134 8973 8186
rect 9025 8134 9037 8186
rect 9089 8134 14002 8186
rect 14054 8134 14066 8186
rect 14118 8134 14130 8186
rect 14182 8134 14194 8186
rect 14246 8134 14258 8186
rect 14310 8134 19223 8186
rect 19275 8134 19287 8186
rect 19339 8134 19351 8186
rect 19403 8134 19415 8186
rect 19467 8134 19479 8186
rect 19531 8134 21988 8186
rect 1104 8112 21988 8134
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 5626 8072 5632 8084
rect 4387 8044 5632 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 7156 8044 7297 8072
rect 7156 8032 7162 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 8386 8072 8392 8084
rect 7285 8035 7343 8041
rect 7852 8044 8392 8072
rect 4617 8007 4675 8013
rect 4617 7973 4629 8007
rect 4663 8004 4675 8007
rect 4706 8004 4712 8016
rect 4663 7976 4712 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 3050 7896 3056 7948
rect 3108 7936 3114 7948
rect 5169 7939 5227 7945
rect 3108 7908 3832 7936
rect 3108 7896 3114 7908
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 2866 7868 2872 7880
rect 1903 7840 2872 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 2866 7828 2872 7840
rect 2924 7868 2930 7880
rect 3510 7868 3516 7880
rect 2924 7840 3516 7868
rect 2924 7828 2930 7840
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3804 7877 3832 7908
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5258 7936 5264 7948
rect 5215 7908 5264 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3789 7831 3847 7837
rect 3896 7840 4077 7868
rect 2124 7803 2182 7809
rect 2124 7769 2136 7803
rect 2170 7800 2182 7803
rect 2222 7800 2228 7812
rect 2170 7772 2228 7800
rect 2170 7769 2182 7772
rect 2124 7763 2182 7769
rect 2222 7760 2228 7772
rect 2280 7760 2286 7812
rect 3142 7760 3148 7812
rect 3200 7800 3206 7812
rect 3896 7800 3924 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4154 7828 4160 7880
rect 4212 7877 4218 7880
rect 4212 7868 4220 7877
rect 5350 7868 5356 7880
rect 4212 7840 5356 7868
rect 4212 7831 4220 7840
rect 4212 7828 4218 7831
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6730 7868 6736 7880
rect 5951 7840 6736 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 7300 7868 7328 8035
rect 7852 7877 7880 8044
rect 8386 8032 8392 8044
rect 8444 8072 8450 8084
rect 9030 8072 9036 8084
rect 8444 8044 9036 8072
rect 8444 8032 8450 8044
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 10134 8032 10140 8084
rect 10192 8032 10198 8084
rect 12342 8072 12348 8084
rect 11992 8044 12348 8072
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7936 9827 7939
rect 10226 7936 10232 7948
rect 9815 7908 10232 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11992 7945 12020 8044
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 13357 8075 13415 8081
rect 13357 8072 13369 8075
rect 12676 8044 13369 8072
rect 12676 8032 12682 8044
rect 13357 8041 13369 8044
rect 13403 8041 13415 8075
rect 13357 8035 13415 8041
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 13872 8044 15117 8072
rect 13872 8032 13878 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 16942 8032 16948 8084
rect 17000 8032 17006 8084
rect 20622 8032 20628 8084
rect 20680 8032 20686 8084
rect 14274 7964 14280 8016
rect 14332 8004 14338 8016
rect 15381 8007 15439 8013
rect 15381 8004 15393 8007
rect 14332 7976 15393 8004
rect 14332 7964 14338 7976
rect 15381 7973 15393 7976
rect 15427 7973 15439 8007
rect 15381 7967 15439 7973
rect 16482 7964 16488 8016
rect 16540 8004 16546 8016
rect 17310 8004 17316 8016
rect 16540 7976 17316 8004
rect 16540 7964 16546 7976
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 20901 8007 20959 8013
rect 20901 7973 20913 8007
rect 20947 8004 20959 8007
rect 21174 8004 21180 8016
rect 20947 7976 21180 8004
rect 20947 7973 20959 7976
rect 20901 7967 20959 7973
rect 21174 7964 21180 7976
rect 21232 7964 21238 8016
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7905 12035 7939
rect 11977 7899 12035 7905
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 16758 7936 16764 7948
rect 14056 7908 16764 7936
rect 14056 7896 14062 7908
rect 16758 7896 16764 7908
rect 16816 7896 16822 7948
rect 18322 7896 18328 7948
rect 18380 7936 18386 7948
rect 19245 7939 19303 7945
rect 19245 7936 19257 7939
rect 18380 7908 19257 7936
rect 18380 7896 18386 7908
rect 19245 7905 19257 7908
rect 19291 7905 19303 7939
rect 19245 7899 19303 7905
rect 21358 7896 21364 7948
rect 21416 7896 21422 7948
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 7300 7840 7757 7868
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 7984 7840 8309 7868
rect 7984 7828 7990 7840
rect 8297 7837 8309 7840
rect 8343 7868 8355 7871
rect 8386 7868 8392 7880
rect 8343 7840 8392 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10496 7871 10554 7877
rect 10496 7837 10508 7871
rect 10542 7868 10554 7871
rect 11514 7868 11520 7880
rect 10542 7840 11520 7868
rect 10542 7837 10554 7840
rect 10496 7831 10554 7837
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 12066 7828 12072 7880
rect 12124 7868 12130 7880
rect 12233 7871 12291 7877
rect 12233 7868 12245 7871
rect 12124 7840 12245 7868
rect 12124 7828 12130 7840
rect 12233 7837 12245 7840
rect 12279 7837 12291 7871
rect 12233 7831 12291 7837
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7868 14887 7871
rect 15010 7868 15016 7880
rect 14875 7840 15016 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 15010 7828 15016 7840
rect 15068 7868 15074 7880
rect 15657 7871 15715 7877
rect 15657 7868 15669 7871
rect 15068 7840 15669 7868
rect 15068 7828 15074 7840
rect 15657 7837 15669 7840
rect 15703 7868 15715 7871
rect 15746 7868 15752 7880
rect 15703 7840 15752 7868
rect 15703 7837 15715 7840
rect 15657 7831 15715 7837
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 17218 7868 17224 7880
rect 15856 7840 17224 7868
rect 15856 7812 15884 7840
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 18230 7828 18236 7880
rect 18288 7868 18294 7880
rect 18601 7871 18659 7877
rect 18601 7868 18613 7871
rect 18288 7840 18613 7868
rect 18288 7828 18294 7840
rect 18601 7837 18613 7840
rect 18647 7837 18659 7871
rect 18601 7831 18659 7837
rect 18874 7828 18880 7880
rect 18932 7828 18938 7880
rect 21082 7828 21088 7880
rect 21140 7868 21146 7880
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 21140 7840 21465 7868
rect 21140 7828 21146 7840
rect 21453 7837 21465 7840
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 3200 7772 3924 7800
rect 3200 7760 3206 7772
rect 3970 7760 3976 7812
rect 4028 7760 4034 7812
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7769 4951 7803
rect 4893 7763 4951 7769
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3237 7735 3295 7741
rect 3237 7732 3249 7735
rect 3108 7704 3249 7732
rect 3108 7692 3114 7704
rect 3237 7701 3249 7704
rect 3283 7701 3295 7735
rect 3237 7695 3295 7701
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 4908 7732 4936 7763
rect 5074 7760 5080 7812
rect 5132 7760 5138 7812
rect 6172 7803 6230 7809
rect 6172 7769 6184 7803
rect 6218 7800 6230 7803
rect 6546 7800 6552 7812
rect 6218 7772 6552 7800
rect 6218 7769 6230 7772
rect 6172 7763 6230 7769
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 8113 7803 8171 7809
rect 8113 7800 8125 7803
rect 7708 7772 8125 7800
rect 7708 7760 7714 7772
rect 8113 7769 8125 7772
rect 8159 7769 8171 7803
rect 8113 7763 8171 7769
rect 8478 7760 8484 7812
rect 8536 7760 8542 7812
rect 8941 7803 8999 7809
rect 8941 7769 8953 7803
rect 8987 7800 8999 7803
rect 9214 7800 9220 7812
rect 8987 7772 9220 7800
rect 8987 7769 8999 7772
rect 8941 7763 8999 7769
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 12710 7760 12716 7812
rect 12768 7800 12774 7812
rect 14553 7803 14611 7809
rect 14553 7800 14565 7803
rect 12768 7772 14565 7800
rect 12768 7760 12774 7772
rect 14553 7769 14565 7772
rect 14599 7769 14611 7803
rect 14553 7763 14611 7769
rect 15838 7760 15844 7812
rect 15896 7760 15902 7812
rect 15933 7803 15991 7809
rect 15933 7769 15945 7803
rect 15979 7800 15991 7803
rect 16022 7800 16028 7812
rect 15979 7772 16028 7800
rect 15979 7769 15991 7772
rect 15933 7763 15991 7769
rect 16022 7760 16028 7772
rect 16080 7760 16086 7812
rect 16206 7760 16212 7812
rect 16264 7760 16270 7812
rect 18080 7803 18138 7809
rect 18080 7769 18092 7803
rect 18126 7800 18138 7803
rect 19512 7803 19570 7809
rect 18126 7772 18460 7800
rect 18126 7769 18138 7772
rect 18080 7763 18138 7769
rect 3844 7704 4936 7732
rect 3844 7692 3850 7704
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7432 7704 7573 7732
rect 7432 7692 7438 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 11609 7735 11667 7741
rect 11609 7732 11621 7735
rect 11296 7704 11621 7732
rect 11296 7692 11302 7704
rect 11609 7701 11621 7704
rect 11655 7732 11667 7735
rect 12342 7732 12348 7744
rect 11655 7704 12348 7732
rect 11655 7701 11667 7704
rect 11609 7695 11667 7701
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 18432 7741 18460 7772
rect 19512 7769 19524 7803
rect 19558 7800 19570 7803
rect 19794 7800 19800 7812
rect 19558 7772 19800 7800
rect 19558 7769 19570 7772
rect 19512 7763 19570 7769
rect 19794 7760 19800 7772
rect 19852 7760 19858 7812
rect 21266 7760 21272 7812
rect 21324 7800 21330 7812
rect 21361 7803 21419 7809
rect 21361 7800 21373 7803
rect 21324 7772 21373 7800
rect 21324 7760 21330 7772
rect 21361 7769 21373 7772
rect 21407 7769 21419 7803
rect 21361 7763 21419 7769
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14424 7704 14657 7732
rect 14424 7692 14430 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 18417 7735 18475 7741
rect 18417 7701 18429 7735
rect 18463 7701 18475 7735
rect 18417 7695 18475 7701
rect 18690 7692 18696 7744
rect 18748 7692 18754 7744
rect 1104 7642 21988 7664
rect 1104 7590 4220 7642
rect 4272 7590 4284 7642
rect 4336 7590 4348 7642
rect 4400 7590 4412 7642
rect 4464 7590 4476 7642
rect 4528 7590 9441 7642
rect 9493 7590 9505 7642
rect 9557 7590 9569 7642
rect 9621 7590 9633 7642
rect 9685 7590 9697 7642
rect 9749 7590 14662 7642
rect 14714 7590 14726 7642
rect 14778 7590 14790 7642
rect 14842 7590 14854 7642
rect 14906 7590 14918 7642
rect 14970 7590 19883 7642
rect 19935 7590 19947 7642
rect 19999 7590 20011 7642
rect 20063 7590 20075 7642
rect 20127 7590 20139 7642
rect 20191 7590 21988 7642
rect 1104 7568 21988 7590
rect 2222 7488 2228 7540
rect 2280 7488 2286 7540
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 5258 7528 5264 7540
rect 4488 7500 5264 7528
rect 4488 7488 4494 7500
rect 5258 7488 5264 7500
rect 5316 7528 5322 7540
rect 5442 7528 5448 7540
rect 5316 7500 5448 7528
rect 5316 7488 5322 7500
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6546 7488 6552 7540
rect 6604 7488 6610 7540
rect 6733 7531 6791 7537
rect 6733 7497 6745 7531
rect 6779 7497 6791 7531
rect 6733 7491 6791 7497
rect 3510 7420 3516 7472
rect 3568 7420 3574 7472
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 5074 7460 5080 7472
rect 4028 7432 5080 7460
rect 4028 7420 4034 7432
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 6086 7420 6092 7472
rect 6144 7460 6150 7472
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 6144 7432 6653 7460
rect 6144 7420 6150 7432
rect 6641 7429 6653 7432
rect 6687 7429 6699 7463
rect 6641 7423 6699 7429
rect 2406 7352 2412 7404
rect 2464 7352 2470 7404
rect 2774 7352 2780 7404
rect 2832 7352 2838 7404
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3292 7364 3801 7392
rect 3292 7352 3298 7364
rect 3789 7361 3801 7364
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4162 7395 4220 7401
rect 4162 7361 4174 7395
rect 4208 7361 4220 7395
rect 4162 7355 4220 7361
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 4080 7324 4108 7355
rect 3108 7296 4108 7324
rect 3108 7284 3114 7296
rect 3878 7216 3884 7268
rect 3936 7256 3942 7268
rect 4062 7256 4068 7268
rect 3936 7228 4068 7256
rect 3936 7216 3942 7228
rect 4062 7216 4068 7228
rect 4120 7256 4126 7268
rect 4172 7256 4200 7355
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5902 7392 5908 7404
rect 5215 7364 5908 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 4985 7327 5043 7333
rect 4985 7293 4997 7327
rect 5031 7293 5043 7327
rect 6748 7324 6776 7491
rect 6822 7488 6828 7540
rect 6880 7488 6886 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 7340 7500 7757 7528
rect 7340 7488 7346 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 8294 7488 8300 7540
rect 8352 7488 8358 7540
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 8481 7531 8539 7537
rect 8481 7528 8493 7531
rect 8444 7500 8493 7528
rect 8444 7488 8450 7500
rect 8481 7497 8493 7500
rect 8527 7497 8539 7531
rect 8481 7491 8539 7497
rect 9306 7488 9312 7540
rect 9364 7528 9370 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9364 7500 9597 7528
rect 9364 7488 9370 7500
rect 9585 7497 9597 7500
rect 9631 7528 9643 7531
rect 10318 7528 10324 7540
rect 9631 7500 10324 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 15654 7528 15660 7540
rect 11900 7500 15660 7528
rect 7009 7463 7067 7469
rect 7009 7429 7021 7463
rect 7055 7460 7067 7463
rect 7374 7460 7380 7472
rect 7055 7432 7380 7460
rect 7055 7429 7067 7432
rect 7009 7423 7067 7429
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 7466 7420 7472 7472
rect 7524 7460 7530 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 7524 7432 7849 7460
rect 7524 7420 7530 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 8312 7460 8340 7488
rect 8941 7463 8999 7469
rect 8941 7460 8953 7463
rect 8312 7432 8953 7460
rect 7837 7423 7895 7429
rect 8941 7429 8953 7432
rect 8987 7429 8999 7463
rect 8941 7423 8999 7429
rect 9030 7420 9036 7472
rect 9088 7460 9094 7472
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 9088 7432 9505 7460
rect 9088 7420 9094 7432
rect 9493 7429 9505 7432
rect 9539 7429 9551 7463
rect 9493 7423 9551 7429
rect 9766 7420 9772 7472
rect 9824 7420 9830 7472
rect 11900 7469 11928 7500
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 15933 7531 15991 7537
rect 15933 7528 15945 7531
rect 15896 7500 15945 7528
rect 15896 7488 15902 7500
rect 15933 7497 15945 7500
rect 15979 7497 15991 7531
rect 15933 7491 15991 7497
rect 16114 7488 16120 7540
rect 16172 7488 16178 7540
rect 16850 7488 16856 7540
rect 16908 7488 16914 7540
rect 17034 7488 17040 7540
rect 17092 7488 17098 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18966 7528 18972 7540
rect 18012 7500 18972 7528
rect 18012 7488 18018 7500
rect 18966 7488 18972 7500
rect 19024 7528 19030 7540
rect 19024 7500 19196 7528
rect 19024 7488 19030 7500
rect 11885 7463 11943 7469
rect 11885 7429 11897 7463
rect 11931 7429 11943 7463
rect 11885 7423 11943 7429
rect 11974 7420 11980 7472
rect 12032 7460 12038 7472
rect 12069 7463 12127 7469
rect 12069 7460 12081 7463
rect 12032 7432 12081 7460
rect 12032 7420 12038 7432
rect 12069 7429 12081 7432
rect 12115 7429 12127 7463
rect 12069 7423 12127 7429
rect 12894 7420 12900 7472
rect 12952 7420 12958 7472
rect 14798 7463 14856 7469
rect 14798 7460 14810 7463
rect 14476 7432 14810 7460
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7650 7392 7656 7404
rect 7607 7364 7656 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 8435 7395 8493 7401
rect 8435 7361 8447 7395
rect 8481 7392 8493 7395
rect 8570 7392 8576 7404
rect 8481 7364 8576 7392
rect 8481 7361 8493 7364
rect 8435 7355 8493 7361
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 6748 7296 7389 7324
rect 4985 7287 5043 7293
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 8312 7324 8340 7355
rect 8570 7352 8576 7364
rect 8628 7352 8634 7404
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8312 7296 8616 7324
rect 7377 7287 7435 7293
rect 4120 7228 4200 7256
rect 4341 7259 4399 7265
rect 4120 7216 4126 7228
rect 4341 7225 4353 7259
rect 4387 7256 4399 7259
rect 5000 7256 5028 7287
rect 4387 7228 5028 7256
rect 5353 7259 5411 7265
rect 4387 7225 4399 7228
rect 4341 7219 4399 7225
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 7742 7256 7748 7268
rect 5399 7228 7748 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 7742 7216 7748 7228
rect 7800 7216 7806 7268
rect 8113 7259 8171 7265
rect 8113 7225 8125 7259
rect 8159 7256 8171 7259
rect 8294 7256 8300 7268
rect 8159 7228 8300 7256
rect 8159 7225 8171 7228
rect 8113 7219 8171 7225
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 4982 7148 4988 7200
rect 5040 7148 5046 7200
rect 8588 7188 8616 7296
rect 8680 7256 8708 7355
rect 9048 7324 9076 7420
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9784 7392 9812 7420
rect 9171 7364 9812 7392
rect 12713 7395 12771 7401
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 12713 7361 12725 7395
rect 12759 7392 12771 7395
rect 13538 7392 13544 7404
rect 12759 7364 13544 7392
rect 12759 7361 12771 7364
rect 12713 7355 12771 7361
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13998 7352 14004 7404
rect 14056 7352 14062 7404
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 9309 7327 9367 7333
rect 9309 7324 9321 7327
rect 9048 7296 9321 7324
rect 9309 7293 9321 7296
rect 9355 7324 9367 7327
rect 9766 7324 9772 7336
rect 9355 7296 9772 7324
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7324 12219 7327
rect 12618 7324 12624 7336
rect 12207 7296 12624 7324
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 12618 7284 12624 7296
rect 12676 7324 12682 7336
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12676 7296 13001 7324
rect 12676 7284 12682 7296
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 9674 7256 9680 7268
rect 8680 7228 9680 7256
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 10045 7259 10103 7265
rect 10045 7256 10057 7259
rect 10008 7228 10057 7256
rect 10008 7216 10014 7228
rect 10045 7225 10057 7228
rect 10091 7225 10103 7259
rect 10045 7219 10103 7225
rect 11606 7216 11612 7268
rect 11664 7216 11670 7268
rect 14476 7265 14504 7432
rect 14798 7429 14810 7432
rect 14844 7429 14856 7463
rect 14798 7423 14856 7429
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 18172 7463 18230 7469
rect 15160 7432 18000 7460
rect 15160 7420 15166 7432
rect 14550 7352 14556 7404
rect 14608 7352 14614 7404
rect 16298 7352 16304 7404
rect 16356 7352 16362 7404
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7392 16727 7395
rect 17586 7392 17592 7404
rect 16715 7364 17592 7392
rect 16715 7361 16727 7364
rect 16669 7355 16727 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17972 7392 18000 7432
rect 18172 7429 18184 7463
rect 18218 7460 18230 7463
rect 18690 7460 18696 7472
rect 18218 7432 18696 7460
rect 18218 7429 18230 7432
rect 18172 7423 18230 7429
rect 18690 7420 18696 7432
rect 18748 7420 18754 7472
rect 18782 7420 18788 7472
rect 18840 7460 18846 7472
rect 19168 7469 19196 7500
rect 19702 7488 19708 7540
rect 19760 7528 19766 7540
rect 19889 7531 19947 7537
rect 19889 7528 19901 7531
rect 19760 7500 19901 7528
rect 19760 7488 19766 7500
rect 19889 7497 19901 7500
rect 19935 7497 19947 7531
rect 19889 7491 19947 7497
rect 20456 7500 20852 7528
rect 19061 7463 19119 7469
rect 19061 7460 19073 7463
rect 18840 7432 19073 7460
rect 18840 7420 18846 7432
rect 19061 7429 19073 7432
rect 19107 7429 19119 7463
rect 19061 7423 19119 7429
rect 19153 7463 19211 7469
rect 19153 7429 19165 7463
rect 19199 7460 19211 7463
rect 20456 7460 20484 7500
rect 20824 7472 20852 7500
rect 20990 7488 20996 7540
rect 21048 7488 21054 7540
rect 19199 7432 20484 7460
rect 19199 7429 19211 7432
rect 19153 7423 19211 7429
rect 20530 7420 20536 7472
rect 20588 7420 20594 7472
rect 20622 7420 20628 7472
rect 20680 7420 20686 7472
rect 20714 7420 20720 7472
rect 20772 7420 20778 7472
rect 20806 7420 20812 7472
rect 20864 7420 20870 7472
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 17972 7364 18889 7392
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 19705 7395 19763 7401
rect 19705 7361 19717 7395
rect 19751 7392 19763 7395
rect 20640 7392 20668 7420
rect 19751 7364 20668 7392
rect 19751 7361 19763 7364
rect 19705 7355 19763 7361
rect 21174 7352 21180 7404
rect 21232 7352 21238 7404
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 14461 7259 14519 7265
rect 14461 7225 14473 7259
rect 14507 7225 14519 7259
rect 18432 7256 18460 7287
rect 19610 7284 19616 7336
rect 19668 7324 19674 7336
rect 19981 7327 20039 7333
rect 19981 7324 19993 7327
rect 19668 7296 19993 7324
rect 19668 7284 19674 7296
rect 19981 7293 19993 7296
rect 20027 7324 20039 7327
rect 20990 7324 20996 7336
rect 20027 7296 20996 7324
rect 20027 7293 20039 7296
rect 19981 7287 20039 7293
rect 20990 7284 20996 7296
rect 21048 7284 21054 7336
rect 19058 7256 19064 7268
rect 18432 7228 19064 7256
rect 14461 7219 14519 7225
rect 19058 7216 19064 7228
rect 19116 7216 19122 7268
rect 19429 7259 19487 7265
rect 19429 7225 19441 7259
rect 19475 7256 19487 7259
rect 19702 7256 19708 7268
rect 19475 7228 19708 7256
rect 19475 7225 19487 7228
rect 19429 7219 19487 7225
rect 19702 7216 19708 7228
rect 19760 7216 19766 7268
rect 9858 7188 9864 7200
rect 8588 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 12434 7148 12440 7200
rect 12492 7148 12498 7200
rect 14185 7191 14243 7197
rect 14185 7157 14197 7191
rect 14231 7188 14243 7191
rect 14826 7188 14832 7200
rect 14231 7160 14832 7188
rect 14231 7157 14243 7160
rect 14185 7151 14243 7157
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 18598 7148 18604 7200
rect 18656 7148 18662 7200
rect 19610 7148 19616 7200
rect 19668 7188 19674 7200
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 19668 7160 20269 7188
rect 19668 7148 19674 7160
rect 20257 7157 20269 7160
rect 20303 7157 20315 7191
rect 20257 7151 20315 7157
rect 1104 7098 21988 7120
rect 1104 7046 3560 7098
rect 3612 7046 3624 7098
rect 3676 7046 3688 7098
rect 3740 7046 3752 7098
rect 3804 7046 3816 7098
rect 3868 7046 8781 7098
rect 8833 7046 8845 7098
rect 8897 7046 8909 7098
rect 8961 7046 8973 7098
rect 9025 7046 9037 7098
rect 9089 7046 14002 7098
rect 14054 7046 14066 7098
rect 14118 7046 14130 7098
rect 14182 7046 14194 7098
rect 14246 7046 14258 7098
rect 14310 7046 19223 7098
rect 19275 7046 19287 7098
rect 19339 7046 19351 7098
rect 19403 7046 19415 7098
rect 19467 7046 19479 7098
rect 19531 7046 21988 7098
rect 1104 7024 21988 7046
rect 1857 6987 1915 6993
rect 1857 6953 1869 6987
rect 1903 6984 1915 6987
rect 2406 6984 2412 6996
rect 1903 6956 2412 6984
rect 1903 6953 1915 6956
rect 1857 6947 1915 6953
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 4948 6956 5181 6984
rect 4948 6944 4954 6956
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 5169 6947 5227 6953
rect 7377 6987 7435 6993
rect 7377 6953 7389 6987
rect 7423 6984 7435 6987
rect 7650 6984 7656 6996
rect 7423 6956 7656 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 7650 6944 7656 6956
rect 7708 6944 7714 6996
rect 17957 6987 18015 6993
rect 17957 6953 17969 6987
rect 18003 6984 18015 6987
rect 18874 6984 18880 6996
rect 18003 6956 18880 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 20714 6944 20720 6996
rect 20772 6944 20778 6996
rect 2685 6919 2743 6925
rect 2685 6916 2697 6919
rect 2663 6888 2697 6916
rect 2685 6885 2697 6888
rect 2731 6885 2743 6919
rect 2685 6879 2743 6885
rect 2792 6888 3096 6916
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 2700 6848 2728 6879
rect 1820 6820 2728 6848
rect 1820 6808 1826 6820
rect 1118 6740 1124 6792
rect 1176 6780 1182 6792
rect 2133 6783 2191 6789
rect 2133 6780 2145 6783
rect 1176 6752 2145 6780
rect 1176 6740 1182 6752
rect 2133 6749 2145 6752
rect 2179 6749 2191 6783
rect 2133 6743 2191 6749
rect 2314 6740 2320 6792
rect 2372 6740 2378 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2792 6780 2820 6888
rect 2958 6848 2964 6860
rect 2455 6752 2820 6780
rect 2884 6820 2964 6848
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2332 6712 2360 6740
rect 2884 6712 2912 6820
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 3068 6848 3096 6888
rect 5902 6876 5908 6928
rect 5960 6916 5966 6928
rect 9122 6916 9128 6928
rect 5960 6888 6960 6916
rect 5960 6876 5966 6888
rect 3237 6851 3295 6857
rect 3237 6848 3249 6851
rect 3068 6820 3249 6848
rect 3237 6817 3249 6820
rect 3283 6848 3295 6851
rect 3326 6848 3332 6860
rect 3283 6820 3332 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3326 6808 3332 6820
rect 3384 6808 3390 6860
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 5258 6848 5264 6860
rect 4387 6820 5264 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 6822 6848 6828 6860
rect 5776 6820 6828 6848
rect 5776 6808 5782 6820
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 6932 6848 6960 6888
rect 8772 6888 9128 6916
rect 6932 6820 7144 6848
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 3863 6783 3921 6789
rect 3863 6780 3875 6783
rect 3651 6752 3875 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 3863 6749 3875 6752
rect 3909 6749 3921 6783
rect 3863 6743 3921 6749
rect 4430 6740 4436 6792
rect 4488 6740 4494 6792
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 4706 6780 4712 6792
rect 4663 6752 4712 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5037 6783 5095 6789
rect 5037 6749 5049 6783
rect 5083 6780 5095 6783
rect 5353 6783 5411 6789
rect 5083 6749 5120 6780
rect 5037 6743 5120 6749
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 6454 6780 6460 6792
rect 5399 6752 6460 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 2332 6684 2912 6712
rect 2958 6672 2964 6724
rect 3016 6672 3022 6724
rect 3142 6672 3148 6724
rect 3200 6672 3206 6724
rect 4798 6672 4804 6724
rect 4856 6672 4862 6724
rect 4893 6715 4951 6721
rect 4893 6681 4905 6715
rect 4939 6681 4951 6715
rect 4893 6675 4951 6681
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 3050 6644 3056 6656
rect 2363 6616 3056 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3418 6604 3424 6656
rect 3476 6604 3482 6656
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 4614 6644 4620 6656
rect 4387 6616 4620 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 4614 6604 4620 6616
rect 4672 6644 4678 6656
rect 4908 6644 4936 6675
rect 4672 6616 4936 6644
rect 5092 6644 5120 6743
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 7116 6780 7144 6820
rect 7190 6808 7196 6860
rect 7248 6808 7254 6860
rect 8772 6857 8800 6888
rect 9122 6876 9128 6888
rect 9180 6876 9186 6928
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9824 6888 10088 6916
rect 9824 6876 9830 6888
rect 10060 6857 10088 6888
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6817 8815 6851
rect 10045 6851 10103 6857
rect 8757 6811 8815 6817
rect 9140 6820 9996 6848
rect 9140 6780 9168 6820
rect 7116 6752 9168 6780
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 9508 6789 9536 6820
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 5166 6672 5172 6724
rect 5224 6712 5230 6724
rect 5537 6715 5595 6721
rect 5537 6712 5549 6715
rect 5224 6684 5549 6712
rect 5224 6672 5230 6684
rect 5537 6681 5549 6684
rect 5583 6681 5595 6715
rect 5537 6675 5595 6681
rect 5905 6715 5963 6721
rect 5905 6681 5917 6715
rect 5951 6712 5963 6715
rect 6825 6715 6883 6721
rect 6825 6712 6837 6715
rect 5951 6684 6837 6712
rect 5951 6681 5963 6684
rect 5905 6675 5963 6681
rect 6825 6681 6837 6684
rect 6871 6681 6883 6715
rect 6825 6675 6883 6681
rect 7926 6672 7932 6724
rect 7984 6712 7990 6724
rect 8490 6715 8548 6721
rect 8490 6712 8502 6715
rect 7984 6684 8502 6712
rect 7984 6672 7990 6684
rect 8490 6681 8502 6684
rect 8536 6681 8548 6715
rect 8490 6675 8548 6681
rect 9582 6672 9588 6724
rect 9640 6712 9646 6724
rect 9876 6712 9904 6743
rect 9640 6684 9904 6712
rect 9968 6712 9996 6820
rect 10045 6817 10057 6851
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6848 13047 6851
rect 13906 6848 13912 6860
rect 13035 6820 13912 6848
rect 13035 6817 13047 6820
rect 12989 6811 13047 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 17034 6808 17040 6860
rect 17092 6848 17098 6860
rect 17497 6851 17555 6857
rect 17497 6848 17509 6851
rect 17092 6820 17509 6848
rect 17092 6808 17098 6820
rect 17497 6817 17509 6820
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 18064 6820 19472 6848
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10042 6712 10048 6724
rect 9968 6684 10048 6712
rect 9640 6672 9646 6684
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 10152 6712 10180 6743
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 10284 6752 10333 6780
rect 10284 6740 10290 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 12434 6780 12440 6792
rect 12391 6752 12440 6780
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 14550 6740 14556 6792
rect 14608 6740 14614 6792
rect 14826 6789 14832 6792
rect 14820 6780 14832 6789
rect 14787 6752 14832 6780
rect 14820 6743 14832 6752
rect 14826 6740 14832 6743
rect 14884 6740 14890 6792
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 16264 6752 16405 6780
rect 16264 6740 16270 6752
rect 16393 6749 16405 6752
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 16807 6752 17417 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 17405 6749 17417 6752
rect 17451 6780 17463 6783
rect 18064 6780 18092 6820
rect 17451 6752 18092 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 18138 6740 18144 6792
rect 18196 6740 18202 6792
rect 19337 6783 19395 6789
rect 19337 6780 19349 6783
rect 19076 6752 19349 6780
rect 19076 6724 19104 6752
rect 19337 6749 19349 6752
rect 19383 6749 19395 6783
rect 19444 6780 19472 6820
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21545 6851 21603 6857
rect 21545 6848 21557 6851
rect 21048 6820 21557 6848
rect 21048 6808 21054 6820
rect 21545 6817 21557 6820
rect 21591 6817 21603 6851
rect 21545 6811 21603 6817
rect 21008 6780 21036 6808
rect 19444 6752 21036 6780
rect 19337 6743 19395 6749
rect 10410 6712 10416 6724
rect 10152 6684 10416 6712
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 10502 6672 10508 6724
rect 10560 6672 10566 6724
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 12989 6715 13047 6721
rect 12989 6712 13001 6715
rect 12952 6684 13001 6712
rect 12952 6672 12958 6684
rect 12989 6681 13001 6684
rect 13035 6681 13047 6715
rect 12989 6675 13047 6681
rect 13081 6715 13139 6721
rect 13081 6681 13093 6715
rect 13127 6712 13139 6715
rect 13170 6712 13176 6724
rect 13127 6684 13176 6712
rect 13127 6681 13139 6684
rect 13081 6675 13139 6681
rect 13170 6672 13176 6684
rect 13228 6672 13234 6724
rect 17034 6712 17040 6724
rect 15948 6684 17040 6712
rect 5350 6644 5356 6656
rect 5092 6616 5356 6644
rect 4672 6604 4678 6616
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5626 6604 5632 6656
rect 5684 6604 5690 6656
rect 5718 6604 5724 6656
rect 5776 6604 5782 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 5997 6647 6055 6653
rect 5997 6644 6009 6647
rect 5868 6616 6009 6644
rect 5868 6604 5874 6616
rect 5997 6613 6009 6616
rect 6043 6613 6055 6647
rect 5997 6607 6055 6613
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 8444 6616 9045 6644
rect 8444 6604 8450 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 9766 6644 9772 6656
rect 9456 6616 9772 6644
rect 9456 6604 9462 6616
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 12158 6604 12164 6656
rect 12216 6604 12222 6656
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 15948 6653 15976 6684
rect 17034 6672 17040 6684
rect 17092 6672 17098 6724
rect 18969 6715 19027 6721
rect 18969 6681 18981 6715
rect 19015 6712 19027 6715
rect 19058 6712 19064 6724
rect 19015 6684 19064 6712
rect 19015 6681 19027 6684
rect 18969 6675 19027 6681
rect 19058 6672 19064 6684
rect 19116 6672 19122 6724
rect 19426 6672 19432 6724
rect 19484 6712 19490 6724
rect 19582 6715 19640 6721
rect 19582 6712 19594 6715
rect 19484 6684 19594 6712
rect 19484 6672 19490 6684
rect 19582 6681 19594 6684
rect 19628 6681 19640 6715
rect 20975 6715 21033 6721
rect 20975 6712 20987 6715
rect 19582 6675 19640 6681
rect 19720 6684 20987 6712
rect 12511 6647 12569 6653
rect 12511 6644 12523 6647
rect 12308 6616 12523 6644
rect 12308 6604 12314 6616
rect 12511 6613 12523 6616
rect 12557 6613 12569 6647
rect 12511 6607 12569 6613
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6613 15991 6647
rect 15933 6607 15991 6613
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17497 6647 17555 6653
rect 17497 6644 17509 6647
rect 17000 6616 17509 6644
rect 17000 6604 17006 6616
rect 17497 6613 17509 6616
rect 17543 6613 17555 6647
rect 17497 6607 17555 6613
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 19720 6644 19748 6684
rect 20975 6681 20987 6684
rect 21021 6681 21033 6715
rect 20975 6675 21033 6681
rect 21082 6672 21088 6724
rect 21140 6712 21146 6724
rect 21269 6715 21327 6721
rect 21269 6712 21281 6715
rect 21140 6684 21281 6712
rect 21140 6672 21146 6684
rect 21269 6681 21281 6684
rect 21315 6681 21327 6715
rect 21269 6675 21327 6681
rect 19208 6616 19748 6644
rect 19208 6604 19214 6616
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 21453 6647 21511 6653
rect 21453 6644 21465 6647
rect 20772 6616 21465 6644
rect 20772 6604 20778 6616
rect 21453 6613 21465 6616
rect 21499 6613 21511 6647
rect 21453 6607 21511 6613
rect 1104 6554 21988 6576
rect 1104 6502 4220 6554
rect 4272 6502 4284 6554
rect 4336 6502 4348 6554
rect 4400 6502 4412 6554
rect 4464 6502 4476 6554
rect 4528 6502 9441 6554
rect 9493 6502 9505 6554
rect 9557 6502 9569 6554
rect 9621 6502 9633 6554
rect 9685 6502 9697 6554
rect 9749 6502 14662 6554
rect 14714 6502 14726 6554
rect 14778 6502 14790 6554
rect 14842 6502 14854 6554
rect 14906 6502 14918 6554
rect 14970 6502 19883 6554
rect 19935 6502 19947 6554
rect 19999 6502 20011 6554
rect 20063 6502 20075 6554
rect 20127 6502 20139 6554
rect 20191 6502 21988 6554
rect 1104 6480 21988 6502
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 2774 6440 2780 6452
rect 2271 6412 2780 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 2774 6400 2780 6412
rect 2832 6440 2838 6452
rect 3234 6440 3240 6452
rect 2832 6412 3240 6440
rect 2832 6400 2838 6412
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4614 6440 4620 6452
rect 4203 6412 4620 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 5350 6440 5356 6452
rect 4816 6412 5356 6440
rect 2041 6375 2099 6381
rect 2041 6341 2053 6375
rect 2087 6372 2099 6375
rect 2087 6344 2636 6372
rect 2087 6341 2099 6344
rect 2041 6335 2099 6341
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 2314 6196 2320 6248
rect 2372 6196 2378 6248
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 2516 6168 2544 6267
rect 1811 6140 2544 6168
rect 2608 6168 2636 6344
rect 2884 6344 4752 6372
rect 2884 6316 2912 6344
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 2866 6304 2872 6316
rect 2823 6276 2872 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 3044 6307 3102 6313
rect 3044 6273 3056 6307
rect 3090 6304 3102 6307
rect 3418 6304 3424 6316
rect 3090 6276 3424 6304
rect 3090 6273 3102 6276
rect 3044 6267 3102 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 4724 6313 4752 6344
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 4816 6236 4844 6412
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 6089 6443 6147 6449
rect 6089 6409 6101 6443
rect 6135 6440 6147 6443
rect 6546 6440 6552 6452
rect 6135 6412 6552 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 7745 6443 7803 6449
rect 7745 6440 7757 6443
rect 7064 6412 7757 6440
rect 7064 6400 7070 6412
rect 7745 6409 7757 6412
rect 7791 6409 7803 6443
rect 7745 6403 7803 6409
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 9272 6412 9413 6440
rect 9272 6400 9278 6412
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 9401 6403 9459 6409
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9916 6412 10057 6440
rect 9916 6400 9922 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 12250 6440 12256 6452
rect 10045 6403 10103 6409
rect 11532 6412 12256 6440
rect 8294 6381 8300 6384
rect 8288 6372 8300 6381
rect 6380 6344 8064 6372
rect 8255 6344 8300 6372
rect 4976 6307 5034 6313
rect 4976 6273 4988 6307
rect 5022 6304 5034 6307
rect 5350 6304 5356 6316
rect 5022 6276 5356 6304
rect 5022 6273 5034 6276
rect 4976 6267 5034 6273
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 6380 6313 6408 6344
rect 8036 6316 8064 6344
rect 8288 6335 8300 6344
rect 8294 6332 8300 6335
rect 8352 6332 8358 6384
rect 10226 6372 10232 6384
rect 9140 6344 10232 6372
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5500 6276 6377 6304
rect 5500 6264 5506 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6621 6307 6679 6313
rect 6621 6304 6633 6307
rect 6512 6276 6633 6304
rect 6512 6264 6518 6276
rect 6621 6273 6633 6276
rect 6667 6273 6679 6307
rect 6621 6267 6679 6273
rect 8018 6264 8024 6316
rect 8076 6264 8082 6316
rect 9140 6304 9168 6344
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 10502 6332 10508 6384
rect 10560 6332 10566 6384
rect 10597 6375 10655 6381
rect 10597 6341 10609 6375
rect 10643 6372 10655 6375
rect 11238 6372 11244 6384
rect 10643 6344 11244 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 11238 6332 11244 6344
rect 11296 6332 11302 6384
rect 8128 6276 9168 6304
rect 4396 6208 4844 6236
rect 4396 6196 4402 6208
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 8128 6236 8156 6276
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9272 6276 9597 6304
rect 9272 6264 9278 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10042 6304 10048 6316
rect 9907 6276 10048 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 7616 6208 8156 6236
rect 9769 6239 9827 6245
rect 7616 6196 7622 6208
rect 9769 6205 9781 6239
rect 9815 6236 9827 6239
rect 10134 6236 10140 6248
rect 9815 6208 10140 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10520 6236 10548 6332
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 10962 6304 10968 6316
rect 10827 6276 10968 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11532 6313 11560 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 12952 6412 13185 6440
rect 12952 6400 12958 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 18598 6440 18604 6452
rect 13173 6403 13231 6409
rect 17236 6412 18604 6440
rect 12060 6375 12118 6381
rect 11624 6344 12020 6372
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 11624 6236 11652 6344
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6304 11851 6307
rect 11882 6304 11888 6316
rect 11839 6276 11888 6304
rect 11839 6273 11851 6276
rect 11793 6267 11851 6273
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 11992 6304 12020 6344
rect 12060 6341 12072 6375
rect 12106 6372 12118 6375
rect 12158 6372 12164 6384
rect 12106 6344 12164 6372
rect 12106 6341 12118 6344
rect 12060 6335 12118 6341
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 13446 6332 13452 6384
rect 13504 6332 13510 6384
rect 15105 6375 15163 6381
rect 15105 6341 15117 6375
rect 15151 6372 15163 6375
rect 15470 6372 15476 6384
rect 15151 6344 15476 6372
rect 15151 6341 15163 6344
rect 15105 6335 15163 6341
rect 15470 6332 15476 6344
rect 15528 6332 15534 6384
rect 12618 6304 12624 6316
rect 11992 6276 12624 6304
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 15562 6264 15568 6316
rect 15620 6264 15626 6316
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17236 6304 17264 6412
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 19337 6443 19395 6449
rect 19337 6409 19349 6443
rect 19383 6409 19395 6443
rect 19337 6403 19395 6409
rect 17954 6372 17960 6384
rect 17328 6344 17960 6372
rect 17328 6313 17356 6344
rect 17954 6332 17960 6344
rect 18012 6372 18018 6384
rect 19058 6372 19064 6384
rect 18012 6344 19064 6372
rect 18012 6332 18018 6344
rect 19058 6332 19064 6344
rect 19116 6332 19122 6384
rect 19352 6372 19380 6403
rect 19426 6400 19432 6452
rect 19484 6400 19490 6452
rect 19950 6375 20008 6381
rect 19950 6372 19962 6375
rect 19352 6344 19962 6372
rect 19950 6341 19962 6344
rect 19996 6341 20008 6375
rect 19950 6335 20008 6341
rect 17083 6276 17264 6304
rect 17313 6307 17371 6313
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17313 6273 17325 6307
rect 17359 6273 17371 6307
rect 17569 6307 17627 6313
rect 17569 6304 17581 6307
rect 17313 6267 17371 6273
rect 17420 6276 17581 6304
rect 10520 6208 11652 6236
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 14185 6239 14243 6245
rect 14185 6236 14197 6239
rect 13872 6208 14197 6236
rect 13872 6196 13878 6208
rect 14185 6205 14197 6208
rect 14231 6236 14243 6239
rect 14550 6236 14556 6248
rect 14231 6208 14556 6236
rect 14231 6205 14243 6208
rect 14185 6199 14243 6205
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 15102 6196 15108 6248
rect 15160 6196 15166 6248
rect 15197 6239 15255 6245
rect 15197 6205 15209 6239
rect 15243 6236 15255 6239
rect 15286 6236 15292 6248
rect 15243 6208 15292 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 15286 6196 15292 6208
rect 15344 6236 15350 6248
rect 16022 6236 16028 6248
rect 15344 6208 16028 6236
rect 15344 6196 15350 6208
rect 16022 6196 16028 6208
rect 16080 6196 16086 6248
rect 17126 6196 17132 6248
rect 17184 6236 17190 6248
rect 17420 6236 17448 6276
rect 17569 6273 17581 6276
rect 17615 6273 17627 6307
rect 17569 6267 17627 6273
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6304 18935 6307
rect 18923 6276 19012 6304
rect 18923 6273 18935 6276
rect 18877 6267 18935 6273
rect 17184 6208 17448 6236
rect 17184 6196 17190 6208
rect 18984 6168 19012 6276
rect 19150 6264 19156 6316
rect 19208 6264 19214 6316
rect 19610 6264 19616 6316
rect 19668 6264 19674 6316
rect 19058 6196 19064 6248
rect 19116 6236 19122 6248
rect 19705 6239 19763 6245
rect 19705 6236 19717 6239
rect 19116 6208 19717 6236
rect 19116 6196 19122 6208
rect 19705 6205 19717 6208
rect 19751 6205 19763 6239
rect 19705 6199 19763 6205
rect 19610 6168 19616 6180
rect 2608 6140 2820 6168
rect 18984 6140 19616 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 2682 6060 2688 6112
rect 2740 6060 2746 6112
rect 2792 6100 2820 6140
rect 19610 6128 19616 6140
rect 19668 6128 19674 6180
rect 21082 6128 21088 6180
rect 21140 6128 21146 6180
rect 3142 6100 3148 6112
rect 2792 6072 3148 6100
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 4890 6100 4896 6112
rect 4764 6072 4896 6100
rect 4764 6060 4770 6072
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 4982 6060 4988 6112
rect 5040 6100 5046 6112
rect 9766 6100 9772 6112
rect 5040 6072 9772 6100
rect 5040 6060 5046 6072
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 11054 6060 11060 6112
rect 11112 6060 11118 6112
rect 11701 6103 11759 6109
rect 11701 6069 11713 6103
rect 11747 6100 11759 6103
rect 12158 6100 12164 6112
rect 11747 6072 12164 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14645 6103 14703 6109
rect 14645 6100 14657 6103
rect 13780 6072 14657 6100
rect 13780 6060 13786 6072
rect 14645 6069 14657 6072
rect 14691 6069 14703 6103
rect 14645 6063 14703 6069
rect 15378 6060 15384 6112
rect 15436 6060 15442 6112
rect 17221 6103 17279 6109
rect 17221 6069 17233 6103
rect 17267 6100 17279 6103
rect 17310 6100 17316 6112
rect 17267 6072 17316 6100
rect 17267 6069 17279 6072
rect 17221 6063 17279 6069
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 18690 6060 18696 6112
rect 18748 6060 18754 6112
rect 19061 6103 19119 6109
rect 19061 6069 19073 6103
rect 19107 6100 19119 6103
rect 19702 6100 19708 6112
rect 19107 6072 19708 6100
rect 19107 6069 19119 6072
rect 19061 6063 19119 6069
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 1104 6010 21988 6032
rect 1104 5958 3560 6010
rect 3612 5958 3624 6010
rect 3676 5958 3688 6010
rect 3740 5958 3752 6010
rect 3804 5958 3816 6010
rect 3868 5958 8781 6010
rect 8833 5958 8845 6010
rect 8897 5958 8909 6010
rect 8961 5958 8973 6010
rect 9025 5958 9037 6010
rect 9089 5958 14002 6010
rect 14054 5958 14066 6010
rect 14118 5958 14130 6010
rect 14182 5958 14194 6010
rect 14246 5958 14258 6010
rect 14310 5958 19223 6010
rect 19275 5958 19287 6010
rect 19339 5958 19351 6010
rect 19403 5958 19415 6010
rect 19467 5958 19479 6010
rect 19531 5958 21988 6010
rect 1104 5936 21988 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 2774 5896 2780 5908
rect 1627 5868 2780 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 4982 5856 4988 5908
rect 5040 5856 5046 5908
rect 5166 5856 5172 5908
rect 5224 5856 5230 5908
rect 5350 5856 5356 5908
rect 5408 5856 5414 5908
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 6273 5899 6331 5905
rect 6273 5896 6285 5899
rect 5684 5868 6285 5896
rect 5684 5856 5690 5868
rect 6273 5865 6285 5868
rect 6319 5865 6331 5899
rect 6273 5859 6331 5865
rect 7926 5856 7932 5908
rect 7984 5856 7990 5908
rect 8570 5896 8576 5908
rect 8036 5868 8576 5896
rect 4525 5831 4583 5837
rect 4525 5797 4537 5831
rect 4571 5797 4583 5831
rect 7558 5828 7564 5840
rect 4525 5791 4583 5797
rect 6012 5800 7564 5828
rect 2682 5652 2688 5704
rect 2740 5701 2746 5704
rect 2740 5692 2752 5701
rect 2740 5664 2785 5692
rect 2740 5655 2752 5664
rect 2740 5652 2746 5655
rect 2866 5652 2872 5704
rect 2924 5692 2930 5704
rect 2961 5695 3019 5701
rect 2961 5692 2973 5695
rect 2924 5664 2973 5692
rect 2924 5652 2930 5664
rect 2961 5661 2973 5664
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 4338 5652 4344 5704
rect 4396 5701 4402 5704
rect 4396 5692 4404 5701
rect 4540 5692 4568 5791
rect 4798 5720 4804 5772
rect 4856 5720 4862 5772
rect 5810 5769 5816 5772
rect 5796 5763 5816 5769
rect 5796 5729 5808 5763
rect 5796 5723 5816 5729
rect 5810 5720 5816 5723
rect 5868 5720 5874 5772
rect 6012 5769 6040 5800
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 7653 5831 7711 5837
rect 7653 5797 7665 5831
rect 7699 5828 7711 5831
rect 8036 5828 8064 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13906 5896 13912 5908
rect 13311 5868 13912 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13906 5856 13912 5868
rect 13964 5896 13970 5908
rect 15102 5896 15108 5908
rect 13964 5868 15108 5896
rect 13964 5856 13970 5868
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15470 5856 15476 5908
rect 15528 5856 15534 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15620 5868 15761 5896
rect 15620 5856 15626 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 19337 5899 19395 5905
rect 19337 5896 19349 5899
rect 15749 5859 15807 5865
rect 16960 5868 19349 5896
rect 7699 5800 8064 5828
rect 8297 5831 8355 5837
rect 7699 5797 7711 5800
rect 7653 5791 7711 5797
rect 8297 5797 8309 5831
rect 8343 5828 8355 5831
rect 8386 5828 8392 5840
rect 8343 5800 8392 5828
rect 8343 5797 8355 5800
rect 8297 5791 8355 5797
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 11425 5831 11483 5837
rect 11425 5797 11437 5831
rect 11471 5828 11483 5831
rect 11882 5828 11888 5840
rect 11471 5800 11888 5828
rect 11471 5797 11483 5800
rect 11425 5791 11483 5797
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5729 6055 5763
rect 7190 5760 7196 5772
rect 5997 5723 6055 5729
rect 6380 5732 7196 5760
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4396 5664 4441 5692
rect 4540 5664 4721 5692
rect 4396 5655 4404 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5692 5043 5695
rect 5902 5692 5908 5704
rect 5031 5664 5908 5692
rect 5031 5661 5043 5664
rect 4985 5655 5043 5661
rect 4396 5652 4402 5655
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6086 5652 6092 5704
rect 6144 5652 6150 5704
rect 4157 5627 4215 5633
rect 4157 5593 4169 5627
rect 4203 5593 4215 5627
rect 4157 5587 4215 5593
rect 4249 5627 4307 5633
rect 4249 5593 4261 5627
rect 4295 5624 4307 5627
rect 4614 5624 4620 5636
rect 4295 5596 4620 5624
rect 4295 5593 4307 5596
rect 4249 5587 4307 5593
rect 4172 5556 4200 5587
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 5537 5627 5595 5633
rect 5537 5593 5549 5627
rect 5583 5624 5595 5627
rect 6380 5624 6408 5732
rect 7190 5720 7196 5732
rect 7248 5760 7254 5772
rect 7248 5732 7604 5760
rect 7248 5720 7254 5732
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 6546 5692 6552 5704
rect 6503 5664 6552 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 7064 5664 7481 5692
rect 7064 5652 7070 5664
rect 7469 5661 7481 5664
rect 7515 5661 7527 5695
rect 7576 5692 7604 5732
rect 8018 5720 8024 5772
rect 8076 5760 8082 5772
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8076 5732 9045 5760
rect 8076 5720 8082 5732
rect 9033 5729 9045 5732
rect 9079 5760 9091 5763
rect 9858 5760 9864 5772
rect 9079 5732 9864 5760
rect 9079 5729 9091 5732
rect 9033 5723 9091 5729
rect 9858 5720 9864 5732
rect 9916 5760 9922 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9916 5732 10057 5760
rect 9916 5720 9922 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 15488 5760 15516 5856
rect 16301 5763 16359 5769
rect 15488 5732 16252 5760
rect 10045 5723 10103 5729
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7576 5664 8125 5692
rect 7469 5655 7527 5661
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8294 5692 8300 5704
rect 8251 5664 8300 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 8478 5692 8484 5704
rect 8435 5664 8484 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11112 5664 11805 5692
rect 11112 5652 11118 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 11974 5692 11980 5704
rect 11931 5664 11980 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12158 5701 12164 5704
rect 12152 5692 12164 5701
rect 12119 5664 12164 5692
rect 12152 5655 12164 5664
rect 12158 5652 12164 5655
rect 12216 5652 12222 5704
rect 13722 5652 13728 5704
rect 13780 5652 13786 5704
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13872 5664 14105 5692
rect 13872 5652 13878 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 5583 5596 6408 5624
rect 6733 5627 6791 5633
rect 5583 5593 5595 5596
rect 5537 5587 5595 5593
rect 6733 5593 6745 5627
rect 6779 5624 6791 5627
rect 7193 5627 7251 5633
rect 7193 5624 7205 5627
rect 6779 5596 7205 5624
rect 6779 5593 6791 5596
rect 6733 5587 6791 5593
rect 7193 5593 7205 5596
rect 7239 5624 7251 5627
rect 7374 5624 7380 5636
rect 7239 5596 7380 5624
rect 7239 5593 7251 5596
rect 7193 5587 7251 5593
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 9861 5627 9919 5633
rect 9861 5593 9873 5627
rect 9907 5624 9919 5627
rect 9950 5624 9956 5636
rect 9907 5596 9956 5624
rect 9907 5593 9919 5596
rect 9861 5587 9919 5593
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10290 5627 10348 5633
rect 10290 5624 10302 5627
rect 10100 5596 10302 5624
rect 10100 5584 10106 5596
rect 10290 5593 10302 5596
rect 10336 5593 10348 5627
rect 14338 5627 14396 5633
rect 14338 5624 14350 5627
rect 10290 5587 10348 5593
rect 13924 5596 14350 5624
rect 4706 5556 4712 5568
rect 4172 5528 4712 5556
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 6641 5559 6699 5565
rect 6641 5556 6653 5559
rect 5951 5528 6653 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 6641 5525 6653 5528
rect 6687 5556 6699 5559
rect 7282 5556 7288 5568
rect 6687 5528 7288 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 11606 5516 11612 5568
rect 11664 5516 11670 5568
rect 13924 5565 13952 5596
rect 14338 5593 14350 5596
rect 14384 5593 14396 5627
rect 14338 5587 14396 5593
rect 16025 5627 16083 5633
rect 16025 5593 16037 5627
rect 16071 5624 16083 5627
rect 16114 5624 16120 5636
rect 16071 5596 16120 5624
rect 16071 5593 16083 5596
rect 16025 5587 16083 5593
rect 16114 5584 16120 5596
rect 16172 5584 16178 5636
rect 16224 5633 16252 5732
rect 16301 5729 16313 5763
rect 16347 5760 16359 5763
rect 16482 5760 16488 5772
rect 16347 5732 16488 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 16960 5701 16988 5868
rect 19337 5865 19349 5868
rect 19383 5865 19395 5899
rect 19337 5859 19395 5865
rect 17126 5788 17132 5840
rect 17184 5788 17190 5840
rect 18601 5831 18659 5837
rect 18601 5797 18613 5831
rect 18647 5828 18659 5831
rect 18782 5828 18788 5840
rect 18647 5800 18788 5828
rect 18647 5797 18659 5800
rect 18601 5791 18659 5797
rect 18782 5788 18788 5800
rect 18840 5788 18846 5840
rect 19518 5788 19524 5840
rect 19576 5828 19582 5840
rect 20165 5831 20223 5837
rect 20165 5828 20177 5831
rect 19576 5800 20177 5828
rect 19576 5788 19582 5800
rect 20165 5797 20177 5800
rect 20211 5797 20223 5831
rect 20165 5791 20223 5797
rect 21542 5788 21548 5840
rect 21600 5788 21606 5840
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 18748 5732 19809 5760
rect 18748 5720 18754 5732
rect 19797 5729 19809 5732
rect 19843 5760 19855 5763
rect 20346 5760 20352 5772
rect 19843 5732 20352 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 20346 5720 20352 5732
rect 20404 5720 20410 5772
rect 20717 5763 20775 5769
rect 20717 5729 20729 5763
rect 20763 5760 20775 5763
rect 20806 5760 20812 5772
rect 20763 5732 20812 5760
rect 20763 5729 20775 5732
rect 20717 5723 20775 5729
rect 20806 5720 20812 5732
rect 20864 5720 20870 5772
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5661 17003 5695
rect 16945 5655 17003 5661
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5692 17279 5695
rect 17954 5692 17960 5704
rect 17267 5664 17960 5692
rect 17267 5661 17279 5664
rect 17221 5655 17279 5661
rect 17954 5652 17960 5664
rect 18012 5652 18018 5704
rect 20438 5652 20444 5704
rect 20496 5652 20502 5704
rect 16209 5627 16267 5633
rect 16209 5593 16221 5627
rect 16255 5593 16267 5627
rect 16209 5587 16267 5593
rect 17310 5584 17316 5636
rect 17368 5624 17374 5636
rect 17466 5627 17524 5633
rect 17466 5624 17478 5627
rect 17368 5596 17478 5624
rect 17368 5584 17374 5596
rect 17466 5593 17478 5596
rect 17512 5593 17524 5627
rect 17466 5587 17524 5593
rect 18782 5584 18788 5636
rect 18840 5624 18846 5636
rect 19797 5627 19855 5633
rect 19797 5624 19809 5627
rect 18840 5596 19809 5624
rect 18840 5584 18846 5596
rect 19797 5593 19809 5596
rect 19843 5593 19855 5627
rect 19797 5587 19855 5593
rect 19889 5627 19947 5633
rect 19889 5593 19901 5627
rect 19935 5624 19947 5627
rect 20990 5624 20996 5636
rect 19935 5596 20996 5624
rect 19935 5593 19947 5596
rect 19889 5587 19947 5593
rect 20990 5584 20996 5596
rect 21048 5584 21054 5636
rect 21269 5627 21327 5633
rect 21269 5593 21281 5627
rect 21315 5624 21327 5627
rect 21450 5624 21456 5636
rect 21315 5596 21456 5624
rect 21315 5593 21327 5596
rect 21269 5587 21327 5593
rect 21450 5584 21456 5596
rect 21508 5584 21514 5636
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5525 13967 5559
rect 13909 5519 13967 5525
rect 20625 5559 20683 5565
rect 20625 5525 20637 5559
rect 20671 5556 20683 5559
rect 21085 5559 21143 5565
rect 21085 5556 21097 5559
rect 20671 5528 21097 5556
rect 20671 5525 20683 5528
rect 20625 5519 20683 5525
rect 21085 5525 21097 5528
rect 21131 5556 21143 5559
rect 21174 5556 21180 5568
rect 21131 5528 21180 5556
rect 21131 5525 21143 5528
rect 21085 5519 21143 5525
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 1104 5466 21988 5488
rect 1104 5414 4220 5466
rect 4272 5414 4284 5466
rect 4336 5414 4348 5466
rect 4400 5414 4412 5466
rect 4464 5414 4476 5466
rect 4528 5414 9441 5466
rect 9493 5414 9505 5466
rect 9557 5414 9569 5466
rect 9621 5414 9633 5466
rect 9685 5414 9697 5466
rect 9749 5414 14662 5466
rect 14714 5414 14726 5466
rect 14778 5414 14790 5466
rect 14842 5414 14854 5466
rect 14906 5414 14918 5466
rect 14970 5414 19883 5466
rect 19935 5414 19947 5466
rect 19999 5414 20011 5466
rect 20063 5414 20075 5466
rect 20127 5414 20139 5466
rect 20191 5414 21988 5466
rect 1104 5392 21988 5414
rect 3142 5312 3148 5364
rect 3200 5352 3206 5364
rect 3329 5355 3387 5361
rect 3329 5352 3341 5355
rect 3200 5324 3341 5352
rect 3200 5312 3206 5324
rect 3329 5321 3341 5324
rect 3375 5352 3387 5355
rect 4614 5352 4620 5364
rect 3375 5324 4620 5352
rect 3375 5321 3387 5324
rect 3329 5315 3387 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 8202 5312 8208 5364
rect 8260 5352 8266 5364
rect 9769 5355 9827 5361
rect 8260 5324 8616 5352
rect 8260 5312 8266 5324
rect 2866 5284 2872 5296
rect 1964 5256 2872 5284
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1854 5216 1860 5228
rect 1719 5188 1860 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 1964 5225 1992 5256
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 3234 5244 3240 5296
rect 3292 5284 3298 5296
rect 4341 5287 4399 5293
rect 4341 5284 4353 5287
rect 3292 5256 4353 5284
rect 3292 5244 3298 5256
rect 4341 5253 4353 5256
rect 4387 5253 4399 5287
rect 4341 5247 4399 5253
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 5592 5256 6592 5284
rect 5592 5244 5598 5256
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 2205 5219 2263 5225
rect 2205 5216 2217 5219
rect 1949 5179 2007 5185
rect 2056 5188 2217 5216
rect 2056 5148 2084 5188
rect 2205 5185 2217 5188
rect 2251 5185 2263 5219
rect 2205 5179 2263 5185
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 1872 5120 2084 5148
rect 3988 5148 4016 5179
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4249 5219 4307 5225
rect 4120 5188 4165 5216
rect 4120 5176 4126 5188
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 4479 5219 4537 5225
rect 4479 5185 4491 5219
rect 4525 5216 4537 5219
rect 4706 5216 4712 5228
rect 4525 5188 4712 5216
rect 4525 5185 4537 5188
rect 4479 5179 4537 5185
rect 4264 5148 4292 5179
rect 4706 5176 4712 5188
rect 4764 5216 4770 5228
rect 5813 5219 5871 5225
rect 4764 5188 5580 5216
rect 4764 5176 4770 5188
rect 5074 5148 5080 5160
rect 3988 5120 4077 5148
rect 4264 5120 5080 5148
rect 1872 5089 1900 5120
rect 1857 5083 1915 5089
rect 1857 5049 1869 5083
rect 1903 5049 1915 5083
rect 4049 5080 4077 5120
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5552 5148 5580 5188
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 6564 5216 6592 5256
rect 6730 5244 6736 5296
rect 6788 5284 6794 5296
rect 6917 5287 6975 5293
rect 6917 5284 6929 5287
rect 6788 5256 6929 5284
rect 6788 5244 6794 5256
rect 6917 5253 6929 5256
rect 6963 5253 6975 5287
rect 6917 5247 6975 5253
rect 7282 5244 7288 5296
rect 7340 5284 7346 5296
rect 7340 5256 8064 5284
rect 7340 5244 7346 5256
rect 5859 5188 6500 5216
rect 6564 5188 6868 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 5552 5120 6215 5148
rect 4522 5080 4528 5092
rect 4049 5052 4528 5080
rect 1857 5043 1915 5049
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 4617 5083 4675 5089
rect 4617 5049 4629 5083
rect 4663 5080 4675 5083
rect 6086 5080 6092 5092
rect 4663 5052 6092 5080
rect 4663 5049 4675 5052
rect 4617 5043 4675 5049
rect 6086 5040 6092 5052
rect 6144 5040 6150 5092
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 6187 5012 6215 5120
rect 6472 5089 6500 5188
rect 6840 5157 6868 5188
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 8036 5225 8064 5256
rect 8386 5244 8392 5296
rect 8444 5284 8450 5296
rect 8481 5287 8539 5293
rect 8481 5284 8493 5287
rect 8444 5256 8493 5284
rect 8444 5244 8450 5256
rect 8481 5253 8493 5256
rect 8527 5253 8539 5287
rect 8481 5247 8539 5253
rect 8588 5225 8616 5324
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10042 5352 10048 5364
rect 9815 5324 10048 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 11238 5312 11244 5364
rect 11296 5352 11302 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11296 5324 12081 5352
rect 11296 5312 11302 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 13170 5352 13176 5364
rect 12069 5315 12127 5321
rect 13004 5324 13176 5352
rect 8849 5287 8907 5293
rect 8849 5253 8861 5287
rect 8895 5284 8907 5287
rect 9306 5284 9312 5296
rect 8895 5256 9312 5284
rect 8895 5253 8907 5256
rect 8849 5247 8907 5253
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 10128 5287 10186 5293
rect 9600 5256 9996 5284
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7524 5188 7849 5216
rect 7524 5176 7530 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8239 5219 8297 5225
rect 8239 5185 8251 5219
rect 8285 5185 8297 5219
rect 8239 5179 8297 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7006 5108 7012 5160
rect 7064 5108 7070 5160
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 8128 5148 8156 5179
rect 7800 5120 8156 5148
rect 8254 5148 8282 5179
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8720 5188 8769 5216
rect 8720 5176 8726 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 8993 5219 9051 5225
rect 8993 5185 9005 5219
rect 9039 5216 9051 5219
rect 9122 5216 9128 5228
rect 9039 5188 9128 5216
rect 9039 5185 9051 5188
rect 8993 5179 9051 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9600 5225 9628 5256
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 9858 5176 9864 5228
rect 9916 5176 9922 5228
rect 9968 5216 9996 5256
rect 10128 5253 10140 5287
rect 10174 5284 10186 5287
rect 11606 5284 11612 5296
rect 10174 5256 11612 5284
rect 10174 5253 10186 5256
rect 10128 5247 10186 5253
rect 11606 5244 11612 5256
rect 11664 5244 11670 5296
rect 11790 5244 11796 5296
rect 11848 5284 11854 5296
rect 12897 5287 12955 5293
rect 12897 5284 12909 5287
rect 11848 5256 12909 5284
rect 11848 5244 11854 5256
rect 12897 5253 12909 5256
rect 12943 5253 12955 5287
rect 12897 5247 12955 5253
rect 9968 5188 11652 5216
rect 8254 5120 8331 5148
rect 7800 5108 7806 5120
rect 6457 5083 6515 5089
rect 6457 5049 6469 5083
rect 6503 5049 6515 5083
rect 8303 5080 8331 5120
rect 11624 5089 11652 5188
rect 11882 5176 11888 5228
rect 11940 5176 11946 5228
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 13004 5216 13032 5324
rect 13170 5312 13176 5324
rect 13228 5352 13234 5364
rect 14366 5352 14372 5364
rect 13228 5324 14372 5352
rect 13228 5312 13234 5324
rect 13081 5287 13139 5293
rect 13081 5253 13093 5287
rect 13127 5284 13139 5287
rect 13446 5284 13452 5296
rect 13127 5256 13452 5284
rect 13127 5253 13139 5256
rect 13081 5247 13139 5253
rect 13446 5244 13452 5256
rect 13504 5284 13510 5296
rect 14016 5293 14044 5324
rect 14366 5312 14372 5324
rect 14424 5352 14430 5364
rect 16482 5352 16488 5364
rect 14424 5324 16488 5352
rect 14424 5312 14430 5324
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5321 19763 5355
rect 19705 5315 19763 5321
rect 13909 5287 13967 5293
rect 13909 5284 13921 5287
rect 13504 5256 13921 5284
rect 13504 5244 13510 5256
rect 13909 5253 13921 5256
rect 13955 5253 13967 5287
rect 13909 5247 13967 5253
rect 14001 5287 14059 5293
rect 14001 5253 14013 5287
rect 14047 5253 14059 5287
rect 14001 5247 14059 5253
rect 14452 5287 14510 5293
rect 14452 5253 14464 5287
rect 14498 5284 14510 5287
rect 15378 5284 15384 5296
rect 14498 5256 15384 5284
rect 14498 5253 14510 5256
rect 14452 5247 14510 5253
rect 15378 5244 15384 5256
rect 15436 5244 15442 5296
rect 17954 5284 17960 5296
rect 16684 5256 17960 5284
rect 12207 5188 13032 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 16684 5225 16712 5256
rect 17954 5244 17960 5256
rect 18012 5244 18018 5296
rect 18046 5244 18052 5296
rect 18104 5284 18110 5296
rect 18601 5287 18659 5293
rect 18601 5284 18613 5287
rect 18104 5256 18613 5284
rect 18104 5244 18110 5256
rect 18601 5253 18613 5256
rect 18647 5253 18659 5287
rect 18601 5247 18659 5253
rect 18785 5287 18843 5293
rect 18785 5253 18797 5287
rect 18831 5253 18843 5287
rect 18785 5247 18843 5253
rect 18877 5287 18935 5293
rect 18877 5253 18889 5287
rect 18923 5284 18935 5287
rect 18966 5284 18972 5296
rect 18923 5256 18972 5284
rect 18923 5253 18935 5256
rect 18877 5247 18935 5253
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16669 5219 16727 5225
rect 16347 5188 16436 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 13173 5151 13231 5157
rect 13173 5148 13185 5151
rect 12676 5120 13185 5148
rect 12676 5108 12682 5120
rect 13173 5117 13185 5120
rect 13219 5117 13231 5151
rect 13173 5111 13231 5117
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5117 14243 5151
rect 14185 5111 14243 5117
rect 9125 5083 9183 5089
rect 9125 5080 9137 5083
rect 8303 5052 9137 5080
rect 6457 5043 6515 5049
rect 9125 5049 9137 5052
rect 9171 5049 9183 5083
rect 9125 5043 9183 5049
rect 11609 5083 11667 5089
rect 11609 5049 11621 5083
rect 11655 5049 11667 5083
rect 11609 5043 11667 5049
rect 11698 5040 11704 5092
rect 11756 5080 11762 5092
rect 13449 5083 13507 5089
rect 13449 5080 13461 5083
rect 11756 5052 13461 5080
rect 11756 5040 11762 5052
rect 13449 5049 13461 5052
rect 13495 5049 13507 5083
rect 14200 5080 14228 5111
rect 13449 5043 13507 5049
rect 13832 5052 14228 5080
rect 13832 5024 13860 5052
rect 6822 5012 6828 5024
rect 6187 4984 6828 5012
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 11848 4984 12633 5012
rect 11848 4972 11854 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 13814 4972 13820 5024
rect 13872 4972 13878 5024
rect 15565 5015 15623 5021
rect 15565 4981 15577 5015
rect 15611 5012 15623 5015
rect 16114 5012 16120 5024
rect 15611 4984 16120 5012
rect 15611 4981 15623 4984
rect 15565 4975 15623 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 16408 5012 16436 5188
rect 16669 5185 16681 5219
rect 16715 5185 16727 5219
rect 16925 5219 16983 5225
rect 16925 5216 16937 5219
rect 16669 5179 16727 5185
rect 16776 5188 16937 5216
rect 16776 5148 16804 5188
rect 16925 5185 16937 5188
rect 16971 5185 16983 5219
rect 16925 5179 16983 5185
rect 16500 5120 16804 5148
rect 16500 5089 16528 5120
rect 16485 5083 16543 5089
rect 16485 5049 16497 5083
rect 16531 5049 16543 5083
rect 18325 5083 18383 5089
rect 18325 5080 18337 5083
rect 16485 5043 16543 5049
rect 17604 5052 18337 5080
rect 17604 5012 17632 5052
rect 18325 5049 18337 5052
rect 18371 5049 18383 5083
rect 18325 5043 18383 5049
rect 16408 4984 17632 5012
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 18800 5012 18828 5247
rect 18966 5244 18972 5256
rect 19024 5244 19030 5296
rect 19720 5284 19748 5315
rect 21174 5312 21180 5364
rect 21232 5312 21238 5364
rect 20042 5287 20100 5293
rect 20042 5284 20054 5287
rect 19720 5256 20054 5284
rect 20042 5253 20054 5256
rect 20088 5253 20100 5287
rect 20042 5247 20100 5253
rect 19518 5176 19524 5228
rect 19576 5176 19582 5228
rect 21542 5176 21548 5228
rect 21600 5176 21606 5228
rect 19058 5108 19064 5160
rect 19116 5148 19122 5160
rect 19797 5151 19855 5157
rect 19797 5148 19809 5151
rect 19116 5120 19809 5148
rect 19116 5108 19122 5120
rect 19797 5117 19809 5120
rect 19843 5117 19855 5151
rect 19797 5111 19855 5117
rect 18104 4984 18828 5012
rect 18104 4972 18110 4984
rect 21358 4972 21364 5024
rect 21416 4972 21422 5024
rect 1104 4922 21988 4944
rect 1104 4870 3560 4922
rect 3612 4870 3624 4922
rect 3676 4870 3688 4922
rect 3740 4870 3752 4922
rect 3804 4870 3816 4922
rect 3868 4870 8781 4922
rect 8833 4870 8845 4922
rect 8897 4870 8909 4922
rect 8961 4870 8973 4922
rect 9025 4870 9037 4922
rect 9089 4870 14002 4922
rect 14054 4870 14066 4922
rect 14118 4870 14130 4922
rect 14182 4870 14194 4922
rect 14246 4870 14258 4922
rect 14310 4870 19223 4922
rect 19275 4870 19287 4922
rect 19339 4870 19351 4922
rect 19403 4870 19415 4922
rect 19467 4870 19479 4922
rect 19531 4870 21988 4922
rect 1104 4848 21988 4870
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 1872 4780 3893 4808
rect 1872 4613 1900 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 3881 4771 3939 4777
rect 4709 4811 4767 4817
rect 4709 4777 4721 4811
rect 4755 4808 4767 4811
rect 4798 4808 4804 4820
rect 4755 4780 4804 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 6730 4768 6736 4820
rect 6788 4768 6794 4820
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4808 7711 4811
rect 9214 4808 9220 4820
rect 7699 4780 9220 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 13446 4768 13452 4820
rect 13504 4768 13510 4820
rect 21542 4768 21548 4820
rect 21600 4768 21606 4820
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4604 2191 4607
rect 2866 4604 2872 4616
rect 2179 4576 2872 4604
rect 2179 4573 2191 4576
rect 2133 4567 2191 4573
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3418 4564 3424 4616
rect 3476 4604 3482 4616
rect 4157 4607 4215 4613
rect 4157 4604 4169 4607
rect 3476 4576 4169 4604
rect 3476 4564 3482 4576
rect 4157 4573 4169 4576
rect 4203 4573 4215 4607
rect 4888 4607 4946 4613
rect 4888 4604 4900 4607
rect 4157 4567 4215 4573
rect 4361 4576 4900 4604
rect 2378 4539 2436 4545
rect 2378 4536 2390 4539
rect 2056 4508 2390 4536
rect 2056 4477 2084 4508
rect 2378 4505 2390 4508
rect 2424 4505 2436 4539
rect 2378 4499 2436 4505
rect 3786 4496 3792 4548
rect 3844 4536 3850 4548
rect 4361 4536 4389 4576
rect 4888 4573 4900 4576
rect 4934 4573 4946 4607
rect 4888 4567 4946 4573
rect 3844 4508 4389 4536
rect 4433 4539 4491 4545
rect 3844 4496 3850 4508
rect 4433 4505 4445 4539
rect 4479 4536 4491 4539
rect 4798 4536 4804 4548
rect 4479 4508 4804 4536
rect 4479 4505 4491 4508
rect 4433 4499 4491 4505
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 2041 4471 2099 4477
rect 2041 4437 2053 4471
rect 2087 4437 2099 4471
rect 2041 4431 2099 4437
rect 3513 4471 3571 4477
rect 3513 4437 3525 4471
rect 3559 4468 3571 4471
rect 4062 4468 4068 4480
rect 3559 4440 4068 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 4062 4428 4068 4440
rect 4120 4468 4126 4480
rect 4341 4471 4399 4477
rect 4341 4468 4353 4471
rect 4120 4440 4353 4468
rect 4120 4428 4126 4440
rect 4341 4437 4353 4440
rect 4387 4437 4399 4471
rect 4903 4468 4931 4567
rect 5074 4564 5080 4616
rect 5132 4564 5138 4616
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5442 4604 5448 4616
rect 5399 4576 5448 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5626 4613 5632 4616
rect 5620 4604 5632 4613
rect 5587 4576 5632 4604
rect 5620 4567 5632 4576
rect 5626 4564 5632 4567
rect 5684 4564 5690 4616
rect 6748 4604 6776 4768
rect 8113 4743 8171 4749
rect 8113 4709 8125 4743
rect 8159 4740 8171 4743
rect 8202 4740 8208 4752
rect 8159 4712 8208 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 16574 4740 16580 4752
rect 16316 4712 16580 4740
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 8478 4672 8484 4684
rect 6880 4644 8484 4672
rect 6880 4632 6886 4644
rect 7536 4613 7564 4644
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 8662 4672 8668 4684
rect 8619 4644 8668 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 6748 4576 7113 4604
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7521 4607 7579 4613
rect 7521 4573 7533 4607
rect 7567 4573 7579 4607
rect 7521 4567 7579 4573
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 9766 4604 9772 4616
rect 8987 4576 9772 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4604 11575 4607
rect 11698 4604 11704 4616
rect 11563 4576 11704 4604
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11790 4564 11796 4616
rect 11848 4564 11854 4616
rect 12066 4564 12072 4616
rect 12124 4564 12130 4616
rect 16316 4613 16344 4712
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4573 16359 4607
rect 16301 4567 16359 4573
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4604 16635 4607
rect 18690 4604 18696 4616
rect 16623 4576 18696 4604
rect 16623 4573 16635 4576
rect 16577 4567 16635 4573
rect 18690 4564 18696 4576
rect 18748 4604 18754 4616
rect 19058 4604 19064 4616
rect 18748 4576 19064 4604
rect 18748 4564 18754 4576
rect 19058 4564 19064 4576
rect 19116 4604 19122 4616
rect 20165 4607 20223 4613
rect 20165 4604 20177 4607
rect 19116 4576 20177 4604
rect 19116 4564 19122 4576
rect 20165 4573 20177 4576
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 20432 4607 20490 4613
rect 20432 4573 20444 4607
rect 20478 4604 20490 4607
rect 21358 4604 21364 4616
rect 20478 4576 21364 4604
rect 20478 4573 20490 4576
rect 20432 4567 20490 4573
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 4982 4496 4988 4548
rect 5040 4496 5046 4548
rect 5092 4536 5120 4564
rect 7282 4536 7288 4548
rect 5092 4508 7288 4536
rect 7282 4496 7288 4508
rect 7340 4496 7346 4548
rect 7377 4539 7435 4545
rect 7377 4505 7389 4539
rect 7423 4505 7435 4539
rect 7377 4499 7435 4505
rect 6822 4468 6828 4480
rect 4903 4440 6828 4468
rect 4341 4431 4399 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7392 4468 7420 4499
rect 8478 4496 8484 4548
rect 8536 4536 8542 4548
rect 8665 4539 8723 4545
rect 8665 4536 8677 4539
rect 8536 4508 8677 4536
rect 8536 4496 8542 4508
rect 8665 4505 8677 4508
rect 8711 4505 8723 4539
rect 8665 4499 8723 4505
rect 8754 4496 8760 4548
rect 8812 4536 8818 4548
rect 9186 4539 9244 4545
rect 9186 4536 9198 4539
rect 8812 4508 9198 4536
rect 8812 4496 8818 4508
rect 9186 4505 9198 4508
rect 9232 4505 9244 4539
rect 12314 4539 12372 4545
rect 12314 4536 12326 4539
rect 9186 4499 9244 4505
rect 11992 4508 12326 4536
rect 7156 4440 7420 4468
rect 8573 4471 8631 4477
rect 7156 4428 7162 4440
rect 8573 4437 8585 4471
rect 8619 4468 8631 4471
rect 9306 4468 9312 4480
rect 8619 4440 9312 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 9306 4428 9312 4440
rect 9364 4468 9370 4480
rect 10321 4471 10379 4477
rect 10321 4468 10333 4471
rect 9364 4440 10333 4468
rect 9364 4428 9370 4440
rect 10321 4437 10333 4440
rect 10367 4437 10379 4471
rect 10321 4431 10379 4437
rect 11698 4428 11704 4480
rect 11756 4428 11762 4480
rect 11992 4477 12020 4508
rect 12314 4505 12326 4508
rect 12360 4505 12372 4539
rect 16822 4539 16880 4545
rect 16822 4536 16834 4539
rect 12314 4499 12372 4505
rect 16500 4508 16834 4536
rect 16500 4477 16528 4508
rect 16822 4505 16834 4508
rect 16868 4505 16880 4539
rect 16822 4499 16880 4505
rect 11977 4471 12035 4477
rect 11977 4437 11989 4471
rect 12023 4437 12035 4471
rect 11977 4431 12035 4437
rect 16485 4471 16543 4477
rect 16485 4437 16497 4471
rect 16531 4437 16543 4471
rect 16485 4431 16543 4437
rect 17954 4428 17960 4480
rect 18012 4428 18018 4480
rect 1104 4378 21988 4400
rect 1104 4326 4220 4378
rect 4272 4326 4284 4378
rect 4336 4326 4348 4378
rect 4400 4326 4412 4378
rect 4464 4326 4476 4378
rect 4528 4326 9441 4378
rect 9493 4326 9505 4378
rect 9557 4326 9569 4378
rect 9621 4326 9633 4378
rect 9685 4326 9697 4378
rect 9749 4326 14662 4378
rect 14714 4326 14726 4378
rect 14778 4326 14790 4378
rect 14842 4326 14854 4378
rect 14906 4326 14918 4378
rect 14970 4326 19883 4378
rect 19935 4326 19947 4378
rect 19999 4326 20011 4378
rect 20063 4326 20075 4378
rect 20127 4326 20139 4378
rect 20191 4326 21988 4378
rect 1104 4304 21988 4326
rect 4525 4267 4583 4273
rect 4525 4233 4537 4267
rect 4571 4264 4583 4267
rect 5258 4264 5264 4276
rect 4571 4236 5264 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 5258 4224 5264 4236
rect 5316 4224 5322 4276
rect 8389 4267 8447 4273
rect 8389 4233 8401 4267
rect 8435 4264 8447 4267
rect 8754 4264 8760 4276
rect 8435 4236 8760 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 13449 4267 13507 4273
rect 13449 4233 13461 4267
rect 13495 4264 13507 4267
rect 13538 4264 13544 4276
rect 13495 4236 13544 4264
rect 13495 4233 13507 4236
rect 13449 4227 13507 4233
rect 13538 4224 13544 4236
rect 13596 4264 13602 4276
rect 13722 4264 13728 4276
rect 13596 4236 13728 4264
rect 13596 4224 13602 4236
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14366 4264 14372 4276
rect 13832 4236 14372 4264
rect 2225 4199 2283 4205
rect 2225 4165 2237 4199
rect 2271 4196 2283 4199
rect 2958 4196 2964 4208
rect 2271 4168 2964 4196
rect 2271 4165 2283 4168
rect 2225 4159 2283 4165
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 3053 4199 3111 4205
rect 3053 4165 3065 4199
rect 3099 4196 3111 4199
rect 3142 4196 3148 4208
rect 3099 4168 3148 4196
rect 3099 4165 3111 4168
rect 3053 4159 3111 4165
rect 3142 4156 3148 4168
rect 3200 4156 3206 4208
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 5353 4199 5411 4205
rect 5353 4196 5365 4199
rect 5132 4168 5365 4196
rect 5132 4156 5138 4168
rect 5353 4165 5365 4168
rect 5399 4165 5411 4199
rect 5353 4159 5411 4165
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 6972 4168 7236 4196
rect 6972 4156 6978 4168
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 1443 4100 1808 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1780 4001 1808 4100
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2832 4100 2881 4128
rect 2832 4088 2838 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 3936 4100 4353 4128
rect 3936 4088 3942 4100
rect 4341 4097 4353 4100
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4764 4100 5181 4128
rect 4764 4088 4770 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 5868 4100 6745 4128
rect 5868 4088 5874 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 7006 4088 7012 4140
rect 7064 4088 7070 4140
rect 7208 4137 7236 4168
rect 7282 4156 7288 4208
rect 7340 4196 7346 4208
rect 7377 4199 7435 4205
rect 7377 4196 7389 4199
rect 7340 4168 7389 4196
rect 7340 4156 7346 4168
rect 7377 4165 7389 4168
rect 7423 4196 7435 4199
rect 10410 4196 10416 4208
rect 7423 4168 10416 4196
rect 7423 4165 7435 4168
rect 7377 4159 7435 4165
rect 10410 4156 10416 4168
rect 10468 4156 10474 4208
rect 11146 4156 11152 4208
rect 11204 4156 11210 4208
rect 11698 4156 11704 4208
rect 11756 4196 11762 4208
rect 12314 4199 12372 4205
rect 12314 4196 12326 4199
rect 11756 4168 12326 4196
rect 11756 4156 11762 4168
rect 12314 4165 12326 4168
rect 12360 4165 12372 4199
rect 13832 4196 13860 4236
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 15286 4264 15292 4276
rect 14844 4236 15292 4264
rect 12314 4159 12372 4165
rect 12406 4168 13860 4196
rect 14016 4168 14688 4196
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7466 4088 7472 4140
rect 7524 4088 7530 4140
rect 7566 4131 7624 4137
rect 7566 4097 7578 4131
rect 7612 4097 7624 4131
rect 7566 4091 7624 4097
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 1765 3995 1823 4001
rect 1765 3961 1777 3995
rect 1811 3961 1823 3995
rect 2240 3992 2268 4023
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 3145 4063 3203 4069
rect 3145 4060 3157 4063
rect 2372 4032 3157 4060
rect 2372 4020 2378 4032
rect 3145 4029 3157 4032
rect 3191 4060 3203 4063
rect 4617 4063 4675 4069
rect 4617 4060 4629 4063
rect 3191 4032 4629 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 4617 4029 4629 4032
rect 4663 4029 4675 4063
rect 4617 4023 4675 4029
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 5626 4060 5632 4072
rect 5491 4032 5632 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 2958 3992 2964 4004
rect 2240 3964 2964 3992
rect 1765 3955 1823 3961
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 3786 3952 3792 4004
rect 3844 3992 3850 4004
rect 3970 3992 3976 4004
rect 3844 3964 3976 3992
rect 3844 3952 3850 3964
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4632 3992 4660 4023
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7581 4060 7609 4091
rect 7926 4088 7932 4140
rect 7984 4088 7990 4140
rect 8202 4088 8208 4140
rect 8260 4088 8266 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8570 4128 8576 4140
rect 8527 4100 8576 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 8901 4131 8959 4137
rect 8901 4097 8913 4131
rect 8947 4128 8959 4131
rect 9122 4128 9128 4140
rect 8947 4100 9128 4128
rect 8947 4097 8959 4100
rect 8901 4091 8959 4097
rect 8680 4060 8708 4091
rect 6880 4032 8708 4060
rect 8772 4060 8800 4091
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 11241 4131 11299 4137
rect 10551 4100 10732 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 9490 4060 9496 4072
rect 8772 4032 9496 4060
rect 6880 4020 6886 4032
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 10134 4020 10140 4072
rect 10192 4020 10198 4072
rect 4798 3992 4804 4004
rect 4632 3964 4804 3992
rect 4798 3952 4804 3964
rect 4856 3992 4862 4004
rect 7006 3992 7012 4004
rect 4856 3964 7012 3992
rect 4856 3952 4862 3964
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 7742 3952 7748 4004
rect 7800 3952 7806 4004
rect 9033 3995 9091 4001
rect 9033 3961 9045 3995
rect 9079 3992 9091 3995
rect 10152 3992 10180 4020
rect 10704 4001 10732 4100
rect 11241 4097 11253 4131
rect 11287 4128 11299 4131
rect 12406 4128 12434 4168
rect 14016 4128 14044 4168
rect 11287 4100 12434 4128
rect 13648 4100 14044 4128
rect 14093 4131 14151 4137
rect 11287 4097 11299 4100
rect 11241 4091 11299 4097
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11057 4063 11115 4069
rect 11057 4060 11069 4063
rect 11020 4032 11069 4060
rect 11020 4020 11026 4032
rect 11057 4029 11069 4032
rect 11103 4029 11115 4063
rect 11057 4023 11115 4029
rect 12066 4020 12072 4072
rect 12124 4020 12130 4072
rect 9079 3964 10180 3992
rect 10689 3995 10747 4001
rect 9079 3961 9091 3964
rect 9033 3955 9091 3961
rect 10689 3961 10701 3995
rect 10735 3961 10747 3995
rect 10689 3955 10747 3961
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 1670 3924 1676 3936
rect 1627 3896 1676 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 1854 3884 1860 3936
rect 1912 3924 1918 3936
rect 2593 3927 2651 3933
rect 2593 3924 2605 3927
rect 1912 3896 2605 3924
rect 1912 3884 1918 3896
rect 2593 3893 2605 3896
rect 2639 3893 2651 3927
rect 2593 3887 2651 3893
rect 3142 3884 3148 3936
rect 3200 3924 3206 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3200 3896 4077 3924
rect 3200 3884 3206 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 4890 3884 4896 3936
rect 4948 3884 4954 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 5960 3896 6469 3924
rect 5960 3884 5966 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 6457 3887 6515 3893
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8294 3924 8300 3936
rect 8159 3896 8300 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10192 3896 10333 3924
rect 10192 3884 10198 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 13648 3924 13676 4100
rect 14093 4097 14105 4131
rect 14139 4128 14151 4131
rect 14550 4128 14556 4140
rect 14139 4100 14556 4128
rect 14139 4097 14151 4100
rect 14093 4091 14151 4097
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 14660 4128 14688 4168
rect 14734 4156 14740 4208
rect 14792 4156 14798 4208
rect 14844 4205 14872 4236
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 17681 4267 17739 4273
rect 17681 4233 17693 4267
rect 17727 4264 17739 4267
rect 18046 4264 18052 4276
rect 17727 4236 18052 4264
rect 17727 4233 17739 4236
rect 17681 4227 17739 4233
rect 18046 4224 18052 4236
rect 18104 4224 18110 4276
rect 18966 4224 18972 4276
rect 19024 4224 19030 4276
rect 14829 4199 14887 4205
rect 14829 4165 14841 4199
rect 14875 4165 14887 4199
rect 15304 4196 15332 4224
rect 15304 4168 15424 4196
rect 14829 4159 14887 4165
rect 15102 4128 15108 4140
rect 14660 4100 15108 4128
rect 13722 4020 13728 4072
rect 13780 4060 13786 4072
rect 14752 4069 14780 4100
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 15286 4137 15292 4140
rect 15280 4091 15292 4137
rect 15286 4088 15292 4091
rect 15344 4088 15350 4140
rect 15396 4128 15424 4168
rect 18230 4156 18236 4208
rect 18288 4196 18294 4208
rect 18509 4199 18567 4205
rect 18509 4196 18521 4199
rect 18288 4168 18521 4196
rect 18288 4156 18294 4168
rect 18509 4165 18521 4168
rect 18555 4165 18567 4199
rect 18984 4196 19012 4224
rect 20073 4199 20131 4205
rect 18984 4168 19748 4196
rect 18509 4159 18567 4165
rect 16298 4128 16304 4140
rect 15396 4100 16304 4128
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 18046 4128 18052 4140
rect 17543 4100 18052 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4097 19027 4131
rect 18969 4091 19027 4097
rect 19245 4131 19303 4137
rect 19245 4097 19257 4131
rect 19291 4128 19303 4131
rect 19595 4131 19653 4137
rect 19595 4128 19607 4131
rect 19291 4100 19607 4128
rect 19291 4097 19303 4100
rect 19245 4091 19303 4097
rect 19595 4097 19607 4100
rect 19641 4097 19653 4131
rect 19720 4128 19748 4168
rect 20073 4165 20085 4199
rect 20119 4196 20131 4199
rect 20622 4196 20628 4208
rect 20119 4168 20628 4196
rect 20119 4165 20131 4168
rect 20073 4159 20131 4165
rect 20622 4156 20628 4168
rect 20680 4156 20686 4208
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 19720 4100 20177 4128
rect 19595 4091 19653 4097
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 14259 4063 14317 4069
rect 14259 4060 14271 4063
rect 13780 4032 14271 4060
rect 13780 4020 13786 4032
rect 14259 4029 14271 4032
rect 14305 4029 14317 4063
rect 14259 4023 14317 4029
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4029 14795 4063
rect 14737 4023 14795 4029
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 17773 4063 17831 4069
rect 17773 4029 17785 4063
rect 17819 4029 17831 4063
rect 17773 4023 17831 4029
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 15028 3992 15056 4023
rect 13872 3964 15056 3992
rect 13872 3952 13878 3964
rect 16574 3952 16580 4004
rect 16632 3992 16638 4004
rect 17221 3995 17279 4001
rect 17221 3992 17233 3995
rect 16632 3964 17233 3992
rect 16632 3952 16638 3964
rect 17221 3961 17233 3964
rect 17267 3961 17279 3995
rect 17788 3992 17816 4023
rect 18506 4020 18512 4072
rect 18564 4020 18570 4072
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4029 18659 4063
rect 18984 4060 19012 4091
rect 18984 4032 19840 4060
rect 18601 4023 18659 4029
rect 18616 3992 18644 4023
rect 19429 3995 19487 4001
rect 17788 3964 19288 3992
rect 17221 3955 17279 3961
rect 11112 3896 13676 3924
rect 11112 3884 11118 3896
rect 13906 3884 13912 3936
rect 13964 3884 13970 3936
rect 16393 3927 16451 3933
rect 16393 3893 16405 3927
rect 16439 3924 16451 3927
rect 16850 3924 16856 3936
rect 16439 3896 16856 3924
rect 16439 3893 16451 3896
rect 16393 3887 16451 3893
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 16942 3884 16948 3936
rect 17000 3924 17006 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17000 3896 18061 3924
rect 17000 3884 17006 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 19153 3927 19211 3933
rect 19153 3924 19165 3927
rect 19116 3896 19165 3924
rect 19116 3884 19122 3896
rect 19153 3893 19165 3896
rect 19199 3893 19211 3927
rect 19260 3924 19288 3964
rect 19429 3961 19441 3995
rect 19475 3992 19487 3995
rect 19702 3992 19708 4004
rect 19475 3964 19708 3992
rect 19475 3961 19487 3964
rect 19429 3955 19487 3961
rect 19702 3952 19708 3964
rect 19760 3952 19766 4004
rect 19812 3992 19840 4032
rect 19886 4020 19892 4072
rect 19944 4060 19950 4072
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19944 4032 19993 4060
rect 19944 4020 19950 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 20898 3992 20904 4004
rect 19812 3964 20904 3992
rect 20898 3952 20904 3964
rect 20956 3952 20962 4004
rect 20990 3924 20996 3936
rect 19260 3896 20996 3924
rect 19153 3887 19211 3893
rect 20990 3884 20996 3896
rect 21048 3884 21054 3936
rect 1104 3834 21988 3856
rect 1104 3782 3560 3834
rect 3612 3782 3624 3834
rect 3676 3782 3688 3834
rect 3740 3782 3752 3834
rect 3804 3782 3816 3834
rect 3868 3782 8781 3834
rect 8833 3782 8845 3834
rect 8897 3782 8909 3834
rect 8961 3782 8973 3834
rect 9025 3782 9037 3834
rect 9089 3782 14002 3834
rect 14054 3782 14066 3834
rect 14118 3782 14130 3834
rect 14182 3782 14194 3834
rect 14246 3782 14258 3834
rect 14310 3782 19223 3834
rect 19275 3782 19287 3834
rect 19339 3782 19351 3834
rect 19403 3782 19415 3834
rect 19467 3782 19479 3834
rect 19531 3782 21988 3834
rect 1104 3760 21988 3782
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5258 3720 5264 3732
rect 5215 3692 5264 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 6825 3723 6883 3729
rect 6825 3689 6837 3723
rect 6871 3720 6883 3723
rect 6914 3720 6920 3732
rect 6871 3692 6920 3720
rect 6871 3689 6883 3692
rect 6825 3683 6883 3689
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 7926 3680 7932 3732
rect 7984 3720 7990 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 7984 3692 9045 3720
rect 7984 3680 7990 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 15010 3720 15016 3732
rect 14792 3692 15016 3720
rect 14792 3680 14798 3692
rect 15010 3680 15016 3692
rect 15068 3720 15074 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15068 3692 15485 3720
rect 15068 3680 15074 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 18966 3720 18972 3732
rect 15473 3683 15531 3689
rect 18248 3692 18972 3720
rect 8110 3612 8116 3664
rect 8168 3612 8174 3664
rect 12069 3655 12127 3661
rect 12069 3621 12081 3655
rect 12115 3621 12127 3655
rect 12069 3615 12127 3621
rect 3694 3584 3700 3596
rect 2884 3556 3700 3584
rect 2884 3528 2912 3556
rect 3694 3544 3700 3556
rect 3752 3584 3758 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 3752 3556 3801 3584
rect 3752 3544 3758 3556
rect 3789 3553 3801 3556
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 5442 3544 5448 3596
rect 5500 3544 5506 3596
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 8680 3556 9597 3584
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 2866 3516 2872 3528
rect 1636 3488 2872 3516
rect 1636 3476 1642 3488
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3142 3476 3148 3528
rect 3200 3476 3206 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 4890 3516 4896 3528
rect 3467 3488 4896 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 6512 3488 7389 3516
rect 6512 3476 6518 3488
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 8478 3516 8484 3528
rect 7377 3479 7435 3485
rect 7668 3488 8484 3516
rect 1848 3451 1906 3457
rect 1848 3417 1860 3451
rect 1894 3448 1906 3451
rect 1946 3448 1952 3460
rect 1894 3420 1952 3448
rect 1894 3417 1906 3420
rect 1848 3411 1906 3417
rect 1946 3408 1952 3420
rect 2004 3408 2010 3460
rect 4034 3451 4092 3457
rect 4034 3448 4046 3451
rect 3344 3420 4046 3448
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3344 3389 3372 3420
rect 4034 3417 4046 3420
rect 4080 3417 4092 3451
rect 4034 3411 4092 3417
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 5350 3448 5356 3460
rect 4212 3420 5356 3448
rect 4212 3408 4218 3420
rect 5350 3408 5356 3420
rect 5408 3408 5414 3460
rect 5718 3457 5724 3460
rect 5712 3411 5724 3457
rect 5718 3408 5724 3411
rect 5776 3408 5782 3460
rect 5994 3408 6000 3460
rect 6052 3448 6058 3460
rect 7083 3451 7141 3457
rect 7083 3448 7095 3451
rect 6052 3420 7095 3448
rect 6052 3408 6058 3420
rect 7083 3417 7095 3420
rect 7129 3417 7141 3451
rect 7083 3411 7141 3417
rect 7466 3408 7472 3460
rect 7524 3448 7530 3460
rect 7668 3457 7696 3488
rect 8478 3476 8484 3488
rect 8536 3516 8542 3528
rect 8680 3525 8708 3556
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9824 3556 9873 3584
rect 9824 3544 9830 3556
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 10134 3525 10140 3528
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 8536 3488 8677 3516
rect 8536 3476 8542 3488
rect 8665 3485 8677 3488
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 10128 3516 10140 3525
rect 9355 3488 9904 3516
rect 10095 3488 10140 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9876 3460 9904 3488
rect 10128 3479 10140 3488
rect 10134 3476 10140 3479
rect 10192 3476 10198 3528
rect 11330 3476 11336 3528
rect 11388 3516 11394 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11388 3488 11621 3516
rect 11388 3476 11394 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 11885 3519 11943 3525
rect 11885 3485 11897 3519
rect 11931 3516 11943 3519
rect 12084 3516 12112 3615
rect 13354 3612 13360 3664
rect 13412 3652 13418 3664
rect 13449 3655 13507 3661
rect 13449 3652 13461 3655
rect 13412 3624 13461 3652
rect 13412 3612 13418 3624
rect 13449 3621 13461 3624
rect 13495 3621 13507 3655
rect 13449 3615 13507 3621
rect 16758 3612 16764 3664
rect 16816 3652 16822 3664
rect 17865 3655 17923 3661
rect 17865 3652 17877 3655
rect 16816 3624 17877 3652
rect 16816 3612 16822 3624
rect 17865 3621 17877 3624
rect 17911 3621 17923 3655
rect 17865 3615 17923 3621
rect 12526 3544 12532 3596
rect 12584 3544 12590 3596
rect 13814 3584 13820 3596
rect 13648 3556 13820 3584
rect 13648 3516 13676 3556
rect 13814 3544 13820 3556
rect 13872 3584 13878 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13872 3556 14105 3584
rect 13872 3544 13878 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 11931 3488 12112 3516
rect 12406 3488 13676 3516
rect 11931 3485 11943 3488
rect 11885 3479 11943 3485
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 7524 3420 7573 3448
rect 7524 3408 7530 3420
rect 7561 3417 7573 3420
rect 7607 3417 7619 3451
rect 7561 3411 7619 3417
rect 7653 3451 7711 3457
rect 7653 3417 7665 3451
rect 7699 3417 7711 3451
rect 7653 3411 7711 3417
rect 2961 3383 3019 3389
rect 2961 3380 2973 3383
rect 2924 3352 2973 3380
rect 2924 3340 2930 3352
rect 2961 3349 2973 3352
rect 3007 3349 3019 3383
rect 2961 3343 3019 3349
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3349 3387 3383
rect 3329 3343 3387 3349
rect 3602 3340 3608 3392
rect 3660 3340 3666 3392
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5626 3380 5632 3392
rect 5040 3352 5632 3380
rect 5040 3340 5046 3352
rect 5626 3340 5632 3352
rect 5684 3380 5690 3392
rect 7668 3380 7696 3411
rect 8386 3408 8392 3460
rect 8444 3408 8450 3460
rect 9490 3408 9496 3460
rect 9548 3408 9554 3460
rect 9858 3408 9864 3460
rect 9916 3408 9922 3460
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 12066 3448 12072 3460
rect 11572 3420 12072 3448
rect 11572 3408 11578 3420
rect 12066 3408 12072 3420
rect 12124 3448 12130 3460
rect 12406 3448 12434 3488
rect 13722 3476 13728 3528
rect 13780 3476 13786 3528
rect 14108 3516 14136 3547
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 15160 3556 15792 3584
rect 15160 3544 15166 3556
rect 15657 3519 15715 3525
rect 15657 3516 15669 3519
rect 14108 3488 15669 3516
rect 15657 3485 15669 3488
rect 15703 3485 15715 3519
rect 15764 3516 15792 3556
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 17402 3584 17408 3596
rect 16908 3556 17408 3584
rect 16908 3544 16914 3556
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 18141 3587 18199 3593
rect 18141 3553 18153 3587
rect 18187 3584 18199 3587
rect 18248 3584 18276 3692
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 20622 3680 20628 3732
rect 20680 3680 20686 3732
rect 20898 3680 20904 3732
rect 20956 3680 20962 3732
rect 18693 3655 18751 3661
rect 18693 3621 18705 3655
rect 18739 3621 18751 3655
rect 18693 3615 18751 3621
rect 18187 3556 18276 3584
rect 18187 3553 18199 3556
rect 18141 3547 18199 3553
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 15764 3488 18429 3516
rect 15657 3479 15715 3485
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18708 3516 18736 3615
rect 21358 3544 21364 3596
rect 21416 3544 21422 3596
rect 19061 3519 19119 3525
rect 19061 3516 19073 3519
rect 18708 3488 19073 3516
rect 18417 3479 18475 3485
rect 19061 3485 19073 3488
rect 19107 3485 19119 3519
rect 19061 3479 19119 3485
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 12124 3420 12434 3448
rect 12124 3408 12130 3420
rect 12618 3408 12624 3460
rect 12676 3408 12682 3460
rect 12897 3451 12955 3457
rect 12897 3417 12909 3451
rect 12943 3448 12955 3451
rect 12943 3420 13124 3448
rect 12943 3417 12955 3420
rect 12897 3411 12955 3417
rect 5684 3352 7696 3380
rect 5684 3340 5690 3352
rect 8570 3340 8576 3392
rect 8628 3340 8634 3392
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 11241 3383 11299 3389
rect 11241 3380 11253 3383
rect 11020 3352 11253 3380
rect 11020 3340 11026 3352
rect 11241 3349 11253 3352
rect 11287 3349 11299 3383
rect 11241 3343 11299 3349
rect 11422 3340 11428 3392
rect 11480 3340 11486 3392
rect 11701 3383 11759 3389
rect 11701 3349 11713 3383
rect 11747 3380 11759 3383
rect 11790 3380 11796 3392
rect 11747 3352 11796 3380
rect 11747 3349 11759 3352
rect 11701 3343 11759 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 12529 3383 12587 3389
rect 12529 3349 12541 3383
rect 12575 3380 12587 3383
rect 12986 3380 12992 3392
rect 12575 3352 12992 3380
rect 12575 3349 12587 3352
rect 12529 3343 12587 3349
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13096 3380 13124 3420
rect 13170 3408 13176 3460
rect 13228 3408 13234 3460
rect 14338 3451 14396 3457
rect 14338 3448 14350 3451
rect 13924 3420 14350 3448
rect 13722 3380 13728 3392
rect 13096 3352 13728 3380
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13924 3389 13952 3420
rect 14338 3417 14350 3420
rect 14384 3417 14396 3451
rect 14338 3411 14396 3417
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 15902 3451 15960 3457
rect 15902 3448 15914 3451
rect 15620 3420 15914 3448
rect 15620 3408 15626 3420
rect 15902 3417 15914 3420
rect 15948 3417 15960 3451
rect 15902 3411 15960 3417
rect 16666 3408 16672 3460
rect 16724 3448 16730 3460
rect 17313 3451 17371 3457
rect 17313 3448 17325 3451
rect 16724 3420 17325 3448
rect 16724 3408 16730 3420
rect 17313 3417 17325 3420
rect 17359 3417 17371 3451
rect 17313 3411 17371 3417
rect 18690 3408 18696 3460
rect 18748 3448 18754 3460
rect 19260 3448 19288 3479
rect 20990 3476 20996 3528
rect 21048 3516 21054 3528
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 21048 3488 21465 3516
rect 21048 3476 21054 3488
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 18748 3420 19288 3448
rect 19512 3451 19570 3457
rect 18748 3408 18754 3420
rect 19512 3417 19524 3451
rect 19558 3448 19570 3451
rect 19702 3448 19708 3460
rect 19558 3420 19708 3448
rect 19558 3417 19570 3420
rect 19512 3411 19570 3417
rect 19702 3408 19708 3420
rect 19760 3408 19766 3460
rect 13909 3383 13967 3389
rect 13909 3349 13921 3383
rect 13955 3349 13967 3383
rect 13909 3343 13967 3349
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 17405 3383 17463 3389
rect 17405 3380 17417 3383
rect 17092 3352 17417 3380
rect 17092 3340 17098 3352
rect 17405 3349 17417 3352
rect 17451 3349 17463 3383
rect 17405 3343 17463 3349
rect 18230 3340 18236 3392
rect 18288 3340 18294 3392
rect 18874 3340 18880 3392
rect 18932 3340 18938 3392
rect 20622 3340 20628 3392
rect 20680 3380 20686 3392
rect 21361 3383 21419 3389
rect 21361 3380 21373 3383
rect 20680 3352 21373 3380
rect 20680 3340 20686 3352
rect 21361 3349 21373 3352
rect 21407 3349 21419 3383
rect 21361 3343 21419 3349
rect 1104 3290 21988 3312
rect 1104 3238 4220 3290
rect 4272 3238 4284 3290
rect 4336 3238 4348 3290
rect 4400 3238 4412 3290
rect 4464 3238 4476 3290
rect 4528 3238 9441 3290
rect 9493 3238 9505 3290
rect 9557 3238 9569 3290
rect 9621 3238 9633 3290
rect 9685 3238 9697 3290
rect 9749 3238 14662 3290
rect 14714 3238 14726 3290
rect 14778 3238 14790 3290
rect 14842 3238 14854 3290
rect 14906 3238 14918 3290
rect 14970 3238 19883 3290
rect 19935 3238 19947 3290
rect 19999 3238 20011 3290
rect 20063 3238 20075 3290
rect 20127 3238 20139 3290
rect 20191 3238 21988 3290
rect 1104 3216 21988 3238
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3050 3176 3056 3188
rect 3007 3148 3056 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 5074 3136 5080 3188
rect 5132 3136 5138 3188
rect 5718 3136 5724 3188
rect 5776 3136 5782 3188
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7524 3148 7757 3176
rect 7524 3136 7530 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9364 3148 9413 3176
rect 9364 3136 9370 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 11146 3136 11152 3188
rect 11204 3136 11210 3188
rect 13173 3179 13231 3185
rect 13173 3176 13185 3179
rect 12406 3148 13185 3176
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 1826 3111 1884 3117
rect 1826 3108 1838 3111
rect 1728 3080 1838 3108
rect 1728 3068 1734 3080
rect 1826 3077 1838 3080
rect 1872 3077 1884 3111
rect 1826 3071 1884 3077
rect 3602 3068 3608 3120
rect 3660 3108 3666 3120
rect 3942 3111 4000 3117
rect 3942 3108 3954 3111
rect 3660 3080 3954 3108
rect 3660 3068 3666 3080
rect 3942 3077 3954 3080
rect 3988 3077 4000 3111
rect 3942 3071 4000 3077
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 7282 3108 7288 3120
rect 5500 3080 7288 3108
rect 5500 3068 5506 3080
rect 1578 3000 1584 3052
rect 1636 3000 1642 3052
rect 3694 3000 3700 3052
rect 3752 3000 3758 3052
rect 5902 3000 5908 3052
rect 5960 3000 5966 3052
rect 5994 3000 6000 3052
rect 6052 3000 6058 3052
rect 6380 3049 6408 3080
rect 7282 3068 7288 3080
rect 7340 3108 7346 3120
rect 8294 3117 8300 3120
rect 8288 3108 8300 3117
rect 7340 3080 8064 3108
rect 8255 3080 8300 3108
rect 7340 3068 7346 3080
rect 8036 3049 8064 3080
rect 8288 3071 8300 3080
rect 8294 3068 8300 3071
rect 8352 3068 8358 3120
rect 10036 3111 10094 3117
rect 10036 3077 10048 3111
rect 10082 3108 10094 3111
rect 11422 3108 11428 3120
rect 10082 3080 11428 3108
rect 10082 3077 10094 3080
rect 10036 3071 10094 3077
rect 11422 3068 11428 3080
rect 11480 3068 11486 3120
rect 11876 3111 11934 3117
rect 11876 3077 11888 3111
rect 11922 3108 11934 3111
rect 12406 3108 12434 3148
rect 13173 3145 13185 3148
rect 13219 3145 13231 3179
rect 13173 3139 13231 3145
rect 13832 3148 14780 3176
rect 11922 3080 12434 3108
rect 11922 3077 11934 3080
rect 11876 3071 11934 3077
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 13832 3108 13860 3148
rect 12584 3080 13860 3108
rect 12584 3068 12590 3080
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 14062 3111 14120 3117
rect 14062 3108 14074 3111
rect 13964 3080 14074 3108
rect 13964 3068 13970 3080
rect 14062 3077 14074 3080
rect 14108 3077 14120 3111
rect 14752 3108 14780 3148
rect 15562 3136 15568 3188
rect 15620 3136 15626 3188
rect 16209 3179 16267 3185
rect 16209 3145 16221 3179
rect 16255 3176 16267 3179
rect 17034 3176 17040 3188
rect 16255 3148 17040 3176
rect 16255 3145 16267 3148
rect 16209 3139 16267 3145
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3176 17371 3179
rect 18230 3176 18236 3188
rect 17359 3148 18236 3176
rect 17359 3145 17371 3148
rect 17313 3139 17371 3145
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 19794 3176 19800 3188
rect 18340 3148 19800 3176
rect 16025 3111 16083 3117
rect 16025 3108 16037 3111
rect 14752 3080 16037 3108
rect 14062 3071 14120 3077
rect 16025 3077 16037 3080
rect 16071 3108 16083 3111
rect 18340 3108 18368 3148
rect 19794 3136 19800 3148
rect 19852 3136 19858 3188
rect 20349 3179 20407 3185
rect 20349 3145 20361 3179
rect 20395 3176 20407 3179
rect 21358 3176 21364 3188
rect 20395 3148 21364 3176
rect 20395 3145 20407 3148
rect 20349 3139 20407 3145
rect 21358 3136 21364 3148
rect 21416 3136 21422 3188
rect 16071 3080 18368 3108
rect 18448 3111 18506 3117
rect 16071 3077 16083 3080
rect 16025 3071 16083 3077
rect 18448 3077 18460 3111
rect 18494 3108 18506 3111
rect 18874 3108 18880 3120
rect 18494 3080 18880 3108
rect 18494 3077 18506 3080
rect 18448 3071 18506 3077
rect 18874 3068 18880 3080
rect 18932 3068 18938 3120
rect 19058 3068 19064 3120
rect 19116 3108 19122 3120
rect 19214 3111 19272 3117
rect 19214 3108 19226 3111
rect 19116 3080 19226 3108
rect 19116 3068 19122 3080
rect 19214 3077 19226 3080
rect 19260 3077 19272 3111
rect 19214 3071 19272 3077
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6621 3043 6679 3049
rect 6621 3040 6633 3043
rect 6365 3003 6423 3009
rect 6472 3012 6633 3040
rect 6472 2972 6500 3012
rect 6621 3009 6633 3012
rect 6667 3009 6679 3043
rect 6621 3003 6679 3009
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 13354 3000 13360 3052
rect 13412 3000 13418 3052
rect 13814 3000 13820 3052
rect 13872 3000 13878 3052
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 15427 3012 15792 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 6380 2944 6500 2972
rect 6181 2907 6239 2913
rect 6181 2873 6193 2907
rect 6227 2904 6239 2907
rect 6380 2904 6408 2944
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 11609 2975 11667 2981
rect 11609 2972 11621 2975
rect 11572 2944 11621 2972
rect 11572 2932 11578 2944
rect 11609 2941 11621 2944
rect 11655 2941 11667 2975
rect 11609 2935 11667 2941
rect 6227 2876 6408 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 12894 2864 12900 2916
rect 12952 2904 12958 2916
rect 12989 2907 13047 2913
rect 12989 2904 13001 2907
rect 12952 2876 13001 2904
rect 12952 2864 12958 2876
rect 12989 2873 13001 2876
rect 13035 2904 13047 2907
rect 13170 2904 13176 2916
rect 13035 2876 13176 2904
rect 13035 2873 13047 2876
rect 12989 2867 13047 2873
rect 13170 2864 13176 2876
rect 13228 2864 13234 2916
rect 15764 2913 15792 3012
rect 16298 3000 16304 3052
rect 16356 3000 16362 3052
rect 16942 3000 16948 3052
rect 17000 3000 17006 3052
rect 18690 2932 18696 2984
rect 18748 2972 18754 2984
rect 18969 2975 19027 2981
rect 18969 2972 18981 2975
rect 18748 2944 18981 2972
rect 18748 2932 18754 2944
rect 18969 2941 18981 2944
rect 19015 2941 19027 2975
rect 18969 2935 19027 2941
rect 15749 2907 15807 2913
rect 15749 2873 15761 2907
rect 15795 2873 15807 2907
rect 15749 2867 15807 2873
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 9122 2836 9128 2848
rect 5408 2808 9128 2836
rect 5408 2796 5414 2808
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 15197 2839 15255 2845
rect 15197 2805 15209 2839
rect 15243 2836 15255 2839
rect 15470 2836 15476 2848
rect 15243 2808 15476 2836
rect 15243 2805 15255 2808
rect 15197 2799 15255 2805
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 17126 2796 17132 2848
rect 17184 2796 17190 2848
rect 1104 2746 21988 2768
rect 1104 2694 3560 2746
rect 3612 2694 3624 2746
rect 3676 2694 3688 2746
rect 3740 2694 3752 2746
rect 3804 2694 3816 2746
rect 3868 2694 8781 2746
rect 8833 2694 8845 2746
rect 8897 2694 8909 2746
rect 8961 2694 8973 2746
rect 9025 2694 9037 2746
rect 9089 2694 14002 2746
rect 14054 2694 14066 2746
rect 14118 2694 14130 2746
rect 14182 2694 14194 2746
rect 14246 2694 14258 2746
rect 14310 2694 19223 2746
rect 19275 2694 19287 2746
rect 19339 2694 19351 2746
rect 19403 2694 19415 2746
rect 19467 2694 19479 2746
rect 19531 2694 21988 2746
rect 1104 2672 21988 2694
rect 1946 2592 1952 2644
rect 2004 2592 2010 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4614 2632 4620 2644
rect 4387 2604 4620 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 8665 2635 8723 2641
rect 8665 2632 8677 2635
rect 8628 2604 8677 2632
rect 8628 2592 8634 2604
rect 8665 2601 8677 2604
rect 8711 2601 8723 2635
rect 8665 2595 8723 2601
rect 10965 2635 11023 2641
rect 10965 2601 10977 2635
rect 11011 2632 11023 2635
rect 11330 2632 11336 2644
rect 11011 2604 11336 2632
rect 11011 2601 11023 2604
rect 10965 2595 11023 2601
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 12618 2632 12624 2644
rect 11532 2604 12624 2632
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2533 2467 2567
rect 4982 2564 4988 2576
rect 2409 2527 2467 2533
rect 2976 2536 4988 2564
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2424 2428 2452 2527
rect 2774 2456 2780 2508
rect 2832 2456 2838 2508
rect 2976 2505 3004 2536
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 11532 2564 11560 2604
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 12897 2635 12955 2641
rect 12897 2601 12909 2635
rect 12943 2632 12955 2635
rect 12986 2632 12992 2644
rect 12943 2604 12992 2632
rect 12943 2601 12955 2604
rect 12897 2595 12955 2601
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 14550 2592 14556 2644
rect 14608 2592 14614 2644
rect 15286 2592 15292 2644
rect 15344 2632 15350 2644
rect 15381 2635 15439 2641
rect 15381 2632 15393 2635
rect 15344 2604 15393 2632
rect 15344 2592 15350 2604
rect 15381 2601 15393 2604
rect 15427 2601 15439 2635
rect 15381 2595 15439 2601
rect 10428 2536 11560 2564
rect 2961 2499 3019 2505
rect 2961 2465 2973 2499
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 3108 2468 4108 2496
rect 3108 2456 3114 2468
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2179 2400 2452 2428
rect 2884 2400 3801 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2884 2372 2912 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 4080 2437 4108 2468
rect 7282 2456 7288 2508
rect 7340 2456 7346 2508
rect 10428 2505 10456 2536
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2465 10471 2499
rect 10413 2459 10471 2465
rect 11514 2456 11520 2508
rect 11572 2456 11578 2508
rect 15013 2499 15071 2505
rect 15013 2465 15025 2499
rect 15059 2496 15071 2499
rect 15470 2496 15476 2508
rect 15059 2468 15476 2496
rect 15059 2465 15071 2468
rect 15013 2459 15071 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 4209 2431 4267 2437
rect 4209 2397 4221 2431
rect 4255 2428 4267 2431
rect 5350 2428 5356 2440
rect 4255 2400 5356 2428
rect 4255 2397 4267 2400
rect 4209 2391 4267 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8110 2428 8116 2440
rect 7055 2400 8116 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 11054 2428 11060 2440
rect 10735 2400 11060 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11790 2437 11796 2440
rect 11784 2428 11796 2437
rect 11751 2400 11796 2428
rect 11784 2391 11796 2400
rect 11790 2388 11796 2391
rect 11848 2388 11854 2440
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 13872 2400 15117 2428
rect 13872 2388 13878 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2428 15623 2431
rect 16758 2428 16764 2440
rect 15611 2400 16764 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 18690 2428 18696 2440
rect 17267 2400 18696 2428
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 18690 2388 18696 2400
rect 18748 2388 18754 2440
rect 2866 2320 2872 2372
rect 2924 2320 2930 2372
rect 7530 2363 7588 2369
rect 7530 2360 7542 2363
rect 7208 2332 7542 2360
rect 7208 2301 7236 2332
rect 7530 2329 7542 2332
rect 7576 2329 7588 2363
rect 7530 2323 7588 2329
rect 15010 2320 15016 2372
rect 15068 2320 15074 2372
rect 17126 2320 17132 2372
rect 17184 2360 17190 2372
rect 17466 2363 17524 2369
rect 17466 2360 17478 2363
rect 17184 2332 17478 2360
rect 17184 2320 17190 2332
rect 17466 2329 17478 2332
rect 17512 2329 17524 2363
rect 17466 2323 17524 2329
rect 7193 2295 7251 2301
rect 7193 2261 7205 2295
rect 7239 2261 7251 2295
rect 7193 2255 7251 2261
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2292 10563 2295
rect 11146 2292 11152 2304
rect 10551 2264 11152 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 18506 2252 18512 2304
rect 18564 2292 18570 2304
rect 18601 2295 18659 2301
rect 18601 2292 18613 2295
rect 18564 2264 18613 2292
rect 18564 2252 18570 2264
rect 18601 2261 18613 2264
rect 18647 2292 18659 2295
rect 18690 2292 18696 2304
rect 18647 2264 18696 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 18690 2252 18696 2264
rect 18748 2252 18754 2304
rect 1104 2202 21988 2224
rect 1104 2150 4220 2202
rect 4272 2150 4284 2202
rect 4336 2150 4348 2202
rect 4400 2150 4412 2202
rect 4464 2150 4476 2202
rect 4528 2150 9441 2202
rect 9493 2150 9505 2202
rect 9557 2150 9569 2202
rect 9621 2150 9633 2202
rect 9685 2150 9697 2202
rect 9749 2150 14662 2202
rect 14714 2150 14726 2202
rect 14778 2150 14790 2202
rect 14842 2150 14854 2202
rect 14906 2150 14918 2202
rect 14970 2150 19883 2202
rect 19935 2150 19947 2202
rect 19999 2150 20011 2202
rect 20063 2150 20075 2202
rect 20127 2150 20139 2202
rect 20191 2150 21988 2202
rect 1104 2128 21988 2150
<< via1 >>
rect 4220 22822 4272 22874
rect 4284 22822 4336 22874
rect 4348 22822 4400 22874
rect 4412 22822 4464 22874
rect 4476 22822 4528 22874
rect 9441 22822 9493 22874
rect 9505 22822 9557 22874
rect 9569 22822 9621 22874
rect 9633 22822 9685 22874
rect 9697 22822 9749 22874
rect 14662 22822 14714 22874
rect 14726 22822 14778 22874
rect 14790 22822 14842 22874
rect 14854 22822 14906 22874
rect 14918 22822 14970 22874
rect 19883 22822 19935 22874
rect 19947 22822 19999 22874
rect 20011 22822 20063 22874
rect 20075 22822 20127 22874
rect 20139 22822 20191 22874
rect 7104 22720 7156 22772
rect 7380 22720 7432 22772
rect 9036 22720 9088 22772
rect 3056 22652 3108 22704
rect 8576 22652 8628 22704
rect 2780 22516 2832 22568
rect 2044 22380 2096 22432
rect 2780 22380 2832 22432
rect 4804 22559 4856 22568
rect 4804 22525 4813 22559
rect 4813 22525 4847 22559
rect 4847 22525 4856 22559
rect 4804 22516 4856 22525
rect 6920 22584 6972 22636
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 9220 22584 9272 22636
rect 11612 22584 11664 22636
rect 13820 22584 13872 22636
rect 17868 22652 17920 22704
rect 16396 22584 16448 22636
rect 19340 22652 19392 22704
rect 19616 22652 19668 22704
rect 18696 22584 18748 22636
rect 21364 22652 21416 22704
rect 7012 22559 7064 22568
rect 7012 22525 7021 22559
rect 7021 22525 7055 22559
rect 7055 22525 7064 22559
rect 7012 22516 7064 22525
rect 9588 22559 9640 22568
rect 9588 22525 9597 22559
rect 9597 22525 9631 22559
rect 9631 22525 9640 22559
rect 9588 22516 9640 22525
rect 16028 22516 16080 22568
rect 16856 22516 16908 22568
rect 21088 22627 21140 22636
rect 21088 22593 21097 22627
rect 21097 22593 21131 22627
rect 21131 22593 21140 22627
rect 21088 22584 21140 22593
rect 16396 22448 16448 22500
rect 19708 22516 19760 22568
rect 20536 22516 20588 22568
rect 20996 22516 21048 22568
rect 18788 22448 18840 22500
rect 5448 22423 5500 22432
rect 5448 22389 5457 22423
rect 5457 22389 5491 22423
rect 5491 22389 5500 22423
rect 5448 22380 5500 22389
rect 5816 22380 5868 22432
rect 8668 22423 8720 22432
rect 8668 22389 8677 22423
rect 8677 22389 8711 22423
rect 8711 22389 8720 22423
rect 8668 22380 8720 22389
rect 9128 22380 9180 22432
rect 11060 22380 11112 22432
rect 12992 22423 13044 22432
rect 12992 22389 13001 22423
rect 13001 22389 13035 22423
rect 13035 22389 13044 22423
rect 12992 22380 13044 22389
rect 16672 22380 16724 22432
rect 17316 22423 17368 22432
rect 17316 22389 17325 22423
rect 17325 22389 17359 22423
rect 17359 22389 17368 22423
rect 17316 22380 17368 22389
rect 18512 22423 18564 22432
rect 18512 22389 18521 22423
rect 18521 22389 18555 22423
rect 18555 22389 18564 22423
rect 18512 22380 18564 22389
rect 20628 22380 20680 22432
rect 3560 22278 3612 22330
rect 3624 22278 3676 22330
rect 3688 22278 3740 22330
rect 3752 22278 3804 22330
rect 3816 22278 3868 22330
rect 8781 22278 8833 22330
rect 8845 22278 8897 22330
rect 8909 22278 8961 22330
rect 8973 22278 9025 22330
rect 9037 22278 9089 22330
rect 14002 22278 14054 22330
rect 14066 22278 14118 22330
rect 14130 22278 14182 22330
rect 14194 22278 14246 22330
rect 14258 22278 14310 22330
rect 19223 22278 19275 22330
rect 19287 22278 19339 22330
rect 19351 22278 19403 22330
rect 19415 22278 19467 22330
rect 19479 22278 19531 22330
rect 3976 22040 4028 22092
rect 7104 22219 7156 22228
rect 7104 22185 7113 22219
rect 7113 22185 7147 22219
rect 7147 22185 7156 22219
rect 7104 22176 7156 22185
rect 9588 22176 9640 22228
rect 13820 22176 13872 22228
rect 7380 22151 7432 22160
rect 7380 22117 7389 22151
rect 7389 22117 7423 22151
rect 7423 22117 7432 22151
rect 7380 22108 7432 22117
rect 8944 22108 8996 22160
rect 9220 22108 9272 22160
rect 9312 22083 9364 22092
rect 2044 22015 2096 22024
rect 2044 21981 2053 22015
rect 2053 21981 2087 22015
rect 2087 21981 2096 22015
rect 2044 21972 2096 21981
rect 2780 21972 2832 22024
rect 4068 21972 4120 22024
rect 5632 22015 5684 22024
rect 5632 21981 5641 22015
rect 5641 21981 5675 22015
rect 5675 21981 5684 22015
rect 5632 21972 5684 21981
rect 5816 21972 5868 22024
rect 9312 22049 9321 22083
rect 9321 22049 9355 22083
rect 9355 22049 9364 22083
rect 9312 22040 9364 22049
rect 8852 21972 8904 22024
rect 10876 21972 10928 22024
rect 2964 21904 3016 21956
rect 1676 21836 1728 21888
rect 3884 21836 3936 21888
rect 4620 21836 4672 21888
rect 8300 21904 8352 21956
rect 9220 21904 9272 21956
rect 10048 21836 10100 21888
rect 10784 21836 10836 21888
rect 11244 21947 11296 21956
rect 11244 21913 11253 21947
rect 11253 21913 11287 21947
rect 11287 21913 11296 21947
rect 11244 21904 11296 21913
rect 11336 21947 11388 21956
rect 11336 21913 11345 21947
rect 11345 21913 11379 21947
rect 11379 21913 11388 21947
rect 11336 21904 11388 21913
rect 15108 22040 15160 22092
rect 18052 22040 18104 22092
rect 19708 22040 19760 22092
rect 12440 22015 12492 22024
rect 12440 21981 12449 22015
rect 12449 21981 12483 22015
rect 12483 21981 12492 22015
rect 12440 21972 12492 21981
rect 12992 21972 13044 22024
rect 13268 21904 13320 21956
rect 12348 21836 12400 21888
rect 15936 22015 15988 22024
rect 15936 21981 15945 22015
rect 15945 21981 15979 22015
rect 15979 21981 15988 22015
rect 15936 21972 15988 21981
rect 16672 22015 16724 22024
rect 16672 21981 16706 22015
rect 16706 21981 16724 22015
rect 16672 21972 16724 21981
rect 19800 22015 19852 22024
rect 19800 21981 19809 22015
rect 19809 21981 19843 22015
rect 19843 21981 19852 22015
rect 19800 21972 19852 21981
rect 14556 21904 14608 21956
rect 15292 21947 15344 21956
rect 15292 21913 15301 21947
rect 15301 21913 15335 21947
rect 15335 21913 15344 21947
rect 15292 21904 15344 21913
rect 15568 21947 15620 21956
rect 15568 21913 15577 21947
rect 15577 21913 15611 21947
rect 15611 21913 15620 21947
rect 15568 21904 15620 21913
rect 17960 21904 18012 21956
rect 18972 21904 19024 21956
rect 20352 21904 20404 21956
rect 13728 21836 13780 21888
rect 13912 21836 13964 21888
rect 15016 21879 15068 21888
rect 15016 21845 15049 21879
rect 15049 21845 15068 21879
rect 15016 21836 15068 21845
rect 15384 21836 15436 21888
rect 15752 21879 15804 21888
rect 15752 21845 15761 21879
rect 15761 21845 15795 21879
rect 15795 21845 15804 21879
rect 15752 21836 15804 21845
rect 18052 21879 18104 21888
rect 18052 21845 18085 21879
rect 18085 21845 18104 21879
rect 18052 21836 18104 21845
rect 21088 21836 21140 21888
rect 4220 21734 4272 21786
rect 4284 21734 4336 21786
rect 4348 21734 4400 21786
rect 4412 21734 4464 21786
rect 4476 21734 4528 21786
rect 9441 21734 9493 21786
rect 9505 21734 9557 21786
rect 9569 21734 9621 21786
rect 9633 21734 9685 21786
rect 9697 21734 9749 21786
rect 14662 21734 14714 21786
rect 14726 21734 14778 21786
rect 14790 21734 14842 21786
rect 14854 21734 14906 21786
rect 14918 21734 14970 21786
rect 19883 21734 19935 21786
rect 19947 21734 19999 21786
rect 20011 21734 20063 21786
rect 20075 21734 20127 21786
rect 20139 21734 20191 21786
rect 2964 21675 3016 21684
rect 2964 21641 2973 21675
rect 2973 21641 3007 21675
rect 3007 21641 3016 21675
rect 2964 21632 3016 21641
rect 5264 21632 5316 21684
rect 5724 21675 5776 21684
rect 5724 21641 5733 21675
rect 5733 21641 5767 21675
rect 5767 21641 5776 21675
rect 5724 21632 5776 21641
rect 6000 21632 6052 21684
rect 2780 21564 2832 21616
rect 1676 21539 1728 21548
rect 1676 21505 1710 21539
rect 1710 21505 1728 21539
rect 1676 21496 1728 21505
rect 4068 21564 4120 21616
rect 4804 21564 4856 21616
rect 5356 21564 5408 21616
rect 5540 21564 5592 21616
rect 6644 21564 6696 21616
rect 8392 21564 8444 21616
rect 8944 21632 8996 21684
rect 9404 21632 9456 21684
rect 10968 21632 11020 21684
rect 11244 21675 11296 21684
rect 11244 21641 11253 21675
rect 11253 21641 11287 21675
rect 11287 21641 11296 21675
rect 11244 21632 11296 21641
rect 12256 21632 12308 21684
rect 13084 21632 13136 21684
rect 3056 21360 3108 21412
rect 5816 21496 5868 21548
rect 3884 21471 3936 21480
rect 3884 21437 3893 21471
rect 3893 21437 3927 21471
rect 3927 21437 3936 21471
rect 3884 21428 3936 21437
rect 3976 21428 4028 21480
rect 6552 21496 6604 21548
rect 7380 21428 7432 21480
rect 5356 21360 5408 21412
rect 6828 21360 6880 21412
rect 7012 21360 7064 21412
rect 8300 21496 8352 21548
rect 8484 21539 8536 21548
rect 8484 21505 8518 21539
rect 8518 21505 8536 21539
rect 8484 21496 8536 21505
rect 9312 21496 9364 21548
rect 10784 21564 10836 21616
rect 11152 21564 11204 21616
rect 12348 21564 12400 21616
rect 12440 21564 12492 21616
rect 11336 21496 11388 21548
rect 11704 21496 11756 21548
rect 12716 21539 12768 21548
rect 12716 21505 12725 21539
rect 12725 21505 12759 21539
rect 12759 21505 12768 21539
rect 12716 21496 12768 21505
rect 15108 21564 15160 21616
rect 16120 21632 16172 21684
rect 17040 21632 17092 21684
rect 19616 21675 19668 21684
rect 19616 21641 19625 21675
rect 19625 21641 19659 21675
rect 19659 21641 19668 21675
rect 19616 21632 19668 21641
rect 8116 21428 8168 21480
rect 14832 21539 14884 21548
rect 14832 21505 14866 21539
rect 14866 21505 14884 21539
rect 14832 21496 14884 21505
rect 15660 21496 15712 21548
rect 16764 21496 16816 21548
rect 19800 21564 19852 21616
rect 20628 21564 20680 21616
rect 18512 21539 18564 21548
rect 18512 21505 18546 21539
rect 18546 21505 18564 21539
rect 18512 21496 18564 21505
rect 5264 21292 5316 21344
rect 6092 21292 6144 21344
rect 6368 21292 6420 21344
rect 6920 21292 6972 21344
rect 8024 21292 8076 21344
rect 11612 21403 11664 21412
rect 11612 21369 11621 21403
rect 11621 21369 11655 21403
rect 11655 21369 11664 21403
rect 11612 21360 11664 21369
rect 19800 21471 19852 21480
rect 19800 21437 19809 21471
rect 19809 21437 19843 21471
rect 19843 21437 19852 21471
rect 19800 21428 19852 21437
rect 16396 21360 16448 21412
rect 10876 21292 10928 21344
rect 14464 21292 14516 21344
rect 15292 21292 15344 21344
rect 16028 21292 16080 21344
rect 21180 21335 21232 21344
rect 21180 21301 21189 21335
rect 21189 21301 21223 21335
rect 21223 21301 21232 21335
rect 21180 21292 21232 21301
rect 3560 21190 3612 21242
rect 3624 21190 3676 21242
rect 3688 21190 3740 21242
rect 3752 21190 3804 21242
rect 3816 21190 3868 21242
rect 8781 21190 8833 21242
rect 8845 21190 8897 21242
rect 8909 21190 8961 21242
rect 8973 21190 9025 21242
rect 9037 21190 9089 21242
rect 14002 21190 14054 21242
rect 14066 21190 14118 21242
rect 14130 21190 14182 21242
rect 14194 21190 14246 21242
rect 14258 21190 14310 21242
rect 19223 21190 19275 21242
rect 19287 21190 19339 21242
rect 19351 21190 19403 21242
rect 19415 21190 19467 21242
rect 19479 21190 19531 21242
rect 1952 21020 2004 21072
rect 5632 21088 5684 21140
rect 5816 21088 5868 21140
rect 2872 21020 2924 21072
rect 5540 21020 5592 21072
rect 4620 20952 4672 21004
rect 6000 20952 6052 21004
rect 2412 20816 2464 20868
rect 2688 20859 2740 20868
rect 2688 20825 2697 20859
rect 2697 20825 2731 20859
rect 2731 20825 2740 20859
rect 3884 20884 3936 20936
rect 4896 20884 4948 20936
rect 5448 20927 5500 20936
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 5632 20927 5684 20936
rect 5632 20893 5641 20927
rect 5641 20893 5675 20927
rect 5675 20893 5684 20927
rect 5632 20884 5684 20893
rect 5724 20927 5776 20936
rect 5724 20893 5733 20927
rect 5733 20893 5767 20927
rect 5767 20893 5776 20927
rect 5724 20884 5776 20893
rect 5908 20927 5960 20936
rect 5908 20893 5911 20927
rect 5911 20893 5960 20927
rect 5908 20884 5960 20893
rect 2688 20816 2740 20825
rect 4528 20816 4580 20868
rect 4988 20816 5040 20868
rect 2596 20791 2648 20800
rect 2596 20757 2605 20791
rect 2605 20757 2639 20791
rect 2639 20757 2648 20791
rect 2596 20748 2648 20757
rect 4620 20748 4672 20800
rect 6644 21088 6696 21140
rect 8484 21088 8536 21140
rect 9220 21088 9272 21140
rect 12256 21088 12308 21140
rect 12716 21088 12768 21140
rect 14832 21088 14884 21140
rect 16856 21088 16908 21140
rect 19616 21088 19668 21140
rect 8392 21020 8444 21072
rect 12900 21020 12952 21072
rect 15108 21020 15160 21072
rect 6368 20952 6420 21004
rect 9312 20952 9364 21004
rect 13912 20995 13964 21004
rect 13912 20961 13921 20995
rect 13921 20961 13955 20995
rect 13955 20961 13964 20995
rect 13912 20952 13964 20961
rect 6092 20816 6144 20868
rect 9128 20927 9180 20936
rect 9128 20893 9137 20927
rect 9137 20893 9171 20927
rect 9171 20893 9180 20927
rect 9128 20884 9180 20893
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 11060 20884 11112 20936
rect 11336 20884 11388 20936
rect 13084 20884 13136 20936
rect 14464 20927 14516 20936
rect 14464 20893 14473 20927
rect 14473 20893 14507 20927
rect 14507 20893 14516 20927
rect 14464 20884 14516 20893
rect 6828 20816 6880 20868
rect 9864 20816 9916 20868
rect 6184 20748 6236 20800
rect 8116 20748 8168 20800
rect 10232 20791 10284 20800
rect 10232 20757 10241 20791
rect 10241 20757 10275 20791
rect 10275 20757 10284 20791
rect 10232 20748 10284 20757
rect 13452 20816 13504 20868
rect 15016 20884 15068 20936
rect 10968 20748 11020 20800
rect 13820 20748 13872 20800
rect 15384 20816 15436 20868
rect 15016 20748 15068 20800
rect 15752 20816 15804 20868
rect 17500 20859 17552 20868
rect 17500 20825 17534 20859
rect 17534 20825 17552 20859
rect 17500 20816 17552 20825
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 19800 20884 19852 20936
rect 21272 20884 21324 20936
rect 17868 20748 17920 20800
rect 20628 20791 20680 20800
rect 20628 20757 20637 20791
rect 20637 20757 20671 20791
rect 20671 20757 20680 20791
rect 20628 20748 20680 20757
rect 21456 20748 21508 20800
rect 4220 20646 4272 20698
rect 4284 20646 4336 20698
rect 4348 20646 4400 20698
rect 4412 20646 4464 20698
rect 4476 20646 4528 20698
rect 9441 20646 9493 20698
rect 9505 20646 9557 20698
rect 9569 20646 9621 20698
rect 9633 20646 9685 20698
rect 9697 20646 9749 20698
rect 14662 20646 14714 20698
rect 14726 20646 14778 20698
rect 14790 20646 14842 20698
rect 14854 20646 14906 20698
rect 14918 20646 14970 20698
rect 19883 20646 19935 20698
rect 19947 20646 19999 20698
rect 20011 20646 20063 20698
rect 20075 20646 20127 20698
rect 20139 20646 20191 20698
rect 2780 20476 2832 20528
rect 4160 20544 4212 20596
rect 4620 20544 4672 20596
rect 5172 20544 5224 20596
rect 1676 20451 1728 20460
rect 1676 20417 1710 20451
rect 1710 20417 1728 20451
rect 1676 20408 1728 20417
rect 3976 20476 4028 20528
rect 4712 20519 4764 20528
rect 4712 20485 4721 20519
rect 4721 20485 4755 20519
rect 4755 20485 4764 20519
rect 4712 20476 4764 20485
rect 5356 20519 5408 20528
rect 5356 20485 5365 20519
rect 5365 20485 5399 20519
rect 5399 20485 5408 20519
rect 5356 20476 5408 20485
rect 5632 20544 5684 20596
rect 5908 20587 5960 20596
rect 5908 20553 5917 20587
rect 5917 20553 5951 20587
rect 5951 20553 5960 20587
rect 5908 20544 5960 20553
rect 6552 20544 6604 20596
rect 6644 20587 6696 20596
rect 6644 20553 6653 20587
rect 6653 20553 6687 20587
rect 6687 20553 6696 20587
rect 6644 20544 6696 20553
rect 8668 20587 8720 20596
rect 8668 20553 8677 20587
rect 8677 20553 8711 20587
rect 8711 20553 8720 20587
rect 8668 20544 8720 20553
rect 9312 20544 9364 20596
rect 5540 20476 5592 20528
rect 6092 20476 6144 20528
rect 2688 20272 2740 20324
rect 4896 20408 4948 20460
rect 4620 20383 4672 20392
rect 4620 20349 4629 20383
rect 4629 20349 4663 20383
rect 4663 20349 4672 20383
rect 4620 20340 4672 20349
rect 4988 20340 5040 20392
rect 5632 20451 5684 20460
rect 5632 20417 5641 20451
rect 5641 20417 5675 20451
rect 5675 20417 5684 20451
rect 5632 20408 5684 20417
rect 7748 20451 7800 20460
rect 8300 20476 8352 20528
rect 8392 20476 8444 20528
rect 10048 20476 10100 20528
rect 12072 20476 12124 20528
rect 7748 20417 7766 20451
rect 7766 20417 7800 20451
rect 7748 20408 7800 20417
rect 8668 20408 8720 20460
rect 5908 20340 5960 20392
rect 8208 20340 8260 20392
rect 11796 20408 11848 20460
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 14464 20544 14516 20596
rect 12992 20476 13044 20528
rect 15292 20476 15344 20528
rect 16856 20544 16908 20596
rect 13084 20451 13136 20460
rect 13084 20417 13093 20451
rect 13093 20417 13127 20451
rect 13127 20417 13136 20451
rect 13084 20408 13136 20417
rect 13268 20451 13320 20460
rect 13268 20417 13282 20451
rect 13282 20417 13316 20451
rect 13316 20417 13320 20451
rect 13268 20408 13320 20417
rect 6828 20272 6880 20324
rect 8576 20272 8628 20324
rect 2044 20204 2096 20256
rect 3976 20204 4028 20256
rect 5080 20247 5132 20256
rect 5080 20213 5089 20247
rect 5089 20213 5123 20247
rect 5123 20213 5132 20247
rect 5080 20204 5132 20213
rect 7380 20204 7432 20256
rect 11704 20315 11756 20324
rect 11704 20281 11713 20315
rect 11713 20281 11747 20315
rect 11747 20281 11756 20315
rect 11704 20272 11756 20281
rect 12256 20383 12308 20392
rect 12256 20349 12265 20383
rect 12265 20349 12299 20383
rect 12299 20349 12308 20383
rect 12256 20340 12308 20349
rect 16028 20408 16080 20460
rect 16396 20476 16448 20528
rect 17040 20519 17092 20528
rect 17040 20485 17049 20519
rect 17049 20485 17083 20519
rect 17083 20485 17092 20519
rect 17040 20476 17092 20485
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 18420 20587 18472 20596
rect 18420 20553 18429 20587
rect 18429 20553 18463 20587
rect 18463 20553 18472 20587
rect 18420 20544 18472 20553
rect 20536 20544 20588 20596
rect 18328 20476 18380 20528
rect 20628 20476 20680 20528
rect 14740 20340 14792 20392
rect 16856 20340 16908 20392
rect 13452 20315 13504 20324
rect 13452 20281 13461 20315
rect 13461 20281 13495 20315
rect 13495 20281 13504 20315
rect 13452 20272 13504 20281
rect 14556 20272 14608 20324
rect 15936 20272 15988 20324
rect 16764 20315 16816 20324
rect 16764 20281 16773 20315
rect 16773 20281 16807 20315
rect 16807 20281 16816 20315
rect 16764 20272 16816 20281
rect 17316 20451 17368 20460
rect 17316 20417 17325 20451
rect 17325 20417 17359 20451
rect 17359 20417 17368 20451
rect 17316 20408 17368 20417
rect 18052 20408 18104 20460
rect 18696 20408 18748 20460
rect 19616 20408 19668 20460
rect 20996 20451 21048 20460
rect 20996 20417 21045 20451
rect 21045 20417 21048 20451
rect 20996 20408 21048 20417
rect 21180 20451 21232 20460
rect 21180 20417 21189 20451
rect 21189 20417 21223 20451
rect 21223 20417 21232 20451
rect 21180 20408 21232 20417
rect 21364 20408 21416 20460
rect 21456 20451 21508 20460
rect 21456 20417 21465 20451
rect 21465 20417 21499 20451
rect 21499 20417 21508 20451
rect 21456 20408 21508 20417
rect 17132 20340 17184 20392
rect 18972 20340 19024 20392
rect 19800 20383 19852 20392
rect 19800 20349 19809 20383
rect 19809 20349 19843 20383
rect 19843 20349 19852 20383
rect 19800 20340 19852 20349
rect 18512 20272 18564 20324
rect 18880 20315 18932 20324
rect 18880 20281 18889 20315
rect 18889 20281 18923 20315
rect 18923 20281 18932 20315
rect 18880 20272 18932 20281
rect 9864 20204 9916 20256
rect 12256 20204 12308 20256
rect 12808 20204 12860 20256
rect 13268 20204 13320 20256
rect 17224 20204 17276 20256
rect 20812 20204 20864 20256
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 3560 20102 3612 20154
rect 3624 20102 3676 20154
rect 3688 20102 3740 20154
rect 3752 20102 3804 20154
rect 3816 20102 3868 20154
rect 8781 20102 8833 20154
rect 8845 20102 8897 20154
rect 8909 20102 8961 20154
rect 8973 20102 9025 20154
rect 9037 20102 9089 20154
rect 14002 20102 14054 20154
rect 14066 20102 14118 20154
rect 14130 20102 14182 20154
rect 14194 20102 14246 20154
rect 14258 20102 14310 20154
rect 19223 20102 19275 20154
rect 19287 20102 19339 20154
rect 19351 20102 19403 20154
rect 19415 20102 19467 20154
rect 19479 20102 19531 20154
rect 1676 20000 1728 20052
rect 4160 20000 4212 20052
rect 5632 20000 5684 20052
rect 7748 20043 7800 20052
rect 7748 20009 7757 20043
rect 7757 20009 7791 20043
rect 7791 20009 7800 20043
rect 7748 20000 7800 20009
rect 8208 20000 8260 20052
rect 10600 20000 10652 20052
rect 11796 20000 11848 20052
rect 12440 20000 12492 20052
rect 13452 20000 13504 20052
rect 18420 20000 18472 20052
rect 20352 20000 20404 20052
rect 21180 20000 21232 20052
rect 5356 19932 5408 19984
rect 8392 19932 8444 19984
rect 14464 19932 14516 19984
rect 5448 19864 5500 19916
rect 9772 19864 9824 19916
rect 13912 19864 13964 19916
rect 1952 19839 2004 19848
rect 1952 19805 1961 19839
rect 1961 19805 1995 19839
rect 1995 19805 2004 19839
rect 1952 19796 2004 19805
rect 2780 19796 2832 19848
rect 3976 19839 4028 19848
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 6092 19796 6144 19848
rect 7932 19839 7984 19848
rect 7932 19805 7941 19839
rect 7941 19805 7975 19839
rect 7975 19805 7984 19839
rect 7932 19796 7984 19805
rect 8024 19796 8076 19848
rect 11152 19796 11204 19848
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 12808 19839 12860 19848
rect 12808 19805 12826 19839
rect 12826 19805 12860 19839
rect 12808 19796 12860 19805
rect 2320 19771 2372 19780
rect 2320 19737 2354 19771
rect 2354 19737 2372 19771
rect 2320 19728 2372 19737
rect 5080 19728 5132 19780
rect 7288 19771 7340 19780
rect 7288 19737 7297 19771
rect 7297 19737 7331 19771
rect 7331 19737 7340 19771
rect 7288 19728 7340 19737
rect 8116 19728 8168 19780
rect 9864 19728 9916 19780
rect 10232 19728 10284 19780
rect 13452 19728 13504 19780
rect 14280 19796 14332 19848
rect 3792 19703 3844 19712
rect 3792 19669 3801 19703
rect 3801 19669 3835 19703
rect 3835 19669 3844 19703
rect 3792 19660 3844 19669
rect 5816 19660 5868 19712
rect 7472 19703 7524 19712
rect 7472 19669 7481 19703
rect 7481 19669 7515 19703
rect 7515 19669 7524 19703
rect 7472 19660 7524 19669
rect 9680 19660 9732 19712
rect 9956 19660 10008 19712
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 11612 19660 11664 19712
rect 11796 19660 11848 19712
rect 13820 19771 13872 19780
rect 13820 19737 13829 19771
rect 13829 19737 13863 19771
rect 13863 19737 13872 19771
rect 15568 19864 15620 19916
rect 13820 19728 13872 19737
rect 14740 19771 14792 19780
rect 14740 19737 14749 19771
rect 14749 19737 14783 19771
rect 14783 19737 14792 19771
rect 14740 19728 14792 19737
rect 15200 19796 15252 19848
rect 17040 19932 17092 19984
rect 18144 19864 18196 19916
rect 18328 19864 18380 19916
rect 15476 19728 15528 19780
rect 16212 19728 16264 19780
rect 16764 19771 16816 19780
rect 16764 19737 16773 19771
rect 16773 19737 16807 19771
rect 16807 19737 16816 19771
rect 16764 19728 16816 19737
rect 17408 19796 17460 19848
rect 18052 19839 18104 19848
rect 18052 19805 18061 19839
rect 18061 19805 18095 19839
rect 18095 19805 18104 19839
rect 18052 19796 18104 19805
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 18604 19839 18656 19848
rect 18604 19805 18613 19839
rect 18613 19805 18647 19839
rect 18647 19805 18656 19839
rect 18604 19796 18656 19805
rect 15108 19660 15160 19712
rect 16856 19660 16908 19712
rect 17132 19728 17184 19780
rect 17592 19771 17644 19780
rect 17592 19737 17601 19771
rect 17601 19737 17635 19771
rect 17635 19737 17644 19771
rect 17592 19728 17644 19737
rect 18972 19728 19024 19780
rect 19708 19864 19760 19916
rect 19800 19796 19852 19848
rect 20904 19796 20956 19848
rect 21272 19728 21324 19780
rect 17224 19660 17276 19712
rect 17868 19660 17920 19712
rect 18328 19660 18380 19712
rect 21456 19660 21508 19712
rect 4220 19558 4272 19610
rect 4284 19558 4336 19610
rect 4348 19558 4400 19610
rect 4412 19558 4464 19610
rect 4476 19558 4528 19610
rect 9441 19558 9493 19610
rect 9505 19558 9557 19610
rect 9569 19558 9621 19610
rect 9633 19558 9685 19610
rect 9697 19558 9749 19610
rect 14662 19558 14714 19610
rect 14726 19558 14778 19610
rect 14790 19558 14842 19610
rect 14854 19558 14906 19610
rect 14918 19558 14970 19610
rect 19883 19558 19935 19610
rect 19947 19558 19999 19610
rect 20011 19558 20063 19610
rect 20075 19558 20127 19610
rect 20139 19558 20191 19610
rect 2320 19456 2372 19508
rect 4620 19456 4672 19508
rect 5448 19456 5500 19508
rect 7656 19456 7708 19508
rect 7932 19456 7984 19508
rect 8024 19456 8076 19508
rect 8668 19456 8720 19508
rect 2780 19388 2832 19440
rect 2044 19363 2096 19372
rect 2044 19329 2053 19363
rect 2053 19329 2087 19363
rect 2087 19329 2096 19363
rect 2044 19320 2096 19329
rect 3056 19320 3108 19372
rect 3792 19388 3844 19440
rect 5816 19431 5868 19440
rect 5816 19397 5825 19431
rect 5825 19397 5859 19431
rect 5859 19397 5868 19431
rect 5816 19388 5868 19397
rect 6920 19388 6972 19440
rect 4712 19320 4764 19372
rect 7288 19320 7340 19372
rect 8208 19388 8260 19440
rect 9128 19388 9180 19440
rect 9680 19456 9732 19508
rect 9864 19499 9916 19508
rect 9864 19465 9873 19499
rect 9873 19465 9907 19499
rect 9907 19465 9916 19499
rect 9864 19456 9916 19465
rect 12072 19456 12124 19508
rect 14556 19456 14608 19508
rect 16212 19499 16264 19508
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 17408 19456 17460 19508
rect 19616 19499 19668 19508
rect 19616 19465 19625 19499
rect 19625 19465 19659 19499
rect 19659 19465 19668 19499
rect 19616 19456 19668 19465
rect 21272 19456 21324 19508
rect 8484 19320 8536 19372
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 7472 19295 7524 19304
rect 7472 19261 7481 19295
rect 7481 19261 7515 19295
rect 7515 19261 7524 19295
rect 7472 19252 7524 19261
rect 10692 19320 10744 19372
rect 11612 19320 11664 19372
rect 12348 19320 12400 19372
rect 13912 19388 13964 19440
rect 15108 19431 15160 19440
rect 15108 19397 15142 19431
rect 15142 19397 15160 19431
rect 15108 19388 15160 19397
rect 13544 19363 13596 19372
rect 13544 19329 13578 19363
rect 13578 19329 13596 19363
rect 13544 19320 13596 19329
rect 16948 19363 17000 19372
rect 16948 19329 16982 19363
rect 16982 19329 17000 19363
rect 16948 19320 17000 19329
rect 18328 19320 18380 19372
rect 19800 19363 19852 19372
rect 19800 19329 19809 19363
rect 19809 19329 19843 19363
rect 19843 19329 19852 19363
rect 19800 19320 19852 19329
rect 21456 19320 21508 19372
rect 8300 19184 8352 19236
rect 6000 19116 6052 19168
rect 6828 19116 6880 19168
rect 7104 19116 7156 19168
rect 9680 19116 9732 19168
rect 10876 19116 10928 19168
rect 11796 19116 11848 19168
rect 15016 19116 15068 19168
rect 18512 19116 18564 19168
rect 20996 19116 21048 19168
rect 3560 19014 3612 19066
rect 3624 19014 3676 19066
rect 3688 19014 3740 19066
rect 3752 19014 3804 19066
rect 3816 19014 3868 19066
rect 8781 19014 8833 19066
rect 8845 19014 8897 19066
rect 8909 19014 8961 19066
rect 8973 19014 9025 19066
rect 9037 19014 9089 19066
rect 14002 19014 14054 19066
rect 14066 19014 14118 19066
rect 14130 19014 14182 19066
rect 14194 19014 14246 19066
rect 14258 19014 14310 19066
rect 19223 19014 19275 19066
rect 19287 19014 19339 19066
rect 19351 19014 19403 19066
rect 19415 19014 19467 19066
rect 19479 19014 19531 19066
rect 1308 18912 1360 18964
rect 4712 18955 4764 18964
rect 4712 18921 4721 18955
rect 4721 18921 4755 18955
rect 4755 18921 4764 18955
rect 4712 18912 4764 18921
rect 7472 18912 7524 18964
rect 10692 18955 10744 18964
rect 10692 18921 10701 18955
rect 10701 18921 10735 18955
rect 10735 18921 10744 18955
rect 10692 18912 10744 18921
rect 14372 18912 14424 18964
rect 15200 18955 15252 18964
rect 15200 18921 15209 18955
rect 15209 18921 15243 18955
rect 15243 18921 15252 18955
rect 15200 18912 15252 18921
rect 17592 18955 17644 18964
rect 17592 18921 17601 18955
rect 17601 18921 17635 18955
rect 17635 18921 17644 18955
rect 17592 18912 17644 18921
rect 18052 18912 18104 18964
rect 2504 18844 2556 18896
rect 8300 18844 8352 18896
rect 2688 18776 2740 18828
rect 4620 18776 4672 18828
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 2780 18708 2832 18760
rect 5540 18708 5592 18760
rect 7104 18708 7156 18760
rect 8392 18708 8444 18760
rect 10140 18708 10192 18760
rect 14280 18844 14332 18896
rect 14740 18844 14792 18896
rect 16120 18887 16172 18896
rect 16120 18853 16129 18887
rect 16129 18853 16163 18887
rect 16163 18853 16172 18887
rect 16120 18844 16172 18853
rect 12348 18819 12400 18828
rect 12348 18785 12357 18819
rect 12357 18785 12391 18819
rect 12391 18785 12400 18819
rect 12348 18776 12400 18785
rect 13912 18776 13964 18828
rect 19616 18912 19668 18964
rect 20628 18955 20680 18964
rect 20628 18921 20637 18955
rect 20637 18921 20671 18955
rect 20671 18921 20680 18955
rect 20628 18912 20680 18921
rect 20996 18912 21048 18964
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 17040 18708 17092 18760
rect 1492 18640 1544 18692
rect 4896 18640 4948 18692
rect 5080 18640 5132 18692
rect 6184 18640 6236 18692
rect 3240 18572 3292 18624
rect 8576 18572 8628 18624
rect 11520 18683 11572 18692
rect 11520 18649 11529 18683
rect 11529 18649 11563 18683
rect 11563 18649 11572 18683
rect 11520 18640 11572 18649
rect 12440 18640 12492 18692
rect 12716 18640 12768 18692
rect 15016 18683 15068 18692
rect 15016 18649 15025 18683
rect 15025 18649 15059 18683
rect 15059 18649 15068 18683
rect 15016 18640 15068 18649
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 11152 18572 11204 18624
rect 11612 18572 11664 18624
rect 15660 18615 15712 18624
rect 15660 18581 15669 18615
rect 15669 18581 15703 18615
rect 15703 18581 15712 18615
rect 15660 18572 15712 18581
rect 16120 18640 16172 18692
rect 16672 18640 16724 18692
rect 19800 18708 19852 18760
rect 18880 18640 18932 18692
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 20628 18640 20680 18692
rect 21180 18708 21232 18760
rect 21364 18640 21416 18692
rect 17132 18572 17184 18624
rect 17868 18572 17920 18624
rect 18420 18572 18472 18624
rect 4220 18470 4272 18522
rect 4284 18470 4336 18522
rect 4348 18470 4400 18522
rect 4412 18470 4464 18522
rect 4476 18470 4528 18522
rect 9441 18470 9493 18522
rect 9505 18470 9557 18522
rect 9569 18470 9621 18522
rect 9633 18470 9685 18522
rect 9697 18470 9749 18522
rect 14662 18470 14714 18522
rect 14726 18470 14778 18522
rect 14790 18470 14842 18522
rect 14854 18470 14906 18522
rect 14918 18470 14970 18522
rect 19883 18470 19935 18522
rect 19947 18470 19999 18522
rect 20011 18470 20063 18522
rect 20075 18470 20127 18522
rect 20139 18470 20191 18522
rect 1492 18411 1544 18420
rect 1492 18377 1501 18411
rect 1501 18377 1535 18411
rect 1535 18377 1544 18411
rect 1492 18368 1544 18377
rect 2688 18411 2740 18420
rect 2688 18377 2697 18411
rect 2697 18377 2731 18411
rect 2731 18377 2740 18411
rect 2688 18368 2740 18377
rect 4344 18411 4396 18420
rect 4344 18377 4353 18411
rect 4353 18377 4387 18411
rect 4387 18377 4396 18411
rect 4344 18368 4396 18377
rect 1308 18300 1360 18352
rect 2780 18300 2832 18352
rect 7656 18368 7708 18420
rect 9956 18368 10008 18420
rect 10876 18368 10928 18420
rect 11152 18368 11204 18420
rect 12716 18411 12768 18420
rect 12716 18377 12725 18411
rect 12725 18377 12759 18411
rect 12759 18377 12768 18411
rect 12716 18368 12768 18377
rect 13544 18368 13596 18420
rect 14556 18368 14608 18420
rect 15660 18368 15712 18420
rect 2504 18232 2556 18284
rect 3976 18232 4028 18284
rect 10324 18300 10376 18352
rect 12440 18300 12492 18352
rect 13176 18300 13228 18352
rect 14372 18300 14424 18352
rect 14464 18343 14516 18352
rect 14464 18309 14473 18343
rect 14473 18309 14507 18343
rect 14507 18309 14516 18343
rect 14464 18300 14516 18309
rect 5632 18232 5684 18284
rect 6000 18275 6052 18284
rect 6000 18241 6009 18275
rect 6009 18241 6043 18275
rect 6043 18241 6052 18275
rect 6000 18232 6052 18241
rect 8300 18232 8352 18284
rect 8576 18232 8628 18284
rect 10600 18232 10652 18284
rect 11612 18232 11664 18284
rect 11796 18232 11848 18284
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 2412 18207 2464 18216
rect 2412 18173 2421 18207
rect 2421 18173 2455 18207
rect 2455 18173 2464 18207
rect 2412 18164 2464 18173
rect 12072 18207 12124 18216
rect 12072 18173 12081 18207
rect 12081 18173 12115 18207
rect 12115 18173 12124 18207
rect 12072 18164 12124 18173
rect 13820 18232 13872 18284
rect 15108 18275 15160 18284
rect 15108 18241 15117 18275
rect 15117 18241 15151 18275
rect 15151 18241 15160 18275
rect 15108 18232 15160 18241
rect 16672 18300 16724 18352
rect 17592 18368 17644 18420
rect 19708 18368 19760 18420
rect 18144 18343 18196 18352
rect 18144 18309 18153 18343
rect 18153 18309 18187 18343
rect 18187 18309 18196 18343
rect 18144 18300 18196 18309
rect 21272 18300 21324 18352
rect 17960 18275 18012 18284
rect 17960 18241 17969 18275
rect 17969 18241 18003 18275
rect 18003 18241 18012 18275
rect 17960 18232 18012 18241
rect 18512 18232 18564 18284
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 10140 18139 10192 18148
rect 10140 18105 10149 18139
rect 10149 18105 10183 18139
rect 10183 18105 10192 18139
rect 10140 18096 10192 18105
rect 11244 18096 11296 18148
rect 6736 18028 6788 18080
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 13176 18028 13228 18080
rect 17316 18207 17368 18216
rect 17316 18173 17325 18207
rect 17325 18173 17359 18207
rect 17359 18173 17368 18207
rect 17316 18164 17368 18173
rect 19064 18164 19116 18216
rect 20352 18207 20404 18216
rect 20352 18173 20361 18207
rect 20361 18173 20395 18207
rect 20395 18173 20404 18207
rect 20352 18164 20404 18173
rect 20996 18207 21048 18216
rect 20996 18173 21005 18207
rect 21005 18173 21039 18207
rect 21039 18173 21048 18207
rect 20996 18164 21048 18173
rect 16764 18139 16816 18148
rect 16764 18105 16773 18139
rect 16773 18105 16807 18139
rect 16807 18105 16816 18139
rect 16764 18096 16816 18105
rect 20444 18096 20496 18148
rect 14372 18028 14424 18080
rect 19616 18028 19668 18080
rect 21640 18071 21692 18080
rect 21640 18037 21649 18071
rect 21649 18037 21683 18071
rect 21683 18037 21692 18071
rect 21640 18028 21692 18037
rect 3560 17926 3612 17978
rect 3624 17926 3676 17978
rect 3688 17926 3740 17978
rect 3752 17926 3804 17978
rect 3816 17926 3868 17978
rect 8781 17926 8833 17978
rect 8845 17926 8897 17978
rect 8909 17926 8961 17978
rect 8973 17926 9025 17978
rect 9037 17926 9089 17978
rect 14002 17926 14054 17978
rect 14066 17926 14118 17978
rect 14130 17926 14182 17978
rect 14194 17926 14246 17978
rect 14258 17926 14310 17978
rect 19223 17926 19275 17978
rect 19287 17926 19339 17978
rect 19351 17926 19403 17978
rect 19415 17926 19467 17978
rect 19479 17926 19531 17978
rect 3240 17867 3292 17876
rect 3240 17833 3249 17867
rect 3249 17833 3283 17867
rect 3283 17833 3292 17867
rect 3240 17824 3292 17833
rect 3976 17824 4028 17876
rect 4344 17824 4396 17876
rect 5632 17824 5684 17876
rect 6184 17824 6236 17876
rect 9772 17824 9824 17876
rect 12532 17824 12584 17876
rect 12992 17824 13044 17876
rect 17960 17824 18012 17876
rect 1860 17663 1912 17672
rect 1860 17629 1869 17663
rect 1869 17629 1903 17663
rect 1903 17629 1912 17663
rect 1860 17620 1912 17629
rect 5816 17756 5868 17808
rect 6552 17756 6604 17808
rect 6828 17756 6880 17808
rect 4620 17688 4672 17740
rect 6000 17688 6052 17740
rect 6920 17688 6972 17740
rect 8484 17799 8536 17808
rect 8484 17765 8493 17799
rect 8493 17765 8527 17799
rect 8527 17765 8536 17799
rect 8484 17756 8536 17765
rect 10784 17688 10836 17740
rect 1952 17552 2004 17604
rect 2872 17552 2924 17604
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 5724 17663 5776 17672
rect 5724 17629 5733 17663
rect 5733 17629 5767 17663
rect 5767 17629 5776 17663
rect 5724 17620 5776 17629
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 5908 17663 5960 17672
rect 5908 17629 5922 17663
rect 5922 17629 5956 17663
rect 5956 17629 5960 17663
rect 5908 17620 5960 17629
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 4988 17552 5040 17604
rect 8668 17620 8720 17672
rect 9864 17620 9916 17672
rect 11520 17756 11572 17808
rect 13084 17756 13136 17808
rect 15200 17799 15252 17808
rect 15200 17765 15209 17799
rect 15209 17765 15243 17799
rect 15243 17765 15252 17799
rect 15200 17756 15252 17765
rect 15844 17756 15896 17808
rect 11336 17731 11388 17740
rect 11336 17697 11345 17731
rect 11345 17697 11379 17731
rect 11379 17697 11388 17731
rect 11336 17688 11388 17697
rect 13820 17688 13872 17740
rect 13636 17620 13688 17672
rect 4712 17484 4764 17536
rect 6920 17595 6972 17604
rect 6920 17561 6929 17595
rect 6929 17561 6963 17595
rect 6963 17561 6972 17595
rect 6920 17552 6972 17561
rect 5356 17484 5408 17536
rect 5540 17484 5592 17536
rect 8208 17552 8260 17604
rect 8116 17484 8168 17536
rect 10324 17484 10376 17536
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 11428 17552 11480 17604
rect 12716 17552 12768 17604
rect 13084 17552 13136 17604
rect 13452 17595 13504 17604
rect 13452 17561 13461 17595
rect 13461 17561 13495 17595
rect 13495 17561 13504 17595
rect 13452 17552 13504 17561
rect 15016 17595 15068 17604
rect 15016 17561 15025 17595
rect 15025 17561 15059 17595
rect 15059 17561 15068 17595
rect 15016 17552 15068 17561
rect 15476 17595 15528 17604
rect 15476 17561 15485 17595
rect 15485 17561 15519 17595
rect 15519 17561 15528 17595
rect 15476 17552 15528 17561
rect 15568 17595 15620 17604
rect 15568 17561 15577 17595
rect 15577 17561 15611 17595
rect 15611 17561 15620 17595
rect 15568 17552 15620 17561
rect 15660 17552 15712 17604
rect 16672 17620 16724 17672
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 17224 17620 17276 17672
rect 20536 17824 20588 17876
rect 21548 17867 21600 17876
rect 21548 17833 21557 17867
rect 21557 17833 21591 17867
rect 21591 17833 21600 17867
rect 21548 17824 21600 17833
rect 18604 17756 18656 17808
rect 18880 17688 18932 17740
rect 19800 17688 19852 17740
rect 18512 17620 18564 17672
rect 18972 17620 19024 17672
rect 19616 17620 19668 17672
rect 20996 17620 21048 17672
rect 12256 17484 12308 17536
rect 12532 17484 12584 17536
rect 13176 17484 13228 17536
rect 13544 17484 13596 17536
rect 13728 17484 13780 17536
rect 16580 17527 16632 17536
rect 16580 17493 16589 17527
rect 16589 17493 16623 17527
rect 16623 17493 16632 17527
rect 16580 17484 16632 17493
rect 16948 17484 17000 17536
rect 18144 17552 18196 17604
rect 21088 17552 21140 17604
rect 19800 17484 19852 17536
rect 20260 17484 20312 17536
rect 4220 17382 4272 17434
rect 4284 17382 4336 17434
rect 4348 17382 4400 17434
rect 4412 17382 4464 17434
rect 4476 17382 4528 17434
rect 9441 17382 9493 17434
rect 9505 17382 9557 17434
rect 9569 17382 9621 17434
rect 9633 17382 9685 17434
rect 9697 17382 9749 17434
rect 14662 17382 14714 17434
rect 14726 17382 14778 17434
rect 14790 17382 14842 17434
rect 14854 17382 14906 17434
rect 14918 17382 14970 17434
rect 19883 17382 19935 17434
rect 19947 17382 19999 17434
rect 20011 17382 20063 17434
rect 20075 17382 20127 17434
rect 20139 17382 20191 17434
rect 1860 17280 1912 17332
rect 2688 17280 2740 17332
rect 2872 17212 2924 17264
rect 3056 17255 3108 17264
rect 3056 17221 3065 17255
rect 3065 17221 3099 17255
rect 3099 17221 3108 17255
rect 3056 17212 3108 17221
rect 6460 17280 6512 17332
rect 6920 17280 6972 17332
rect 1952 17051 2004 17060
rect 1952 17017 1961 17051
rect 1961 17017 1995 17051
rect 1995 17017 2004 17051
rect 1952 17008 2004 17017
rect 3240 17144 3292 17196
rect 4896 17212 4948 17264
rect 6000 17212 6052 17264
rect 8208 17280 8260 17332
rect 7932 17212 7984 17264
rect 8024 17255 8076 17264
rect 8024 17221 8033 17255
rect 8033 17221 8067 17255
rect 8067 17221 8076 17255
rect 8024 17212 8076 17221
rect 10508 17212 10560 17264
rect 11428 17280 11480 17332
rect 11796 17280 11848 17332
rect 13360 17280 13412 17332
rect 13452 17280 13504 17332
rect 15476 17280 15528 17332
rect 17960 17280 18012 17332
rect 18972 17280 19024 17332
rect 19708 17280 19760 17332
rect 20168 17280 20220 17332
rect 21272 17280 21324 17332
rect 11704 17212 11756 17264
rect 4068 17076 4120 17128
rect 4712 17076 4764 17128
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 5908 17144 5960 17196
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 7840 17144 7892 17196
rect 9588 17144 9640 17196
rect 11796 17144 11848 17196
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 12808 17212 12860 17264
rect 13728 17212 13780 17264
rect 13820 17212 13872 17264
rect 15200 17255 15252 17264
rect 15200 17221 15234 17255
rect 15234 17221 15252 17255
rect 15200 17212 15252 17221
rect 17040 17212 17092 17264
rect 17408 17212 17460 17264
rect 13636 17144 13688 17196
rect 17316 17187 17368 17196
rect 6828 17076 6880 17128
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 8116 17076 8168 17128
rect 9312 17076 9364 17128
rect 11060 17076 11112 17128
rect 11612 17076 11664 17128
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 6276 17008 6328 17060
rect 6552 17008 6604 17060
rect 9588 17008 9640 17060
rect 13544 17008 13596 17060
rect 14648 17119 14700 17128
rect 14648 17085 14657 17119
rect 14657 17085 14691 17119
rect 14691 17085 14700 17119
rect 17316 17153 17325 17187
rect 17325 17153 17359 17187
rect 17359 17153 17368 17187
rect 17316 17144 17368 17153
rect 17960 17144 18012 17196
rect 19064 17212 19116 17264
rect 18604 17144 18656 17196
rect 21456 17212 21508 17264
rect 20260 17144 20312 17196
rect 20444 17187 20496 17196
rect 20444 17153 20478 17187
rect 20478 17153 20496 17187
rect 20444 17144 20496 17153
rect 14648 17076 14700 17085
rect 15936 17076 15988 17128
rect 19064 17076 19116 17128
rect 5540 16940 5592 16992
rect 6460 16940 6512 16992
rect 6920 16983 6972 16992
rect 6920 16949 6929 16983
rect 6929 16949 6963 16983
rect 6963 16949 6972 16983
rect 6920 16940 6972 16949
rect 9680 16940 9732 16992
rect 12256 16940 12308 16992
rect 14464 16940 14516 16992
rect 14556 16940 14608 16992
rect 15660 16940 15712 16992
rect 16764 16983 16816 16992
rect 16764 16949 16773 16983
rect 16773 16949 16807 16983
rect 16807 16949 16816 16983
rect 16764 16940 16816 16949
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 19616 16983 19668 16992
rect 19616 16949 19625 16983
rect 19625 16949 19659 16983
rect 19659 16949 19668 16983
rect 19616 16940 19668 16949
rect 19708 16940 19760 16992
rect 3560 16838 3612 16890
rect 3624 16838 3676 16890
rect 3688 16838 3740 16890
rect 3752 16838 3804 16890
rect 3816 16838 3868 16890
rect 8781 16838 8833 16890
rect 8845 16838 8897 16890
rect 8909 16838 8961 16890
rect 8973 16838 9025 16890
rect 9037 16838 9089 16890
rect 14002 16838 14054 16890
rect 14066 16838 14118 16890
rect 14130 16838 14182 16890
rect 14194 16838 14246 16890
rect 14258 16838 14310 16890
rect 19223 16838 19275 16890
rect 19287 16838 19339 16890
rect 19351 16838 19403 16890
rect 19415 16838 19467 16890
rect 19479 16838 19531 16890
rect 5356 16779 5408 16788
rect 5356 16745 5365 16779
rect 5365 16745 5399 16779
rect 5399 16745 5408 16779
rect 5356 16736 5408 16745
rect 6552 16736 6604 16788
rect 4068 16600 4120 16652
rect 2688 16532 2740 16584
rect 1676 16507 1728 16516
rect 1676 16473 1710 16507
rect 1710 16473 1728 16507
rect 1676 16464 1728 16473
rect 2780 16439 2832 16448
rect 2780 16405 2789 16439
rect 2789 16405 2823 16439
rect 2823 16405 2832 16439
rect 2780 16396 2832 16405
rect 2964 16439 3016 16448
rect 2964 16405 2973 16439
rect 2973 16405 3007 16439
rect 3007 16405 3016 16439
rect 2964 16396 3016 16405
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 3884 16532 3936 16584
rect 4620 16600 4672 16652
rect 4712 16600 4764 16652
rect 5632 16600 5684 16652
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 9312 16736 9364 16788
rect 9588 16736 9640 16788
rect 7932 16668 7984 16720
rect 8392 16668 8444 16720
rect 11520 16736 11572 16788
rect 11888 16736 11940 16788
rect 13820 16779 13872 16788
rect 13820 16745 13829 16779
rect 13829 16745 13863 16779
rect 13863 16745 13872 16779
rect 13820 16736 13872 16745
rect 6736 16600 6788 16609
rect 9312 16600 9364 16652
rect 15660 16668 15712 16720
rect 20536 16736 20588 16788
rect 17408 16643 17460 16652
rect 17408 16609 17417 16643
rect 17417 16609 17451 16643
rect 17451 16609 17460 16643
rect 17408 16600 17460 16609
rect 19064 16600 19116 16652
rect 21456 16779 21508 16788
rect 21456 16745 21465 16779
rect 21465 16745 21499 16779
rect 21499 16745 21508 16779
rect 21456 16736 21508 16745
rect 6460 16575 6512 16584
rect 6460 16541 6478 16575
rect 6478 16541 6512 16575
rect 6460 16532 6512 16541
rect 6920 16532 6972 16584
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 8668 16532 8720 16584
rect 9680 16532 9732 16584
rect 4712 16396 4764 16448
rect 8944 16396 8996 16448
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 13636 16532 13688 16584
rect 14372 16575 14424 16584
rect 14372 16541 14406 16575
rect 14406 16541 14424 16575
rect 14372 16532 14424 16541
rect 16580 16532 16632 16584
rect 17684 16575 17736 16584
rect 17684 16541 17718 16575
rect 17718 16541 17736 16575
rect 17684 16532 17736 16541
rect 19340 16532 19392 16584
rect 9956 16507 10008 16516
rect 9956 16473 9965 16507
rect 9965 16473 9999 16507
rect 9999 16473 10008 16507
rect 9956 16464 10008 16473
rect 18880 16464 18932 16516
rect 19616 16464 19668 16516
rect 16580 16396 16632 16448
rect 17224 16439 17276 16448
rect 17224 16405 17233 16439
rect 17233 16405 17267 16439
rect 17267 16405 17276 16439
rect 17224 16396 17276 16405
rect 18604 16396 18656 16448
rect 20352 16396 20404 16448
rect 20904 16396 20956 16448
rect 4220 16294 4272 16346
rect 4284 16294 4336 16346
rect 4348 16294 4400 16346
rect 4412 16294 4464 16346
rect 4476 16294 4528 16346
rect 9441 16294 9493 16346
rect 9505 16294 9557 16346
rect 9569 16294 9621 16346
rect 9633 16294 9685 16346
rect 9697 16294 9749 16346
rect 14662 16294 14714 16346
rect 14726 16294 14778 16346
rect 14790 16294 14842 16346
rect 14854 16294 14906 16346
rect 14918 16294 14970 16346
rect 19883 16294 19935 16346
rect 19947 16294 19999 16346
rect 20011 16294 20063 16346
rect 20075 16294 20127 16346
rect 20139 16294 20191 16346
rect 1676 16235 1728 16244
rect 1676 16201 1685 16235
rect 1685 16201 1719 16235
rect 1719 16201 1728 16235
rect 1676 16192 1728 16201
rect 2780 16192 2832 16244
rect 4252 16192 4304 16244
rect 4804 16192 4856 16244
rect 7564 16192 7616 16244
rect 8484 16235 8536 16244
rect 8484 16201 8493 16235
rect 8493 16201 8527 16235
rect 8527 16201 8536 16235
rect 8484 16192 8536 16201
rect 9864 16192 9916 16244
rect 3424 16124 3476 16176
rect 5540 16167 5592 16176
rect 5540 16133 5558 16167
rect 5558 16133 5592 16167
rect 5540 16124 5592 16133
rect 2872 16056 2924 16108
rect 5724 16056 5776 16108
rect 5908 16099 5960 16108
rect 5908 16065 5917 16099
rect 5917 16065 5951 16099
rect 5951 16065 5960 16099
rect 5908 16056 5960 16065
rect 6736 16124 6788 16176
rect 7932 16124 7984 16176
rect 9312 16124 9364 16176
rect 11888 16192 11940 16244
rect 2412 15988 2464 16040
rect 2688 15988 2740 16040
rect 9036 16056 9088 16108
rect 12256 16124 12308 16176
rect 13452 16167 13504 16176
rect 13452 16133 13461 16167
rect 13461 16133 13495 16167
rect 13495 16133 13504 16167
rect 13452 16124 13504 16133
rect 15844 16167 15896 16176
rect 15844 16133 15853 16167
rect 15853 16133 15887 16167
rect 15887 16133 15896 16167
rect 15844 16124 15896 16133
rect 16764 16192 16816 16244
rect 20996 16192 21048 16244
rect 12072 16056 12124 16108
rect 4804 15920 4856 15972
rect 7840 15920 7892 15972
rect 4896 15852 4948 15904
rect 11336 15920 11388 15972
rect 13084 16056 13136 16108
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 16580 16056 16632 16108
rect 17224 16124 17276 16176
rect 17408 16124 17460 16176
rect 18604 16167 18656 16176
rect 18604 16133 18613 16167
rect 18613 16133 18647 16167
rect 18647 16133 18656 16167
rect 18604 16124 18656 16133
rect 16948 16099 17000 16108
rect 16948 16065 16982 16099
rect 16982 16065 17000 16099
rect 16948 16056 17000 16065
rect 18052 16056 18104 16108
rect 19340 16056 19392 16108
rect 19800 16124 19852 16176
rect 21548 16124 21600 16176
rect 19524 16056 19576 16108
rect 21180 16099 21232 16108
rect 21180 16065 21229 16099
rect 21229 16065 21232 16099
rect 21180 16056 21232 16065
rect 21456 16099 21508 16108
rect 21456 16065 21465 16099
rect 21465 16065 21499 16099
rect 21499 16065 21508 16099
rect 21456 16056 21508 16065
rect 21640 16099 21692 16108
rect 21640 16065 21649 16099
rect 21649 16065 21683 16099
rect 21683 16065 21692 16099
rect 21640 16056 21692 16065
rect 10876 15852 10928 15904
rect 11060 15852 11112 15904
rect 11704 15852 11756 15904
rect 13636 15988 13688 16040
rect 18880 16031 18932 16040
rect 18880 15997 18889 16031
rect 18889 15997 18923 16031
rect 18923 15997 18932 16031
rect 18880 15988 18932 15997
rect 15936 15920 15988 15972
rect 16672 15920 16724 15972
rect 17960 15920 18012 15972
rect 21088 15963 21140 15972
rect 21088 15929 21097 15963
rect 21097 15929 21131 15963
rect 21131 15929 21140 15963
rect 21088 15920 21140 15929
rect 14464 15852 14516 15904
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 17040 15852 17092 15904
rect 3560 15750 3612 15802
rect 3624 15750 3676 15802
rect 3688 15750 3740 15802
rect 3752 15750 3804 15802
rect 3816 15750 3868 15802
rect 8781 15750 8833 15802
rect 8845 15750 8897 15802
rect 8909 15750 8961 15802
rect 8973 15750 9025 15802
rect 9037 15750 9089 15802
rect 14002 15750 14054 15802
rect 14066 15750 14118 15802
rect 14130 15750 14182 15802
rect 14194 15750 14246 15802
rect 14258 15750 14310 15802
rect 19223 15750 19275 15802
rect 19287 15750 19339 15802
rect 19351 15750 19403 15802
rect 19415 15750 19467 15802
rect 19479 15750 19531 15802
rect 3884 15691 3936 15700
rect 3884 15657 3893 15691
rect 3893 15657 3927 15691
rect 3927 15657 3936 15691
rect 3884 15648 3936 15657
rect 5908 15648 5960 15700
rect 4620 15580 4672 15632
rect 4252 15555 4304 15564
rect 4252 15521 4261 15555
rect 4261 15521 4295 15555
rect 4295 15521 4304 15555
rect 4252 15512 4304 15521
rect 4988 15512 5040 15564
rect 5632 15512 5684 15564
rect 2688 15444 2740 15496
rect 6000 15444 6052 15496
rect 2964 15376 3016 15428
rect 4712 15376 4764 15428
rect 8484 15648 8536 15700
rect 9956 15648 10008 15700
rect 10508 15648 10560 15700
rect 10600 15648 10652 15700
rect 12164 15648 12216 15700
rect 15108 15648 15160 15700
rect 16856 15648 16908 15700
rect 7564 15444 7616 15496
rect 8668 15444 8720 15496
rect 10968 15580 11020 15632
rect 13820 15512 13872 15564
rect 15660 15580 15712 15632
rect 18880 15580 18932 15632
rect 20260 15580 20312 15632
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 17040 15555 17092 15564
rect 17040 15521 17049 15555
rect 17049 15521 17083 15555
rect 17083 15521 17092 15555
rect 17040 15512 17092 15521
rect 17132 15555 17184 15564
rect 17132 15521 17141 15555
rect 17141 15521 17175 15555
rect 17175 15521 17184 15555
rect 17132 15512 17184 15521
rect 21548 15512 21600 15564
rect 4988 15308 5040 15360
rect 10048 15376 10100 15428
rect 11244 15444 11296 15496
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 13360 15444 13412 15496
rect 15936 15487 15988 15496
rect 10600 15419 10652 15428
rect 10600 15385 10609 15419
rect 10609 15385 10643 15419
rect 10643 15385 10652 15419
rect 10600 15376 10652 15385
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 18236 15444 18288 15496
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 10232 15351 10284 15360
rect 10232 15317 10266 15351
rect 10266 15317 10284 15351
rect 10232 15308 10284 15317
rect 10508 15308 10560 15360
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 12808 15308 12860 15360
rect 13452 15308 13504 15360
rect 18052 15376 18104 15428
rect 21456 15376 21508 15428
rect 17684 15351 17736 15360
rect 17684 15317 17693 15351
rect 17693 15317 17727 15351
rect 17727 15317 17736 15351
rect 17684 15308 17736 15317
rect 21180 15351 21232 15360
rect 21180 15317 21189 15351
rect 21189 15317 21223 15351
rect 21223 15317 21232 15351
rect 21180 15308 21232 15317
rect 4220 15206 4272 15258
rect 4284 15206 4336 15258
rect 4348 15206 4400 15258
rect 4412 15206 4464 15258
rect 4476 15206 4528 15258
rect 9441 15206 9493 15258
rect 9505 15206 9557 15258
rect 9569 15206 9621 15258
rect 9633 15206 9685 15258
rect 9697 15206 9749 15258
rect 14662 15206 14714 15258
rect 14726 15206 14778 15258
rect 14790 15206 14842 15258
rect 14854 15206 14906 15258
rect 14918 15206 14970 15258
rect 19883 15206 19935 15258
rect 19947 15206 19999 15258
rect 20011 15206 20063 15258
rect 20075 15206 20127 15258
rect 20139 15206 20191 15258
rect 4620 15104 4672 15156
rect 4068 15036 4120 15088
rect 3424 14968 3476 15020
rect 9312 15104 9364 15156
rect 15476 15104 15528 15156
rect 9036 15036 9088 15088
rect 10232 15036 10284 15088
rect 10508 15079 10560 15088
rect 10508 15045 10517 15079
rect 10517 15045 10551 15079
rect 10551 15045 10560 15079
rect 10508 15036 10560 15045
rect 10876 15079 10928 15088
rect 10876 15045 10885 15079
rect 10885 15045 10919 15079
rect 10919 15045 10928 15079
rect 10876 15036 10928 15045
rect 11244 15079 11296 15088
rect 11244 15045 11253 15079
rect 11253 15045 11287 15079
rect 11287 15045 11296 15079
rect 11244 15036 11296 15045
rect 12072 15079 12124 15088
rect 12072 15045 12081 15079
rect 12081 15045 12115 15079
rect 12115 15045 12124 15079
rect 12072 15036 12124 15045
rect 11980 14968 12032 15020
rect 15844 15036 15896 15088
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 17960 15036 18012 15088
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 17316 14968 17368 15020
rect 5080 14900 5132 14952
rect 5356 14900 5408 14952
rect 7748 14900 7800 14952
rect 12624 14900 12676 14952
rect 13544 14900 13596 14952
rect 16580 14900 16632 14952
rect 2872 14832 2924 14884
rect 2964 14807 3016 14816
rect 2964 14773 2973 14807
rect 2973 14773 3007 14807
rect 3007 14773 3016 14807
rect 2964 14764 3016 14773
rect 5816 14764 5868 14816
rect 10692 14832 10744 14884
rect 11612 14875 11664 14884
rect 11612 14841 11621 14875
rect 11621 14841 11655 14875
rect 11655 14841 11664 14875
rect 11612 14832 11664 14841
rect 14740 14832 14792 14884
rect 20260 14968 20312 15020
rect 19800 14900 19852 14952
rect 19892 14832 19944 14884
rect 10416 14764 10468 14816
rect 10600 14764 10652 14816
rect 12992 14807 13044 14816
rect 12992 14773 13001 14807
rect 13001 14773 13035 14807
rect 13035 14773 13044 14807
rect 12992 14764 13044 14773
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 18604 14807 18656 14816
rect 18604 14773 18613 14807
rect 18613 14773 18647 14807
rect 18647 14773 18656 14807
rect 18604 14764 18656 14773
rect 19616 14764 19668 14816
rect 21548 14807 21600 14816
rect 21548 14773 21557 14807
rect 21557 14773 21591 14807
rect 21591 14773 21600 14807
rect 21548 14764 21600 14773
rect 3560 14662 3612 14714
rect 3624 14662 3676 14714
rect 3688 14662 3740 14714
rect 3752 14662 3804 14714
rect 3816 14662 3868 14714
rect 8781 14662 8833 14714
rect 8845 14662 8897 14714
rect 8909 14662 8961 14714
rect 8973 14662 9025 14714
rect 9037 14662 9089 14714
rect 14002 14662 14054 14714
rect 14066 14662 14118 14714
rect 14130 14662 14182 14714
rect 14194 14662 14246 14714
rect 14258 14662 14310 14714
rect 19223 14662 19275 14714
rect 19287 14662 19339 14714
rect 19351 14662 19403 14714
rect 19415 14662 19467 14714
rect 19479 14662 19531 14714
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 2596 14424 2648 14476
rect 3332 14424 3384 14476
rect 5080 14492 5132 14544
rect 5632 14492 5684 14544
rect 7656 14560 7708 14612
rect 10324 14560 10376 14612
rect 10600 14560 10652 14612
rect 11980 14603 12032 14612
rect 11980 14569 11989 14603
rect 11989 14569 12023 14603
rect 12023 14569 12032 14603
rect 11980 14560 12032 14569
rect 12900 14560 12952 14612
rect 16028 14560 16080 14612
rect 16580 14560 16632 14612
rect 2964 14356 3016 14408
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4988 14424 5040 14476
rect 1584 14288 1636 14340
rect 3240 14288 3292 14340
rect 2872 14220 2924 14272
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 4620 14356 4672 14408
rect 5172 14356 5224 14408
rect 5540 14356 5592 14408
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 7748 14467 7800 14476
rect 7748 14433 7757 14467
rect 7757 14433 7791 14467
rect 7791 14433 7800 14467
rect 7748 14424 7800 14433
rect 10416 14492 10468 14544
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 18236 14603 18288 14612
rect 18236 14569 18245 14603
rect 18245 14569 18279 14603
rect 18279 14569 18288 14603
rect 18236 14560 18288 14569
rect 19524 14560 19576 14612
rect 19892 14560 19944 14612
rect 9312 14424 9364 14476
rect 13636 14424 13688 14476
rect 14372 14424 14424 14476
rect 21364 14467 21416 14476
rect 21364 14433 21373 14467
rect 21373 14433 21407 14467
rect 21407 14433 21416 14467
rect 21364 14424 21416 14433
rect 21456 14467 21508 14476
rect 21456 14433 21465 14467
rect 21465 14433 21499 14467
rect 21499 14433 21508 14467
rect 21456 14424 21508 14433
rect 4712 14288 4764 14340
rect 5264 14288 5316 14340
rect 6828 14288 6880 14340
rect 11428 14356 11480 14408
rect 12256 14356 12308 14408
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15292 14399 15344 14408
rect 15292 14365 15326 14399
rect 15326 14365 15344 14399
rect 15292 14356 15344 14365
rect 17224 14356 17276 14408
rect 18696 14356 18748 14408
rect 4896 14220 4948 14272
rect 6000 14220 6052 14272
rect 7012 14220 7064 14272
rect 7840 14220 7892 14272
rect 9220 14288 9272 14340
rect 10232 14331 10284 14340
rect 10232 14297 10241 14331
rect 10241 14297 10275 14331
rect 10275 14297 10284 14331
rect 10232 14288 10284 14297
rect 12440 14331 12492 14340
rect 12440 14297 12474 14331
rect 12474 14297 12492 14331
rect 12440 14288 12492 14297
rect 8668 14220 8720 14272
rect 9128 14220 9180 14272
rect 9772 14220 9824 14272
rect 13544 14263 13596 14272
rect 13544 14229 13553 14263
rect 13553 14229 13587 14263
rect 13587 14229 13596 14263
rect 13544 14220 13596 14229
rect 13912 14263 13964 14272
rect 13912 14229 13921 14263
rect 13921 14229 13955 14263
rect 13955 14229 13964 14263
rect 13912 14220 13964 14229
rect 19340 14356 19392 14408
rect 19800 14356 19852 14408
rect 15844 14220 15896 14272
rect 18236 14220 18288 14272
rect 18604 14220 18656 14272
rect 19616 14288 19668 14340
rect 20720 14220 20772 14272
rect 20812 14220 20864 14272
rect 4220 14118 4272 14170
rect 4284 14118 4336 14170
rect 4348 14118 4400 14170
rect 4412 14118 4464 14170
rect 4476 14118 4528 14170
rect 9441 14118 9493 14170
rect 9505 14118 9557 14170
rect 9569 14118 9621 14170
rect 9633 14118 9685 14170
rect 9697 14118 9749 14170
rect 14662 14118 14714 14170
rect 14726 14118 14778 14170
rect 14790 14118 14842 14170
rect 14854 14118 14906 14170
rect 14918 14118 14970 14170
rect 19883 14118 19935 14170
rect 19947 14118 19999 14170
rect 20011 14118 20063 14170
rect 20075 14118 20127 14170
rect 20139 14118 20191 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2688 14016 2740 14068
rect 2044 13991 2096 14000
rect 2044 13957 2053 13991
rect 2053 13957 2087 13991
rect 2087 13957 2096 13991
rect 2044 13948 2096 13957
rect 2872 13948 2924 14000
rect 5724 14016 5776 14068
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 3240 13991 3292 14000
rect 3240 13957 3249 13991
rect 3249 13957 3283 13991
rect 3283 13957 3292 13991
rect 3240 13948 3292 13957
rect 4528 13948 4580 14000
rect 4620 13948 4672 14000
rect 5632 13991 5684 14000
rect 5632 13957 5641 13991
rect 5641 13957 5675 13991
rect 5675 13957 5684 13991
rect 5632 13948 5684 13957
rect 6736 13948 6788 14000
rect 4712 13855 4764 13864
rect 4712 13821 4721 13855
rect 4721 13821 4755 13855
rect 4755 13821 4764 13855
rect 4712 13812 4764 13821
rect 5080 13812 5132 13864
rect 5172 13744 5224 13796
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 9312 14016 9364 14068
rect 12348 14016 12400 14068
rect 7840 13991 7892 14000
rect 7840 13957 7849 13991
rect 7849 13957 7883 13991
rect 7883 13957 7892 13991
rect 7840 13948 7892 13957
rect 8576 13948 8628 14000
rect 10508 13948 10560 14000
rect 9772 13923 9824 13932
rect 5632 13744 5684 13796
rect 5264 13676 5316 13728
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 7472 13855 7524 13864
rect 7472 13821 7481 13855
rect 7481 13821 7515 13855
rect 7515 13821 7524 13855
rect 7472 13812 7524 13821
rect 8300 13812 8352 13864
rect 9772 13889 9781 13923
rect 9781 13889 9815 13923
rect 9815 13889 9824 13923
rect 9772 13880 9824 13889
rect 10140 13880 10192 13932
rect 10692 13923 10744 13932
rect 10692 13889 10701 13923
rect 10701 13889 10735 13923
rect 10735 13889 10744 13923
rect 10692 13880 10744 13889
rect 10876 13948 10928 14000
rect 12900 14016 12952 14068
rect 13544 14016 13596 14068
rect 12624 13948 12676 14000
rect 13176 13948 13228 14000
rect 10416 13812 10468 13864
rect 13452 13880 13504 13932
rect 13912 13991 13964 14000
rect 17316 14016 17368 14068
rect 18696 14059 18748 14068
rect 18696 14025 18705 14059
rect 18705 14025 18739 14059
rect 18739 14025 18748 14059
rect 18696 14016 18748 14025
rect 18788 14016 18840 14068
rect 13912 13957 13930 13991
rect 13930 13957 13964 13991
rect 13912 13948 13964 13957
rect 14832 13991 14884 14000
rect 14832 13957 14841 13991
rect 14841 13957 14875 13991
rect 14875 13957 14884 13991
rect 14832 13948 14884 13957
rect 15844 13991 15896 14000
rect 15844 13957 15853 13991
rect 15853 13957 15887 13991
rect 15887 13957 15896 13991
rect 15844 13948 15896 13957
rect 16028 13991 16080 14000
rect 16028 13957 16037 13991
rect 16037 13957 16071 13991
rect 16071 13957 16080 13991
rect 16028 13948 16080 13957
rect 17684 13948 17736 14000
rect 15660 13880 15712 13932
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 17224 13880 17276 13932
rect 19340 13948 19392 14000
rect 18972 13880 19024 13932
rect 20260 14016 20312 14068
rect 20628 13991 20680 14000
rect 20628 13957 20637 13991
rect 20637 13957 20671 13991
rect 20671 13957 20680 13991
rect 20628 13948 20680 13957
rect 20812 13991 20864 14000
rect 20812 13957 20821 13991
rect 20821 13957 20855 13991
rect 20855 13957 20864 13991
rect 20812 13948 20864 13957
rect 12624 13812 12676 13864
rect 14372 13812 14424 13864
rect 15476 13812 15528 13864
rect 11796 13744 11848 13796
rect 15936 13812 15988 13864
rect 20536 13855 20588 13864
rect 20536 13821 20545 13855
rect 20545 13821 20579 13855
rect 20579 13821 20588 13855
rect 20536 13812 20588 13821
rect 20720 13880 20772 13932
rect 20904 13812 20956 13864
rect 19892 13744 19944 13796
rect 8484 13676 8536 13728
rect 9220 13676 9272 13728
rect 10232 13676 10284 13728
rect 13268 13676 13320 13728
rect 13820 13676 13872 13728
rect 20812 13676 20864 13728
rect 3560 13574 3612 13626
rect 3624 13574 3676 13626
rect 3688 13574 3740 13626
rect 3752 13574 3804 13626
rect 3816 13574 3868 13626
rect 8781 13574 8833 13626
rect 8845 13574 8897 13626
rect 8909 13574 8961 13626
rect 8973 13574 9025 13626
rect 9037 13574 9089 13626
rect 14002 13574 14054 13626
rect 14066 13574 14118 13626
rect 14130 13574 14182 13626
rect 14194 13574 14246 13626
rect 14258 13574 14310 13626
rect 19223 13574 19275 13626
rect 19287 13574 19339 13626
rect 19351 13574 19403 13626
rect 19415 13574 19467 13626
rect 19479 13574 19531 13626
rect 2780 13472 2832 13524
rect 2688 13336 2740 13388
rect 4528 13515 4580 13524
rect 4528 13481 4537 13515
rect 4537 13481 4571 13515
rect 4571 13481 4580 13515
rect 4528 13472 4580 13481
rect 4804 13472 4856 13524
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 3332 13268 3384 13320
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 4712 13336 4764 13388
rect 7104 13472 7156 13524
rect 7380 13472 7432 13524
rect 8300 13472 8352 13524
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 10048 13472 10100 13524
rect 12440 13472 12492 13524
rect 13452 13472 13504 13524
rect 17040 13472 17092 13524
rect 18972 13472 19024 13524
rect 21180 13472 21232 13524
rect 5632 13379 5684 13388
rect 5632 13345 5641 13379
rect 5641 13345 5675 13379
rect 5675 13345 5684 13379
rect 5632 13336 5684 13345
rect 5724 13379 5776 13388
rect 5724 13345 5733 13379
rect 5733 13345 5767 13379
rect 5767 13345 5776 13379
rect 5724 13336 5776 13345
rect 6000 13379 6052 13388
rect 6000 13345 6009 13379
rect 6009 13345 6043 13379
rect 6043 13345 6052 13379
rect 6000 13336 6052 13345
rect 6092 13336 6144 13388
rect 7380 13336 7432 13388
rect 10140 13404 10192 13456
rect 16856 13404 16908 13456
rect 8576 13336 8628 13388
rect 9956 13336 10008 13388
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 15936 13379 15988 13388
rect 15936 13345 15945 13379
rect 15945 13345 15979 13379
rect 15979 13345 15988 13379
rect 15936 13336 15988 13345
rect 4528 13268 4580 13320
rect 2044 13243 2096 13252
rect 2044 13209 2053 13243
rect 2053 13209 2087 13243
rect 2087 13209 2096 13243
rect 2044 13200 2096 13209
rect 3056 13200 3108 13252
rect 3424 13200 3476 13252
rect 4988 13268 5040 13320
rect 5356 13200 5408 13252
rect 6092 13200 6144 13252
rect 7012 13200 7064 13252
rect 3976 13175 4028 13184
rect 3976 13141 3985 13175
rect 3985 13141 4019 13175
rect 4019 13141 4028 13175
rect 3976 13132 4028 13141
rect 6736 13132 6788 13184
rect 8300 13268 8352 13320
rect 8668 13268 8720 13320
rect 9220 13311 9272 13320
rect 9220 13277 9230 13311
rect 9230 13277 9264 13311
rect 9264 13277 9272 13311
rect 9220 13268 9272 13277
rect 10048 13268 10100 13320
rect 10232 13268 10284 13320
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10692 13268 10744 13320
rect 13820 13268 13872 13320
rect 18236 13379 18288 13388
rect 18236 13345 18245 13379
rect 18245 13345 18279 13379
rect 18279 13345 18288 13379
rect 18236 13336 18288 13345
rect 19800 13336 19852 13388
rect 19892 13268 19944 13320
rect 20260 13311 20312 13320
rect 20260 13277 20294 13311
rect 20294 13277 20312 13311
rect 20260 13268 20312 13277
rect 10876 13200 10928 13252
rect 12348 13200 12400 13252
rect 14464 13200 14516 13252
rect 9864 13132 9916 13184
rect 10416 13132 10468 13184
rect 14556 13132 14608 13184
rect 16304 13243 16356 13252
rect 16304 13209 16313 13243
rect 16313 13209 16347 13243
rect 16347 13209 16356 13243
rect 16304 13200 16356 13209
rect 16488 13243 16540 13252
rect 16488 13209 16497 13243
rect 16497 13209 16531 13243
rect 16531 13209 16540 13243
rect 16488 13200 16540 13209
rect 18144 13200 18196 13252
rect 20536 13200 20588 13252
rect 16580 13132 16632 13184
rect 17316 13132 17368 13184
rect 18236 13175 18288 13184
rect 18236 13141 18245 13175
rect 18245 13141 18279 13175
rect 18279 13141 18288 13175
rect 18236 13132 18288 13141
rect 18420 13132 18472 13184
rect 4220 13030 4272 13082
rect 4284 13030 4336 13082
rect 4348 13030 4400 13082
rect 4412 13030 4464 13082
rect 4476 13030 4528 13082
rect 9441 13030 9493 13082
rect 9505 13030 9557 13082
rect 9569 13030 9621 13082
rect 9633 13030 9685 13082
rect 9697 13030 9749 13082
rect 14662 13030 14714 13082
rect 14726 13030 14778 13082
rect 14790 13030 14842 13082
rect 14854 13030 14906 13082
rect 14918 13030 14970 13082
rect 19883 13030 19935 13082
rect 19947 13030 19999 13082
rect 20011 13030 20063 13082
rect 20075 13030 20127 13082
rect 20139 13030 20191 13082
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 3424 12792 3476 12844
rect 4712 12928 4764 12980
rect 5632 12928 5684 12980
rect 6460 12971 6512 12980
rect 6460 12937 6469 12971
rect 6469 12937 6503 12971
rect 6503 12937 6512 12971
rect 6460 12928 6512 12937
rect 6920 12928 6972 12980
rect 7104 12928 7156 12980
rect 4620 12860 4672 12912
rect 5816 12860 5868 12912
rect 6552 12860 6604 12912
rect 7288 12903 7340 12912
rect 7288 12869 7297 12903
rect 7297 12869 7331 12903
rect 7331 12869 7340 12903
rect 7288 12860 7340 12869
rect 7472 12860 7524 12912
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 5908 12835 5960 12844
rect 5908 12801 5917 12835
rect 5917 12801 5951 12835
rect 5951 12801 5960 12835
rect 5908 12792 5960 12801
rect 4896 12724 4948 12776
rect 6276 12792 6328 12844
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 6736 12792 6788 12844
rect 7012 12724 7064 12776
rect 7380 12724 7432 12776
rect 7656 12792 7708 12844
rect 8668 12792 8720 12844
rect 9312 12860 9364 12912
rect 10140 12860 10192 12912
rect 10876 12860 10928 12912
rect 6552 12656 6604 12708
rect 3792 12588 3844 12640
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 8576 12656 8628 12708
rect 9864 12767 9916 12776
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 9864 12724 9916 12733
rect 10232 12724 10284 12776
rect 10784 12792 10836 12844
rect 12716 12860 12768 12912
rect 13176 12903 13228 12912
rect 13176 12869 13185 12903
rect 13185 12869 13219 12903
rect 13219 12869 13228 12903
rect 13176 12860 13228 12869
rect 16304 12928 16356 12980
rect 18052 12971 18104 12980
rect 18052 12937 18061 12971
rect 18061 12937 18095 12971
rect 18095 12937 18104 12971
rect 18052 12928 18104 12937
rect 20352 12928 20404 12980
rect 11796 12792 11848 12844
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 18144 12903 18196 12912
rect 18144 12869 18153 12903
rect 18153 12869 18187 12903
rect 18187 12869 18196 12903
rect 18144 12860 18196 12869
rect 12992 12724 13044 12776
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 14372 12724 14424 12776
rect 10048 12656 10100 12708
rect 10140 12656 10192 12708
rect 10324 12656 10376 12708
rect 10600 12656 10652 12708
rect 13636 12656 13688 12708
rect 13728 12699 13780 12708
rect 13728 12665 13737 12699
rect 13737 12665 13771 12699
rect 13771 12665 13780 12699
rect 13728 12656 13780 12665
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18512 12860 18564 12912
rect 21180 12860 21232 12912
rect 18604 12792 18656 12844
rect 20352 12792 20404 12844
rect 20536 12792 20588 12844
rect 18972 12767 19024 12776
rect 18972 12733 18981 12767
rect 18981 12733 19015 12767
rect 19015 12733 19024 12767
rect 18972 12724 19024 12733
rect 18236 12656 18288 12708
rect 20720 12699 20772 12708
rect 20720 12665 20729 12699
rect 20729 12665 20763 12699
rect 20763 12665 20772 12699
rect 20720 12656 20772 12665
rect 9220 12588 9272 12640
rect 10232 12631 10284 12640
rect 10232 12597 10241 12631
rect 10241 12597 10275 12631
rect 10275 12597 10284 12631
rect 10232 12588 10284 12597
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12440 12588 12492 12597
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 16856 12588 16908 12640
rect 18420 12631 18472 12640
rect 18420 12597 18429 12631
rect 18429 12597 18463 12631
rect 18463 12597 18472 12631
rect 18420 12588 18472 12597
rect 3560 12486 3612 12538
rect 3624 12486 3676 12538
rect 3688 12486 3740 12538
rect 3752 12486 3804 12538
rect 3816 12486 3868 12538
rect 8781 12486 8833 12538
rect 8845 12486 8897 12538
rect 8909 12486 8961 12538
rect 8973 12486 9025 12538
rect 9037 12486 9089 12538
rect 14002 12486 14054 12538
rect 14066 12486 14118 12538
rect 14130 12486 14182 12538
rect 14194 12486 14246 12538
rect 14258 12486 14310 12538
rect 19223 12486 19275 12538
rect 19287 12486 19339 12538
rect 19351 12486 19403 12538
rect 19415 12486 19467 12538
rect 19479 12486 19531 12538
rect 6644 12384 6696 12436
rect 9128 12384 9180 12436
rect 2872 12291 2924 12300
rect 2872 12257 2881 12291
rect 2881 12257 2915 12291
rect 2915 12257 2924 12291
rect 2872 12248 2924 12257
rect 4620 12248 4672 12300
rect 5724 12248 5776 12300
rect 7380 12248 7432 12300
rect 2780 12180 2832 12232
rect 7196 12180 7248 12232
rect 8208 12180 8260 12232
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 9864 12316 9916 12368
rect 10416 12316 10468 12368
rect 10600 12384 10652 12436
rect 12440 12384 12492 12436
rect 12992 12384 13044 12436
rect 16488 12384 16540 12436
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9312 12180 9364 12232
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 13268 12291 13320 12300
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 11060 12180 11112 12232
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13728 12180 13780 12232
rect 15016 12180 15068 12232
rect 18420 12384 18472 12436
rect 18604 12316 18656 12368
rect 18972 12316 19024 12368
rect 16856 12223 16908 12232
rect 16856 12189 16865 12223
rect 16865 12189 16899 12223
rect 16899 12189 16908 12223
rect 16856 12180 16908 12189
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 21272 12316 21324 12368
rect 19708 12248 19760 12300
rect 20444 12248 20496 12300
rect 20536 12180 20588 12232
rect 3056 12112 3108 12164
rect 4896 12112 4948 12164
rect 6552 12112 6604 12164
rect 10324 12112 10376 12164
rect 12624 12112 12676 12164
rect 13176 12112 13228 12164
rect 16672 12112 16724 12164
rect 1860 12044 1912 12096
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 3332 12044 3384 12096
rect 4988 12044 5040 12096
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 9956 12087 10008 12096
rect 9956 12053 9965 12087
rect 9965 12053 9999 12087
rect 9999 12053 10008 12087
rect 9956 12044 10008 12053
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 11336 12044 11388 12096
rect 12440 12044 12492 12096
rect 12716 12044 12768 12096
rect 13452 12044 13504 12096
rect 20812 12112 20864 12164
rect 21364 12112 21416 12164
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 19248 12044 19300 12096
rect 20720 12087 20772 12096
rect 20720 12053 20729 12087
rect 20729 12053 20763 12087
rect 20763 12053 20772 12087
rect 20720 12044 20772 12053
rect 4220 11942 4272 11994
rect 4284 11942 4336 11994
rect 4348 11942 4400 11994
rect 4412 11942 4464 11994
rect 4476 11942 4528 11994
rect 9441 11942 9493 11994
rect 9505 11942 9557 11994
rect 9569 11942 9621 11994
rect 9633 11942 9685 11994
rect 9697 11942 9749 11994
rect 14662 11942 14714 11994
rect 14726 11942 14778 11994
rect 14790 11942 14842 11994
rect 14854 11942 14906 11994
rect 14918 11942 14970 11994
rect 19883 11942 19935 11994
rect 19947 11942 19999 11994
rect 20011 11942 20063 11994
rect 20075 11942 20127 11994
rect 20139 11942 20191 11994
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 10048 11840 10100 11892
rect 10600 11840 10652 11892
rect 1860 11747 1912 11756
rect 1860 11713 1894 11747
rect 1894 11713 1912 11747
rect 1860 11704 1912 11713
rect 7748 11772 7800 11824
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 5080 11704 5132 11756
rect 10324 11772 10376 11824
rect 11152 11815 11204 11824
rect 11152 11781 11161 11815
rect 11161 11781 11195 11815
rect 11195 11781 11204 11815
rect 11152 11772 11204 11781
rect 11336 11772 11388 11824
rect 13268 11840 13320 11892
rect 13728 11840 13780 11892
rect 15936 11840 15988 11892
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 2964 11543 3016 11552
rect 2964 11509 2973 11543
rect 2973 11509 3007 11543
rect 3007 11509 3016 11543
rect 2964 11500 3016 11509
rect 4988 11611 5040 11620
rect 4988 11577 4997 11611
rect 4997 11577 5031 11611
rect 5031 11577 5040 11611
rect 4988 11568 5040 11577
rect 6092 11568 6144 11620
rect 4620 11500 4672 11552
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 8576 11636 8628 11688
rect 9588 11636 9640 11688
rect 9864 11636 9916 11688
rect 11060 11568 11112 11620
rect 10508 11500 10560 11552
rect 11612 11636 11664 11688
rect 13452 11747 13504 11756
rect 13452 11713 13470 11747
rect 13470 11713 13504 11747
rect 13452 11704 13504 11713
rect 13820 11747 13872 11756
rect 13820 11713 13829 11747
rect 13829 11713 13863 11747
rect 13863 11713 13872 11747
rect 13820 11704 13872 11713
rect 16028 11815 16080 11824
rect 16028 11781 16037 11815
rect 16037 11781 16071 11815
rect 16071 11781 16080 11815
rect 16028 11772 16080 11781
rect 17040 11772 17092 11824
rect 20720 11840 20772 11892
rect 15660 11704 15712 11756
rect 16488 11747 16540 11756
rect 16488 11713 16497 11747
rect 16497 11713 16531 11747
rect 16531 11713 16540 11747
rect 16488 11704 16540 11713
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 12532 11636 12584 11688
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 19064 11636 19116 11688
rect 11888 11543 11940 11552
rect 11888 11509 11897 11543
rect 11897 11509 11931 11543
rect 11931 11509 11940 11543
rect 11888 11500 11940 11509
rect 15108 11568 15160 11620
rect 12624 11500 12676 11552
rect 13084 11500 13136 11552
rect 14372 11500 14424 11552
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 21088 11543 21140 11552
rect 21088 11509 21097 11543
rect 21097 11509 21131 11543
rect 21131 11509 21140 11543
rect 21088 11500 21140 11509
rect 3560 11398 3612 11450
rect 3624 11398 3676 11450
rect 3688 11398 3740 11450
rect 3752 11398 3804 11450
rect 3816 11398 3868 11450
rect 8781 11398 8833 11450
rect 8845 11398 8897 11450
rect 8909 11398 8961 11450
rect 8973 11398 9025 11450
rect 9037 11398 9089 11450
rect 14002 11398 14054 11450
rect 14066 11398 14118 11450
rect 14130 11398 14182 11450
rect 14194 11398 14246 11450
rect 14258 11398 14310 11450
rect 19223 11398 19275 11450
rect 19287 11398 19339 11450
rect 19351 11398 19403 11450
rect 19415 11398 19467 11450
rect 19479 11398 19531 11450
rect 4804 11296 4856 11348
rect 4896 11296 4948 11348
rect 7104 11296 7156 11348
rect 8300 11296 8352 11348
rect 6644 11271 6696 11280
rect 6644 11237 6653 11271
rect 6653 11237 6687 11271
rect 6687 11237 6696 11271
rect 6644 11228 6696 11237
rect 7288 11271 7340 11280
rect 7288 11237 7297 11271
rect 7297 11237 7331 11271
rect 7331 11237 7340 11271
rect 7288 11228 7340 11237
rect 9220 11228 9272 11280
rect 11612 11296 11664 11348
rect 11888 11296 11940 11348
rect 1676 11092 1728 11144
rect 2964 11092 3016 11144
rect 3332 11024 3384 11076
rect 3792 10956 3844 11008
rect 4620 11092 4672 11144
rect 5172 11092 5224 11144
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 5356 11024 5408 11076
rect 6920 11160 6972 11212
rect 9128 11160 9180 11212
rect 9956 11160 10008 11212
rect 10232 11203 10284 11212
rect 10232 11169 10241 11203
rect 10241 11169 10275 11203
rect 10275 11169 10284 11203
rect 10232 11160 10284 11169
rect 10600 11160 10652 11212
rect 4896 10956 4948 11008
rect 5540 10956 5592 11008
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 10324 11092 10376 11144
rect 10508 11092 10560 11144
rect 11244 11135 11296 11144
rect 11244 11101 11278 11135
rect 11278 11101 11296 11135
rect 11244 11092 11296 11101
rect 13360 11296 13412 11348
rect 12808 11228 12860 11280
rect 13636 11228 13688 11280
rect 13820 11296 13872 11348
rect 16488 11296 16540 11348
rect 16120 11228 16172 11280
rect 17592 11228 17644 11280
rect 13268 11160 13320 11212
rect 16580 11160 16632 11212
rect 17224 11203 17276 11212
rect 17224 11169 17233 11203
rect 17233 11169 17267 11203
rect 17267 11169 17276 11203
rect 17224 11160 17276 11169
rect 20720 11296 20772 11348
rect 21364 11339 21416 11348
rect 21364 11305 21373 11339
rect 21373 11305 21407 11339
rect 21407 11305 21416 11339
rect 21364 11296 21416 11305
rect 19064 11160 19116 11212
rect 15108 11135 15160 11144
rect 15108 11101 15117 11135
rect 15117 11101 15151 11135
rect 15151 11101 15160 11135
rect 15108 11092 15160 11101
rect 16304 11092 16356 11144
rect 8208 10956 8260 11008
rect 8484 10956 8536 11008
rect 10784 11024 10836 11076
rect 12440 11024 12492 11076
rect 9128 10956 9180 11008
rect 12624 10956 12676 11008
rect 13084 11024 13136 11076
rect 13452 11067 13504 11076
rect 13452 11033 13461 11067
rect 13461 11033 13495 11067
rect 13495 11033 13504 11067
rect 13452 11024 13504 11033
rect 16028 11024 16080 11076
rect 14464 10956 14516 11008
rect 15016 10956 15068 11008
rect 16580 11024 16632 11076
rect 17316 11067 17368 11076
rect 17316 11033 17325 11067
rect 17325 11033 17359 11067
rect 17359 11033 17368 11067
rect 17316 11024 17368 11033
rect 17960 11067 18012 11076
rect 17960 11033 17969 11067
rect 17969 11033 18003 11067
rect 18003 11033 18012 11067
rect 17960 11024 18012 11033
rect 21088 11092 21140 11144
rect 20904 11024 20956 11076
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 19800 10956 19852 11008
rect 4220 10854 4272 10906
rect 4284 10854 4336 10906
rect 4348 10854 4400 10906
rect 4412 10854 4464 10906
rect 4476 10854 4528 10906
rect 9441 10854 9493 10906
rect 9505 10854 9557 10906
rect 9569 10854 9621 10906
rect 9633 10854 9685 10906
rect 9697 10854 9749 10906
rect 14662 10854 14714 10906
rect 14726 10854 14778 10906
rect 14790 10854 14842 10906
rect 14854 10854 14906 10906
rect 14918 10854 14970 10906
rect 19883 10854 19935 10906
rect 19947 10854 19999 10906
rect 20011 10854 20063 10906
rect 20075 10854 20127 10906
rect 20139 10854 20191 10906
rect 3792 10795 3844 10804
rect 3792 10761 3801 10795
rect 3801 10761 3835 10795
rect 3835 10761 3844 10795
rect 3792 10752 3844 10761
rect 4160 10752 4212 10804
rect 5264 10752 5316 10804
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 3240 10684 3292 10736
rect 4712 10684 4764 10736
rect 5448 10684 5500 10736
rect 11796 10752 11848 10804
rect 12532 10752 12584 10804
rect 13452 10752 13504 10804
rect 16028 10752 16080 10804
rect 1952 10659 2004 10668
rect 1952 10625 1986 10659
rect 1986 10625 2004 10659
rect 1952 10616 2004 10625
rect 5908 10616 5960 10668
rect 6828 10616 6880 10668
rect 7012 10616 7064 10668
rect 7932 10616 7984 10668
rect 8116 10659 8168 10668
rect 8116 10625 8125 10659
rect 8125 10625 8159 10659
rect 8159 10625 8168 10659
rect 8116 10616 8168 10625
rect 8484 10659 8536 10668
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9220 10616 9272 10668
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 14372 10727 14424 10736
rect 14372 10693 14390 10727
rect 14390 10693 14424 10727
rect 14372 10684 14424 10693
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 4160 10548 4212 10600
rect 4804 10548 4856 10600
rect 3332 10523 3384 10532
rect 3332 10489 3341 10523
rect 3341 10489 3375 10523
rect 3375 10489 3384 10523
rect 3332 10480 3384 10489
rect 5448 10548 5500 10600
rect 2872 10412 2924 10464
rect 5080 10523 5132 10532
rect 5080 10489 5089 10523
rect 5089 10489 5123 10523
rect 5123 10489 5132 10523
rect 5080 10480 5132 10489
rect 5264 10480 5316 10532
rect 10416 10591 10468 10600
rect 10416 10557 10425 10591
rect 10425 10557 10459 10591
rect 10459 10557 10468 10591
rect 10416 10548 10468 10557
rect 10324 10480 10376 10532
rect 10692 10480 10744 10532
rect 11244 10616 11296 10668
rect 12072 10616 12124 10668
rect 16120 10684 16172 10736
rect 17132 10684 17184 10736
rect 15108 10616 15160 10668
rect 15292 10659 15344 10668
rect 15292 10625 15326 10659
rect 15326 10625 15344 10659
rect 15292 10616 15344 10625
rect 21364 10684 21416 10736
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 13268 10523 13320 10532
rect 13268 10489 13277 10523
rect 13277 10489 13311 10523
rect 13311 10489 13320 10523
rect 13268 10480 13320 10489
rect 19064 10548 19116 10600
rect 20812 10548 20864 10600
rect 20996 10591 21048 10600
rect 20996 10557 21005 10591
rect 21005 10557 21039 10591
rect 21039 10557 21048 10591
rect 20996 10548 21048 10557
rect 5816 10412 5868 10464
rect 6000 10412 6052 10464
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 7748 10412 7800 10421
rect 14372 10412 14424 10464
rect 17960 10412 18012 10464
rect 3560 10310 3612 10362
rect 3624 10310 3676 10362
rect 3688 10310 3740 10362
rect 3752 10310 3804 10362
rect 3816 10310 3868 10362
rect 8781 10310 8833 10362
rect 8845 10310 8897 10362
rect 8909 10310 8961 10362
rect 8973 10310 9025 10362
rect 9037 10310 9089 10362
rect 14002 10310 14054 10362
rect 14066 10310 14118 10362
rect 14130 10310 14182 10362
rect 14194 10310 14246 10362
rect 14258 10310 14310 10362
rect 19223 10310 19275 10362
rect 19287 10310 19339 10362
rect 19351 10310 19403 10362
rect 19415 10310 19467 10362
rect 19479 10310 19531 10362
rect 1952 10208 2004 10260
rect 3148 10208 3200 10260
rect 6092 10208 6144 10260
rect 4160 10140 4212 10192
rect 5448 10140 5500 10192
rect 7748 10208 7800 10260
rect 3056 10004 3108 10056
rect 3332 10004 3384 10056
rect 4160 10004 4212 10056
rect 5080 10004 5132 10056
rect 1308 9936 1360 9988
rect 2964 9979 3016 9988
rect 2964 9945 2973 9979
rect 2973 9945 3007 9979
rect 3007 9945 3016 9979
rect 2964 9936 3016 9945
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 4620 9936 4672 9988
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 7380 10140 7432 10192
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 8484 10208 8536 10260
rect 11244 10208 11296 10260
rect 8208 10183 8260 10192
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 8208 10140 8260 10149
rect 12072 10208 12124 10260
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 15292 10208 15344 10260
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 17316 10208 17368 10260
rect 18144 10208 18196 10260
rect 8300 10047 8352 10056
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 9220 10004 9272 10056
rect 12532 10072 12584 10124
rect 12900 10115 12952 10124
rect 12900 10081 12909 10115
rect 12909 10081 12943 10115
rect 12943 10081 12952 10115
rect 12900 10072 12952 10081
rect 17132 10115 17184 10124
rect 17132 10081 17141 10115
rect 17141 10081 17175 10115
rect 17175 10081 17184 10115
rect 17132 10072 17184 10081
rect 12348 10004 12400 10056
rect 10324 9936 10376 9988
rect 10784 9936 10836 9988
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 12808 9979 12860 9988
rect 12808 9945 12817 9979
rect 12817 9945 12851 9979
rect 12851 9945 12860 9979
rect 12808 9936 12860 9945
rect 4252 9868 4304 9920
rect 4804 9868 4856 9920
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 7012 9911 7064 9920
rect 7012 9877 7021 9911
rect 7021 9877 7055 9911
rect 7055 9877 7064 9911
rect 7012 9868 7064 9877
rect 7380 9868 7432 9920
rect 7932 9868 7984 9920
rect 12440 9868 12492 9920
rect 13176 9868 13228 9920
rect 14372 10004 14424 10056
rect 15384 10004 15436 10056
rect 15568 10047 15620 10056
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 19064 10004 19116 10056
rect 19892 10004 19944 10056
rect 20628 10004 20680 10056
rect 16212 9936 16264 9988
rect 17408 9979 17460 9988
rect 17408 9945 17442 9979
rect 17442 9945 17460 9979
rect 17408 9936 17460 9945
rect 20260 9936 20312 9988
rect 21272 9868 21324 9920
rect 4220 9766 4272 9818
rect 4284 9766 4336 9818
rect 4348 9766 4400 9818
rect 4412 9766 4464 9818
rect 4476 9766 4528 9818
rect 9441 9766 9493 9818
rect 9505 9766 9557 9818
rect 9569 9766 9621 9818
rect 9633 9766 9685 9818
rect 9697 9766 9749 9818
rect 14662 9766 14714 9818
rect 14726 9766 14778 9818
rect 14790 9766 14842 9818
rect 14854 9766 14906 9818
rect 14918 9766 14970 9818
rect 19883 9766 19935 9818
rect 19947 9766 19999 9818
rect 20011 9766 20063 9818
rect 20075 9766 20127 9818
rect 20139 9766 20191 9818
rect 1308 9596 1360 9648
rect 2872 9596 2924 9648
rect 3056 9528 3108 9580
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 3884 9596 3936 9648
rect 5632 9596 5684 9648
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 6552 9596 6604 9648
rect 9680 9664 9732 9716
rect 10416 9664 10468 9716
rect 17408 9707 17460 9716
rect 17408 9673 17417 9707
rect 17417 9673 17451 9707
rect 17451 9673 17460 9707
rect 17408 9664 17460 9673
rect 18144 9664 18196 9716
rect 21364 9707 21416 9716
rect 21364 9673 21373 9707
rect 21373 9673 21407 9707
rect 21407 9673 21416 9707
rect 21364 9664 21416 9673
rect 3976 9571 4028 9580
rect 3976 9537 3985 9571
rect 3985 9537 4019 9571
rect 4019 9537 4028 9571
rect 3976 9528 4028 9537
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 4988 9528 5040 9580
rect 6092 9528 6144 9580
rect 8484 9596 8536 9648
rect 6736 9528 6788 9580
rect 7564 9528 7616 9580
rect 7656 9528 7708 9580
rect 2964 9460 3016 9512
rect 4712 9392 4764 9444
rect 4804 9435 4856 9444
rect 4804 9401 4813 9435
rect 4813 9401 4847 9435
rect 4847 9401 4856 9435
rect 4804 9392 4856 9401
rect 5632 9435 5684 9444
rect 5632 9401 5641 9435
rect 5641 9401 5675 9435
rect 5675 9401 5684 9435
rect 5632 9392 5684 9401
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 3976 9324 4028 9376
rect 6000 9324 6052 9376
rect 7932 9460 7984 9512
rect 9128 9528 9180 9580
rect 10600 9596 10652 9648
rect 12624 9596 12676 9648
rect 10784 9528 10836 9580
rect 8024 9392 8076 9444
rect 8668 9392 8720 9444
rect 14372 9639 14424 9648
rect 14372 9605 14381 9639
rect 14381 9605 14415 9639
rect 14415 9605 14424 9639
rect 14372 9596 14424 9605
rect 15752 9596 15804 9648
rect 17040 9596 17092 9648
rect 19064 9596 19116 9648
rect 20444 9596 20496 9648
rect 20536 9596 20588 9648
rect 13820 9460 13872 9512
rect 15384 9528 15436 9580
rect 15476 9460 15528 9512
rect 15660 9528 15712 9580
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 18144 9528 18196 9580
rect 21180 9528 21232 9580
rect 15844 9460 15896 9512
rect 17316 9460 17368 9512
rect 8300 9324 8352 9376
rect 8392 9324 8444 9376
rect 10048 9324 10100 9376
rect 12164 9324 12216 9376
rect 13728 9367 13780 9376
rect 13728 9333 13737 9367
rect 13737 9333 13771 9367
rect 13771 9333 13780 9367
rect 13728 9324 13780 9333
rect 16304 9324 16356 9376
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 18880 9392 18932 9444
rect 19892 9392 19944 9444
rect 21364 9503 21416 9512
rect 21364 9469 21373 9503
rect 21373 9469 21407 9503
rect 21407 9469 21416 9503
rect 21364 9460 21416 9469
rect 20352 9392 20404 9444
rect 20628 9435 20680 9444
rect 20628 9401 20637 9435
rect 20637 9401 20671 9435
rect 20671 9401 20680 9435
rect 20628 9392 20680 9401
rect 20904 9435 20956 9444
rect 20904 9401 20913 9435
rect 20913 9401 20947 9435
rect 20947 9401 20956 9435
rect 20904 9392 20956 9401
rect 20536 9324 20588 9376
rect 3560 9222 3612 9274
rect 3624 9222 3676 9274
rect 3688 9222 3740 9274
rect 3752 9222 3804 9274
rect 3816 9222 3868 9274
rect 8781 9222 8833 9274
rect 8845 9222 8897 9274
rect 8909 9222 8961 9274
rect 8973 9222 9025 9274
rect 9037 9222 9089 9274
rect 14002 9222 14054 9274
rect 14066 9222 14118 9274
rect 14130 9222 14182 9274
rect 14194 9222 14246 9274
rect 14258 9222 14310 9274
rect 19223 9222 19275 9274
rect 19287 9222 19339 9274
rect 19351 9222 19403 9274
rect 19415 9222 19467 9274
rect 19479 9222 19531 9274
rect 7656 9120 7708 9172
rect 17040 9163 17092 9172
rect 17040 9129 17049 9163
rect 17049 9129 17083 9163
rect 17083 9129 17092 9163
rect 17040 9120 17092 9129
rect 18236 9120 18288 9172
rect 20812 9120 20864 9172
rect 4896 9052 4948 9104
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 1952 8959 2004 8968
rect 1952 8925 1986 8959
rect 1986 8925 2004 8959
rect 1952 8916 2004 8925
rect 4712 8916 4764 8968
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 7564 9095 7616 9104
rect 7564 9061 7573 9095
rect 7573 9061 7607 9095
rect 7607 9061 7616 9095
rect 7564 9052 7616 9061
rect 7840 9052 7892 9104
rect 11704 9052 11756 9104
rect 13912 9052 13964 9104
rect 7288 8984 7340 9036
rect 5540 8916 5592 8968
rect 6736 8916 6788 8968
rect 7012 8916 7064 8968
rect 8024 8916 8076 8968
rect 8484 8959 8536 8968
rect 8484 8925 8493 8959
rect 8493 8925 8527 8959
rect 8527 8925 8536 8959
rect 8484 8916 8536 8925
rect 3884 8848 3936 8900
rect 4620 8891 4672 8900
rect 4620 8857 4629 8891
rect 4629 8857 4663 8891
rect 4663 8857 4672 8891
rect 4620 8848 4672 8857
rect 4804 8848 4856 8900
rect 5080 8891 5132 8900
rect 5080 8857 5089 8891
rect 5089 8857 5123 8891
rect 5123 8857 5132 8891
rect 5080 8848 5132 8857
rect 5172 8891 5224 8900
rect 5172 8857 5181 8891
rect 5181 8857 5215 8891
rect 5215 8857 5224 8891
rect 5172 8848 5224 8857
rect 5632 8848 5684 8900
rect 8392 8848 8444 8900
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 11520 8984 11572 9036
rect 14096 9027 14148 9036
rect 9128 8916 9180 8968
rect 11612 8916 11664 8968
rect 14096 8993 14105 9027
rect 14105 8993 14139 9027
rect 14139 8993 14148 9027
rect 14096 8984 14148 8993
rect 17132 8984 17184 9036
rect 9680 8848 9732 8900
rect 10140 8848 10192 8900
rect 11244 8891 11296 8900
rect 11244 8857 11253 8891
rect 11253 8857 11287 8891
rect 11287 8857 11296 8891
rect 11244 8848 11296 8857
rect 12164 8891 12216 8900
rect 12164 8857 12198 8891
rect 12198 8857 12216 8891
rect 3056 8823 3108 8832
rect 3056 8789 3065 8823
rect 3065 8789 3099 8823
rect 3099 8789 3108 8823
rect 3056 8780 3108 8789
rect 4068 8780 4120 8832
rect 5816 8780 5868 8832
rect 6552 8780 6604 8832
rect 6828 8780 6880 8832
rect 7932 8823 7984 8832
rect 7932 8789 7941 8823
rect 7941 8789 7975 8823
rect 7975 8789 7984 8823
rect 7932 8780 7984 8789
rect 9312 8780 9364 8832
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 11428 8823 11480 8832
rect 11428 8789 11437 8823
rect 11437 8789 11471 8823
rect 11471 8789 11480 8823
rect 11428 8780 11480 8789
rect 12164 8848 12216 8857
rect 12348 8848 12400 8900
rect 13728 8916 13780 8968
rect 15108 8916 15160 8968
rect 18328 8916 18380 8968
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 13820 8848 13872 8900
rect 16120 8848 16172 8900
rect 16856 8848 16908 8900
rect 19708 8848 19760 8900
rect 20996 8848 21048 8900
rect 13176 8780 13228 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 18420 8780 18472 8832
rect 18880 8780 18932 8832
rect 20536 8780 20588 8832
rect 20904 8780 20956 8832
rect 21364 8780 21416 8832
rect 4220 8678 4272 8730
rect 4284 8678 4336 8730
rect 4348 8678 4400 8730
rect 4412 8678 4464 8730
rect 4476 8678 4528 8730
rect 9441 8678 9493 8730
rect 9505 8678 9557 8730
rect 9569 8678 9621 8730
rect 9633 8678 9685 8730
rect 9697 8678 9749 8730
rect 14662 8678 14714 8730
rect 14726 8678 14778 8730
rect 14790 8678 14842 8730
rect 14854 8678 14906 8730
rect 14918 8678 14970 8730
rect 19883 8678 19935 8730
rect 19947 8678 19999 8730
rect 20011 8678 20063 8730
rect 20075 8678 20127 8730
rect 20139 8678 20191 8730
rect 5172 8576 5224 8628
rect 7288 8619 7340 8628
rect 7288 8585 7297 8619
rect 7297 8585 7331 8619
rect 7331 8585 7340 8619
rect 7288 8576 7340 8585
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 7932 8619 7984 8628
rect 7932 8585 7941 8619
rect 7941 8585 7975 8619
rect 7975 8585 7984 8619
rect 7932 8576 7984 8585
rect 14372 8576 14424 8628
rect 17040 8576 17092 8628
rect 1676 8508 1728 8560
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 4620 8508 4672 8560
rect 6092 8508 6144 8560
rect 7380 8551 7432 8560
rect 7380 8517 7389 8551
rect 7389 8517 7423 8551
rect 7423 8517 7432 8551
rect 7380 8508 7432 8517
rect 4160 8440 4212 8492
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 8300 8440 8352 8492
rect 10232 8508 10284 8560
rect 10508 8508 10560 8560
rect 12624 8551 12676 8560
rect 12624 8517 12633 8551
rect 12633 8517 12667 8551
rect 12667 8517 12676 8551
rect 12624 8508 12676 8517
rect 13452 8508 13504 8560
rect 14096 8508 14148 8560
rect 14556 8508 14608 8560
rect 15108 8508 15160 8560
rect 15844 8551 15896 8560
rect 15844 8517 15853 8551
rect 15853 8517 15887 8551
rect 15887 8517 15896 8551
rect 15844 8508 15896 8517
rect 16948 8508 17000 8560
rect 17224 8551 17276 8560
rect 17224 8517 17233 8551
rect 17233 8517 17267 8551
rect 17267 8517 17276 8551
rect 17224 8508 17276 8517
rect 19616 8576 19668 8628
rect 21180 8576 21232 8628
rect 20260 8551 20312 8560
rect 6736 8372 6788 8424
rect 3148 8236 3200 8288
rect 4988 8236 5040 8288
rect 5448 8236 5500 8288
rect 6092 8279 6144 8288
rect 6092 8245 6101 8279
rect 6101 8245 6135 8279
rect 6135 8245 6144 8279
rect 6092 8236 6144 8245
rect 10600 8440 10652 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 9128 8236 9180 8288
rect 11428 8304 11480 8356
rect 11888 8304 11940 8356
rect 12348 8440 12400 8492
rect 12532 8372 12584 8424
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 14464 8483 14516 8492
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 17960 8440 18012 8492
rect 15108 8372 15160 8424
rect 15752 8372 15804 8424
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17316 8415 17368 8424
rect 17316 8381 17325 8415
rect 17325 8381 17359 8415
rect 17359 8381 17368 8415
rect 17316 8372 17368 8381
rect 18236 8440 18288 8492
rect 18328 8483 18380 8492
rect 18328 8449 18337 8483
rect 18337 8449 18371 8483
rect 18371 8449 18380 8483
rect 18328 8440 18380 8449
rect 18880 8440 18932 8492
rect 20260 8517 20294 8551
rect 20294 8517 20312 8551
rect 20260 8508 20312 8517
rect 13912 8304 13964 8356
rect 14464 8304 14516 8356
rect 18236 8304 18288 8356
rect 9588 8279 9640 8288
rect 9588 8245 9597 8279
rect 9597 8245 9631 8279
rect 9631 8245 9640 8279
rect 9588 8236 9640 8245
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 12072 8236 12124 8288
rect 16764 8279 16816 8288
rect 16764 8245 16773 8279
rect 16773 8245 16807 8279
rect 16807 8245 16816 8279
rect 16764 8236 16816 8245
rect 17592 8279 17644 8288
rect 17592 8245 17601 8279
rect 17601 8245 17635 8279
rect 17635 8245 17644 8279
rect 17592 8236 17644 8245
rect 19708 8279 19760 8288
rect 19708 8245 19717 8279
rect 19717 8245 19751 8279
rect 19751 8245 19760 8279
rect 19708 8236 19760 8245
rect 3560 8134 3612 8186
rect 3624 8134 3676 8186
rect 3688 8134 3740 8186
rect 3752 8134 3804 8186
rect 3816 8134 3868 8186
rect 8781 8134 8833 8186
rect 8845 8134 8897 8186
rect 8909 8134 8961 8186
rect 8973 8134 9025 8186
rect 9037 8134 9089 8186
rect 14002 8134 14054 8186
rect 14066 8134 14118 8186
rect 14130 8134 14182 8186
rect 14194 8134 14246 8186
rect 14258 8134 14310 8186
rect 19223 8134 19275 8186
rect 19287 8134 19339 8186
rect 19351 8134 19403 8186
rect 19415 8134 19467 8186
rect 19479 8134 19531 8186
rect 5632 8032 5684 8084
rect 7104 8032 7156 8084
rect 4712 7964 4764 8016
rect 3056 7896 3108 7948
rect 2872 7828 2924 7880
rect 3516 7828 3568 7880
rect 5264 7896 5316 7948
rect 2228 7760 2280 7812
rect 3148 7760 3200 7812
rect 4160 7871 4212 7880
rect 4160 7837 4174 7871
rect 4174 7837 4208 7871
rect 4208 7837 4212 7871
rect 4160 7828 4212 7837
rect 5356 7828 5408 7880
rect 6736 7828 6788 7880
rect 8392 8032 8444 8084
rect 9036 8032 9088 8084
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 10232 7939 10284 7948
rect 10232 7905 10241 7939
rect 10241 7905 10275 7939
rect 10275 7905 10284 7939
rect 10232 7896 10284 7905
rect 12348 8032 12400 8084
rect 12624 8032 12676 8084
rect 13820 8032 13872 8084
rect 16948 8075 17000 8084
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 20628 8075 20680 8084
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 14280 7964 14332 8016
rect 16488 8007 16540 8016
rect 16488 7973 16497 8007
rect 16497 7973 16531 8007
rect 16531 7973 16540 8007
rect 16488 7964 16540 7973
rect 17316 7964 17368 8016
rect 21180 7964 21232 8016
rect 14004 7896 14056 7948
rect 16764 7896 16816 7948
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 21364 7939 21416 7948
rect 21364 7905 21373 7939
rect 21373 7905 21407 7939
rect 21407 7905 21416 7939
rect 21364 7896 21416 7905
rect 7932 7828 7984 7880
rect 8392 7828 8444 7880
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 11520 7828 11572 7880
rect 12072 7828 12124 7880
rect 15016 7828 15068 7880
rect 15752 7828 15804 7880
rect 17224 7828 17276 7880
rect 18236 7828 18288 7880
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 21088 7828 21140 7880
rect 3976 7803 4028 7812
rect 3976 7769 3985 7803
rect 3985 7769 4019 7803
rect 4019 7769 4028 7803
rect 3976 7760 4028 7769
rect 3056 7692 3108 7744
rect 3792 7692 3844 7744
rect 5080 7803 5132 7812
rect 5080 7769 5089 7803
rect 5089 7769 5123 7803
rect 5123 7769 5132 7803
rect 5080 7760 5132 7769
rect 6552 7760 6604 7812
rect 7656 7760 7708 7812
rect 8484 7803 8536 7812
rect 8484 7769 8493 7803
rect 8493 7769 8527 7803
rect 8527 7769 8536 7803
rect 8484 7760 8536 7769
rect 9220 7760 9272 7812
rect 12716 7760 12768 7812
rect 15844 7803 15896 7812
rect 15844 7769 15853 7803
rect 15853 7769 15887 7803
rect 15887 7769 15896 7803
rect 15844 7760 15896 7769
rect 16028 7760 16080 7812
rect 16212 7803 16264 7812
rect 16212 7769 16221 7803
rect 16221 7769 16255 7803
rect 16255 7769 16264 7803
rect 16212 7760 16264 7769
rect 7380 7692 7432 7744
rect 11244 7692 11296 7744
rect 12348 7692 12400 7744
rect 14372 7692 14424 7744
rect 19800 7760 19852 7812
rect 21272 7760 21324 7812
rect 18696 7735 18748 7744
rect 18696 7701 18705 7735
rect 18705 7701 18739 7735
rect 18739 7701 18748 7735
rect 18696 7692 18748 7701
rect 4220 7590 4272 7642
rect 4284 7590 4336 7642
rect 4348 7590 4400 7642
rect 4412 7590 4464 7642
rect 4476 7590 4528 7642
rect 9441 7590 9493 7642
rect 9505 7590 9557 7642
rect 9569 7590 9621 7642
rect 9633 7590 9685 7642
rect 9697 7590 9749 7642
rect 14662 7590 14714 7642
rect 14726 7590 14778 7642
rect 14790 7590 14842 7642
rect 14854 7590 14906 7642
rect 14918 7590 14970 7642
rect 19883 7590 19935 7642
rect 19947 7590 19999 7642
rect 20011 7590 20063 7642
rect 20075 7590 20127 7642
rect 20139 7590 20191 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 4436 7488 4488 7540
rect 5264 7488 5316 7540
rect 5448 7488 5500 7540
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 3516 7463 3568 7472
rect 3516 7429 3525 7463
rect 3525 7429 3559 7463
rect 3559 7429 3568 7463
rect 3516 7420 3568 7429
rect 3976 7463 4028 7472
rect 3976 7429 3985 7463
rect 3985 7429 4019 7463
rect 4019 7429 4028 7463
rect 3976 7420 4028 7429
rect 5080 7420 5132 7472
rect 6092 7420 6144 7472
rect 2412 7395 2464 7404
rect 2412 7361 2421 7395
rect 2421 7361 2455 7395
rect 2455 7361 2464 7395
rect 2412 7352 2464 7361
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 3240 7352 3292 7404
rect 3056 7284 3108 7336
rect 3884 7216 3936 7268
rect 4068 7216 4120 7268
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5908 7352 5960 7404
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 7288 7488 7340 7540
rect 8300 7488 8352 7540
rect 8392 7488 8444 7540
rect 9312 7488 9364 7540
rect 10324 7488 10376 7540
rect 7380 7420 7432 7472
rect 7472 7420 7524 7472
rect 9036 7420 9088 7472
rect 9772 7463 9824 7472
rect 9772 7429 9781 7463
rect 9781 7429 9815 7463
rect 9815 7429 9824 7463
rect 9772 7420 9824 7429
rect 15660 7488 15712 7540
rect 15844 7488 15896 7540
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 16856 7531 16908 7540
rect 16856 7497 16865 7531
rect 16865 7497 16899 7531
rect 16899 7497 16908 7531
rect 16856 7488 16908 7497
rect 17040 7531 17092 7540
rect 17040 7497 17049 7531
rect 17049 7497 17083 7531
rect 17083 7497 17092 7531
rect 17040 7488 17092 7497
rect 17960 7488 18012 7540
rect 18972 7488 19024 7540
rect 11980 7420 12032 7472
rect 12900 7463 12952 7472
rect 12900 7429 12909 7463
rect 12909 7429 12943 7463
rect 12943 7429 12952 7463
rect 12900 7420 12952 7429
rect 7656 7352 7708 7404
rect 8576 7352 8628 7404
rect 7748 7216 7800 7268
rect 8300 7216 8352 7268
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 13544 7352 13596 7404
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 9772 7284 9824 7336
rect 12624 7284 12676 7336
rect 9680 7216 9732 7268
rect 9956 7216 10008 7268
rect 11612 7259 11664 7268
rect 11612 7225 11621 7259
rect 11621 7225 11655 7259
rect 11655 7225 11664 7259
rect 11612 7216 11664 7225
rect 15108 7420 15160 7472
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 17592 7352 17644 7404
rect 18696 7420 18748 7472
rect 18788 7420 18840 7472
rect 19708 7488 19760 7540
rect 20996 7531 21048 7540
rect 20996 7497 21005 7531
rect 21005 7497 21039 7531
rect 21039 7497 21048 7531
rect 20996 7488 21048 7497
rect 20536 7463 20588 7472
rect 20536 7429 20545 7463
rect 20545 7429 20579 7463
rect 20579 7429 20588 7463
rect 20536 7420 20588 7429
rect 20628 7420 20680 7472
rect 20720 7463 20772 7472
rect 20720 7429 20729 7463
rect 20729 7429 20763 7463
rect 20763 7429 20772 7463
rect 20720 7420 20772 7429
rect 20812 7463 20864 7472
rect 20812 7429 20821 7463
rect 20821 7429 20855 7463
rect 20855 7429 20864 7463
rect 20812 7420 20864 7429
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 19616 7284 19668 7336
rect 20996 7284 21048 7336
rect 19064 7216 19116 7268
rect 19708 7216 19760 7268
rect 9864 7148 9916 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 14832 7148 14884 7200
rect 18604 7191 18656 7200
rect 18604 7157 18613 7191
rect 18613 7157 18647 7191
rect 18647 7157 18656 7191
rect 18604 7148 18656 7157
rect 19616 7148 19668 7200
rect 3560 7046 3612 7098
rect 3624 7046 3676 7098
rect 3688 7046 3740 7098
rect 3752 7046 3804 7098
rect 3816 7046 3868 7098
rect 8781 7046 8833 7098
rect 8845 7046 8897 7098
rect 8909 7046 8961 7098
rect 8973 7046 9025 7098
rect 9037 7046 9089 7098
rect 14002 7046 14054 7098
rect 14066 7046 14118 7098
rect 14130 7046 14182 7098
rect 14194 7046 14246 7098
rect 14258 7046 14310 7098
rect 19223 7046 19275 7098
rect 19287 7046 19339 7098
rect 19351 7046 19403 7098
rect 19415 7046 19467 7098
rect 19479 7046 19531 7098
rect 2412 6944 2464 6996
rect 4896 6944 4948 6996
rect 7656 6944 7708 6996
rect 18880 6944 18932 6996
rect 20720 6987 20772 6996
rect 20720 6953 20729 6987
rect 20729 6953 20763 6987
rect 20763 6953 20772 6987
rect 20720 6944 20772 6953
rect 1768 6808 1820 6860
rect 1124 6740 1176 6792
rect 2320 6740 2372 6792
rect 2964 6808 3016 6860
rect 5908 6876 5960 6928
rect 3332 6808 3384 6860
rect 5264 6808 5316 6860
rect 5724 6808 5776 6860
rect 6828 6808 6880 6860
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 4712 6740 4764 6792
rect 2964 6715 3016 6724
rect 2964 6681 2973 6715
rect 2973 6681 3007 6715
rect 3007 6681 3016 6715
rect 2964 6672 3016 6681
rect 3148 6715 3200 6724
rect 3148 6681 3157 6715
rect 3157 6681 3191 6715
rect 3191 6681 3200 6715
rect 3148 6672 3200 6681
rect 4804 6715 4856 6724
rect 4804 6681 4813 6715
rect 4813 6681 4847 6715
rect 4847 6681 4856 6715
rect 4804 6672 4856 6681
rect 3056 6604 3108 6656
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 4620 6604 4672 6656
rect 6460 6740 6512 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 7196 6851 7248 6860
rect 7196 6817 7205 6851
rect 7205 6817 7239 6851
rect 7239 6817 7248 6851
rect 7196 6808 7248 6817
rect 9128 6876 9180 6928
rect 9772 6876 9824 6928
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 5172 6672 5224 6724
rect 7932 6672 7984 6724
rect 9588 6672 9640 6724
rect 13912 6808 13964 6860
rect 17040 6808 17092 6860
rect 10048 6672 10100 6724
rect 10232 6740 10284 6792
rect 12440 6740 12492 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 14832 6783 14884 6792
rect 14832 6749 14866 6783
rect 14866 6749 14884 6783
rect 14832 6740 14884 6749
rect 16212 6740 16264 6792
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 20996 6808 21048 6860
rect 10416 6672 10468 6724
rect 10508 6715 10560 6724
rect 10508 6681 10517 6715
rect 10517 6681 10551 6715
rect 10551 6681 10560 6715
rect 10508 6672 10560 6681
rect 12900 6672 12952 6724
rect 13176 6672 13228 6724
rect 5356 6604 5408 6656
rect 5632 6647 5684 6656
rect 5632 6613 5641 6647
rect 5641 6613 5675 6647
rect 5675 6613 5684 6647
rect 5632 6604 5684 6613
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 5816 6604 5868 6656
rect 8392 6604 8444 6656
rect 9404 6604 9456 6656
rect 9772 6604 9824 6656
rect 12164 6647 12216 6656
rect 12164 6613 12173 6647
rect 12173 6613 12207 6647
rect 12207 6613 12216 6647
rect 12164 6604 12216 6613
rect 12256 6604 12308 6656
rect 17040 6672 17092 6724
rect 19064 6672 19116 6724
rect 19432 6672 19484 6724
rect 16948 6604 17000 6656
rect 19156 6604 19208 6656
rect 21088 6672 21140 6724
rect 20720 6604 20772 6656
rect 4220 6502 4272 6554
rect 4284 6502 4336 6554
rect 4348 6502 4400 6554
rect 4412 6502 4464 6554
rect 4476 6502 4528 6554
rect 9441 6502 9493 6554
rect 9505 6502 9557 6554
rect 9569 6502 9621 6554
rect 9633 6502 9685 6554
rect 9697 6502 9749 6554
rect 14662 6502 14714 6554
rect 14726 6502 14778 6554
rect 14790 6502 14842 6554
rect 14854 6502 14906 6554
rect 14918 6502 14970 6554
rect 19883 6502 19935 6554
rect 19947 6502 19999 6554
rect 20011 6502 20063 6554
rect 20075 6502 20127 6554
rect 20139 6502 20191 6554
rect 2780 6400 2832 6452
rect 3240 6400 3292 6452
rect 4620 6400 4672 6452
rect 2320 6239 2372 6248
rect 2320 6205 2329 6239
rect 2329 6205 2363 6239
rect 2363 6205 2372 6239
rect 2320 6196 2372 6205
rect 2872 6264 2924 6316
rect 3424 6264 3476 6316
rect 4344 6196 4396 6248
rect 5356 6400 5408 6452
rect 6552 6400 6604 6452
rect 7012 6400 7064 6452
rect 9220 6400 9272 6452
rect 9864 6400 9916 6452
rect 8300 6375 8352 6384
rect 5356 6264 5408 6316
rect 5448 6264 5500 6316
rect 8300 6341 8334 6375
rect 8334 6341 8352 6375
rect 8300 6332 8352 6341
rect 6460 6264 6512 6316
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 10232 6332 10284 6384
rect 10508 6375 10560 6384
rect 10508 6341 10517 6375
rect 10517 6341 10551 6375
rect 10551 6341 10560 6375
rect 10508 6332 10560 6341
rect 11244 6332 11296 6384
rect 7564 6196 7616 6248
rect 9220 6264 9272 6316
rect 10048 6264 10100 6316
rect 10140 6196 10192 6248
rect 10968 6264 11020 6316
rect 12256 6400 12308 6452
rect 12900 6400 12952 6452
rect 11888 6264 11940 6316
rect 12164 6332 12216 6384
rect 13452 6375 13504 6384
rect 13452 6341 13461 6375
rect 13461 6341 13495 6375
rect 13495 6341 13504 6375
rect 13452 6332 13504 6341
rect 15476 6332 15528 6384
rect 12624 6264 12676 6316
rect 15568 6307 15620 6316
rect 15568 6273 15577 6307
rect 15577 6273 15611 6307
rect 15611 6273 15620 6307
rect 15568 6264 15620 6273
rect 18604 6400 18656 6452
rect 17960 6332 18012 6384
rect 19064 6332 19116 6384
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 13820 6196 13872 6248
rect 14556 6196 14608 6248
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 15292 6196 15344 6248
rect 16028 6196 16080 6248
rect 17132 6196 17184 6248
rect 19156 6307 19208 6316
rect 19156 6273 19165 6307
rect 19165 6273 19199 6307
rect 19199 6273 19208 6307
rect 19156 6264 19208 6273
rect 19616 6307 19668 6316
rect 19616 6273 19625 6307
rect 19625 6273 19659 6307
rect 19659 6273 19668 6307
rect 19616 6264 19668 6273
rect 19064 6196 19116 6248
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 19616 6128 19668 6180
rect 21088 6171 21140 6180
rect 21088 6137 21097 6171
rect 21097 6137 21131 6171
rect 21131 6137 21140 6171
rect 21088 6128 21140 6137
rect 3148 6060 3200 6112
rect 4712 6060 4764 6112
rect 4896 6060 4948 6112
rect 4988 6060 5040 6112
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 12164 6060 12216 6112
rect 13728 6060 13780 6112
rect 15384 6103 15436 6112
rect 15384 6069 15393 6103
rect 15393 6069 15427 6103
rect 15427 6069 15436 6103
rect 15384 6060 15436 6069
rect 17316 6060 17368 6112
rect 18696 6103 18748 6112
rect 18696 6069 18705 6103
rect 18705 6069 18739 6103
rect 18739 6069 18748 6103
rect 18696 6060 18748 6069
rect 19708 6060 19760 6112
rect 3560 5958 3612 6010
rect 3624 5958 3676 6010
rect 3688 5958 3740 6010
rect 3752 5958 3804 6010
rect 3816 5958 3868 6010
rect 8781 5958 8833 6010
rect 8845 5958 8897 6010
rect 8909 5958 8961 6010
rect 8973 5958 9025 6010
rect 9037 5958 9089 6010
rect 14002 5958 14054 6010
rect 14066 5958 14118 6010
rect 14130 5958 14182 6010
rect 14194 5958 14246 6010
rect 14258 5958 14310 6010
rect 19223 5958 19275 6010
rect 19287 5958 19339 6010
rect 19351 5958 19403 6010
rect 19415 5958 19467 6010
rect 19479 5958 19531 6010
rect 2780 5856 2832 5908
rect 4988 5899 5040 5908
rect 4988 5865 4997 5899
rect 4997 5865 5031 5899
rect 5031 5865 5040 5899
rect 4988 5856 5040 5865
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 5632 5856 5684 5908
rect 7932 5899 7984 5908
rect 7932 5865 7941 5899
rect 7941 5865 7975 5899
rect 7975 5865 7984 5899
rect 7932 5856 7984 5865
rect 2688 5695 2740 5704
rect 2688 5661 2706 5695
rect 2706 5661 2740 5695
rect 2688 5652 2740 5661
rect 2872 5652 2924 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4344 5695 4396 5704
rect 4344 5661 4358 5695
rect 4358 5661 4392 5695
rect 4392 5661 4396 5695
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 5816 5763 5868 5772
rect 5816 5729 5842 5763
rect 5842 5729 5868 5763
rect 5816 5720 5868 5729
rect 7564 5788 7616 5840
rect 8576 5856 8628 5908
rect 13912 5856 13964 5908
rect 15108 5856 15160 5908
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 15568 5856 15620 5908
rect 8392 5788 8444 5840
rect 11888 5788 11940 5840
rect 4344 5652 4396 5661
rect 5908 5652 5960 5704
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 4620 5584 4672 5636
rect 7196 5720 7248 5772
rect 6552 5652 6604 5704
rect 7012 5652 7064 5704
rect 8024 5720 8076 5772
rect 9864 5720 9916 5772
rect 8300 5652 8352 5704
rect 8484 5652 8536 5704
rect 11060 5652 11112 5704
rect 11980 5652 12032 5704
rect 12164 5695 12216 5704
rect 12164 5661 12198 5695
rect 12198 5661 12216 5695
rect 12164 5652 12216 5661
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 13820 5652 13872 5704
rect 7380 5584 7432 5636
rect 9956 5584 10008 5636
rect 10048 5584 10100 5636
rect 4712 5516 4764 5568
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 11612 5559 11664 5568
rect 11612 5525 11621 5559
rect 11621 5525 11655 5559
rect 11655 5525 11664 5559
rect 11612 5516 11664 5525
rect 16120 5584 16172 5636
rect 16488 5720 16540 5772
rect 17132 5831 17184 5840
rect 17132 5797 17141 5831
rect 17141 5797 17175 5831
rect 17175 5797 17184 5831
rect 17132 5788 17184 5797
rect 18788 5788 18840 5840
rect 19524 5788 19576 5840
rect 21548 5831 21600 5840
rect 21548 5797 21557 5831
rect 21557 5797 21591 5831
rect 21591 5797 21600 5831
rect 21548 5788 21600 5797
rect 18696 5720 18748 5772
rect 20352 5720 20404 5772
rect 20812 5720 20864 5772
rect 17960 5652 18012 5704
rect 20444 5695 20496 5704
rect 20444 5661 20453 5695
rect 20453 5661 20487 5695
rect 20487 5661 20496 5695
rect 20444 5652 20496 5661
rect 17316 5584 17368 5636
rect 18788 5584 18840 5636
rect 20996 5627 21048 5636
rect 20996 5593 21005 5627
rect 21005 5593 21039 5627
rect 21039 5593 21048 5627
rect 20996 5584 21048 5593
rect 21456 5584 21508 5636
rect 21180 5516 21232 5568
rect 4220 5414 4272 5466
rect 4284 5414 4336 5466
rect 4348 5414 4400 5466
rect 4412 5414 4464 5466
rect 4476 5414 4528 5466
rect 9441 5414 9493 5466
rect 9505 5414 9557 5466
rect 9569 5414 9621 5466
rect 9633 5414 9685 5466
rect 9697 5414 9749 5466
rect 14662 5414 14714 5466
rect 14726 5414 14778 5466
rect 14790 5414 14842 5466
rect 14854 5414 14906 5466
rect 14918 5414 14970 5466
rect 19883 5414 19935 5466
rect 19947 5414 19999 5466
rect 20011 5414 20063 5466
rect 20075 5414 20127 5466
rect 20139 5414 20191 5466
rect 3148 5312 3200 5364
rect 4620 5312 4672 5364
rect 8208 5312 8260 5364
rect 1860 5176 1912 5228
rect 2872 5244 2924 5296
rect 3240 5244 3292 5296
rect 5540 5244 5592 5296
rect 4068 5219 4120 5228
rect 4068 5185 4078 5219
rect 4078 5185 4112 5219
rect 4112 5185 4120 5219
rect 4068 5176 4120 5185
rect 4712 5176 4764 5228
rect 5080 5108 5132 5160
rect 6736 5244 6788 5296
rect 7288 5244 7340 5296
rect 4528 5040 4580 5092
rect 6092 5040 6144 5092
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 7472 5176 7524 5228
rect 8392 5244 8444 5296
rect 10048 5312 10100 5364
rect 11244 5355 11296 5364
rect 11244 5321 11253 5355
rect 11253 5321 11287 5355
rect 11287 5321 11296 5355
rect 11244 5312 11296 5321
rect 9312 5244 9364 5296
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 7748 5108 7800 5160
rect 8668 5176 8720 5228
rect 9128 5176 9180 5228
rect 9864 5219 9916 5228
rect 9864 5185 9873 5219
rect 9873 5185 9907 5219
rect 9907 5185 9916 5219
rect 9864 5176 9916 5185
rect 11612 5244 11664 5296
rect 11796 5244 11848 5296
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 13176 5312 13228 5364
rect 13452 5244 13504 5296
rect 14372 5312 14424 5364
rect 16488 5312 16540 5364
rect 15384 5244 15436 5296
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 17960 5244 18012 5296
rect 18052 5244 18104 5296
rect 12624 5108 12676 5160
rect 11704 5040 11756 5092
rect 6828 4972 6880 5024
rect 11796 4972 11848 5024
rect 13820 4972 13872 5024
rect 16120 4972 16172 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18972 5244 19024 5296
rect 21180 5355 21232 5364
rect 21180 5321 21189 5355
rect 21189 5321 21223 5355
rect 21223 5321 21232 5355
rect 21180 5312 21232 5321
rect 19524 5219 19576 5228
rect 19524 5185 19533 5219
rect 19533 5185 19567 5219
rect 19567 5185 19576 5219
rect 19524 5176 19576 5185
rect 21548 5219 21600 5228
rect 21548 5185 21557 5219
rect 21557 5185 21591 5219
rect 21591 5185 21600 5219
rect 21548 5176 21600 5185
rect 19064 5108 19116 5160
rect 18052 4972 18104 4981
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 3560 4870 3612 4922
rect 3624 4870 3676 4922
rect 3688 4870 3740 4922
rect 3752 4870 3804 4922
rect 3816 4870 3868 4922
rect 8781 4870 8833 4922
rect 8845 4870 8897 4922
rect 8909 4870 8961 4922
rect 8973 4870 9025 4922
rect 9037 4870 9089 4922
rect 14002 4870 14054 4922
rect 14066 4870 14118 4922
rect 14130 4870 14182 4922
rect 14194 4870 14246 4922
rect 14258 4870 14310 4922
rect 19223 4870 19275 4922
rect 19287 4870 19339 4922
rect 19351 4870 19403 4922
rect 19415 4870 19467 4922
rect 19479 4870 19531 4922
rect 4804 4768 4856 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 9220 4768 9272 4820
rect 13452 4811 13504 4820
rect 13452 4777 13461 4811
rect 13461 4777 13495 4811
rect 13495 4777 13504 4811
rect 13452 4768 13504 4777
rect 21548 4811 21600 4820
rect 21548 4777 21557 4811
rect 21557 4777 21591 4811
rect 21591 4777 21600 4811
rect 21548 4768 21600 4777
rect 2872 4564 2924 4616
rect 3424 4564 3476 4616
rect 3792 4496 3844 4548
rect 4804 4496 4856 4548
rect 4068 4428 4120 4480
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 5264 4607 5316 4616
rect 5264 4573 5273 4607
rect 5273 4573 5307 4607
rect 5307 4573 5316 4607
rect 5264 4564 5316 4573
rect 5448 4564 5500 4616
rect 5632 4607 5684 4616
rect 5632 4573 5666 4607
rect 5666 4573 5684 4607
rect 5632 4564 5684 4573
rect 8208 4700 8260 4752
rect 6828 4632 6880 4684
rect 8484 4632 8536 4684
rect 8668 4632 8720 4684
rect 9772 4564 9824 4616
rect 11704 4564 11756 4616
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 16580 4700 16632 4752
rect 18696 4564 18748 4616
rect 19064 4564 19116 4616
rect 21364 4564 21416 4616
rect 4988 4539 5040 4548
rect 4988 4505 4997 4539
rect 4997 4505 5031 4539
rect 5031 4505 5040 4539
rect 4988 4496 5040 4505
rect 7288 4539 7340 4548
rect 7288 4505 7297 4539
rect 7297 4505 7331 4539
rect 7331 4505 7340 4539
rect 7288 4496 7340 4505
rect 6828 4428 6880 4480
rect 7104 4428 7156 4480
rect 8484 4496 8536 4548
rect 8760 4496 8812 4548
rect 9312 4428 9364 4480
rect 11704 4471 11756 4480
rect 11704 4437 11713 4471
rect 11713 4437 11747 4471
rect 11747 4437 11756 4471
rect 11704 4428 11756 4437
rect 17960 4471 18012 4480
rect 17960 4437 17969 4471
rect 17969 4437 18003 4471
rect 18003 4437 18012 4471
rect 17960 4428 18012 4437
rect 4220 4326 4272 4378
rect 4284 4326 4336 4378
rect 4348 4326 4400 4378
rect 4412 4326 4464 4378
rect 4476 4326 4528 4378
rect 9441 4326 9493 4378
rect 9505 4326 9557 4378
rect 9569 4326 9621 4378
rect 9633 4326 9685 4378
rect 9697 4326 9749 4378
rect 14662 4326 14714 4378
rect 14726 4326 14778 4378
rect 14790 4326 14842 4378
rect 14854 4326 14906 4378
rect 14918 4326 14970 4378
rect 19883 4326 19935 4378
rect 19947 4326 19999 4378
rect 20011 4326 20063 4378
rect 20075 4326 20127 4378
rect 20139 4326 20191 4378
rect 5264 4224 5316 4276
rect 8760 4224 8812 4276
rect 13544 4224 13596 4276
rect 13728 4224 13780 4276
rect 2964 4156 3016 4208
rect 3148 4156 3200 4208
rect 5080 4156 5132 4208
rect 6920 4199 6972 4208
rect 6920 4165 6929 4199
rect 6929 4165 6963 4199
rect 6963 4165 6972 4199
rect 6920 4156 6972 4165
rect 2780 4088 2832 4140
rect 3884 4088 3936 4140
rect 4712 4088 4764 4140
rect 5816 4088 5868 4140
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 7288 4156 7340 4208
rect 10416 4156 10468 4208
rect 11152 4199 11204 4208
rect 11152 4165 11161 4199
rect 11161 4165 11195 4199
rect 11195 4165 11204 4199
rect 11152 4156 11204 4165
rect 11704 4156 11756 4208
rect 14372 4224 14424 4276
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 2320 4063 2372 4072
rect 2320 4029 2329 4063
rect 2329 4029 2363 4063
rect 2363 4029 2372 4063
rect 2320 4020 2372 4029
rect 2964 3952 3016 4004
rect 3792 3952 3844 4004
rect 3976 3952 4028 4004
rect 5632 4020 5684 4072
rect 6828 4020 6880 4072
rect 7932 4131 7984 4140
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 8576 4088 8628 4140
rect 9128 4088 9180 4140
rect 9496 4020 9548 4072
rect 10140 4020 10192 4072
rect 4804 3952 4856 4004
rect 7012 3952 7064 4004
rect 7748 3995 7800 4004
rect 7748 3961 7757 3995
rect 7757 3961 7791 3995
rect 7791 3961 7800 3995
rect 7748 3952 7800 3961
rect 10968 4020 11020 4072
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 1676 3884 1728 3936
rect 1860 3884 1912 3936
rect 3148 3884 3200 3936
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5908 3884 5960 3936
rect 8300 3884 8352 3936
rect 10140 3884 10192 3936
rect 11060 3884 11112 3936
rect 14556 4088 14608 4140
rect 14740 4199 14792 4208
rect 14740 4165 14749 4199
rect 14749 4165 14783 4199
rect 14783 4165 14792 4199
rect 14740 4156 14792 4165
rect 15292 4224 15344 4276
rect 18052 4224 18104 4276
rect 18972 4224 19024 4276
rect 13728 4020 13780 4072
rect 15108 4088 15160 4140
rect 15292 4131 15344 4140
rect 15292 4097 15326 4131
rect 15326 4097 15344 4131
rect 15292 4088 15344 4097
rect 18236 4156 18288 4208
rect 16304 4088 16356 4140
rect 18052 4088 18104 4140
rect 20628 4156 20680 4208
rect 13820 3952 13872 4004
rect 16580 3952 16632 4004
rect 18512 4063 18564 4072
rect 18512 4029 18521 4063
rect 18521 4029 18555 4063
rect 18555 4029 18564 4063
rect 18512 4020 18564 4029
rect 13912 3927 13964 3936
rect 13912 3893 13921 3927
rect 13921 3893 13955 3927
rect 13955 3893 13964 3927
rect 13912 3884 13964 3893
rect 16856 3884 16908 3936
rect 16948 3884 17000 3936
rect 19064 3884 19116 3936
rect 19708 3952 19760 4004
rect 19892 4020 19944 4072
rect 20904 3952 20956 4004
rect 20996 3884 21048 3936
rect 3560 3782 3612 3834
rect 3624 3782 3676 3834
rect 3688 3782 3740 3834
rect 3752 3782 3804 3834
rect 3816 3782 3868 3834
rect 8781 3782 8833 3834
rect 8845 3782 8897 3834
rect 8909 3782 8961 3834
rect 8973 3782 9025 3834
rect 9037 3782 9089 3834
rect 14002 3782 14054 3834
rect 14066 3782 14118 3834
rect 14130 3782 14182 3834
rect 14194 3782 14246 3834
rect 14258 3782 14310 3834
rect 19223 3782 19275 3834
rect 19287 3782 19339 3834
rect 19351 3782 19403 3834
rect 19415 3782 19467 3834
rect 19479 3782 19531 3834
rect 5264 3680 5316 3732
rect 6920 3680 6972 3732
rect 7932 3680 7984 3732
rect 14740 3680 14792 3732
rect 15016 3680 15068 3732
rect 8116 3655 8168 3664
rect 8116 3621 8125 3655
rect 8125 3621 8159 3655
rect 8159 3621 8168 3655
rect 8116 3612 8168 3621
rect 3700 3544 3752 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 2872 3476 2924 3528
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 4896 3476 4948 3528
rect 6460 3476 6512 3528
rect 1952 3408 2004 3460
rect 2872 3340 2924 3392
rect 4160 3408 4212 3460
rect 5356 3408 5408 3460
rect 5724 3451 5776 3460
rect 5724 3417 5758 3451
rect 5758 3417 5776 3451
rect 5724 3408 5776 3417
rect 6000 3408 6052 3460
rect 7472 3408 7524 3460
rect 8484 3476 8536 3528
rect 9772 3544 9824 3596
rect 10140 3519 10192 3528
rect 10140 3485 10174 3519
rect 10174 3485 10192 3519
rect 10140 3476 10192 3485
rect 11336 3476 11388 3528
rect 13360 3612 13412 3664
rect 16764 3612 16816 3664
rect 12532 3587 12584 3596
rect 12532 3553 12541 3587
rect 12541 3553 12575 3587
rect 12575 3553 12584 3587
rect 12532 3544 12584 3553
rect 13820 3544 13872 3596
rect 3608 3383 3660 3392
rect 3608 3349 3617 3383
rect 3617 3349 3651 3383
rect 3651 3349 3660 3383
rect 3608 3340 3660 3349
rect 4988 3340 5040 3392
rect 5632 3340 5684 3392
rect 8392 3451 8444 3460
rect 8392 3417 8401 3451
rect 8401 3417 8435 3451
rect 8435 3417 8444 3451
rect 8392 3408 8444 3417
rect 9496 3451 9548 3460
rect 9496 3417 9505 3451
rect 9505 3417 9539 3451
rect 9539 3417 9548 3451
rect 9496 3408 9548 3417
rect 9864 3408 9916 3460
rect 11520 3408 11572 3460
rect 12072 3408 12124 3460
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 15108 3544 15160 3596
rect 16856 3544 16908 3596
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 18972 3680 19024 3732
rect 20628 3723 20680 3732
rect 20628 3689 20637 3723
rect 20637 3689 20671 3723
rect 20671 3689 20680 3723
rect 20628 3680 20680 3689
rect 20904 3723 20956 3732
rect 20904 3689 20913 3723
rect 20913 3689 20947 3723
rect 20947 3689 20956 3723
rect 20904 3680 20956 3689
rect 21364 3587 21416 3596
rect 21364 3553 21373 3587
rect 21373 3553 21407 3587
rect 21407 3553 21416 3587
rect 21364 3544 21416 3553
rect 12624 3451 12676 3460
rect 12624 3417 12633 3451
rect 12633 3417 12667 3451
rect 12667 3417 12676 3451
rect 12624 3408 12676 3417
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 10968 3340 11020 3392
rect 11428 3383 11480 3392
rect 11428 3349 11437 3383
rect 11437 3349 11471 3383
rect 11471 3349 11480 3383
rect 11428 3340 11480 3349
rect 11796 3340 11848 3392
rect 12992 3383 13044 3392
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 13176 3451 13228 3460
rect 13176 3417 13185 3451
rect 13185 3417 13219 3451
rect 13219 3417 13228 3451
rect 13176 3408 13228 3417
rect 13728 3340 13780 3392
rect 15568 3408 15620 3460
rect 16672 3408 16724 3460
rect 18696 3408 18748 3460
rect 20996 3476 21048 3528
rect 19708 3408 19760 3460
rect 17040 3383 17092 3392
rect 17040 3349 17049 3383
rect 17049 3349 17083 3383
rect 17083 3349 17092 3383
rect 17040 3340 17092 3349
rect 18236 3383 18288 3392
rect 18236 3349 18245 3383
rect 18245 3349 18279 3383
rect 18279 3349 18288 3383
rect 18236 3340 18288 3349
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 20628 3340 20680 3392
rect 4220 3238 4272 3290
rect 4284 3238 4336 3290
rect 4348 3238 4400 3290
rect 4412 3238 4464 3290
rect 4476 3238 4528 3290
rect 9441 3238 9493 3290
rect 9505 3238 9557 3290
rect 9569 3238 9621 3290
rect 9633 3238 9685 3290
rect 9697 3238 9749 3290
rect 14662 3238 14714 3290
rect 14726 3238 14778 3290
rect 14790 3238 14842 3290
rect 14854 3238 14906 3290
rect 14918 3238 14970 3290
rect 19883 3238 19935 3290
rect 19947 3238 19999 3290
rect 20011 3238 20063 3290
rect 20075 3238 20127 3290
rect 20139 3238 20191 3290
rect 3056 3136 3108 3188
rect 5080 3179 5132 3188
rect 5080 3145 5089 3179
rect 5089 3145 5123 3179
rect 5123 3145 5132 3179
rect 5080 3136 5132 3145
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 7472 3136 7524 3188
rect 9312 3136 9364 3188
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 1676 3068 1728 3120
rect 3608 3068 3660 3120
rect 5448 3068 5500 3120
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 7288 3068 7340 3120
rect 8300 3111 8352 3120
rect 8300 3077 8334 3111
rect 8334 3077 8352 3111
rect 8300 3068 8352 3077
rect 11428 3068 11480 3120
rect 12532 3068 12584 3120
rect 13912 3068 13964 3120
rect 15568 3179 15620 3188
rect 15568 3145 15577 3179
rect 15577 3145 15611 3179
rect 15611 3145 15620 3179
rect 15568 3136 15620 3145
rect 17040 3136 17092 3188
rect 18236 3136 18288 3188
rect 19800 3136 19852 3188
rect 21364 3136 21416 3188
rect 18880 3068 18932 3120
rect 19064 3068 19116 3120
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 13360 3043 13412 3052
rect 13360 3009 13369 3043
rect 13369 3009 13403 3043
rect 13403 3009 13412 3043
rect 13360 3000 13412 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 11520 2932 11572 2984
rect 12900 2864 12952 2916
rect 13176 2864 13228 2916
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 5356 2796 5408 2848
rect 9128 2796 9180 2848
rect 15476 2796 15528 2848
rect 17132 2839 17184 2848
rect 17132 2805 17141 2839
rect 17141 2805 17175 2839
rect 17175 2805 17184 2839
rect 17132 2796 17184 2805
rect 3560 2694 3612 2746
rect 3624 2694 3676 2746
rect 3688 2694 3740 2746
rect 3752 2694 3804 2746
rect 3816 2694 3868 2746
rect 8781 2694 8833 2746
rect 8845 2694 8897 2746
rect 8909 2694 8961 2746
rect 8973 2694 9025 2746
rect 9037 2694 9089 2746
rect 14002 2694 14054 2746
rect 14066 2694 14118 2746
rect 14130 2694 14182 2746
rect 14194 2694 14246 2746
rect 14258 2694 14310 2746
rect 19223 2694 19275 2746
rect 19287 2694 19339 2746
rect 19351 2694 19403 2746
rect 19415 2694 19467 2746
rect 19479 2694 19531 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 4620 2592 4672 2644
rect 8576 2592 8628 2644
rect 11336 2592 11388 2644
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 4988 2524 5040 2576
rect 12624 2592 12676 2644
rect 12992 2592 13044 2644
rect 14556 2635 14608 2644
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 15292 2592 15344 2644
rect 3056 2456 3108 2508
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 7288 2499 7340 2508
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 11520 2499 11572 2508
rect 11520 2465 11529 2499
rect 11529 2465 11563 2499
rect 11563 2465 11572 2499
rect 11520 2456 11572 2465
rect 15476 2456 15528 2508
rect 5356 2388 5408 2440
rect 8116 2388 8168 2440
rect 11060 2388 11112 2440
rect 11796 2431 11848 2440
rect 11796 2397 11830 2431
rect 11830 2397 11848 2431
rect 11796 2388 11848 2397
rect 13820 2388 13872 2440
rect 16764 2388 16816 2440
rect 18696 2388 18748 2440
rect 2872 2363 2924 2372
rect 2872 2329 2881 2363
rect 2881 2329 2915 2363
rect 2915 2329 2924 2363
rect 2872 2320 2924 2329
rect 15016 2363 15068 2372
rect 15016 2329 15025 2363
rect 15025 2329 15059 2363
rect 15059 2329 15068 2363
rect 15016 2320 15068 2329
rect 17132 2320 17184 2372
rect 11152 2252 11204 2304
rect 18512 2252 18564 2304
rect 18696 2252 18748 2304
rect 4220 2150 4272 2202
rect 4284 2150 4336 2202
rect 4348 2150 4400 2202
rect 4412 2150 4464 2202
rect 4476 2150 4528 2202
rect 9441 2150 9493 2202
rect 9505 2150 9557 2202
rect 9569 2150 9621 2202
rect 9633 2150 9685 2202
rect 9697 2150 9749 2202
rect 14662 2150 14714 2202
rect 14726 2150 14778 2202
rect 14790 2150 14842 2202
rect 14854 2150 14906 2202
rect 14918 2150 14970 2202
rect 19883 2150 19935 2202
rect 19947 2150 19999 2202
rect 20011 2150 20063 2202
rect 20075 2150 20127 2202
rect 20139 2150 20191 2202
<< metal2 >>
rect 5170 24475 5226 25275
rect 5814 24475 5870 25275
rect 7102 24475 7158 25275
rect 7746 24475 7802 25275
rect 9034 24475 9090 25275
rect 9678 24475 9734 25275
rect 10966 24475 11022 25275
rect 11348 24534 11560 24562
rect 4220 22876 4528 22885
rect 4220 22874 4226 22876
rect 4282 22874 4306 22876
rect 4362 22874 4386 22876
rect 4442 22874 4466 22876
rect 4522 22874 4528 22876
rect 4282 22822 4284 22874
rect 4464 22822 4466 22874
rect 4220 22820 4226 22822
rect 4282 22820 4306 22822
rect 4362 22820 4386 22822
rect 4442 22820 4466 22822
rect 4522 22820 4528 22822
rect 4220 22811 4528 22820
rect 3056 22704 3108 22710
rect 3056 22646 3108 22652
rect 2780 22568 2832 22574
rect 2832 22528 2912 22556
rect 2780 22510 2832 22516
rect 2044 22432 2096 22438
rect 2044 22374 2096 22380
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2056 22030 2084 22374
rect 2792 22114 2820 22374
rect 2700 22086 2820 22114
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1688 21554 1716 21830
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1952 21072 2004 21078
rect 1952 21014 2004 21020
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1688 20058 1716 20402
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1964 19854 1992 21014
rect 2700 20874 2728 22086
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2792 21622 2820 21966
rect 2780 21616 2832 21622
rect 2780 21558 2832 21564
rect 2412 20868 2464 20874
rect 2412 20810 2464 20816
rect 2688 20868 2740 20874
rect 2688 20810 2740 20816
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 1952 19848 2004 19854
rect 1952 19790 2004 19796
rect 2056 19378 2084 20198
rect 2320 19780 2372 19786
rect 2320 19722 2372 19728
rect 2332 19514 2360 19722
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 1306 19136 1362 19145
rect 1306 19071 1362 19080
rect 1320 18970 1348 19071
rect 1308 18964 1360 18970
rect 1308 18906 1360 18912
rect 1320 18358 1348 18906
rect 1492 18692 1544 18698
rect 1492 18634 1544 18640
rect 1504 18426 1532 18634
rect 1492 18420 1544 18426
rect 1492 18362 1544 18368
rect 1308 18352 1360 18358
rect 1308 18294 1360 18300
rect 2424 18222 2452 20810
rect 2596 20800 2648 20806
rect 2596 20742 2648 20748
rect 2608 20482 2636 20742
rect 2792 20534 2820 21558
rect 2884 21078 2912 22528
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2976 21690 3004 21898
rect 3068 21865 3096 22646
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 3560 22332 3868 22341
rect 3560 22330 3566 22332
rect 3622 22330 3646 22332
rect 3702 22330 3726 22332
rect 3782 22330 3806 22332
rect 3862 22330 3868 22332
rect 3622 22278 3624 22330
rect 3804 22278 3806 22330
rect 3560 22276 3566 22278
rect 3622 22276 3646 22278
rect 3702 22276 3726 22278
rect 3782 22276 3806 22278
rect 3862 22276 3868 22278
rect 3560 22267 3868 22276
rect 3976 22092 4028 22098
rect 4816 22094 4844 22510
rect 3976 22034 4028 22040
rect 4632 22066 4844 22094
rect 3884 21888 3936 21894
rect 3054 21856 3110 21865
rect 3884 21830 3936 21836
rect 3054 21791 3110 21800
rect 2964 21684 3016 21690
rect 2964 21626 3016 21632
rect 3068 21418 3096 21791
rect 3896 21486 3924 21830
rect 3988 21486 4016 22034
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4080 21622 4108 21966
rect 4632 21894 4660 22066
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4220 21788 4528 21797
rect 4220 21786 4226 21788
rect 4282 21786 4306 21788
rect 4362 21786 4386 21788
rect 4442 21786 4466 21788
rect 4522 21786 4528 21788
rect 4282 21734 4284 21786
rect 4464 21734 4466 21786
rect 4220 21732 4226 21734
rect 4282 21732 4306 21734
rect 4362 21732 4386 21734
rect 4442 21732 4466 21734
rect 4522 21732 4528 21734
rect 4220 21723 4528 21732
rect 4068 21616 4120 21622
rect 4068 21558 4120 21564
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 3056 21412 3108 21418
rect 3056 21354 3108 21360
rect 3560 21244 3868 21253
rect 3560 21242 3566 21244
rect 3622 21242 3646 21244
rect 3702 21242 3726 21244
rect 3782 21242 3806 21244
rect 3862 21242 3868 21244
rect 3622 21190 3624 21242
rect 3804 21190 3806 21242
rect 3560 21188 3566 21190
rect 3622 21188 3646 21190
rect 3702 21188 3726 21190
rect 3782 21188 3806 21190
rect 3862 21188 3868 21190
rect 3560 21179 3868 21188
rect 2872 21072 2924 21078
rect 2872 21014 2924 21020
rect 3896 20942 3924 21422
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3988 20534 4016 21422
rect 4632 21010 4660 21830
rect 4804 21616 4856 21622
rect 4804 21558 4856 21564
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4540 20874 4752 20890
rect 4528 20868 4752 20874
rect 4580 20862 4752 20868
rect 4724 20856 4752 20862
rect 4816 20856 4844 21558
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4724 20828 4844 20856
rect 4528 20810 4580 20816
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 4220 20700 4528 20709
rect 4220 20698 4226 20700
rect 4282 20698 4306 20700
rect 4362 20698 4386 20700
rect 4442 20698 4466 20700
rect 4522 20698 4528 20700
rect 4282 20646 4284 20698
rect 4464 20646 4466 20698
rect 4220 20644 4226 20646
rect 4282 20644 4306 20646
rect 4362 20644 4386 20646
rect 4442 20644 4466 20646
rect 4522 20644 4528 20646
rect 4220 20635 4528 20644
rect 4632 20602 4660 20742
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 2780 20528 2832 20534
rect 2686 20496 2742 20505
rect 2608 20454 2686 20482
rect 2780 20470 2832 20476
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 2686 20431 2742 20440
rect 2700 20330 2728 20431
rect 2688 20324 2740 20330
rect 2688 20266 2740 20272
rect 2792 19854 2820 20470
rect 3988 20346 4016 20470
rect 3988 20318 4108 20346
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3560 20156 3868 20165
rect 3560 20154 3566 20156
rect 3622 20154 3646 20156
rect 3702 20154 3726 20156
rect 3782 20154 3806 20156
rect 3862 20154 3868 20156
rect 3622 20102 3624 20154
rect 3804 20102 3806 20154
rect 3560 20100 3566 20102
rect 3622 20100 3646 20102
rect 3702 20100 3726 20102
rect 3782 20100 3806 20102
rect 3862 20100 3868 20102
rect 3560 20091 3868 20100
rect 3988 19854 4016 20198
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 2792 19446 2820 19790
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3804 19446 3832 19654
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 2504 18896 2556 18902
rect 2504 18838 2556 18844
rect 2516 18290 2544 18838
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2700 18426 2728 18770
rect 2792 18766 2820 19382
rect 3056 19372 3108 19378
rect 3056 19314 3108 19320
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2792 18358 2820 18702
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1872 17338 1900 17614
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1964 17066 1992 17546
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1676 16516 1728 16522
rect 1676 16458 1728 16464
rect 1688 16250 1716 16458
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 2424 16046 2452 18158
rect 2778 17776 2834 17785
rect 2778 17711 2834 17720
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2700 16590 2728 17274
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2700 16046 2728 16526
rect 2792 16454 2820 17711
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2884 17270 2912 17546
rect 3068 17270 3096 19314
rect 3560 19068 3868 19077
rect 3560 19066 3566 19068
rect 3622 19066 3646 19068
rect 3702 19066 3726 19068
rect 3782 19066 3806 19068
rect 3862 19066 3868 19068
rect 3622 19014 3624 19066
rect 3804 19014 3806 19066
rect 3560 19012 3566 19014
rect 3622 19012 3646 19014
rect 3702 19012 3726 19014
rect 3782 19012 3806 19014
rect 3862 19012 3868 19014
rect 3560 19003 3868 19012
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 17882 3280 18566
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3560 17980 3868 17989
rect 3560 17978 3566 17980
rect 3622 17978 3646 17980
rect 3702 17978 3726 17980
rect 3782 17978 3806 17980
rect 3862 17978 3868 17980
rect 3622 17926 3624 17978
rect 3804 17926 3806 17978
rect 3560 17924 3566 17926
rect 3622 17924 3646 17926
rect 3702 17924 3726 17926
rect 3782 17924 3806 17926
rect 3862 17924 3868 17926
rect 3560 17915 3868 17924
rect 3988 17882 4016 18226
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 2872 17264 2924 17270
rect 3056 17264 3108 17270
rect 2872 17206 2924 17212
rect 3054 17232 3056 17241
rect 3108 17232 3110 17241
rect 3252 17202 3280 17818
rect 3054 17167 3110 17176
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 4080 17134 4108 20318
rect 4172 20058 4200 20538
rect 4712 20528 4764 20534
rect 4712 20470 4764 20476
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4220 19612 4528 19621
rect 4220 19610 4226 19612
rect 4282 19610 4306 19612
rect 4362 19610 4386 19612
rect 4442 19610 4466 19612
rect 4522 19610 4528 19612
rect 4282 19558 4284 19610
rect 4464 19558 4466 19610
rect 4220 19556 4226 19558
rect 4282 19556 4306 19558
rect 4362 19556 4386 19558
rect 4442 19556 4466 19558
rect 4522 19556 4528 19558
rect 4220 19547 4528 19556
rect 4632 19514 4660 20334
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4724 19378 4752 20470
rect 4816 20346 4844 20828
rect 4908 20466 4936 20878
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 5000 20398 5028 20810
rect 5184 20602 5212 24475
rect 5828 22522 5856 24475
rect 7116 22778 7144 24475
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 5736 22494 5856 22522
rect 5448 22432 5500 22438
rect 5448 22374 5500 22380
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5276 21350 5304 21626
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 5368 21418 5396 21558
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5460 20942 5488 22374
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5552 21078 5580 21558
rect 5644 21146 5672 21966
rect 5736 21690 5764 22494
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5828 22030 5856 22374
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5540 21072 5592 21078
rect 5540 21014 5592 21020
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 5552 20534 5580 21014
rect 5736 20942 5764 21626
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5828 21146 5856 21490
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 6012 21010 6040 21626
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6000 21004 6052 21010
rect 6104 20992 6132 21286
rect 6380 21010 6408 21286
rect 6368 21004 6420 21010
rect 6104 20964 6224 20992
rect 6000 20946 6052 20952
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5644 20618 5672 20878
rect 5644 20602 5764 20618
rect 5920 20602 5948 20878
rect 6092 20868 6144 20874
rect 6092 20810 6144 20816
rect 5632 20596 5764 20602
rect 5684 20590 5764 20596
rect 5632 20538 5684 20544
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 4988 20392 5040 20398
rect 4816 20318 4936 20346
rect 4988 20334 5040 20340
rect 4802 19816 4858 19825
rect 4802 19751 4858 19760
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4724 18970 4752 19314
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4220 18524 4528 18533
rect 4220 18522 4226 18524
rect 4282 18522 4306 18524
rect 4362 18522 4386 18524
rect 4442 18522 4466 18524
rect 4522 18522 4528 18524
rect 4282 18470 4284 18522
rect 4464 18470 4466 18522
rect 4220 18468 4226 18470
rect 4282 18468 4306 18470
rect 4362 18468 4386 18470
rect 4442 18468 4466 18470
rect 4522 18468 4528 18470
rect 4220 18459 4528 18468
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4356 18329 4384 18362
rect 4342 18320 4398 18329
rect 4342 18255 4398 18264
rect 4356 17882 4384 18255
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4632 17746 4660 18770
rect 4816 17762 4844 19751
rect 4908 18698 4936 20318
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4724 17734 4844 17762
rect 4724 17542 4752 17734
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4220 17436 4528 17445
rect 4220 17434 4226 17436
rect 4282 17434 4306 17436
rect 4362 17434 4386 17436
rect 4442 17434 4466 17436
rect 4522 17434 4528 17436
rect 4282 17382 4284 17434
rect 4464 17382 4466 17434
rect 4220 17380 4226 17382
rect 4282 17380 4306 17382
rect 4362 17380 4386 17382
rect 4442 17380 4466 17382
rect 4522 17380 4528 17382
rect 4220 17371 4528 17380
rect 4724 17134 4752 17478
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 3560 16892 3868 16901
rect 3560 16890 3566 16892
rect 3622 16890 3646 16892
rect 3702 16890 3726 16892
rect 3782 16890 3806 16892
rect 3862 16890 3868 16892
rect 3622 16838 3624 16890
rect 3804 16838 3806 16890
rect 3560 16836 3566 16838
rect 3622 16836 3646 16838
rect 3702 16836 3726 16838
rect 3782 16836 3806 16838
rect 3862 16836 3868 16838
rect 3560 16827 3868 16836
rect 4080 16658 4108 17070
rect 4724 16658 4752 17070
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 2792 16250 2820 16390
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2700 15502 2728 15982
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2700 14498 2728 15438
rect 2884 14890 2912 16050
rect 2976 15434 3004 16390
rect 3436 16182 3464 16390
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3560 15804 3868 15813
rect 3560 15802 3566 15804
rect 3622 15802 3646 15804
rect 3702 15802 3726 15804
rect 3782 15802 3806 15804
rect 3862 15802 3868 15804
rect 3622 15750 3624 15802
rect 3804 15750 3806 15802
rect 3560 15748 3566 15750
rect 3622 15748 3646 15750
rect 3702 15748 3726 15750
rect 3782 15748 3806 15750
rect 3862 15748 3868 15750
rect 3146 15736 3202 15745
rect 3560 15739 3868 15748
rect 3896 15706 3924 16526
rect 4220 16348 4528 16357
rect 4220 16346 4226 16348
rect 4282 16346 4306 16348
rect 4362 16346 4386 16348
rect 4442 16346 4466 16348
rect 4522 16346 4528 16348
rect 4282 16294 4284 16346
rect 4464 16294 4466 16346
rect 4220 16292 4226 16294
rect 4282 16292 4306 16294
rect 4362 16292 4386 16294
rect 4442 16292 4466 16294
rect 4522 16292 4528 16294
rect 4220 16283 4528 16292
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 3146 15671 3202 15680
rect 3884 15700 3936 15706
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2872 14884 2924 14890
rect 2872 14826 2924 14832
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2608 14482 2728 14498
rect 2596 14476 2728 14482
rect 2648 14470 2728 14476
rect 2596 14418 2648 14424
rect 1584 14340 1636 14346
rect 1584 14282 1636 14288
rect 1596 14074 1624 14282
rect 2700 14074 2728 14470
rect 2976 14414 3004 14758
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2044 14000 2096 14006
rect 2044 13942 2096 13948
rect 2056 13258 2084 13942
rect 2700 13394 2728 14010
rect 2884 14006 2912 14214
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13530 2820 13874
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 2870 13016 2926 13025
rect 3068 12986 3096 13194
rect 2870 12951 2926 12960
rect 3056 12980 3108 12986
rect 2778 12336 2834 12345
rect 2884 12306 2912 12951
rect 3056 12922 3108 12928
rect 2778 12271 2834 12280
rect 2872 12300 2924 12306
rect 2792 12238 2820 12271
rect 2872 12242 2924 12248
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 2872 12096 2924 12102
rect 2924 12056 3004 12084
rect 2872 12038 2924 12044
rect 1872 11762 1900 12038
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 2976 11558 3004 12056
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 11150 3004 11494
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 1688 10606 1716 11086
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1306 10296 1362 10305
rect 1306 10231 1362 10240
rect 1320 9994 1348 10231
rect 1308 9988 1360 9994
rect 1308 9930 1360 9936
rect 1308 9648 1360 9654
rect 1308 9590 1360 9596
rect 1320 8945 1348 9590
rect 1688 8974 1716 10542
rect 1964 10266 1992 10610
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2884 9926 2912 10406
rect 3068 10062 3096 12106
rect 3160 10266 3188 15671
rect 3884 15642 3936 15648
rect 4264 15570 4292 16186
rect 4632 15638 4660 16594
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4264 15348 4292 15506
rect 4080 15320 4292 15348
rect 4080 15094 4108 15320
rect 4220 15260 4528 15269
rect 4220 15258 4226 15260
rect 4282 15258 4306 15260
rect 4362 15258 4386 15260
rect 4442 15258 4466 15260
rect 4522 15258 4528 15260
rect 4282 15206 4284 15258
rect 4464 15206 4466 15258
rect 4220 15204 4226 15206
rect 4282 15204 4306 15206
rect 4362 15204 4386 15206
rect 4442 15204 4466 15206
rect 4522 15204 4528 15206
rect 4220 15195 4528 15204
rect 4632 15162 4660 15574
rect 4724 15434 4752 16390
rect 4816 16250 4844 17614
rect 5000 17610 5028 20334
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5092 19786 5120 20198
rect 5368 19990 5396 20470
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5644 20058 5672 20402
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 5460 19514 5488 19858
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 4988 17604 5040 17610
rect 4988 17546 5040 17552
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4908 16561 4936 17206
rect 4894 16552 4950 16561
rect 4894 16487 4950 16496
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3252 14006 3280 14282
rect 3344 14278 3372 14418
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 3344 13326 3372 14214
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3436 13258 3464 14962
rect 3560 14716 3868 14725
rect 3560 14714 3566 14716
rect 3622 14714 3646 14716
rect 3702 14714 3726 14716
rect 3782 14714 3806 14716
rect 3862 14714 3868 14716
rect 3622 14662 3624 14714
rect 3804 14662 3806 14714
rect 3560 14660 3566 14662
rect 3622 14660 3646 14662
rect 3702 14660 3726 14662
rect 3782 14660 3806 14662
rect 3862 14660 3868 14662
rect 3560 14651 3868 14660
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 3560 13628 3868 13637
rect 3560 13626 3566 13628
rect 3622 13626 3646 13628
rect 3702 13626 3726 13628
rect 3782 13626 3806 13628
rect 3862 13626 3868 13628
rect 3622 13574 3624 13626
rect 3804 13574 3806 13626
rect 3560 13572 3566 13574
rect 3622 13572 3646 13574
rect 3702 13572 3726 13574
rect 3782 13572 3806 13574
rect 3862 13572 3868 13574
rect 3560 13563 3868 13572
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3436 12850 3464 13194
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3804 12646 3832 13262
rect 3988 13190 4016 14350
rect 4220 14172 4528 14181
rect 4220 14170 4226 14172
rect 4282 14170 4306 14172
rect 4362 14170 4386 14172
rect 4442 14170 4466 14172
rect 4522 14170 4528 14172
rect 4282 14118 4284 14170
rect 4464 14118 4466 14170
rect 4220 14116 4226 14118
rect 4282 14116 4306 14118
rect 4362 14116 4386 14118
rect 4442 14116 4466 14118
rect 4522 14116 4528 14118
rect 4220 14107 4528 14116
rect 4632 14006 4660 14350
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4540 13530 4568 13942
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4528 13320 4580 13326
rect 4632 13274 4660 13942
rect 4724 13870 4752 14282
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4724 13394 4752 13806
rect 4816 13530 4844 15914
rect 4908 15910 4936 16487
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 5000 15570 5028 17546
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 5000 15366 5028 15506
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5092 14958 5120 18634
rect 5552 17678 5580 18702
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 17882 5672 18226
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 5736 17678 5764 20590
rect 5908 20596 5960 20602
rect 5908 20538 5960 20544
rect 5920 20398 5948 20538
rect 6104 20534 6132 20810
rect 6196 20806 6224 20964
rect 6368 20946 6420 20952
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6092 20528 6144 20534
rect 6092 20470 6144 20476
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5828 19446 5856 19654
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5828 17678 5856 17750
rect 5920 17678 5948 20334
rect 6104 19854 6132 20470
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18290 6040 19110
rect 6104 18834 6132 19790
rect 6196 19553 6224 20742
rect 6564 20602 6592 21490
rect 6656 21146 6684 21558
rect 6828 21412 6880 21418
rect 6828 21354 6880 21360
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6656 20602 6684 21082
rect 6840 20874 6868 21354
rect 6932 21350 6960 22578
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 7024 21418 7052 22510
rect 7116 22234 7144 22714
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 7392 22166 7420 22714
rect 7380 22160 7432 22166
rect 7380 22102 7432 22108
rect 7760 22094 7788 24475
rect 9048 22778 9076 24475
rect 9692 23066 9720 24475
rect 9692 23038 9812 23066
rect 9441 22876 9749 22885
rect 9441 22874 9447 22876
rect 9503 22874 9527 22876
rect 9583 22874 9607 22876
rect 9663 22874 9687 22876
rect 9743 22874 9749 22876
rect 9503 22822 9505 22874
rect 9685 22822 9687 22874
rect 9441 22820 9447 22822
rect 9503 22820 9527 22822
rect 9583 22820 9607 22822
rect 9663 22820 9687 22822
rect 9743 22820 9749 22822
rect 9441 22811 9749 22820
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 7668 22066 7788 22094
rect 8404 22094 8432 22578
rect 8404 22066 8524 22094
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6828 20868 6880 20874
rect 6828 20810 6880 20816
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6828 20324 6880 20330
rect 6828 20266 6880 20272
rect 6182 19544 6238 19553
rect 6182 19479 6238 19488
rect 6196 19334 6224 19479
rect 6196 19306 6316 19334
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6184 18692 6236 18698
rect 6184 18634 6236 18640
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 6196 17882 6224 18634
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5356 17536 5408 17542
rect 5540 17536 5592 17542
rect 5356 17478 5408 17484
rect 5460 17496 5540 17524
rect 5368 17202 5396 17478
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5354 17096 5410 17105
rect 5460 17082 5488 17496
rect 5540 17478 5592 17484
rect 5736 17218 5764 17614
rect 5552 17202 5764 17218
rect 5920 17202 5948 17614
rect 6012 17270 6040 17682
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 5540 17196 5764 17202
rect 5592 17190 5764 17196
rect 5908 17196 5960 17202
rect 5540 17138 5592 17144
rect 5908 17138 5960 17144
rect 5410 17054 5488 17082
rect 5354 17031 5410 17040
rect 5368 16794 5396 17031
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5552 16182 5580 16934
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5644 15570 5672 16594
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4580 13268 4660 13274
rect 4528 13262 4660 13268
rect 4540 13246 4660 13262
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 4220 13084 4528 13093
rect 4220 13082 4226 13084
rect 4282 13082 4306 13084
rect 4362 13082 4386 13084
rect 4442 13082 4466 13084
rect 4522 13082 4528 13084
rect 4282 13030 4284 13082
rect 4464 13030 4466 13082
rect 4220 13028 4226 13030
rect 4282 13028 4306 13030
rect 4362 13028 4386 13030
rect 4442 13028 4466 13030
rect 4522 13028 4528 13030
rect 4220 13019 4528 13028
rect 4632 12918 4660 13246
rect 4724 12986 4752 13330
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4908 12782 4936 14214
rect 5000 13326 5028 14418
rect 5092 13870 5120 14486
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5184 13802 5212 14350
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 5184 13530 5212 13738
rect 5276 13734 5304 14282
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5276 13530 5304 13670
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5368 13258 5396 14894
rect 5644 14550 5672 15506
rect 5632 14544 5684 14550
rect 5552 14492 5632 14498
rect 5552 14486 5684 14492
rect 5552 14470 5672 14486
rect 5552 14414 5580 14470
rect 5540 14408 5592 14414
rect 5446 14376 5502 14385
rect 5540 14350 5592 14356
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5446 14311 5502 14320
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5368 12850 5396 13194
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 3560 12540 3868 12549
rect 3560 12538 3566 12540
rect 3622 12538 3646 12540
rect 3702 12538 3726 12540
rect 3782 12538 3806 12540
rect 3862 12538 3868 12540
rect 3622 12486 3624 12538
rect 3804 12486 3806 12538
rect 3560 12484 3566 12486
rect 3622 12484 3646 12486
rect 3702 12484 3726 12486
rect 3782 12484 3806 12486
rect 3862 12484 3868 12486
rect 3560 12475 3868 12484
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11762 3372 12038
rect 4220 11996 4528 12005
rect 4220 11994 4226 11996
rect 4282 11994 4306 11996
rect 4362 11994 4386 11996
rect 4442 11994 4466 11996
rect 4522 11994 4528 11996
rect 4282 11942 4284 11994
rect 4464 11942 4466 11994
rect 4220 11940 4226 11942
rect 4282 11940 4306 11942
rect 4362 11940 4386 11942
rect 4442 11940 4466 11942
rect 4522 11940 4528 11942
rect 4220 11931 4528 11940
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3238 11656 3294 11665
rect 3238 11591 3294 11600
rect 3252 10742 3280 11591
rect 4632 11558 4660 12242
rect 4908 12170 4936 12582
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11626 5028 12038
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 3560 11452 3868 11461
rect 3560 11450 3566 11452
rect 3622 11450 3646 11452
rect 3702 11450 3726 11452
rect 3782 11450 3806 11452
rect 3862 11450 3868 11452
rect 3622 11398 3624 11450
rect 3804 11398 3806 11450
rect 3560 11396 3566 11398
rect 3622 11396 3646 11398
rect 3702 11396 3726 11398
rect 3782 11396 3806 11398
rect 3862 11396 3868 11398
rect 3560 11387 3868 11396
rect 4632 11150 4660 11494
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 3344 10538 3372 11018
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 4066 10976 4122 10985
rect 3804 10810 3832 10950
rect 4066 10911 4122 10920
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3560 10364 3868 10373
rect 3560 10362 3566 10364
rect 3622 10362 3646 10364
rect 3702 10362 3726 10364
rect 3782 10362 3806 10364
rect 3862 10362 3868 10364
rect 3622 10310 3624 10362
rect 3804 10310 3806 10362
rect 3560 10308 3566 10310
rect 3622 10308 3646 10310
rect 3702 10308 3726 10310
rect 3782 10308 3806 10310
rect 3862 10308 3868 10310
rect 3560 10299 3868 10308
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9654 2912 9862
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2976 9518 3004 9930
rect 3344 9586 3372 9998
rect 3884 9648 3936 9654
rect 3882 9616 3884 9625
rect 3936 9616 3938 9625
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3332 9580 3384 9586
rect 4080 9586 4108 10911
rect 4220 10908 4528 10917
rect 4220 10906 4226 10908
rect 4282 10906 4306 10908
rect 4362 10906 4386 10908
rect 4442 10906 4466 10908
rect 4522 10906 4528 10908
rect 4282 10854 4284 10906
rect 4464 10854 4466 10906
rect 4220 10852 4226 10854
rect 4282 10852 4306 10854
rect 4362 10852 4386 10854
rect 4442 10852 4466 10854
rect 4522 10852 4528 10854
rect 4220 10843 4528 10852
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4172 10606 4200 10746
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4172 10198 4200 10542
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9908 4200 9998
rect 4632 9994 4660 11086
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4252 9920 4304 9926
rect 4172 9880 4252 9908
rect 4252 9862 4304 9868
rect 4220 9820 4528 9829
rect 4220 9818 4226 9820
rect 4282 9818 4306 9820
rect 4362 9818 4386 9820
rect 4442 9818 4466 9820
rect 4522 9818 4528 9820
rect 4282 9766 4284 9818
rect 4464 9766 4466 9818
rect 4220 9764 4226 9766
rect 4282 9764 4306 9766
rect 4362 9764 4386 9766
rect 4442 9764 4466 9766
rect 4522 9764 4528 9766
rect 4220 9755 4528 9764
rect 3882 9551 3938 9560
rect 3976 9580 4028 9586
rect 3332 9522 3384 9528
rect 3976 9522 4028 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1964 8974 1992 9318
rect 1676 8968 1728 8974
rect 1306 8936 1362 8945
rect 1676 8910 1728 8916
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1306 8871 1362 8880
rect 1688 8566 1716 8910
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1122 6896 1178 6905
rect 1780 6866 1808 8434
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2228 7812 2280 7818
rect 2228 7754 2280 7760
rect 2240 7546 2268 7754
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2778 7440 2834 7449
rect 2412 7404 2464 7410
rect 2778 7375 2780 7384
rect 2412 7346 2464 7352
rect 2832 7375 2834 7384
rect 2780 7346 2832 7352
rect 2424 7002 2452 7346
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 1122 6831 1178 6840
rect 1768 6860 1820 6866
rect 1136 6798 1164 6831
rect 1768 6802 1820 6808
rect 1124 6792 1176 6798
rect 1124 6734 1176 6740
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2332 6254 2360 6734
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1872 3942 1900 5170
rect 2332 4078 2360 6190
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2700 5710 2728 6054
rect 2792 5914 2820 6394
rect 2884 6322 2912 7822
rect 2976 6866 3004 9454
rect 3068 8838 3096 9522
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 7954 3096 8774
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 3160 7818 3188 8230
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7342 3096 7686
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2884 5710 2912 6258
rect 2976 6225 3004 6666
rect 3068 6662 3096 7278
rect 3160 6730 3188 7754
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3252 6458 3280 7346
rect 3344 6866 3372 9522
rect 3988 9382 4016 9522
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3560 9276 3868 9285
rect 3560 9274 3566 9276
rect 3622 9274 3646 9276
rect 3702 9274 3726 9276
rect 3782 9274 3806 9276
rect 3862 9274 3868 9276
rect 3622 9222 3624 9274
rect 3804 9222 3806 9274
rect 3560 9220 3566 9222
rect 3622 9220 3646 9222
rect 3702 9220 3726 9222
rect 3782 9220 3806 9222
rect 3862 9220 3868 9222
rect 3560 9211 3868 9220
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3560 8188 3868 8197
rect 3560 8186 3566 8188
rect 3622 8186 3646 8188
rect 3702 8186 3726 8188
rect 3782 8186 3806 8188
rect 3862 8186 3868 8188
rect 3622 8134 3624 8186
rect 3804 8134 3806 8186
rect 3560 8132 3566 8134
rect 3622 8132 3646 8134
rect 3702 8132 3726 8134
rect 3782 8132 3806 8134
rect 3862 8132 3868 8134
rect 3560 8123 3868 8132
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3528 7478 3556 7822
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7585 3832 7686
rect 3790 7576 3846 7585
rect 3790 7511 3846 7520
rect 3516 7472 3568 7478
rect 3896 7449 3924 8842
rect 3988 7818 4016 9318
rect 4632 8906 4660 9930
rect 4724 9450 4752 10678
rect 4816 10606 4844 11290
rect 4908 11014 4936 11290
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 9450 4844 9862
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4908 9110 4936 10950
rect 5092 10538 5120 11698
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11150 5212 11494
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5276 10538 5304 10746
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 9580 5040 9586
rect 5092 9568 5120 9998
rect 5040 9540 5120 9568
rect 4988 9522 5040 9528
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4080 8514 4108 8774
rect 4220 8732 4528 8741
rect 4220 8730 4226 8732
rect 4282 8730 4306 8732
rect 4362 8730 4386 8732
rect 4442 8730 4466 8732
rect 4522 8730 4528 8732
rect 4282 8678 4284 8730
rect 4464 8678 4466 8730
rect 4220 8676 4226 8678
rect 4282 8676 4306 8678
rect 4362 8676 4386 8678
rect 4442 8676 4466 8678
rect 4522 8676 4528 8678
rect 4220 8667 4528 8676
rect 4632 8566 4660 8842
rect 4620 8560 4672 8566
rect 4080 8498 4200 8514
rect 4620 8502 4672 8508
rect 4080 8492 4212 8498
rect 4080 8486 4160 8492
rect 4160 8434 4212 8440
rect 4724 8022 4752 8910
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4160 7880 4212 7886
rect 4080 7840 4160 7868
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7478 4016 7754
rect 3976 7472 4028 7478
rect 3516 7414 3568 7420
rect 3882 7440 3938 7449
rect 3976 7414 4028 7420
rect 3882 7375 3938 7384
rect 4080 7274 4108 7840
rect 4160 7822 4212 7828
rect 4220 7644 4528 7653
rect 4220 7642 4226 7644
rect 4282 7642 4306 7644
rect 4362 7642 4386 7644
rect 4442 7642 4466 7644
rect 4522 7642 4528 7644
rect 4282 7590 4284 7642
rect 4464 7590 4466 7642
rect 4220 7588 4226 7590
rect 4282 7588 4306 7590
rect 4362 7588 4386 7590
rect 4442 7588 4466 7590
rect 4522 7588 4528 7590
rect 4220 7579 4528 7588
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3560 7100 3868 7109
rect 3560 7098 3566 7100
rect 3622 7098 3646 7100
rect 3702 7098 3726 7100
rect 3782 7098 3806 7100
rect 3862 7098 3868 7100
rect 3622 7046 3624 7098
rect 3804 7046 3806 7098
rect 3560 7044 3566 7046
rect 3622 7044 3646 7046
rect 3702 7044 3726 7046
rect 3782 7044 3806 7046
rect 3862 7044 3868 7046
rect 3560 7035 3868 7044
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3436 6322 3464 6598
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 2962 6216 3018 6225
rect 2962 6151 3018 6160
rect 3148 6112 3200 6118
rect 3200 6072 3372 6100
rect 3148 6054 3200 6060
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5302 2912 5646
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2884 4622 2912 5238
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2778 4176 2834 4185
rect 2778 4111 2780 4120
rect 2832 4111 2834 4120
rect 2780 4082 2832 4088
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 3058 1624 3470
rect 1688 3126 1716 3878
rect 2884 3534 2912 4558
rect 3160 4214 3188 5306
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 2964 4208 3016 4214
rect 3148 4208 3200 4214
rect 3016 4156 3096 4162
rect 2964 4150 3096 4156
rect 3148 4150 3200 4156
rect 2976 4134 3096 4150
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1964 2650 1992 3402
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2778 2816 2834 2825
rect 2778 2751 2834 2760
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2792 2514 2820 2751
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2884 2378 2912 3334
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2976 2145 3004 3946
rect 3068 3194 3096 4134
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3160 3534 3188 3878
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3068 2514 3096 3130
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 2962 2136 3018 2145
rect 2962 2071 3018 2080
rect 3252 800 3280 5238
rect 3344 2774 3372 6072
rect 3560 6012 3868 6021
rect 3560 6010 3566 6012
rect 3622 6010 3646 6012
rect 3702 6010 3726 6012
rect 3782 6010 3806 6012
rect 3862 6010 3868 6012
rect 3622 5958 3624 6010
rect 3804 5958 3806 6010
rect 3560 5956 3566 5958
rect 3622 5956 3646 5958
rect 3702 5956 3726 5958
rect 3782 5956 3806 5958
rect 3862 5956 3868 5958
rect 3560 5947 3868 5956
rect 3560 4924 3868 4933
rect 3560 4922 3566 4924
rect 3622 4922 3646 4924
rect 3702 4922 3726 4924
rect 3782 4922 3806 4924
rect 3862 4922 3868 4924
rect 3622 4870 3624 4922
rect 3804 4870 3806 4922
rect 3560 4868 3566 4870
rect 3622 4868 3646 4870
rect 3702 4868 3726 4870
rect 3782 4868 3806 4870
rect 3862 4868 3868 4870
rect 3422 4856 3478 4865
rect 3560 4859 3868 4868
rect 3422 4791 3478 4800
rect 3436 4622 3464 4791
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3792 4548 3844 4554
rect 3896 4536 3924 7210
rect 4448 6798 4476 7482
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4220 6556 4528 6565
rect 4220 6554 4226 6556
rect 4282 6554 4306 6556
rect 4362 6554 4386 6556
rect 4442 6554 4466 6556
rect 4522 6554 4528 6556
rect 4282 6502 4284 6554
rect 4464 6502 4466 6554
rect 4220 6500 4226 6502
rect 4282 6500 4306 6502
rect 4362 6500 4386 6502
rect 4442 6500 4466 6502
rect 4522 6500 4528 6502
rect 4220 6491 4528 6500
rect 4632 6458 4660 6598
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4356 5710 4384 6190
rect 4724 6118 4752 6734
rect 4816 6730 4844 8842
rect 4908 7993 4936 8910
rect 5092 8906 5120 9540
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 8634 5212 8842
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 4988 8288 5040 8294
rect 5184 8242 5212 8570
rect 4988 8230 5040 8236
rect 4894 7984 4950 7993
rect 4894 7919 4950 7928
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4908 7002 4936 7346
rect 5000 7206 5028 8230
rect 5092 8214 5212 8242
rect 5092 7818 5120 8214
rect 5276 7954 5304 10474
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5276 7546 5304 7890
rect 5368 7886 5396 11018
rect 5460 10742 5488 14311
rect 5644 14006 5672 14350
rect 5736 14074 5764 16050
rect 5920 15706 5948 16050
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 6012 15502 6040 17206
rect 6288 17066 6316 19306
rect 6840 19174 6868 20266
rect 6932 19446 6960 21286
rect 7392 20262 7420 21422
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6472 17338 6500 17614
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6564 17202 6592 17750
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6472 16590 6500 16934
rect 6564 16794 6592 17002
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6748 16658 6776 18022
rect 6840 17814 6868 19110
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6840 17134 6868 17750
rect 6932 17746 6960 19382
rect 7300 19378 7328 19722
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7484 19310 7512 19654
rect 7668 19514 7696 22066
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8312 21554 8340 21898
rect 8496 21706 8524 22066
rect 8588 21842 8616 22646
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 8680 22094 8708 22374
rect 8781 22332 9089 22341
rect 8781 22330 8787 22332
rect 8843 22330 8867 22332
rect 8923 22330 8947 22332
rect 9003 22330 9027 22332
rect 9083 22330 9089 22332
rect 8843 22278 8845 22330
rect 9025 22278 9027 22330
rect 8781 22276 8787 22278
rect 8843 22276 8867 22278
rect 8923 22276 8947 22278
rect 9003 22276 9027 22278
rect 9083 22276 9089 22278
rect 8781 22267 9089 22276
rect 8944 22160 8996 22166
rect 8944 22102 8996 22108
rect 8680 22066 8892 22094
rect 8864 22030 8892 22066
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8588 21814 8708 21842
rect 8496 21678 8616 21706
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7760 20058 7788 20402
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 8036 19854 8064 21286
rect 8128 20806 8156 21422
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 7944 19514 7972 19790
rect 8128 19786 8156 20742
rect 8312 20534 8340 21490
rect 8404 21078 8432 21558
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 8496 21146 8524 21490
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8392 21072 8444 21078
rect 8392 21014 8444 21020
rect 8404 20534 8432 21014
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8220 20058 8248 20334
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 8022 19544 8078 19553
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7932 19508 7984 19514
rect 8022 19479 8024 19488
rect 7932 19450 7984 19456
rect 8076 19479 8078 19488
rect 8024 19450 8076 19456
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7116 18766 7144 19110
rect 7484 18970 7512 19246
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7668 18426 7696 19450
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6932 17338 6960 17546
rect 8128 17542 8156 19722
rect 8220 19446 8248 19994
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8312 19242 8340 20470
rect 8588 20330 8616 21678
rect 8680 20754 8708 21814
rect 8956 21690 8984 22102
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 8781 21244 9089 21253
rect 8781 21242 8787 21244
rect 8843 21242 8867 21244
rect 8923 21242 8947 21244
rect 9003 21242 9027 21244
rect 9083 21242 9089 21244
rect 8843 21190 8845 21242
rect 9025 21190 9027 21242
rect 8781 21188 8787 21190
rect 8843 21188 8867 21190
rect 8923 21188 8947 21190
rect 9003 21188 9027 21190
rect 9083 21188 9089 21190
rect 8781 21179 9089 21188
rect 9140 20942 9168 22374
rect 9232 22166 9260 22578
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9600 22234 9628 22510
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9220 22160 9272 22166
rect 9220 22102 9272 22108
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9232 21146 9260 21898
rect 9324 21554 9352 22034
rect 9441 21788 9749 21797
rect 9441 21786 9447 21788
rect 9503 21786 9527 21788
rect 9583 21786 9607 21788
rect 9663 21786 9687 21788
rect 9743 21786 9749 21788
rect 9503 21734 9505 21786
rect 9685 21734 9687 21786
rect 9441 21732 9447 21734
rect 9503 21732 9527 21734
rect 9583 21732 9607 21734
rect 9663 21732 9687 21734
rect 9743 21732 9749 21734
rect 9441 21723 9749 21732
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9324 21010 9352 21490
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9416 20856 9444 21626
rect 9324 20828 9444 20856
rect 8680 20726 9168 20754
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8680 20466 8708 20538
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8576 20324 8628 20330
rect 8576 20266 8628 20272
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8312 18902 8340 19178
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 8312 18290 8340 18838
rect 8404 18766 8432 19926
rect 8680 19514 8708 20402
rect 8781 20156 9089 20165
rect 8781 20154 8787 20156
rect 8843 20154 8867 20156
rect 8923 20154 8947 20156
rect 9003 20154 9027 20156
rect 9083 20154 9089 20156
rect 8843 20102 8845 20154
rect 9025 20102 9027 20154
rect 8781 20100 8787 20102
rect 8843 20100 8867 20102
rect 8923 20100 8947 20102
rect 9003 20100 9027 20102
rect 9083 20100 9089 20102
rect 8781 20091 9089 20100
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 9140 19446 9168 20726
rect 9324 20602 9352 20828
rect 9441 20700 9749 20709
rect 9441 20698 9447 20700
rect 9503 20698 9527 20700
rect 9583 20698 9607 20700
rect 9663 20698 9687 20700
rect 9743 20698 9749 20700
rect 9503 20646 9505 20698
rect 9685 20646 9687 20698
rect 9441 20644 9447 20646
rect 9503 20644 9527 20646
rect 9583 20644 9607 20646
rect 9663 20644 9687 20646
rect 9743 20644 9749 20646
rect 9441 20635 9749 20644
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9784 20040 9812 23038
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10060 20942 10088 21830
rect 10796 21622 10824 21830
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 10888 21350 10916 21966
rect 10980 21690 11008 24475
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 11072 20942 11100 22374
rect 11348 22094 11376 24534
rect 11532 24426 11560 24534
rect 11610 24475 11666 25275
rect 12254 24475 12310 25275
rect 12898 24475 12954 25275
rect 13542 24475 13598 25275
rect 13924 24534 14136 24562
rect 11624 24426 11652 24475
rect 11532 24398 11652 24426
rect 11612 22636 11664 22642
rect 11612 22578 11664 22584
rect 11348 22066 11468 22094
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11256 21690 11284 21898
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9876 20262 9904 20810
rect 10060 20534 10088 20878
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10048 20528 10100 20534
rect 10048 20470 10100 20476
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9692 20012 9812 20040
rect 9692 19718 9720 20012
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9441 19612 9749 19621
rect 9441 19610 9447 19612
rect 9503 19610 9527 19612
rect 9583 19610 9607 19612
rect 9663 19610 9687 19612
rect 9743 19610 9749 19612
rect 9503 19558 9505 19610
rect 9685 19558 9687 19610
rect 9441 19556 9447 19558
rect 9503 19556 9527 19558
rect 9583 19556 9607 19558
rect 9663 19556 9687 19558
rect 9743 19556 9749 19558
rect 9441 19547 9749 19556
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9128 19440 9180 19446
rect 8574 19408 8630 19417
rect 8484 19372 8536 19378
rect 9128 19382 9180 19388
rect 8574 19343 8576 19352
rect 8484 19314 8536 19320
rect 8628 19343 8630 19352
rect 8576 19314 8628 19320
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8496 18578 8524 19314
rect 9692 19174 9720 19450
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 8781 19068 9089 19077
rect 8781 19066 8787 19068
rect 8843 19066 8867 19068
rect 8923 19066 8947 19068
rect 9003 19066 9027 19068
rect 9083 19066 9089 19068
rect 8843 19014 8845 19066
rect 9025 19014 9027 19066
rect 8781 19012 8787 19014
rect 8843 19012 8867 19014
rect 8923 19012 8947 19014
rect 9003 19012 9027 19014
rect 9083 19012 9089 19014
rect 8781 19003 9089 19012
rect 8404 18550 8524 18578
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7932 17264 7984 17270
rect 8024 17264 8076 17270
rect 7932 17206 7984 17212
rect 8022 17232 8024 17241
rect 8076 17232 8078 17241
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6748 16182 6776 16594
rect 6932 16590 6960 16934
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 7576 16250 7604 17070
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 7576 15502 7604 16186
rect 7852 15978 7880 17138
rect 7944 16726 7972 17206
rect 8022 17167 8078 17176
rect 8128 17134 8156 17478
rect 8220 17338 8248 17546
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 8404 16726 8432 18550
rect 8588 18290 8616 18566
rect 9441 18524 9749 18533
rect 9441 18522 9447 18524
rect 9503 18522 9527 18524
rect 9583 18522 9607 18524
rect 9663 18522 9687 18524
rect 9743 18522 9749 18524
rect 9503 18470 9505 18522
rect 9685 18470 9687 18522
rect 9441 18468 9447 18470
rect 9503 18468 9527 18470
rect 9583 18468 9607 18470
rect 9663 18468 9687 18470
rect 9743 18468 9749 18470
rect 9441 18459 9749 18468
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8781 17980 9089 17989
rect 8781 17978 8787 17980
rect 8843 17978 8867 17980
rect 8923 17978 8947 17980
rect 9003 17978 9027 17980
rect 9083 17978 9089 17980
rect 8843 17926 8845 17978
rect 9025 17926 9027 17978
rect 8781 17924 8787 17926
rect 8843 17924 8867 17926
rect 8923 17924 8947 17926
rect 9003 17924 9027 17926
rect 9083 17924 9089 17926
rect 8781 17915 9089 17924
rect 9784 17882 9812 19858
rect 10244 19786 10272 20742
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 9876 19514 9904 19722
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 8484 17808 8536 17814
rect 8484 17750 8536 17756
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 7944 16182 7972 16662
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 5906 15056 5962 15065
rect 5906 14991 5962 15000
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5828 14618 5856 14758
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5644 13394 5672 13738
rect 5736 13394 5764 14010
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5644 12986 5672 13330
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5828 12918 5856 14010
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5920 12850 5948 14991
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6012 13394 6040 14214
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6458 13424 6514 13433
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6092 13388 6144 13394
rect 6458 13359 6514 13368
rect 6092 13330 6144 13336
rect 6104 13258 6132 13330
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6472 12986 6500 13359
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6564 12918 6592 14010
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6748 13190 6776 13942
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6748 12850 6776 13126
rect 5908 12844 5960 12850
rect 6276 12844 6328 12850
rect 5960 12804 6276 12832
rect 5908 12786 5960 12792
rect 6276 12786 6328 12792
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12306 5764 12582
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 6564 12170 6592 12650
rect 6656 12442 6684 12786
rect 6840 12646 6868 14282
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 12986 6960 13806
rect 7024 13258 7052 14214
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7392 13530 7420 13874
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7116 12986 7144 13466
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7288 12912 7340 12918
rect 7288 12854 7340 12860
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6104 11150 6132 11562
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10810 5580 10950
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5460 10198 5488 10542
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5460 8294 5488 10134
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9654 5672 9862
rect 5828 9654 5856 10406
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5552 8106 5580 8910
rect 5644 8906 5672 9386
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8498 5856 8774
rect 5920 8498 5948 10610
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 10062 6040 10406
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6104 10062 6132 10202
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6012 9382 6040 9998
rect 6564 9654 6592 12106
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6656 10130 6684 11222
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6932 11082 6960 11154
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 7024 10674 7052 12718
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7116 11082 7144 11290
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6840 10062 6868 10610
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6104 8566 6132 9522
rect 6564 8838 6592 9590
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 8974 6776 9522
rect 7024 8974 7052 9862
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5460 8078 5580 8106
rect 5644 8090 5672 8434
rect 5632 8084 5684 8090
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5460 7698 5488 8078
rect 5632 8026 5684 8032
rect 5368 7670 5488 7698
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4816 5930 4844 6666
rect 5000 6118 5028 7142
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4724 5902 4844 5930
rect 3976 5704 4028 5710
rect 4344 5704 4396 5710
rect 3976 5646 4028 5652
rect 4080 5652 4344 5658
rect 4080 5646 4396 5652
rect 3988 5545 4016 5646
rect 4080 5630 4384 5646
rect 4620 5636 4672 5642
rect 3974 5536 4030 5545
rect 3974 5471 4030 5480
rect 4080 5386 4108 5630
rect 4620 5578 4672 5584
rect 4220 5468 4528 5477
rect 4220 5466 4226 5468
rect 4282 5466 4306 5468
rect 4362 5466 4386 5468
rect 4442 5466 4466 5468
rect 4522 5466 4528 5468
rect 4282 5414 4284 5466
rect 4464 5414 4466 5466
rect 4220 5412 4226 5414
rect 4282 5412 4306 5414
rect 4362 5412 4386 5414
rect 4442 5412 4466 5414
rect 4522 5412 4528 5414
rect 4220 5403 4528 5412
rect 3844 4508 3924 4536
rect 3988 5358 4108 5386
rect 4632 5370 4660 5578
rect 4724 5574 4752 5902
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4620 5364 4672 5370
rect 3792 4490 3844 4496
rect 3804 4010 3832 4490
rect 3988 4162 4016 5358
rect 4620 5306 4672 5312
rect 4724 5234 4752 5510
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4080 4486 4108 5170
rect 4528 5092 4580 5098
rect 4580 5052 4660 5080
rect 4528 5034 4580 5040
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4220 4380 4528 4389
rect 4220 4378 4226 4380
rect 4282 4378 4306 4380
rect 4362 4378 4386 4380
rect 4442 4378 4466 4380
rect 4522 4378 4528 4380
rect 4282 4326 4284 4378
rect 4464 4326 4466 4378
rect 4220 4324 4226 4326
rect 4282 4324 4306 4326
rect 4362 4324 4386 4326
rect 4442 4324 4466 4326
rect 4522 4324 4528 4326
rect 4220 4315 4528 4324
rect 3884 4140 3936 4146
rect 3988 4134 4200 4162
rect 3884 4082 3936 4088
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3560 3836 3868 3845
rect 3560 3834 3566 3836
rect 3622 3834 3646 3836
rect 3702 3834 3726 3836
rect 3782 3834 3806 3836
rect 3862 3834 3868 3836
rect 3622 3782 3624 3834
rect 3804 3782 3806 3834
rect 3560 3780 3566 3782
rect 3622 3780 3646 3782
rect 3702 3780 3726 3782
rect 3782 3780 3806 3782
rect 3862 3780 3868 3782
rect 3560 3771 3868 3780
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 3126 3648 3334
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3712 3058 3740 3538
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3344 2746 3464 2774
rect 3436 921 3464 2746
rect 3560 2748 3868 2757
rect 3560 2746 3566 2748
rect 3622 2746 3646 2748
rect 3702 2746 3726 2748
rect 3782 2746 3806 2748
rect 3862 2746 3868 2748
rect 3622 2694 3624 2746
rect 3804 2694 3806 2746
rect 3560 2692 3566 2694
rect 3622 2692 3646 2694
rect 3702 2692 3726 2694
rect 3782 2692 3806 2694
rect 3862 2692 3868 2694
rect 3560 2683 3868 2692
rect 3422 912 3478 921
rect 3422 847 3478 856
rect 3896 800 3924 4082
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3988 2446 4016 3946
rect 4172 3466 4200 4134
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4220 3292 4528 3301
rect 4220 3290 4226 3292
rect 4282 3290 4306 3292
rect 4362 3290 4386 3292
rect 4442 3290 4466 3292
rect 4522 3290 4528 3292
rect 4282 3238 4284 3290
rect 4464 3238 4466 3290
rect 4220 3236 4226 3238
rect 4282 3236 4306 3238
rect 4362 3236 4386 3238
rect 4442 3236 4466 3238
rect 4522 3236 4528 3238
rect 4220 3227 4528 3236
rect 4632 2650 4660 5052
rect 4816 4826 4844 5714
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4220 2204 4528 2213
rect 4220 2202 4226 2204
rect 4282 2202 4306 2204
rect 4362 2202 4386 2204
rect 4442 2202 4466 2204
rect 4522 2202 4528 2204
rect 4282 2150 4284 2202
rect 4464 2150 4466 2202
rect 4220 2148 4226 2150
rect 4282 2148 4306 2150
rect 4362 2148 4386 2150
rect 4442 2148 4466 2150
rect 4522 2148 4528 2150
rect 4220 2139 4528 2148
rect 4724 1986 4752 4082
rect 4816 4010 4844 4490
rect 4908 4026 4936 6054
rect 5000 5914 5028 6054
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 5092 5166 5120 7414
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5184 5914 5212 6666
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5092 4622 5120 5102
rect 5276 4706 5304 6802
rect 5368 6662 5396 7670
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6458 5396 6598
rect 5460 6474 5488 7482
rect 5920 7410 5948 8434
rect 6748 8430 6776 8910
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 7478 6132 8230
rect 6748 7886 6776 8366
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6564 7546 6592 7754
rect 6840 7546 6868 8774
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7116 8090 7144 8434
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 6934 5948 7346
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5736 6662 5764 6802
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5356 6452 5408 6458
rect 5460 6446 5580 6474
rect 5356 6394 5408 6400
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5368 5914 5396 6258
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5184 4678 5304 4706
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5000 4298 5028 4490
rect 5000 4270 5120 4298
rect 5092 4214 5120 4270
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 4804 4004 4856 4010
rect 4908 3998 5028 4026
rect 4804 3946 4856 3952
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3534 4936 3878
rect 4896 3528 4948 3534
rect 5000 3505 5028 3998
rect 4896 3470 4948 3476
rect 4986 3496 5042 3505
rect 4986 3431 5042 3440
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 2582 5028 3334
rect 5092 3194 5120 4150
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 4540 1958 4752 1986
rect 4540 800 4568 1958
rect 5184 1465 5212 4678
rect 5460 4622 5488 6258
rect 5552 5522 5580 6446
rect 5644 5914 5672 6598
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5828 5778 5856 6598
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5920 5710 5948 6870
rect 6840 6866 6868 7482
rect 7208 6866 7236 12174
rect 7300 11286 7328 12854
rect 7392 12782 7420 13330
rect 7484 12918 7512 13806
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7668 12850 7696 14554
rect 7760 14482 7788 14894
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 14006 7880 14214
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8312 13530 8340 13806
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7392 12306 7420 12718
rect 8312 12434 8340 13262
rect 8220 12406 8340 12434
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 8220 12238 8248 12406
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7760 11830 7788 12038
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 8128 10674 8156 12038
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7392 10198 7420 10406
rect 7760 10266 7788 10406
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7944 10062 7972 10610
rect 8220 10198 8248 10950
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8312 10062 8340 11290
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 8634 7328 8978
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7300 7546 7328 8570
rect 7392 8566 7420 9862
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7576 9110 7604 9522
rect 7668 9178 7696 9522
rect 7944 9518 7972 9862
rect 8404 9738 8432 16662
rect 8496 16590 8524 17750
rect 9876 17678 9904 19450
rect 9968 18426 9996 19654
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 10152 18154 10180 18702
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18358 10364 18566
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10140 18148 10192 18154
rect 10140 18090 10192 18096
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 8680 16590 8708 17614
rect 10336 17542 10364 18294
rect 10612 18290 10640 19994
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10704 18970 10732 19314
rect 10888 19174 10916 19654
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10888 18426 10916 19110
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 9441 17436 9749 17445
rect 9441 17434 9447 17436
rect 9503 17434 9527 17436
rect 9583 17434 9607 17436
rect 9663 17434 9687 17436
rect 9743 17434 9749 17436
rect 9503 17382 9505 17434
rect 9685 17382 9687 17434
rect 9441 17380 9447 17382
rect 9503 17380 9527 17382
rect 9583 17380 9607 17382
rect 9663 17380 9687 17382
rect 9743 17380 9749 17382
rect 9441 17371 9749 17380
rect 10520 17270 10548 17478
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 8781 16892 9089 16901
rect 8781 16890 8787 16892
rect 8843 16890 8867 16892
rect 8923 16890 8947 16892
rect 9003 16890 9027 16892
rect 9083 16890 9089 16892
rect 8843 16838 8845 16890
rect 9025 16838 9027 16890
rect 8781 16836 8787 16838
rect 8843 16836 8867 16838
rect 8923 16836 8947 16838
rect 9003 16836 9027 16838
rect 9083 16836 9089 16838
rect 8781 16827 9089 16836
rect 9324 16794 9352 17070
rect 9600 17066 9628 17138
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9600 16794 9628 17002
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9324 16658 9352 16730
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8496 15706 8524 16186
rect 8956 16130 8984 16390
rect 9324 16182 9352 16594
rect 9692 16590 9720 16934
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9441 16348 9749 16357
rect 9441 16346 9447 16348
rect 9503 16346 9527 16348
rect 9583 16346 9607 16348
rect 9663 16346 9687 16348
rect 9743 16346 9749 16348
rect 9503 16294 9505 16346
rect 9685 16294 9687 16346
rect 9441 16292 9447 16294
rect 9503 16292 9527 16294
rect 9583 16292 9607 16294
rect 9663 16292 9687 16294
rect 9743 16292 9749 16294
rect 9441 16283 9749 16292
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9312 16176 9364 16182
rect 8956 16114 9076 16130
rect 9312 16118 9364 16124
rect 8956 16108 9088 16114
rect 8956 16102 9036 16108
rect 9036 16050 9088 16056
rect 8781 15804 9089 15813
rect 8781 15802 8787 15804
rect 8843 15802 8867 15804
rect 8923 15802 8947 15804
rect 9003 15802 9027 15804
rect 9083 15802 9089 15804
rect 8843 15750 8845 15802
rect 9025 15750 9027 15802
rect 8781 15748 8787 15750
rect 8843 15748 8867 15750
rect 8923 15748 8947 15750
rect 9003 15748 9027 15750
rect 9083 15748 9089 15750
rect 8781 15739 9089 15748
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8680 14278 8708 15438
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9048 15094 9076 15302
rect 9324 15162 9352 16118
rect 9441 15260 9749 15269
rect 9441 15258 9447 15260
rect 9503 15258 9527 15260
rect 9583 15258 9607 15260
rect 9663 15258 9687 15260
rect 9743 15258 9749 15260
rect 9503 15206 9505 15258
rect 9685 15206 9687 15258
rect 9441 15204 9447 15206
rect 9503 15204 9527 15206
rect 9583 15204 9607 15206
rect 9663 15204 9687 15206
rect 9743 15204 9749 15206
rect 9441 15195 9749 15204
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 8781 14716 9089 14725
rect 8781 14714 8787 14716
rect 8843 14714 8867 14716
rect 8923 14714 8947 14716
rect 9003 14714 9027 14716
rect 9083 14714 9089 14716
rect 8843 14662 8845 14714
rect 9025 14662 9027 14714
rect 8781 14660 8787 14662
rect 8843 14660 8867 14662
rect 8923 14660 8947 14662
rect 9003 14660 9027 14662
rect 9083 14660 9089 14662
rect 8781 14651 9089 14660
rect 9324 14482 9352 15098
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13376 8524 13670
rect 8588 13530 8616 13942
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8576 13388 8628 13394
rect 8496 13348 8576 13376
rect 8496 12238 8524 13348
rect 8576 13330 8628 13336
rect 8680 13326 8708 14214
rect 8781 13628 9089 13637
rect 8781 13626 8787 13628
rect 8843 13626 8867 13628
rect 8923 13626 8947 13628
rect 9003 13626 9027 13628
rect 9083 13626 9089 13628
rect 8843 13574 8845 13626
rect 9025 13574 9027 13626
rect 8781 13572 8787 13574
rect 8843 13572 8867 13574
rect 8923 13572 8947 13574
rect 9003 13572 9027 13574
rect 9083 13572 9089 13574
rect 8781 13563 9089 13572
rect 9140 13530 9168 14214
rect 9232 13734 9260 14282
rect 9324 14074 9352 14418
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9441 14172 9749 14181
rect 9441 14170 9447 14172
rect 9503 14170 9527 14172
rect 9583 14170 9607 14172
rect 9663 14170 9687 14172
rect 9743 14170 9749 14172
rect 9503 14118 9505 14170
rect 9685 14118 9687 14170
rect 9441 14116 9447 14118
rect 9503 14116 9527 14118
rect 9583 14116 9607 14118
rect 9663 14116 9687 14118
rect 9743 14116 9749 14118
rect 9441 14107 9749 14116
rect 9312 14068 9364 14074
rect 9784 14056 9812 14214
rect 9312 14010 9364 14016
rect 9416 14028 9812 14056
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8588 11694 8616 12650
rect 8680 12238 8708 12786
rect 9232 12646 9260 13262
rect 9416 13240 9444 14028
rect 9876 13977 9904 16186
rect 9968 15706 9996 16458
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 9862 13968 9918 13977
rect 9772 13932 9824 13938
rect 9862 13903 9918 13912
rect 9772 13874 9824 13880
rect 9324 13212 9444 13240
rect 9324 12918 9352 13212
rect 9441 13084 9749 13093
rect 9441 13082 9447 13084
rect 9503 13082 9527 13084
rect 9583 13082 9607 13084
rect 9663 13082 9687 13084
rect 9743 13082 9749 13084
rect 9503 13030 9505 13082
rect 9685 13030 9687 13082
rect 9441 13028 9447 13030
rect 9503 13028 9527 13030
rect 9583 13028 9607 13030
rect 9663 13028 9687 13030
rect 9743 13028 9749 13030
rect 9441 13019 9749 13028
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 8781 12540 9089 12549
rect 8781 12538 8787 12540
rect 8843 12538 8867 12540
rect 8923 12538 8947 12540
rect 9003 12538 9027 12540
rect 9083 12538 9089 12540
rect 8843 12486 8845 12538
rect 9025 12486 9027 12538
rect 8781 12484 8787 12486
rect 8843 12484 8867 12486
rect 8923 12484 8947 12486
rect 9003 12484 9027 12486
rect 9083 12484 9089 12486
rect 8781 12475 9089 12484
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8781 11452 9089 11461
rect 8781 11450 8787 11452
rect 8843 11450 8867 11452
rect 8923 11450 8947 11452
rect 9003 11450 9027 11452
rect 9083 11450 9089 11452
rect 8843 11398 8845 11450
rect 9025 11398 9027 11450
rect 8781 11396 8787 11398
rect 8843 11396 8867 11398
rect 8923 11396 8947 11398
rect 9003 11396 9027 11398
rect 9083 11396 9089 11398
rect 8781 11387 9089 11396
rect 9140 11218 9168 12378
rect 9232 11286 9260 12582
rect 9784 12238 9812 13874
rect 10060 13530 10088 15370
rect 10520 15366 10548 15642
rect 10612 15434 10640 15642
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10244 15094 10272 15302
rect 10520 15094 10548 15302
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10244 14346 10272 15030
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10152 13462 10180 13874
rect 10244 13734 10272 14282
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10140 13456 10192 13462
rect 10060 13404 10140 13410
rect 10060 13398 10192 13404
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10060 13382 10180 13398
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9876 12782 9904 13126
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9324 11898 9352 12174
rect 9441 11996 9749 12005
rect 9441 11994 9447 11996
rect 9503 11994 9527 11996
rect 9583 11994 9607 11996
rect 9663 11994 9687 11996
rect 9743 11994 9749 11996
rect 9503 11942 9505 11994
rect 9685 11942 9687 11994
rect 9441 11940 9447 11942
rect 9503 11940 9527 11942
rect 9583 11940 9607 11942
rect 9663 11940 9687 11942
rect 9743 11940 9749 11942
rect 9441 11931 9749 11940
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9876 11778 9904 12310
rect 9968 12102 9996 13330
rect 10060 13326 10088 13382
rect 10244 13326 10272 13670
rect 10336 13326 10364 14554
rect 10428 14550 10456 14758
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10428 13870 10456 14486
rect 10520 14006 10548 15030
rect 10612 14822 10640 15370
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14618 10640 14758
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10704 13938 10732 14826
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10060 12714 10088 13262
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10152 12714 10180 12854
rect 10244 12782 10272 13262
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10336 12714 10364 13262
rect 10428 13190 10456 13806
rect 10704 13326 10732 13874
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10060 12238 10088 12650
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9692 11750 9904 11778
rect 9588 11688 9640 11694
rect 9692 11676 9720 11750
rect 9640 11648 9720 11676
rect 9864 11688 9916 11694
rect 9588 11630 9640 11636
rect 9864 11630 9916 11636
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9140 11098 9168 11154
rect 9140 11070 9260 11098
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8496 10674 8524 10950
rect 9140 10674 9168 10950
rect 9232 10674 9260 11070
rect 9441 10908 9749 10917
rect 9441 10906 9447 10908
rect 9503 10906 9527 10908
rect 9583 10906 9607 10908
rect 9663 10906 9687 10908
rect 9743 10906 9749 10908
rect 9503 10854 9505 10906
rect 9685 10854 9687 10906
rect 9441 10852 9447 10854
rect 9503 10852 9527 10854
rect 9583 10852 9607 10854
rect 9663 10852 9687 10854
rect 9743 10852 9749 10854
rect 9441 10843 9749 10852
rect 9876 10674 9904 11630
rect 9968 11218 9996 12038
rect 10060 11898 10088 12174
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10244 11218 10272 12582
rect 10428 12374 10456 13126
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10612 12442 10640 12650
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10428 12238 10456 12310
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10336 11830 10364 12106
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10520 11150 10548 11494
rect 10612 11218 10640 11834
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 8496 10266 8524 10610
rect 8781 10364 9089 10373
rect 8781 10362 8787 10364
rect 8843 10362 8867 10364
rect 8923 10362 8947 10364
rect 9003 10362 9027 10364
rect 9083 10362 9089 10364
rect 8843 10310 8845 10362
rect 9025 10310 9027 10362
rect 8781 10308 8787 10310
rect 8843 10308 8867 10310
rect 8923 10308 8947 10310
rect 9003 10308 9027 10310
rect 9083 10308 9089 10310
rect 8781 10299 9089 10308
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 9232 10062 9260 10610
rect 10336 10538 10364 11086
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 10336 9994 10364 10474
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 9441 9820 9749 9829
rect 9441 9818 9447 9820
rect 9503 9818 9527 9820
rect 9583 9818 9607 9820
rect 9663 9818 9687 9820
rect 9743 9818 9749 9820
rect 9503 9766 9505 9818
rect 9685 9766 9687 9818
rect 9441 9764 9447 9766
rect 9503 9764 9527 9766
rect 9583 9764 9607 9766
rect 9663 9764 9687 9766
rect 9743 9764 9749 9766
rect 9441 9755 9749 9764
rect 8404 9710 8708 9738
rect 7932 9512 7984 9518
rect 8404 9466 8432 9710
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 7932 9454 7984 9460
rect 8024 9444 8076 9450
rect 8024 9386 8076 9392
rect 8312 9438 8432 9466
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7852 8634 7880 9046
rect 8036 8974 8064 9386
rect 8312 9382 8340 9438
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7944 8634 7972 8774
rect 8312 8650 8340 9318
rect 8404 8906 8432 9318
rect 8496 8974 8524 9590
rect 8680 9450 8708 9710
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8781 9276 9089 9285
rect 8781 9274 8787 9276
rect 8843 9274 8867 9276
rect 8923 9274 8947 9276
rect 9003 9274 9027 9276
rect 9083 9274 9089 9276
rect 8843 9222 8845 9274
rect 9025 9222 9027 9274
rect 8781 9220 8787 9222
rect 8843 9220 8867 9222
rect 8923 9220 8947 9222
rect 9003 9220 9027 9222
rect 9083 9220 9089 9222
rect 8781 9211 9089 9220
rect 9140 8974 9168 9522
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9692 8906 9720 9658
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7932 8628 7984 8634
rect 8312 8622 8432 8650
rect 7932 8570 7984 8576
rect 7380 8560 7432 8566
rect 7432 8520 7512 8548
rect 7380 8502 7432 8508
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6472 6322 6500 6734
rect 6564 6458 6592 6734
rect 7024 6458 7052 6734
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6564 5710 6592 6394
rect 7024 5710 7052 6394
rect 7208 5778 7236 6802
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 5552 5494 5764 5522
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5276 4282 5304 4558
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5276 3738 5304 4218
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5460 3602 5488 4558
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5368 2854 5396 3402
rect 5460 3126 5488 3538
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5368 2446 5396 2790
rect 5552 2774 5580 5238
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4622 5672 4966
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5632 4072 5684 4078
rect 5736 4060 5764 5494
rect 6104 5098 6132 5646
rect 7300 5574 7328 7482
rect 7392 7478 7420 7686
rect 7484 7478 7512 8520
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7484 5658 7512 7414
rect 7668 7410 7696 7754
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7668 7002 7696 7346
rect 7760 7274 7788 8434
rect 7944 7886 7972 8570
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 8312 7546 8340 8434
rect 8404 8090 8432 8622
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8781 8188 9089 8197
rect 8781 8186 8787 8188
rect 8843 8186 8867 8188
rect 8923 8186 8947 8188
rect 9003 8186 9027 8188
rect 9083 8186 9089 8188
rect 8843 8134 8845 8186
rect 9025 8134 9027 8186
rect 8781 8132 8787 8134
rect 8843 8132 8867 8134
rect 8923 8132 8947 8134
rect 9003 8132 9027 8134
rect 9083 8132 9089 8134
rect 8781 8123 9089 8132
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7546 8432 7822
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7576 5846 7604 6190
rect 7944 5914 7972 6666
rect 8312 6390 8340 7210
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 8036 5778 8064 6258
rect 8404 5846 8432 6598
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 8496 5710 8524 7754
rect 9048 7478 9076 8026
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8588 5914 8616 7346
rect 8781 7100 9089 7109
rect 8781 7098 8787 7100
rect 8843 7098 8867 7100
rect 8923 7098 8947 7100
rect 9003 7098 9027 7100
rect 9083 7098 9089 7100
rect 8843 7046 8845 7098
rect 9025 7046 9027 7098
rect 8781 7044 8787 7046
rect 8843 7044 8867 7046
rect 8923 7044 8947 7046
rect 9003 7044 9027 7046
rect 9083 7044 9089 7046
rect 8781 7035 9089 7044
rect 9140 6934 9168 8230
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9232 7449 9260 7754
rect 9324 7546 9352 8774
rect 9441 8732 9749 8741
rect 9441 8730 9447 8732
rect 9503 8730 9527 8732
rect 9583 8730 9607 8732
rect 9663 8730 9687 8732
rect 9743 8730 9749 8732
rect 9503 8678 9505 8730
rect 9685 8678 9687 8730
rect 9441 8676 9447 8678
rect 9503 8676 9527 8678
rect 9583 8676 9607 8678
rect 9663 8676 9687 8678
rect 9743 8676 9749 8678
rect 9441 8667 9749 8676
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 7834 9628 8230
rect 9956 7880 10008 7886
rect 9600 7806 9812 7834
rect 9956 7822 10008 7828
rect 9441 7644 9749 7653
rect 9441 7642 9447 7644
rect 9503 7642 9527 7644
rect 9583 7642 9607 7644
rect 9663 7642 9687 7644
rect 9743 7642 9749 7644
rect 9503 7590 9505 7642
rect 9685 7590 9687 7642
rect 9441 7588 9447 7590
rect 9503 7588 9527 7590
rect 9583 7588 9607 7590
rect 9663 7588 9687 7590
rect 9743 7588 9749 7590
rect 9441 7579 9749 7588
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9784 7478 9812 7806
rect 9772 7472 9824 7478
rect 9218 7440 9274 7449
rect 9772 7414 9824 7420
rect 9218 7375 9274 7384
rect 9232 7041 9260 7375
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9218 7032 9274 7041
rect 9218 6967 9274 6976
rect 9128 6928 9180 6934
rect 9128 6870 9180 6876
rect 9324 6854 9628 6882
rect 9220 6792 9272 6798
rect 9324 6780 9352 6854
rect 9272 6752 9352 6780
rect 9404 6792 9456 6798
rect 9220 6734 9272 6740
rect 9404 6734 9456 6740
rect 9232 6458 9260 6734
rect 9416 6662 9444 6734
rect 9600 6730 9628 6854
rect 9692 6798 9720 7210
rect 9784 6934 9812 7278
rect 9968 7274 9996 7822
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9441 6556 9749 6565
rect 9441 6554 9447 6556
rect 9503 6554 9527 6556
rect 9583 6554 9607 6556
rect 9663 6554 9687 6556
rect 9743 6554 9749 6556
rect 9503 6502 9505 6554
rect 9685 6502 9687 6554
rect 9441 6500 9447 6502
rect 9503 6500 9527 6502
rect 9583 6500 9607 6502
rect 9663 6500 9687 6502
rect 9743 6500 9749 6502
rect 9441 6491 9749 6500
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 8781 6012 9089 6021
rect 8781 6010 8787 6012
rect 8843 6010 8867 6012
rect 8923 6010 8947 6012
rect 9003 6010 9027 6012
rect 9083 6010 9089 6012
rect 8843 5958 8845 6010
rect 9025 5958 9027 6010
rect 8781 5956 8787 5958
rect 8843 5956 8867 5958
rect 8923 5956 8947 5958
rect 9003 5956 9027 5958
rect 9083 5956 9089 5958
rect 8781 5947 9089 5956
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 7392 5642 7512 5658
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 7380 5636 7512 5642
rect 7432 5630 7512 5636
rect 7380 5578 7432 5584
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5302 7328 5510
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6748 4826 6776 5238
rect 7484 5234 7512 5630
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6840 4690 6868 4966
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5684 4032 5764 4060
rect 5632 4014 5684 4020
rect 5644 3398 5672 4014
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5736 3194 5764 3402
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5460 2746 5580 2774
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5170 1456 5226 1465
rect 5170 1391 5226 1400
rect 5184 870 5304 898
rect 5184 800 5212 870
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5276 762 5304 870
rect 5460 762 5488 2746
rect 5828 800 5856 4082
rect 6840 4078 6868 4422
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5920 3058 5948 3878
rect 6932 3738 6960 4150
rect 7024 4146 7052 5102
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7024 4010 7052 4082
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 6012 3058 6040 3402
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6472 800 6500 3470
rect 7116 800 7144 4422
rect 7300 4214 7328 4490
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 3466 7512 4082
rect 7760 4010 7788 5102
rect 8220 4842 8248 5306
rect 8312 5284 8340 5646
rect 8392 5296 8444 5302
rect 8312 5256 8392 5284
rect 8392 5238 8444 5244
rect 8668 5228 8720 5234
rect 7852 4814 8248 4842
rect 8496 5188 8668 5216
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7484 3194 7512 3402
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7300 2514 7328 3062
rect 7852 2666 7880 4814
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8220 4146 8248 4694
rect 8496 4690 8524 5188
rect 8668 5170 8720 5176
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 8781 4924 9089 4933
rect 8781 4922 8787 4924
rect 8843 4922 8867 4924
rect 8923 4922 8947 4924
rect 9003 4922 9027 4924
rect 9083 4922 9089 4924
rect 8843 4870 8845 4922
rect 9025 4870 9027 4922
rect 8781 4868 8787 4870
rect 8843 4868 8867 4870
rect 8923 4868 8947 4870
rect 9003 4868 9027 4870
rect 9083 4868 9089 4870
rect 8781 4859 9089 4868
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7944 3738 7972 4082
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7760 2638 7880 2666
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7760 800 7788 2638
rect 8128 2446 8156 3606
rect 8312 3126 8340 3878
rect 8496 3534 8524 4490
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8404 800 8432 3402
rect 8588 3398 8616 4082
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8588 2650 8616 3334
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 5276 734 5488 762
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 8680 762 8708 4626
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8772 4282 8800 4490
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 9140 4146 9168 5170
rect 9232 4826 9260 6258
rect 9784 6118 9812 6598
rect 9876 6458 9904 7142
rect 9954 7032 10010 7041
rect 9954 6967 10010 6976
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9968 6225 9996 6967
rect 10060 6730 10088 9318
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10152 8090 10180 8842
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10244 7954 10272 8502
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10336 7834 10364 9930
rect 10428 9722 10456 10542
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10520 9042 10548 11086
rect 10612 10674 10640 11154
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10612 9654 10640 10610
rect 10704 10538 10732 13262
rect 10796 12850 10824 17682
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 15094 10916 15846
rect 10980 15638 11008 20742
rect 11164 19854 11192 21558
rect 11348 21554 11376 21898
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11348 20942 11376 21490
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 18426 11192 18566
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 15910 11100 17070
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10888 13258 10916 13942
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12918 10916 13194
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 11626 11100 12174
rect 11164 11830 11192 18362
rect 11256 18154 11284 19790
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11348 15978 11376 17682
rect 11440 17610 11468 22066
rect 11624 21418 11652 22578
rect 12268 21690 12296 24475
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11612 21412 11664 21418
rect 11612 21354 11664 21360
rect 11716 20330 11744 21490
rect 12268 21146 12296 21626
rect 12360 21622 12388 21830
rect 12452 21622 12480 21966
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12728 21146 12756 21490
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12912 21078 12940 24475
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 13004 22030 13032 22374
rect 13556 22094 13584 24475
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13832 22234 13860 22578
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 13556 22066 13676 22094
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13268 21956 13320 21962
rect 13268 21898 13320 21904
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 12072 20528 12124 20534
rect 12912 20516 12940 21014
rect 13096 20942 13124 21626
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 12992 20528 13044 20534
rect 12912 20488 12992 20516
rect 12072 20470 12124 20476
rect 12992 20470 13044 20476
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11808 20058 11836 20402
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11808 19718 11836 19994
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11624 19378 11652 19654
rect 12084 19514 12112 20470
rect 13096 20466 13124 20878
rect 13280 20466 13308 21898
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12268 20262 12296 20334
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12452 20058 12480 20402
rect 13280 20262 13308 20402
rect 13464 20330 13492 20810
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12820 19854 12848 20198
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 13464 19786 13492 19994
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11532 17814 11560 18634
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11624 18290 11652 18566
rect 11808 18290 11836 19110
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11440 17338 11468 17546
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11532 16794 11560 17750
rect 11624 17134 11652 18226
rect 11808 17338 11836 18226
rect 12084 18222 12112 19450
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 12360 18834 12388 19314
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12452 18358 12480 18634
rect 12728 18426 12756 18634
rect 13556 18426 13584 19314
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12544 17882 12572 18226
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11716 15910 11744 17206
rect 11808 17202 11836 17274
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11900 16794 11928 17138
rect 12268 16998 12296 17478
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12544 17082 12572 17478
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11900 16250 11928 16730
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11256 15094 11284 15438
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11440 14414 11468 15302
rect 11624 14890 11652 15438
rect 11612 14884 11664 14890
rect 11612 14826 11664 14832
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11518 12336 11574 12345
rect 11518 12271 11574 12280
rect 11532 12238 11560 12271
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10796 10674 10824 11018
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10796 9994 10824 10610
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10796 9586 10824 9930
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8566 10548 8978
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10612 8498 10640 8774
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10244 7806 10364 7834
rect 10244 6798 10272 7806
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10060 6322 10088 6666
rect 10244 6390 10272 6734
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10140 6248 10192 6254
rect 9954 6216 10010 6225
rect 10140 6190 10192 6196
rect 9954 6151 10010 6160
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9441 5468 9749 5477
rect 9441 5466 9447 5468
rect 9503 5466 9527 5468
rect 9583 5466 9607 5468
rect 9663 5466 9687 5468
rect 9743 5466 9749 5468
rect 9503 5414 9505 5466
rect 9685 5414 9687 5466
rect 9441 5412 9447 5414
rect 9503 5412 9527 5414
rect 9583 5412 9607 5414
rect 9663 5412 9687 5414
rect 9743 5412 9749 5414
rect 9441 5403 9749 5412
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9324 4486 9352 5238
rect 9876 5234 9904 5714
rect 9968 5642 9996 6151
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10060 5370 10088 5578
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9876 4706 9904 5170
rect 9784 4678 9904 4706
rect 9784 4622 9812 4678
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9441 4380 9749 4389
rect 9441 4378 9447 4380
rect 9503 4378 9527 4380
rect 9583 4378 9607 4380
rect 9663 4378 9687 4380
rect 9743 4378 9749 4380
rect 9503 4326 9505 4378
rect 9685 4326 9687 4378
rect 9441 4324 9447 4326
rect 9503 4324 9527 4326
rect 9583 4324 9607 4326
rect 9663 4324 9687 4326
rect 9743 4324 9749 4326
rect 9441 4315 9749 4324
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8781 3836 9089 3845
rect 8781 3834 8787 3836
rect 8843 3834 8867 3836
rect 8923 3834 8947 3836
rect 9003 3834 9027 3836
rect 9083 3834 9089 3836
rect 8843 3782 8845 3834
rect 9025 3782 9027 3834
rect 8781 3780 8787 3782
rect 8843 3780 8867 3782
rect 8923 3780 8947 3782
rect 9003 3780 9027 3782
rect 9083 3780 9089 3782
rect 8781 3771 9089 3780
rect 9140 2854 9168 4082
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9508 3466 9536 4014
rect 9784 3602 9812 4558
rect 10152 4078 10180 6190
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9496 3460 9548 3466
rect 9324 3420 9496 3448
rect 9324 3194 9352 3420
rect 9496 3402 9548 3408
rect 9441 3292 9749 3301
rect 9441 3290 9447 3292
rect 9503 3290 9527 3292
rect 9583 3290 9607 3292
rect 9663 3290 9687 3292
rect 9743 3290 9749 3292
rect 9503 3238 9505 3290
rect 9685 3238 9687 3290
rect 9441 3236 9447 3238
rect 9503 3236 9527 3238
rect 9583 3236 9607 3238
rect 9663 3236 9687 3238
rect 9743 3236 9749 3238
rect 9441 3227 9749 3236
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9784 3058 9812 3538
rect 10152 3534 10180 3878
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 8781 2748 9089 2757
rect 8781 2746 8787 2748
rect 8843 2746 8867 2748
rect 8923 2746 8947 2748
rect 9003 2746 9027 2748
rect 9083 2746 9089 2748
rect 8843 2694 8845 2746
rect 9025 2694 9027 2746
rect 8781 2692 8787 2694
rect 8843 2692 8867 2694
rect 8923 2692 8947 2694
rect 9003 2692 9027 2694
rect 9083 2692 9089 2694
rect 8781 2683 9089 2692
rect 9441 2204 9749 2213
rect 9441 2202 9447 2204
rect 9503 2202 9527 2204
rect 9583 2202 9607 2204
rect 9663 2202 9687 2204
rect 9743 2202 9749 2204
rect 9503 2150 9505 2202
rect 9685 2150 9687 2202
rect 9441 2148 9447 2150
rect 9503 2148 9527 2150
rect 9583 2148 9607 2150
rect 9663 2148 9687 2150
rect 9743 2148 9749 2150
rect 9441 2139 9749 2148
rect 9876 1714 9904 3402
rect 9692 1686 9904 1714
rect 8956 870 9076 898
rect 8956 762 8984 870
rect 9048 800 9076 870
rect 9692 800 9720 1686
rect 10336 800 10364 7482
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10428 4214 10456 6666
rect 10520 6390 10548 6666
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10966 6352 11022 6361
rect 10966 6287 10968 6296
rect 11020 6287 11022 6296
rect 10968 6258 11020 6264
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5710 11100 6054
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11164 5522 11192 11766
rect 11256 11150 11284 12038
rect 11348 11830 11376 12038
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11624 11354 11652 11630
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11256 10266 11284 10610
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11532 9042 11560 10542
rect 11716 9194 11744 15846
rect 12084 15094 12112 16050
rect 12176 15706 12204 16526
rect 12268 16182 12296 16934
rect 12452 16590 12480 17070
rect 12544 17054 12664 17082
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12636 15042 12664 17054
rect 12728 15450 12756 17546
rect 12820 17270 12848 18022
rect 13004 17882 13032 18226
rect 13188 18086 13216 18294
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 13096 17610 13124 17750
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 13096 16114 13124 17546
rect 13188 17542 13216 18022
rect 13648 17762 13676 22066
rect 13924 21894 13952 24534
rect 14108 24426 14136 24534
rect 14186 24475 14242 25275
rect 14384 24534 14780 24562
rect 14200 24426 14228 24475
rect 14108 24398 14228 24426
rect 14002 22332 14310 22341
rect 14002 22330 14008 22332
rect 14064 22330 14088 22332
rect 14144 22330 14168 22332
rect 14224 22330 14248 22332
rect 14304 22330 14310 22332
rect 14064 22278 14066 22330
rect 14246 22278 14248 22330
rect 14002 22276 14008 22278
rect 14064 22276 14088 22278
rect 14144 22276 14168 22278
rect 14224 22276 14248 22278
rect 14304 22276 14310 22278
rect 14002 22267 14310 22276
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13740 19360 13768 21830
rect 14002 21244 14310 21253
rect 14002 21242 14008 21244
rect 14064 21242 14088 21244
rect 14144 21242 14168 21244
rect 14224 21242 14248 21244
rect 14304 21242 14310 21244
rect 14064 21190 14066 21242
rect 14246 21190 14248 21242
rect 14002 21188 14008 21190
rect 14064 21188 14088 21190
rect 14144 21188 14168 21190
rect 14224 21188 14248 21190
rect 14304 21188 14310 21190
rect 14002 21179 14310 21188
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13832 19786 13860 20742
rect 13924 19922 13952 20946
rect 14002 20156 14310 20165
rect 14002 20154 14008 20156
rect 14064 20154 14088 20156
rect 14144 20154 14168 20156
rect 14224 20154 14248 20156
rect 14304 20154 14310 20156
rect 14064 20102 14066 20154
rect 14246 20102 14248 20154
rect 14002 20100 14008 20102
rect 14064 20100 14088 20102
rect 14144 20100 14168 20102
rect 14224 20100 14248 20102
rect 14304 20100 14310 20102
rect 14002 20091 14310 20100
rect 14384 20074 14412 24534
rect 14752 24426 14780 24534
rect 14830 24475 14886 25275
rect 16118 24475 16174 25275
rect 16762 24475 16818 25275
rect 17406 24475 17462 25275
rect 18050 24475 18106 25275
rect 19338 24475 19394 25275
rect 14844 24426 14872 24475
rect 14752 24398 14872 24426
rect 14662 22876 14970 22885
rect 14662 22874 14668 22876
rect 14724 22874 14748 22876
rect 14804 22874 14828 22876
rect 14884 22874 14908 22876
rect 14964 22874 14970 22876
rect 14724 22822 14726 22874
rect 14906 22822 14908 22874
rect 14662 22820 14668 22822
rect 14724 22820 14748 22822
rect 14804 22820 14828 22822
rect 14884 22820 14908 22822
rect 14964 22820 14970 22822
rect 14662 22811 14970 22820
rect 16028 22568 16080 22574
rect 16028 22510 16080 22516
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14476 20942 14504 21286
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14476 20602 14504 20878
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14568 20330 14596 21898
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 14662 21788 14970 21797
rect 14662 21786 14668 21788
rect 14724 21786 14748 21788
rect 14804 21786 14828 21788
rect 14884 21786 14908 21788
rect 14964 21786 14970 21788
rect 14724 21734 14726 21786
rect 14906 21734 14908 21786
rect 14662 21732 14668 21734
rect 14724 21732 14748 21734
rect 14804 21732 14828 21734
rect 14884 21732 14908 21734
rect 14964 21732 14970 21734
rect 14662 21723 14970 21732
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14844 21146 14872 21490
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 15028 20942 15056 21830
rect 15120 21622 15148 22034
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 15120 21078 15148 21558
rect 15304 21350 15332 21898
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15108 21072 15160 21078
rect 15108 21014 15160 21020
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 14662 20700 14970 20709
rect 14662 20698 14668 20700
rect 14724 20698 14748 20700
rect 14804 20698 14828 20700
rect 14884 20698 14908 20700
rect 14964 20698 14970 20700
rect 14724 20646 14726 20698
rect 14906 20646 14908 20698
rect 14662 20644 14668 20646
rect 14724 20644 14748 20646
rect 14804 20644 14828 20646
rect 14884 20644 14908 20646
rect 14964 20644 14970 20646
rect 14662 20635 14970 20644
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14556 20324 14608 20330
rect 14556 20266 14608 20272
rect 14384 20046 14596 20074
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13924 19446 13952 19858
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13740 19332 13860 19360
rect 13832 18290 13860 19332
rect 13924 18834 13952 19382
rect 14292 19156 14320 19790
rect 14292 19128 14412 19156
rect 14002 19068 14310 19077
rect 14002 19066 14008 19068
rect 14064 19066 14088 19068
rect 14144 19066 14168 19068
rect 14224 19066 14248 19068
rect 14304 19066 14310 19068
rect 14064 19014 14066 19066
rect 14246 19014 14248 19066
rect 14002 19012 14008 19014
rect 14064 19012 14088 19014
rect 14144 19012 14168 19014
rect 14224 19012 14248 19014
rect 14304 19012 14310 19014
rect 14002 19003 14310 19012
rect 14384 18970 14412 19128
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14280 18896 14332 18902
rect 14280 18838 14332 18844
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13556 17734 13676 17762
rect 13832 17746 13860 18226
rect 14292 18204 14320 18838
rect 14384 18358 14412 18906
rect 14476 18358 14504 19926
rect 14568 19514 14596 20046
rect 14752 19825 14780 20334
rect 14738 19816 14794 19825
rect 14738 19751 14740 19760
rect 14792 19751 14794 19760
rect 14740 19722 14792 19728
rect 14662 19612 14970 19621
rect 14662 19610 14668 19612
rect 14724 19610 14748 19612
rect 14804 19610 14828 19612
rect 14884 19610 14908 19612
rect 14964 19610 14970 19612
rect 14724 19558 14726 19610
rect 14906 19558 14908 19610
rect 14662 19556 14668 19558
rect 14724 19556 14748 19558
rect 14804 19556 14828 19558
rect 14884 19556 14908 19558
rect 14964 19556 14970 19558
rect 14662 19547 14970 19556
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14568 18426 14596 19450
rect 14738 19408 14794 19417
rect 14738 19343 14794 19352
rect 14752 18902 14780 19343
rect 15028 19174 15056 20742
rect 15304 20534 15332 21286
rect 15396 20874 15424 21830
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15580 19922 15608 21898
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15200 19848 15252 19854
rect 15672 19802 15700 21490
rect 15764 20874 15792 21830
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15948 20330 15976 21966
rect 16040 21350 16068 22510
rect 16132 21690 16160 24475
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16408 22506 16436 22578
rect 16396 22500 16448 22506
rect 16396 22442 16448 22448
rect 16120 21684 16172 21690
rect 16120 21626 16172 21632
rect 16408 21418 16436 22442
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16684 22030 16712 22374
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16776 21672 16804 24475
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16684 21644 16804 21672
rect 16396 21412 16448 21418
rect 16396 21354 16448 21360
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 16408 20534 16436 21354
rect 16396 20528 16448 20534
rect 16396 20470 16448 20476
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15936 20324 15988 20330
rect 15936 20266 15988 20272
rect 15200 19790 15252 19796
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15120 19446 15148 19654
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15212 18970 15240 19790
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15580 19774 15700 19802
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 15488 18766 15516 19722
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 14662 18524 14970 18533
rect 14662 18522 14668 18524
rect 14724 18522 14748 18524
rect 14804 18522 14828 18524
rect 14884 18522 14908 18524
rect 14964 18522 14970 18524
rect 14724 18470 14726 18522
rect 14906 18470 14908 18522
rect 14662 18468 14668 18470
rect 14724 18468 14748 18470
rect 14804 18468 14828 18470
rect 14884 18468 14908 18470
rect 14964 18468 14970 18470
rect 14662 18459 14970 18468
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14464 18352 14516 18358
rect 15028 18329 15056 18634
rect 14464 18294 14516 18300
rect 15014 18320 15070 18329
rect 15014 18255 15070 18264
rect 15108 18284 15160 18290
rect 14292 18176 14504 18204
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14002 17980 14310 17989
rect 14002 17978 14008 17980
rect 14064 17978 14088 17980
rect 14144 17978 14168 17980
rect 14224 17978 14248 17980
rect 14304 17978 14310 17980
rect 14064 17926 14066 17978
rect 14246 17926 14248 17978
rect 14002 17924 14008 17926
rect 14064 17924 14088 17926
rect 14144 17924 14168 17926
rect 14224 17924 14248 17926
rect 14304 17924 14310 17926
rect 14002 17915 14310 17924
rect 13820 17740 13872 17746
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13464 17338 13492 17546
rect 13556 17542 13584 17734
rect 13820 17682 13872 17688
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 13372 15502 13400 17274
rect 13556 17066 13584 17478
rect 13648 17202 13676 17614
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13740 17270 13768 17478
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13648 16590 13676 17138
rect 13832 16794 13860 17206
rect 14002 16892 14310 16901
rect 14002 16890 14008 16892
rect 14064 16890 14088 16892
rect 14144 16890 14168 16892
rect 14224 16890 14248 16892
rect 14304 16890 14310 16892
rect 14064 16838 14066 16890
rect 14246 16838 14248 16890
rect 14002 16836 14008 16838
rect 14064 16836 14088 16838
rect 14144 16836 14168 16838
rect 14224 16836 14248 16838
rect 14304 16836 14310 16838
rect 14002 16827 14310 16836
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13360 15496 13412 15502
rect 12728 15422 12848 15450
rect 13360 15438 13412 15444
rect 12820 15366 12848 15422
rect 13464 15366 13492 16118
rect 13648 16046 13676 16526
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 11980 15020 12032 15026
rect 12636 15014 12756 15042
rect 11980 14962 12032 14968
rect 11992 14618 12020 14962
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11808 12850 11836 13738
rect 12268 13394 12296 14350
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12360 13258 12388 14010
rect 12452 13530 12480 14282
rect 12636 14006 12664 14894
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12636 13870 12664 13942
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12728 13682 12756 15014
rect 12636 13654 12756 13682
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 11808 10810 11836 12786
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12442 12480 12582
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11900 11354 11928 11494
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 12452 11098 12480 12038
rect 12544 11812 12572 12786
rect 12636 12170 12664 13654
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12728 12102 12756 12854
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12544 11784 12664 11812
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12360 11082 12480 11098
rect 12360 11076 12492 11082
rect 12360 11070 12440 11076
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 10266 12112 10610
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12360 10062 12388 11070
rect 12440 11018 12492 11024
rect 12544 10810 12572 11630
rect 12636 11558 12664 11784
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12820 11370 12848 15302
rect 13176 15020 13228 15026
rect 13228 14980 13308 15008
rect 13176 14962 13228 14968
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12912 14074 12940 14554
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13004 12782 13032 14758
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13188 12918 13216 13942
rect 13280 13734 13308 14980
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 13938 13492 14758
rect 13556 14278 13584 14894
rect 13648 14482 13676 15982
rect 13832 15570 13860 16730
rect 14384 16590 14412 18022
rect 14476 17082 14504 18176
rect 15028 17610 15056 18255
rect 15108 18226 15160 18232
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 14662 17436 14970 17445
rect 14662 17434 14668 17436
rect 14724 17434 14748 17436
rect 14804 17434 14828 17436
rect 14884 17434 14908 17436
rect 14964 17434 14970 17436
rect 14724 17382 14726 17434
rect 14906 17382 14908 17434
rect 14662 17380 14668 17382
rect 14724 17380 14748 17382
rect 14804 17380 14828 17382
rect 14884 17380 14908 17382
rect 14964 17380 14970 17382
rect 14662 17371 14970 17380
rect 15028 17241 15056 17546
rect 15014 17232 15070 17241
rect 15014 17167 15070 17176
rect 14648 17128 14700 17134
rect 14476 17076 14648 17082
rect 14476 17070 14700 17076
rect 14476 17054 14688 17070
rect 14476 16998 14504 17054
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14462 16144 14518 16153
rect 14462 16079 14518 16088
rect 14476 15910 14504 16079
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14002 15804 14310 15813
rect 14002 15802 14008 15804
rect 14064 15802 14088 15804
rect 14144 15802 14168 15804
rect 14224 15802 14248 15804
rect 14304 15802 14310 15804
rect 14064 15750 14066 15802
rect 14246 15750 14248 15802
rect 14002 15748 14008 15750
rect 14064 15748 14088 15750
rect 14144 15748 14168 15750
rect 14224 15748 14248 15750
rect 14304 15748 14310 15750
rect 14002 15739 14310 15748
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 14002 14716 14310 14725
rect 14002 14714 14008 14716
rect 14064 14714 14088 14716
rect 14144 14714 14168 14716
rect 14224 14714 14248 14716
rect 14304 14714 14310 14716
rect 14064 14662 14066 14714
rect 14246 14662 14248 14714
rect 14002 14660 14008 14662
rect 14064 14660 14088 14662
rect 14144 14660 14168 14662
rect 14224 14660 14248 14662
rect 14304 14660 14310 14662
rect 14002 14651 14310 14660
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 14074 13584 14214
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13542 13968 13598 13977
rect 13452 13932 13504 13938
rect 13542 13903 13598 13912
rect 13452 13874 13504 13880
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13280 12782 13308 13670
rect 13464 13530 13492 13874
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 12992 12776 13044 12782
rect 12636 11342 12848 11370
rect 12912 12724 12992 12730
rect 12912 12718 13044 12724
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 12912 12702 13032 12718
rect 12636 11014 12664 11342
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12544 10130 12572 10746
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12348 10056 12400 10062
rect 12636 10010 12664 10950
rect 12348 9998 12400 10004
rect 12544 9982 12664 10010
rect 12820 9994 12848 11222
rect 12912 10130 12940 12702
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13004 10266 13032 12378
rect 13266 12336 13322 12345
rect 13266 12271 13268 12280
rect 13320 12271 13322 12280
rect 13268 12242 13320 12248
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11082 13124 11494
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 13096 10062 13124 11018
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12808 9988 12860 9994
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 11716 9166 11836 9194
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11256 7750 11284 8842
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11440 8362 11468 8774
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 7886 11560 8230
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11624 7274 11652 8910
rect 11716 8498 11744 9046
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11072 5494 11192 5522
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10980 3398 11008 4014
rect 11072 3942 11100 5494
rect 11256 5370 11284 6326
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11624 5302 11652 5510
rect 11808 5302 11836 9166
rect 12176 8906 12204 9318
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12360 8498 12388 8842
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11900 8242 11928 8298
rect 12072 8288 12124 8294
rect 11900 8214 12020 8242
rect 12072 8230 12124 8236
rect 11992 7478 12020 8214
rect 12084 7886 12112 8230
rect 12360 8090 12388 8434
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12176 6390 12204 6598
rect 12268 6458 12296 6598
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 11888 6316 11940 6322
rect 11940 6276 12020 6304
rect 11888 6258 11940 6264
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11900 5234 11928 5782
rect 11992 5710 12020 6276
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12176 5710 12204 6054
rect 11980 5704 12032 5710
rect 12164 5704 12216 5710
rect 12032 5664 12112 5692
rect 11980 5646 12032 5652
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 11716 4622 11744 5034
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4622 11836 4966
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 4214 11744 4422
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10980 800 11008 3334
rect 11072 2446 11100 3878
rect 11164 3194 11192 4150
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11164 2310 11192 3130
rect 11348 2650 11376 3470
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11440 3126 11468 3334
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11532 2990 11560 3402
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11532 2514 11560 2926
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11808 2446 11836 3334
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11624 870 11744 898
rect 11624 800 11652 870
rect 8680 734 8984 762
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 11716 762 11744 870
rect 11900 762 11928 5170
rect 12084 4622 12112 5664
rect 12164 5646 12216 5652
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 4078 12112 4558
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12084 3466 12112 4014
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12360 2774 12388 7686
rect 12452 7290 12480 9862
rect 12544 8430 12572 9982
rect 12808 9930 12860 9936
rect 13188 9926 13216 12106
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13280 11218 13308 11834
rect 13372 11354 13400 12174
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13464 11762 13492 12038
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 10538 13308 11154
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13464 10810 13492 11018
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12636 8566 12664 9590
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12636 8090 12664 8502
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12728 7818 12756 8366
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12728 7426 12756 7754
rect 12636 7398 12756 7426
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12636 7342 12664 7398
rect 12624 7336 12676 7342
rect 12452 7262 12572 7290
rect 12624 7278 12676 7284
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6798 12480 7142
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12544 3602 12572 7262
rect 12636 6322 12664 7278
rect 12912 6730 12940 7414
rect 13188 6730 13216 8774
rect 13464 8566 13492 8774
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13556 7410 13584 13903
rect 13740 12714 13768 14350
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13924 14006 13952 14214
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 14384 13870 14412 14418
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13326 13860 13670
rect 14002 13628 14310 13637
rect 14002 13626 14008 13628
rect 14064 13626 14088 13628
rect 14144 13626 14168 13628
rect 14224 13626 14248 13628
rect 14304 13626 14310 13628
rect 14064 13574 14066 13626
rect 14246 13574 14248 13626
rect 14002 13572 14008 13574
rect 14064 13572 14088 13574
rect 14144 13572 14168 13574
rect 14224 13572 14248 13574
rect 14304 13572 14310 13574
rect 14002 13563 14310 13572
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 14384 12782 14412 13806
rect 14476 13258 14504 15846
rect 14568 15570 14596 16934
rect 14662 16348 14970 16357
rect 14662 16346 14668 16348
rect 14724 16346 14748 16348
rect 14804 16346 14828 16348
rect 14884 16346 14908 16348
rect 14964 16346 14970 16348
rect 14724 16294 14726 16346
rect 14906 16294 14908 16346
rect 14662 16292 14668 16294
rect 14724 16292 14748 16294
rect 14804 16292 14828 16294
rect 14884 16292 14908 16294
rect 14964 16292 14970 16294
rect 14662 16283 14970 16292
rect 15120 15706 15148 18226
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15212 17270 15240 17750
rect 15580 17610 15608 19774
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15672 18426 15700 18566
rect 15660 18420 15712 18426
rect 15660 18362 15712 18368
rect 15844 17808 15896 17814
rect 15844 17750 15896 17756
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15488 17338 15516 17546
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15580 16572 15608 17546
rect 15672 16998 15700 17546
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15672 16726 15700 16934
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15580 16544 15792 16572
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14662 15260 14970 15269
rect 14662 15258 14668 15260
rect 14724 15258 14748 15260
rect 14804 15258 14828 15260
rect 14884 15258 14908 15260
rect 14964 15258 14970 15260
rect 14724 15206 14726 15258
rect 14906 15206 14908 15258
rect 14662 15204 14668 15206
rect 14724 15204 14748 15206
rect 14804 15204 14828 15206
rect 14884 15204 14908 15206
rect 14964 15204 14970 15206
rect 14662 15195 14970 15204
rect 15488 15162 15516 16050
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15638 15700 15846
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14752 14414 14780 14826
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 14414 15332 14758
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14662 14172 14970 14181
rect 14662 14170 14668 14172
rect 14724 14170 14748 14172
rect 14804 14170 14828 14172
rect 14884 14170 14908 14172
rect 14964 14170 14970 14172
rect 14724 14118 14726 14170
rect 14906 14118 14908 14170
rect 14662 14116 14668 14118
rect 14724 14116 14748 14118
rect 14804 14116 14828 14118
rect 14884 14116 14908 14118
rect 14964 14116 14970 14118
rect 14662 14107 14970 14116
rect 14832 14000 14884 14006
rect 14830 13968 14832 13977
rect 14884 13968 14886 13977
rect 14830 13903 14886 13912
rect 15488 13870 15516 14962
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13648 11286 13676 12650
rect 14002 12540 14310 12549
rect 14002 12538 14008 12540
rect 14064 12538 14088 12540
rect 14144 12538 14168 12540
rect 14224 12538 14248 12540
rect 14304 12538 14310 12540
rect 14064 12486 14066 12538
rect 14246 12486 14248 12538
rect 14002 12484 14008 12486
rect 14064 12484 14088 12486
rect 14144 12484 14168 12486
rect 14224 12484 14248 12486
rect 14304 12484 14310 12486
rect 14002 12475 14310 12484
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11898 13768 12174
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13832 11354 13860 11698
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14002 11452 14310 11461
rect 14002 11450 14008 11452
rect 14064 11450 14088 11452
rect 14144 11450 14168 11452
rect 14224 11450 14248 11452
rect 14304 11450 14310 11452
rect 14064 11398 14066 11450
rect 14246 11398 14248 11450
rect 14002 11396 14008 11398
rect 14064 11396 14088 11398
rect 14144 11396 14168 11398
rect 14224 11396 14248 11398
rect 14304 11396 14310 11398
rect 14002 11387 14310 11396
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 14384 10742 14412 11494
rect 14476 11014 14504 13194
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12850 14596 13126
rect 14662 13084 14970 13093
rect 14662 13082 14668 13084
rect 14724 13082 14748 13084
rect 14804 13082 14828 13084
rect 14884 13082 14908 13084
rect 14964 13082 14970 13084
rect 14724 13030 14726 13082
rect 14906 13030 14908 13082
rect 14662 13028 14668 13030
rect 14724 13028 14748 13030
rect 14804 13028 14828 13030
rect 14884 13028 14908 13030
rect 14964 13028 14970 13030
rect 14662 13019 14970 13028
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 15016 12232 15068 12238
rect 15068 12180 15148 12186
rect 15016 12174 15148 12180
rect 15028 12158 15148 12174
rect 14662 11996 14970 12005
rect 14662 11994 14668 11996
rect 14724 11994 14748 11996
rect 14804 11994 14828 11996
rect 14884 11994 14908 11996
rect 14964 11994 14970 11996
rect 14724 11942 14726 11994
rect 14906 11942 14908 11994
rect 14662 11940 14668 11942
rect 14724 11940 14748 11942
rect 14804 11940 14828 11942
rect 14884 11940 14908 11942
rect 14964 11940 14970 11942
rect 14662 11931 14970 11940
rect 15120 11626 15148 12158
rect 15672 11762 15700 13874
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 15120 11150 15148 11562
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 14662 10908 14970 10917
rect 14662 10906 14668 10908
rect 14724 10906 14748 10908
rect 14804 10906 14828 10908
rect 14884 10906 14908 10908
rect 14964 10906 14970 10908
rect 14724 10854 14726 10906
rect 14906 10854 14908 10906
rect 14662 10852 14668 10854
rect 14724 10852 14748 10854
rect 14804 10852 14828 10854
rect 14884 10852 14908 10854
rect 14964 10852 14970 10854
rect 14662 10843 14970 10852
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14002 10364 14310 10373
rect 14002 10362 14008 10364
rect 14064 10362 14088 10364
rect 14144 10362 14168 10364
rect 14224 10362 14248 10364
rect 14304 10362 14310 10364
rect 14064 10310 14066 10362
rect 14246 10310 14248 10362
rect 14002 10308 14008 10310
rect 14064 10308 14088 10310
rect 14144 10308 14168 10310
rect 14224 10308 14248 10310
rect 14304 10308 14310 10310
rect 14002 10299 14310 10308
rect 14384 10062 14412 10406
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14662 9820 14970 9829
rect 14662 9818 14668 9820
rect 14724 9818 14748 9820
rect 14804 9818 14828 9820
rect 14884 9818 14908 9820
rect 14964 9818 14970 9820
rect 14724 9766 14726 9818
rect 14906 9766 14908 9818
rect 14662 9764 14668 9766
rect 14724 9764 14748 9766
rect 14804 9764 14828 9766
rect 14884 9764 14908 9766
rect 14964 9764 14970 9766
rect 14662 9755 14970 9764
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 13820 9512 13872 9518
rect 13872 9460 13952 9466
rect 13820 9454 13952 9460
rect 13832 9438 13952 9454
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 8974 13768 9318
rect 13924 9110 13952 9438
rect 14002 9276 14310 9285
rect 14002 9274 14008 9276
rect 14064 9274 14088 9276
rect 14144 9274 14168 9276
rect 14224 9274 14248 9276
rect 14304 9274 14310 9276
rect 14064 9222 14066 9274
rect 14246 9222 14248 9274
rect 14002 9220 14008 9222
rect 14064 9220 14088 9222
rect 14144 9220 14168 9222
rect 14224 9220 14248 9222
rect 14304 9220 14310 9222
rect 14002 9211 14310 9220
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13832 8090 13860 8842
rect 13924 8362 13952 9046
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 8566 14136 8978
rect 14384 8634 14412 9590
rect 14662 8732 14970 8741
rect 14662 8730 14668 8732
rect 14724 8730 14748 8732
rect 14804 8730 14828 8732
rect 14884 8730 14908 8732
rect 14964 8730 14970 8732
rect 14724 8678 14726 8730
rect 14906 8678 14908 8730
rect 14662 8676 14668 8678
rect 14724 8676 14748 8678
rect 14804 8676 14828 8678
rect 14884 8676 14908 8678
rect 14964 8676 14970 8678
rect 14662 8667 14970 8676
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 14002 8188 14310 8197
rect 14002 8186 14008 8188
rect 14064 8186 14088 8188
rect 14144 8186 14168 8188
rect 14224 8186 14248 8188
rect 14304 8186 14310 8188
rect 14064 8134 14066 8186
rect 14246 8134 14248 8186
rect 14002 8132 14008 8134
rect 14064 8132 14088 8134
rect 14144 8132 14168 8134
rect 14224 8132 14248 8134
rect 14304 8132 14310 8134
rect 14002 8123 14310 8132
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14016 7410 14044 7890
rect 14292 7410 14320 7958
rect 14384 7750 14412 8570
rect 14556 8560 14608 8566
rect 14462 8528 14518 8537
rect 14556 8502 14608 8508
rect 14462 8463 14464 8472
rect 14516 8463 14518 8472
rect 14464 8434 14516 8440
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14002 7100 14310 7109
rect 14002 7098 14008 7100
rect 14064 7098 14088 7100
rect 14144 7098 14168 7100
rect 14224 7098 14248 7100
rect 14304 7098 14310 7100
rect 14064 7046 14066 7098
rect 14246 7046 14248 7098
rect 14002 7044 14008 7046
rect 14064 7044 14088 7046
rect 14144 7044 14168 7046
rect 14224 7044 14248 7046
rect 14304 7044 14310 7046
rect 14002 7035 14310 7044
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 12912 6458 12940 6666
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12636 5166 12664 6258
rect 13188 5370 13216 6666
rect 13450 6488 13506 6497
rect 13450 6423 13506 6432
rect 13464 6390 13492 6423
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13464 6225 13492 6326
rect 13820 6248 13872 6254
rect 13450 6216 13506 6225
rect 13820 6190 13872 6196
rect 13450 6151 13506 6160
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5710 13768 6054
rect 13832 5710 13860 6190
rect 13924 5914 13952 6802
rect 14002 6012 14310 6021
rect 14002 6010 14008 6012
rect 14064 6010 14088 6012
rect 14144 6010 14168 6012
rect 14224 6010 14248 6012
rect 14304 6010 14310 6012
rect 14064 5958 14066 6010
rect 14246 5958 14248 6010
rect 14002 5956 14008 5958
rect 14064 5956 14088 5958
rect 14144 5956 14168 5958
rect 14224 5956 14248 5958
rect 14304 5956 14310 5958
rect 14002 5947 14310 5956
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12544 3126 12572 3538
rect 12636 3466 12664 5102
rect 13464 4826 13492 5238
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13740 4282 13768 5170
rect 13832 5030 13860 5646
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12268 2746 12388 2774
rect 12268 800 12296 2746
rect 12636 2650 12664 3402
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12912 800 12940 2858
rect 13004 2650 13032 3334
rect 13188 2922 13216 3402
rect 13372 3058 13400 3606
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13556 800 13584 4218
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13740 3534 13768 4014
rect 13832 4010 13860 4966
rect 14002 4924 14310 4933
rect 14002 4922 14008 4924
rect 14064 4922 14088 4924
rect 14144 4922 14168 4924
rect 14224 4922 14248 4924
rect 14304 4922 14310 4924
rect 14064 4870 14066 4922
rect 14246 4870 14248 4922
rect 14002 4868 14008 4870
rect 14064 4868 14088 4870
rect 14144 4868 14168 4870
rect 14224 4868 14248 4870
rect 14304 4868 14310 4870
rect 14002 4859 14310 4868
rect 14384 4282 14412 5306
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13832 3602 13860 3946
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 2938 13768 3334
rect 13832 3058 13860 3538
rect 13924 3126 13952 3878
rect 14002 3836 14310 3845
rect 14002 3834 14008 3836
rect 14064 3834 14088 3836
rect 14144 3834 14168 3836
rect 14224 3834 14248 3836
rect 14304 3834 14310 3836
rect 14064 3782 14066 3834
rect 14246 3782 14248 3834
rect 14002 3780 14008 3782
rect 14064 3780 14088 3782
rect 14144 3780 14168 3782
rect 14224 3780 14248 3782
rect 14304 3780 14310 3782
rect 14002 3771 14310 3780
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14384 2938 14412 4218
rect 13740 2910 14412 2938
rect 13832 2446 13860 2910
rect 14002 2748 14310 2757
rect 14002 2746 14008 2748
rect 14064 2746 14088 2748
rect 14144 2746 14168 2748
rect 14224 2746 14248 2748
rect 14304 2746 14310 2748
rect 14064 2694 14066 2746
rect 14246 2694 14248 2746
rect 14002 2692 14008 2694
rect 14064 2692 14088 2694
rect 14144 2692 14168 2694
rect 14224 2692 14248 2694
rect 14304 2692 14310 2694
rect 14002 2683 14310 2692
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14200 870 14320 898
rect 14200 800 14228 870
rect 11716 734 11928 762
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14292 762 14320 870
rect 14476 762 14504 8298
rect 14568 7410 14596 8502
rect 15028 7886 15056 10950
rect 15120 10674 15148 11086
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15120 8974 15148 10610
rect 15304 10266 15332 10610
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15580 10062 15608 11494
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15396 9586 15424 9998
rect 15672 9586 15700 11698
rect 15764 10266 15792 16544
rect 15856 16182 15884 17750
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 15948 15978 15976 17070
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15948 15502 15976 15914
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15856 14278 15884 15030
rect 16040 14618 16068 20402
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 16224 19514 16252 19722
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16120 18896 16172 18902
rect 16120 18838 16172 18844
rect 16132 18698 16160 18838
rect 16684 18698 16712 21644
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 16776 20330 16804 21490
rect 16868 21146 16896 22510
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16868 20602 16896 21082
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 17052 20534 17080 21626
rect 17040 20528 17092 20534
rect 17040 20470 17092 20476
rect 17328 20466 17356 22374
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 16856 20392 16908 20398
rect 17132 20392 17184 20398
rect 16908 20352 17132 20380
rect 16856 20334 16908 20340
rect 17132 20334 17184 20340
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16684 18358 16712 18634
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16776 18154 16804 19722
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16868 19360 16896 19654
rect 16948 19372 17000 19378
rect 16868 19332 16948 19360
rect 16948 19314 17000 19320
rect 17052 18766 17080 19926
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17144 18630 17172 19722
rect 17236 19718 17264 20198
rect 17420 19854 17448 24475
rect 17868 22704 17920 22710
rect 18064 22658 18092 24475
rect 19352 22710 19380 24475
rect 19883 22876 20191 22885
rect 19883 22874 19889 22876
rect 19945 22874 19969 22876
rect 20025 22874 20049 22876
rect 20105 22874 20129 22876
rect 20185 22874 20191 22876
rect 19945 22822 19947 22874
rect 20127 22822 20129 22874
rect 19883 22820 19889 22822
rect 19945 22820 19969 22822
rect 20025 22820 20049 22822
rect 20105 22820 20129 22822
rect 20185 22820 20191 22822
rect 19883 22811 20191 22820
rect 17920 22652 18092 22658
rect 17868 22646 18092 22652
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19616 22704 19668 22710
rect 19616 22646 19668 22652
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 17880 22630 18092 22646
rect 18064 22098 18092 22630
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18708 22488 18736 22578
rect 18788 22500 18840 22506
rect 18708 22460 18788 22488
rect 18788 22442 18840 22448
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17512 20602 17540 20810
rect 17868 20800 17920 20806
rect 17972 20754 18000 21898
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 17920 20748 18000 20754
rect 17868 20742 18000 20748
rect 17880 20726 18000 20742
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 16590 16620 17478
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16592 16114 16620 16390
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16684 15978 16712 17614
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16776 16250 16804 16934
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16868 15706 16896 17614
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16960 16114 16988 17478
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 17052 15910 17080 17206
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 17052 15570 17080 15846
rect 17144 15570 17172 18566
rect 17236 17678 17264 19654
rect 17420 19514 17448 19790
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17604 18970 17632 19722
rect 17880 19718 17908 20726
rect 18064 20466 18092 21830
rect 18524 21554 18552 22374
rect 19223 22332 19531 22341
rect 19223 22330 19229 22332
rect 19285 22330 19309 22332
rect 19365 22330 19389 22332
rect 19445 22330 19469 22332
rect 19525 22330 19531 22332
rect 19285 22278 19287 22330
rect 19467 22278 19469 22330
rect 19223 22276 19229 22278
rect 19285 22276 19309 22278
rect 19365 22276 19389 22278
rect 19445 22276 19469 22278
rect 19525 22276 19531 22278
rect 19223 22267 19531 22276
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18602 21040 18658 21049
rect 18602 20975 18658 20984
rect 18420 20596 18472 20602
rect 18420 20538 18472 20544
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 18340 19922 18368 20470
rect 18432 20058 18460 20538
rect 18512 20324 18564 20330
rect 18512 20266 18564 20272
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17604 18426 17632 18906
rect 17880 18630 17908 19654
rect 18064 18970 18092 19790
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17868 18624 17920 18630
rect 17866 18592 17868 18601
rect 17920 18592 17922 18601
rect 17866 18527 17922 18536
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 18156 18358 18184 19858
rect 18524 19854 18552 20266
rect 18616 19854 18644 20975
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18340 19378 18368 19654
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18524 19174 18552 19790
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17328 17202 17356 18158
rect 17972 17882 18000 18226
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17958 17776 18014 17785
rect 17958 17711 18014 17720
rect 17972 17338 18000 17711
rect 18156 17610 18184 18294
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17420 16658 17448 17206
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17222 16552 17278 16561
rect 17222 16487 17278 16496
rect 17236 16454 17264 16487
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17420 16182 17448 16594
rect 17696 16590 17724 16934
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17236 15026 17264 16118
rect 17972 15978 18000 17138
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17958 15600 18014 15609
rect 17958 15535 18014 15544
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16592 14618 16620 14894
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 14006 15884 14214
rect 16040 14006 16068 14554
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15948 13394 15976 13806
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15948 11898 15976 13330
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16316 12986 16344 13194
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16500 12889 16528 13194
rect 16592 13190 16620 14554
rect 17236 14414 17264 14962
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17236 13938 17264 14350
rect 17328 14074 17356 14962
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17696 14006 17724 15302
rect 17972 15094 18000 15535
rect 18064 15434 18092 16050
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18052 15428 18104 15434
rect 18052 15370 18104 15376
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17972 14618 18000 15030
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17052 13530 17080 13874
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16486 12880 16542 12889
rect 16868 12850 16896 13398
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 16486 12815 16542 12824
rect 16856 12844 16908 12850
rect 16500 12442 16528 12815
rect 16856 12786 16908 12792
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16684 12170 16712 12582
rect 16868 12238 16896 12582
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 17052 11830 17080 12038
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 16040 11082 16068 11766
rect 17144 11762 17172 12174
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16132 11286 16160 11630
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 16040 10810 16068 11018
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16132 10742 16160 11222
rect 16316 11150 16344 11494
rect 16500 11354 16528 11698
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16592 11082 16620 11154
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 17144 10742 17172 11698
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 17132 10736 17184 10742
rect 17236 10713 17264 11154
rect 17328 11082 17356 13126
rect 18064 12986 18092 15370
rect 18248 14618 18276 15438
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 13394 18276 14214
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18156 12918 18184 13194
rect 18432 13190 18460 18566
rect 18524 18290 18552 19110
rect 18708 18329 18736 20402
rect 18892 20330 18920 20878
rect 18984 20398 19012 21898
rect 19628 21690 19656 22646
rect 21088 22636 21140 22642
rect 21140 22596 21220 22624
rect 21088 22578 21140 22584
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 19720 22098 19748 22510
rect 19708 22092 19760 22098
rect 19708 22034 19760 22040
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19223 21244 19531 21253
rect 19223 21242 19229 21244
rect 19285 21242 19309 21244
rect 19365 21242 19389 21244
rect 19445 21242 19469 21244
rect 19525 21242 19531 21244
rect 19285 21190 19287 21242
rect 19467 21190 19469 21242
rect 19223 21188 19229 21190
rect 19285 21188 19309 21190
rect 19365 21188 19389 21190
rect 19445 21188 19469 21190
rect 19525 21188 19531 21190
rect 19223 21179 19531 21188
rect 19616 21140 19668 21146
rect 19720 21128 19748 22034
rect 19800 22024 19852 22030
rect 19800 21966 19852 21972
rect 19812 21622 19840 21966
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 19883 21788 20191 21797
rect 19883 21786 19889 21788
rect 19945 21786 19969 21788
rect 20025 21786 20049 21788
rect 20105 21786 20129 21788
rect 20185 21786 20191 21788
rect 19945 21734 19947 21786
rect 20127 21734 20129 21786
rect 19883 21732 19889 21734
rect 19945 21732 19969 21734
rect 20025 21732 20049 21734
rect 20105 21732 20129 21734
rect 20185 21732 20191 21734
rect 19883 21723 20191 21732
rect 19800 21616 19852 21622
rect 19800 21558 19852 21564
rect 19812 21486 19840 21558
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 19668 21100 19748 21128
rect 19616 21082 19668 21088
rect 19812 20942 19840 21422
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 18984 19786 19012 20334
rect 19223 20156 19531 20165
rect 19223 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19469 20156
rect 19525 20154 19531 20156
rect 19285 20102 19287 20154
rect 19467 20102 19469 20154
rect 19223 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19469 20102
rect 19525 20100 19531 20102
rect 19223 20091 19531 20100
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18984 19334 19012 19722
rect 19628 19514 19656 20402
rect 19812 20398 19840 20878
rect 19883 20700 20191 20709
rect 19883 20698 19889 20700
rect 19945 20698 19969 20700
rect 20025 20698 20049 20700
rect 20105 20698 20129 20700
rect 20185 20698 20191 20700
rect 19945 20646 19947 20698
rect 20127 20646 20129 20698
rect 19883 20644 19889 20646
rect 19945 20644 19969 20646
rect 20025 20644 20049 20646
rect 20105 20644 20129 20646
rect 20185 20644 20191 20646
rect 19883 20635 20191 20644
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 18892 19306 19012 19334
rect 18892 18698 18920 19306
rect 19223 19068 19531 19077
rect 19223 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19469 19068
rect 19525 19066 19531 19068
rect 19285 19014 19287 19066
rect 19467 19014 19469 19066
rect 19223 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19469 19014
rect 19525 19012 19531 19014
rect 19223 19003 19531 19012
rect 19628 18970 19656 19450
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 18970 18864 19026 18873
rect 18970 18799 19026 18808
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18694 18320 18750 18329
rect 18512 18284 18564 18290
rect 18694 18255 18696 18264
rect 18512 18226 18564 18232
rect 18748 18255 18750 18264
rect 18696 18226 18748 18232
rect 18524 17678 18552 18226
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18616 17202 18644 17750
rect 18892 17746 18920 18634
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18892 16522 18920 17682
rect 18984 17678 19012 18799
rect 19720 18426 19748 19858
rect 19812 19854 19840 20334
rect 20364 20058 20392 21898
rect 20548 21434 20576 22510
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20640 21622 20668 22374
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20548 21406 20668 21434
rect 20640 20806 20668 21406
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19812 19378 19840 19790
rect 19883 19612 20191 19621
rect 19883 19610 19889 19612
rect 19945 19610 19969 19612
rect 20025 19610 20049 19612
rect 20105 19610 20129 19612
rect 20185 19610 20191 19612
rect 19945 19558 19947 19610
rect 20127 19558 20129 19610
rect 19883 19556 19889 19558
rect 19945 19556 19969 19558
rect 20025 19556 20049 19558
rect 20105 19556 20129 19558
rect 20185 19556 20191 19558
rect 19883 19547 20191 19556
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19812 18766 19840 19314
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18984 17338 19012 17614
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19076 17270 19104 18158
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19223 17980 19531 17989
rect 19223 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19469 17980
rect 19525 17978 19531 17980
rect 19285 17926 19287 17978
rect 19467 17926 19469 17978
rect 19223 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19469 17926
rect 19525 17924 19531 17926
rect 19223 17915 19531 17924
rect 19628 17678 19656 18022
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19720 17338 19748 18362
rect 19812 17746 19840 18702
rect 20548 18578 20576 20538
rect 20640 20534 20668 20742
rect 20628 20528 20680 20534
rect 20628 20470 20680 20476
rect 21008 20466 21036 22510
rect 21088 21888 21140 21894
rect 21086 21856 21088 21865
rect 21140 21856 21142 21865
rect 21086 21791 21142 21800
rect 21100 21049 21128 21791
rect 21192 21350 21220 22596
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21192 21185 21220 21286
rect 21178 21176 21234 21185
rect 21178 21111 21234 21120
rect 21086 21040 21142 21049
rect 21086 20975 21142 20984
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21178 20496 21234 20505
rect 20996 20460 21048 20466
rect 21178 20431 21180 20440
rect 20996 20402 21048 20408
rect 21232 20431 21234 20440
rect 21180 20402 21232 20408
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20626 19816 20682 19825
rect 20626 19751 20682 19760
rect 20640 18970 20668 19751
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20640 18698 20668 18906
rect 20824 18766 20852 20198
rect 20916 19854 20944 20198
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 21008 19174 21036 20402
rect 21192 20058 21220 20402
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21284 19786 21312 20878
rect 21376 20466 21404 22646
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21468 20466 21496 20742
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21284 19514 21312 19722
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21008 18970 21036 19110
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20548 18550 20668 18578
rect 19883 18524 20191 18533
rect 19883 18522 19889 18524
rect 19945 18522 19969 18524
rect 20025 18522 20049 18524
rect 20105 18522 20129 18524
rect 20185 18522 20191 18524
rect 19945 18470 19947 18522
rect 20127 18470 20129 18522
rect 19883 18468 19889 18470
rect 19945 18468 19969 18470
rect 20025 18468 20049 18470
rect 20105 18468 20129 18470
rect 20185 18468 20191 18470
rect 19883 18459 20191 18468
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 19076 17134 19104 17206
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 19076 16658 19104 17070
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19223 16892 19531 16901
rect 19223 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19469 16892
rect 19525 16890 19531 16892
rect 19285 16838 19287 16890
rect 19467 16838 19469 16890
rect 19223 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19469 16838
rect 19525 16836 19531 16838
rect 19223 16827 19531 16836
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 16182 18644 16390
rect 18604 16176 18656 16182
rect 18604 16118 18656 16124
rect 18892 16046 18920 16458
rect 19352 16114 19380 16526
rect 19628 16522 19656 16934
rect 19616 16516 19668 16522
rect 19616 16458 19668 16464
rect 19720 16402 19748 16934
rect 19536 16374 19748 16402
rect 19536 16114 19564 16374
rect 19812 16266 19840 17478
rect 19883 17436 20191 17445
rect 19883 17434 19889 17436
rect 19945 17434 19969 17436
rect 20025 17434 20049 17436
rect 20105 17434 20129 17436
rect 20185 17434 20191 17436
rect 19945 17382 19947 17434
rect 20127 17382 20129 17434
rect 19883 17380 19889 17382
rect 19945 17380 19969 17382
rect 20025 17380 20049 17382
rect 20105 17380 20129 17382
rect 20185 17380 20191 17382
rect 19883 17371 20191 17380
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20180 17082 20208 17274
rect 20272 17202 20300 17478
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20180 17054 20300 17082
rect 19883 16348 20191 16357
rect 19883 16346 19889 16348
rect 19945 16346 19969 16348
rect 20025 16346 20049 16348
rect 20105 16346 20129 16348
rect 20185 16346 20191 16348
rect 19945 16294 19947 16346
rect 20127 16294 20129 16346
rect 19883 16292 19889 16294
rect 19945 16292 19969 16294
rect 20025 16292 20049 16294
rect 20105 16292 20129 16294
rect 20185 16292 20191 16294
rect 19883 16283 20191 16292
rect 19628 16238 19840 16266
rect 20272 16266 20300 17054
rect 20364 16454 20392 18158
rect 20444 18148 20496 18154
rect 20444 18090 20496 18096
rect 20456 17202 20484 18090
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20548 16794 20576 17818
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20272 16238 20392 16266
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18892 15638 18920 15982
rect 19223 15804 19531 15813
rect 19223 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19469 15804
rect 19525 15802 19531 15804
rect 19285 15750 19287 15802
rect 19467 15750 19469 15802
rect 19223 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19469 15750
rect 19525 15748 19531 15750
rect 19223 15739 19531 15748
rect 19628 15722 19656 16238
rect 19800 16176 19852 16182
rect 19800 16118 19852 16124
rect 19628 15694 19748 15722
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 18616 14278 18644 14758
rect 19223 14716 19531 14725
rect 19223 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19469 14716
rect 19525 14714 19531 14716
rect 19285 14662 19287 14714
rect 19467 14662 19469 14714
rect 19223 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19469 14662
rect 19525 14660 19531 14662
rect 19223 14651 19531 14660
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19536 14521 19564 14554
rect 19522 14512 19578 14521
rect 19522 14447 19578 14456
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18708 14074 18736 14350
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18800 13977 18828 14010
rect 19352 14006 19380 14350
rect 19628 14346 19656 14758
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 19340 14000 19392 14006
rect 18786 13968 18842 13977
rect 19340 13942 19392 13948
rect 18786 13903 18842 13912
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18984 13530 19012 13874
rect 19223 13628 19531 13637
rect 19223 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19469 13628
rect 19525 13626 19531 13628
rect 19285 13574 19287 13626
rect 19467 13574 19469 13626
rect 19223 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19469 13574
rect 19525 13572 19531 13574
rect 19223 13563 19531 13572
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18248 12714 18276 13126
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18248 12434 18276 12650
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18432 12442 18460 12582
rect 17972 12406 18276 12434
rect 18420 12436 18472 12442
rect 17592 11280 17644 11286
rect 17592 11222 17644 11228
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17132 10678 17184 10684
rect 17222 10704 17278 10713
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15764 9654 15792 10202
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15120 8566 15148 8910
rect 15488 8838 15516 9454
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14662 7644 14970 7653
rect 14662 7642 14668 7644
rect 14724 7642 14748 7644
rect 14804 7642 14828 7644
rect 14884 7642 14908 7644
rect 14964 7642 14970 7644
rect 14724 7590 14726 7642
rect 14906 7590 14908 7642
rect 14662 7588 14668 7590
rect 14724 7588 14748 7590
rect 14804 7588 14828 7590
rect 14884 7588 14908 7590
rect 14964 7588 14970 7590
rect 14662 7579 14970 7588
rect 15120 7478 15148 8366
rect 15672 7546 15700 9522
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15856 8566 15884 9454
rect 16132 9058 16160 10678
rect 17144 10130 17172 10678
rect 17222 10639 17278 10648
rect 17328 10266 17356 11018
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16040 9030 16160 9058
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15764 7886 15792 8366
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 16040 7818 16068 9030
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 15856 7546 15884 7754
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14844 6798 14872 7142
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14568 6254 14596 6734
rect 14662 6556 14970 6565
rect 14662 6554 14668 6556
rect 14724 6554 14748 6556
rect 14804 6554 14828 6556
rect 14884 6554 14908 6556
rect 14964 6554 14970 6556
rect 14724 6502 14726 6554
rect 14906 6502 14908 6554
rect 14662 6500 14668 6502
rect 14724 6500 14748 6502
rect 14804 6500 14828 6502
rect 14884 6500 14908 6502
rect 14964 6500 14970 6502
rect 14662 6491 14970 6500
rect 15120 6254 15148 7414
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 14662 5468 14970 5477
rect 14662 5466 14668 5468
rect 14724 5466 14748 5468
rect 14804 5466 14828 5468
rect 14884 5466 14908 5468
rect 14964 5466 14970 5468
rect 14724 5414 14726 5466
rect 14906 5414 14908 5466
rect 14662 5412 14668 5414
rect 14724 5412 14748 5414
rect 14804 5412 14828 5414
rect 14884 5412 14908 5414
rect 14964 5412 14970 5414
rect 14662 5403 14970 5412
rect 14662 4380 14970 4389
rect 14662 4378 14668 4380
rect 14724 4378 14748 4380
rect 14804 4378 14828 4380
rect 14884 4378 14908 4380
rect 14964 4378 14970 4380
rect 14724 4326 14726 4378
rect 14906 4326 14908 4378
rect 14662 4324 14668 4326
rect 14724 4324 14748 4326
rect 14804 4324 14828 4326
rect 14884 4324 14908 4326
rect 14964 4324 14970 4326
rect 14662 4315 14970 4324
rect 15120 4298 15148 5850
rect 15120 4270 15240 4298
rect 15304 4282 15332 6190
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15396 5302 15424 6054
rect 15488 5914 15516 6326
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15580 5914 15608 6258
rect 16040 6254 16068 7754
rect 16132 7546 16160 8842
rect 16224 7818 16252 9930
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16224 6798 16252 7754
rect 16316 7410 16344 9318
rect 17052 9178 17080 9590
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 16500 5778 16528 7958
rect 16776 7954 16804 8230
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16868 7546 16896 8842
rect 17052 8634 17080 9114
rect 17144 9042 17172 10066
rect 17328 9518 17356 10202
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17420 9722 17448 9930
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17604 9586 17632 11222
rect 17972 11082 18000 12406
rect 18420 12378 18472 12384
rect 18524 11898 18552 12854
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18616 12374 18644 12786
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18984 12374 19012 12718
rect 19223 12540 19531 12549
rect 19223 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19469 12540
rect 19525 12538 19531 12540
rect 19285 12486 19287 12538
rect 19467 12486 19469 12538
rect 19223 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19469 12486
rect 19525 12484 19531 12486
rect 19223 12475 19531 12484
rect 18604 12368 18656 12374
rect 18602 12336 18604 12345
rect 18972 12368 19024 12374
rect 18656 12336 18658 12345
rect 18972 12310 19024 12316
rect 19720 12306 19748 15694
rect 19812 14958 19840 16118
rect 20260 15632 20312 15638
rect 20260 15574 20312 15580
rect 19883 15260 20191 15269
rect 19883 15258 19889 15260
rect 19945 15258 19969 15260
rect 20025 15258 20049 15260
rect 20105 15258 20129 15260
rect 20185 15258 20191 15260
rect 19945 15206 19947 15258
rect 20127 15206 20129 15258
rect 19883 15204 19889 15206
rect 19945 15204 19969 15206
rect 20025 15204 20049 15206
rect 20105 15204 20129 15206
rect 20185 15204 20191 15206
rect 19883 15195 20191 15204
rect 20272 15026 20300 15574
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19812 14414 19840 14894
rect 19892 14884 19944 14890
rect 19892 14826 19944 14832
rect 19904 14618 19932 14826
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19812 13394 19840 14350
rect 19883 14172 20191 14181
rect 19883 14170 19889 14172
rect 19945 14170 19969 14172
rect 20025 14170 20049 14172
rect 20105 14170 20129 14172
rect 20185 14170 20191 14172
rect 19945 14118 19947 14170
rect 20127 14118 20129 14170
rect 19883 14116 19889 14118
rect 19945 14116 19969 14118
rect 20025 14116 20049 14118
rect 20105 14116 20129 14118
rect 20185 14116 20191 14118
rect 19883 14107 20191 14116
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 19892 13796 19944 13802
rect 19892 13738 19944 13744
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19904 13326 19932 13738
rect 20272 13326 20300 14010
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 19883 13084 20191 13093
rect 19883 13082 19889 13084
rect 19945 13082 19969 13084
rect 20025 13082 20049 13084
rect 20105 13082 20129 13084
rect 20185 13082 20191 13084
rect 19945 13030 19947 13082
rect 20127 13030 20129 13082
rect 19883 13028 19889 13030
rect 19945 13028 19969 13030
rect 20025 13028 20049 13030
rect 20105 13028 20129 13030
rect 20185 13028 20191 13030
rect 19883 13019 20191 13028
rect 20364 12986 20392 16238
rect 20640 14006 20668 18550
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 21008 17678 21036 18158
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20718 15056 20774 15065
rect 20718 14991 20774 15000
rect 20732 14278 20760 14991
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20824 14006 20852 14214
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20548 13258 20576 13806
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20548 12850 20576 13194
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 18602 12271 18658 12280
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 19260 11762 19288 12038
rect 19883 11996 20191 12005
rect 19883 11994 19889 11996
rect 19945 11994 19969 11996
rect 20025 11994 20049 11996
rect 20105 11994 20129 11996
rect 20185 11994 20191 11996
rect 19945 11942 19947 11994
rect 20127 11942 20129 11994
rect 19883 11940 19889 11942
rect 19945 11940 19969 11942
rect 20025 11940 20049 11942
rect 20105 11940 20129 11942
rect 20185 11940 20191 11942
rect 19883 11931 20191 11940
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19076 11218 19104 11630
rect 19223 11452 19531 11461
rect 19223 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19469 11452
rect 19525 11450 19531 11452
rect 19285 11398 19287 11450
rect 19467 11398 19469 11450
rect 19223 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19469 11398
rect 19525 11396 19531 11398
rect 19223 11387 19531 11396
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17972 10554 18000 11018
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 17880 10526 18000 10554
rect 17880 10044 17908 10526
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 10146 18000 10406
rect 18156 10266 18184 10950
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18050 10160 18106 10169
rect 17972 10118 18050 10146
rect 18050 10095 18106 10104
rect 17880 10016 18000 10044
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17972 8786 18000 10016
rect 18064 9518 18092 10095
rect 18156 9722 18184 10202
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17972 8758 18092 8786
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 16960 8090 16988 8502
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16960 6662 16988 8026
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 17052 7449 17080 7482
rect 17038 7440 17094 7449
rect 17038 7375 17094 7384
rect 17052 6866 17080 7375
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17144 6746 17172 8366
rect 17236 7886 17264 8502
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17328 8022 17356 8366
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17604 7410 17632 8230
rect 17972 7546 18000 8434
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17052 6730 17172 6746
rect 17040 6724 17172 6730
rect 17092 6718 17172 6724
rect 17040 6666 17092 6672
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 16132 5030 16160 5578
rect 16500 5370 16528 5714
rect 17052 5692 17080 6666
rect 17960 6384 18012 6390
rect 18064 6361 18092 8758
rect 18156 8537 18184 9522
rect 18892 9450 18920 10610
rect 19076 10606 19104 11154
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19076 10062 19104 10542
rect 19223 10364 19531 10373
rect 19223 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19469 10364
rect 19525 10362 19531 10364
rect 19285 10310 19287 10362
rect 19467 10310 19469 10362
rect 19223 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19469 10310
rect 19525 10308 19531 10310
rect 19223 10299 19531 10308
rect 19064 10056 19116 10062
rect 19812 10044 19840 10950
rect 19883 10908 20191 10917
rect 19883 10906 19889 10908
rect 19945 10906 19969 10908
rect 20025 10906 20049 10908
rect 20105 10906 20129 10908
rect 20185 10906 20191 10908
rect 19945 10854 19947 10906
rect 20127 10854 20129 10906
rect 19883 10852 19889 10854
rect 19945 10852 19969 10854
rect 20025 10852 20049 10854
rect 20105 10852 20129 10854
rect 20185 10852 20191 10854
rect 19883 10843 20191 10852
rect 19892 10056 19944 10062
rect 19812 10016 19892 10044
rect 19064 9998 19116 10004
rect 19892 9998 19944 10004
rect 19076 9654 19104 9998
rect 20260 9988 20312 9994
rect 20260 9930 20312 9936
rect 19883 9820 20191 9829
rect 19883 9818 19889 9820
rect 19945 9818 19969 9820
rect 20025 9818 20049 9820
rect 20105 9818 20129 9820
rect 20185 9818 20191 9820
rect 19945 9766 19947 9818
rect 20127 9766 20129 9818
rect 19883 9764 19889 9766
rect 19945 9764 19969 9766
rect 20025 9764 20049 9766
rect 20105 9764 20129 9766
rect 20185 9764 20191 9766
rect 19883 9755 20191 9764
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 18880 9444 18932 9450
rect 18880 9386 18932 9392
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19223 9276 19531 9285
rect 19223 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19469 9276
rect 19525 9274 19531 9276
rect 19285 9222 19287 9274
rect 19467 9222 19469 9274
rect 19223 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19469 9222
rect 19525 9220 19531 9222
rect 19223 9211 19531 9220
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18142 8528 18198 8537
rect 18248 8498 18276 9114
rect 19904 8974 19932 9386
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 18340 8498 18368 8910
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18142 8463 18198 8472
rect 18236 8492 18288 8498
rect 18156 6798 18184 8463
rect 18236 8434 18288 8440
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18248 7886 18276 8298
rect 18340 7954 18368 8434
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 17960 6326 18012 6332
rect 18050 6352 18106 6361
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17144 5846 17172 6190
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17052 5664 17172 5692
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14568 2650 14596 4082
rect 14752 3738 14780 4150
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14662 3292 14970 3301
rect 14662 3290 14668 3292
rect 14724 3290 14748 3292
rect 14804 3290 14828 3292
rect 14884 3290 14908 3292
rect 14964 3290 14970 3292
rect 14724 3238 14726 3290
rect 14906 3238 14908 3290
rect 14662 3236 14668 3238
rect 14724 3236 14748 3238
rect 14804 3236 14828 3238
rect 14884 3236 14908 3238
rect 14964 3236 14970 3238
rect 14662 3227 14970 3236
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 15028 2378 15056 3674
rect 15120 3602 15148 4082
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15212 3482 15240 4270
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15120 3454 15240 3482
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 14662 2204 14970 2213
rect 14662 2202 14668 2204
rect 14724 2202 14748 2204
rect 14804 2202 14828 2204
rect 14884 2202 14908 2204
rect 14964 2202 14970 2204
rect 14724 2150 14726 2202
rect 14906 2150 14908 2202
rect 14662 2148 14668 2150
rect 14724 2148 14748 2150
rect 14804 2148 14828 2150
rect 14884 2148 14908 2150
rect 14964 2148 14970 2150
rect 14662 2139 14970 2148
rect 14844 870 14964 898
rect 14844 800 14872 870
rect 14292 734 14504 762
rect 14830 0 14886 800
rect 14936 762 14964 870
rect 15120 762 15148 3454
rect 15304 2650 15332 4082
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15580 3194 15608 3402
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15488 2514 15516 2790
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15488 800 15516 2450
rect 16132 800 16160 4966
rect 16500 4842 16528 5306
rect 16500 4814 16712 4842
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16316 3058 16344 4082
rect 16592 4010 16620 4694
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16684 3466 16712 4814
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16776 2446 16804 3606
rect 16868 3602 16896 3878
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16960 3058 16988 3878
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17052 3194 17080 3334
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17144 3074 17172 5664
rect 17328 5642 17356 6054
rect 17972 5710 18000 6326
rect 18050 6287 18106 6296
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 17972 5302 18000 5646
rect 18064 5302 18092 6287
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17972 4162 18000 4422
rect 18064 4282 18092 4966
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18236 4208 18288 4214
rect 17972 4146 18092 4162
rect 18432 4185 18460 8774
rect 18892 8498 18920 8774
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 19223 8188 19531 8197
rect 19223 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19469 8188
rect 19525 8186 19531 8188
rect 19285 8134 19287 8186
rect 19467 8134 19469 8186
rect 19223 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19469 8134
rect 19525 8132 19531 8134
rect 19223 8123 19531 8132
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18708 7478 18736 7686
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18616 6458 18644 7142
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18708 5778 18736 6054
rect 18800 5846 18828 7414
rect 18892 7002 18920 7822
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18788 5840 18840 5846
rect 18788 5782 18840 5788
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18800 5642 18828 5782
rect 18788 5636 18840 5642
rect 18788 5578 18840 5584
rect 18984 5302 19012 7482
rect 19628 7342 19656 8570
rect 19720 8294 19748 8842
rect 19883 8732 20191 8741
rect 19883 8730 19889 8732
rect 19945 8730 19969 8732
rect 20025 8730 20049 8732
rect 20105 8730 20129 8732
rect 20185 8730 20191 8732
rect 19945 8678 19947 8730
rect 20127 8678 20129 8730
rect 19883 8676 19889 8678
rect 19945 8676 19969 8678
rect 20025 8676 20049 8678
rect 20105 8676 20129 8678
rect 20185 8676 20191 8678
rect 19883 8667 20191 8676
rect 20272 8566 20300 9930
rect 20364 9450 20392 12786
rect 20732 12714 20760 13874
rect 20824 13734 20852 13942
rect 20916 13870 20944 16390
rect 21008 16250 21036 17614
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 21100 15978 21128 17546
rect 21192 16114 21220 18702
rect 21376 18698 21404 20402
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21468 19378 21496 19654
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 21284 17338 21312 18294
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21284 17105 21312 17274
rect 21270 17096 21326 17105
rect 21270 17031 21326 17040
rect 21180 16108 21232 16114
rect 21376 16096 21404 18634
rect 21546 18456 21602 18465
rect 21546 18391 21602 18400
rect 21560 17882 21588 18391
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21456 17264 21508 17270
rect 21456 17206 21508 17212
rect 21468 16794 21496 17206
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21560 16182 21588 17818
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21652 16114 21680 18022
rect 21456 16108 21508 16114
rect 21376 16068 21456 16096
rect 21180 16050 21232 16056
rect 21456 16050 21508 16056
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20916 12434 20944 13806
rect 21192 13530 21220 15302
rect 21468 14521 21496 15370
rect 21560 14822 21588 15506
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21454 14512 21510 14521
rect 21364 14476 21416 14482
rect 21454 14447 21456 14456
rect 21364 14418 21416 14424
rect 21508 14447 21510 14456
rect 21456 14418 21508 14424
rect 21376 14385 21404 14418
rect 21362 14376 21418 14385
rect 21362 14311 21418 14320
rect 21560 13705 21588 14758
rect 21546 13696 21602 13705
rect 21546 13631 21602 13640
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21192 12918 21220 13466
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 20916 12406 21036 12434
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20456 9654 20484 12242
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20548 9654 20576 12174
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11898 20760 12038
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20824 11370 20852 12106
rect 20732 11354 20852 11370
rect 20720 11348 20852 11354
rect 20772 11342 20852 11348
rect 20720 11290 20772 11296
rect 20824 10606 20852 11342
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19720 7546 19748 8230
rect 19800 7812 19852 7818
rect 19800 7754 19852 7760
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19076 6730 19104 7210
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19223 7100 19531 7109
rect 19223 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19469 7100
rect 19525 7098 19531 7100
rect 19285 7046 19287 7098
rect 19467 7046 19469 7098
rect 19223 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19469 7046
rect 19525 7044 19531 7046
rect 19223 7035 19531 7044
rect 19064 6724 19116 6730
rect 19064 6666 19116 6672
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 19076 6390 19104 6666
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19076 6254 19104 6326
rect 19168 6322 19196 6598
rect 19444 6458 19472 6666
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19628 6322 19656 7142
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19064 6248 19116 6254
rect 19720 6202 19748 7210
rect 19064 6190 19116 6196
rect 18972 5296 19024 5302
rect 18972 5238 19024 5244
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18236 4150 18288 4156
rect 18418 4176 18474 4185
rect 17972 4140 18104 4146
rect 17972 4134 18052 4140
rect 18052 4082 18104 4088
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 17052 3046 17172 3074
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16776 870 16896 898
rect 16776 800 16804 870
rect 14936 734 15148 762
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 16868 762 16896 870
rect 17052 762 17080 3046
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 17144 2378 17172 2790
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17420 800 17448 3538
rect 18064 800 18092 4082
rect 18248 3398 18276 4150
rect 18418 4111 18474 4120
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18248 3194 18276 3334
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18524 2310 18552 4014
rect 18708 3466 18736 4558
rect 18984 4282 19012 5238
rect 19076 5166 19104 6190
rect 19628 6186 19748 6202
rect 19616 6180 19748 6186
rect 19668 6174 19748 6180
rect 19616 6122 19668 6128
rect 19708 6112 19760 6118
rect 19812 6100 19840 7754
rect 19883 7644 20191 7653
rect 19883 7642 19889 7644
rect 19945 7642 19969 7644
rect 20025 7642 20049 7644
rect 20105 7642 20129 7644
rect 20185 7642 20191 7644
rect 19945 7590 19947 7642
rect 20127 7590 20129 7642
rect 19883 7588 19889 7590
rect 19945 7588 19969 7590
rect 20025 7588 20049 7590
rect 20105 7588 20129 7590
rect 20185 7588 20191 7590
rect 19883 7579 20191 7588
rect 19883 6556 20191 6565
rect 19883 6554 19889 6556
rect 19945 6554 19969 6556
rect 20025 6554 20049 6556
rect 20105 6554 20129 6556
rect 20185 6554 20191 6556
rect 19945 6502 19947 6554
rect 20127 6502 20129 6554
rect 19883 6500 19889 6502
rect 19945 6500 19969 6502
rect 20025 6500 20049 6502
rect 20105 6500 20129 6502
rect 20185 6500 20191 6502
rect 19883 6491 20191 6500
rect 19760 6072 19840 6100
rect 19708 6054 19760 6060
rect 19223 6012 19531 6021
rect 19223 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19469 6012
rect 19525 6010 19531 6012
rect 19285 5958 19287 6010
rect 19467 5958 19469 6010
rect 19223 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19469 5958
rect 19525 5956 19531 5958
rect 19223 5947 19531 5956
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19536 5234 19564 5782
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20364 5545 20392 5714
rect 20456 5710 20484 9590
rect 20548 9382 20576 9590
rect 20640 9450 20668 9998
rect 20916 9450 20944 11018
rect 21008 10606 21036 12406
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21284 11762 21312 12310
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21376 11665 21404 12106
rect 21362 11656 21418 11665
rect 21362 11591 21418 11600
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21100 11150 21128 11494
rect 21376 11354 21404 11591
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20824 8945 20852 9114
rect 21008 9058 21036 10542
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21284 9602 21312 9862
rect 21376 9722 21404 10678
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21362 9616 21418 9625
rect 21180 9580 21232 9586
rect 21284 9574 21362 9602
rect 21362 9551 21418 9560
rect 21180 9522 21232 9528
rect 20916 9030 21036 9058
rect 20810 8936 20866 8945
rect 20810 8871 20866 8880
rect 20916 8838 20944 9030
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20548 7478 20576 8774
rect 20626 8256 20682 8265
rect 20626 8191 20682 8200
rect 20640 8090 20668 8191
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20640 7478 20668 8026
rect 21008 7546 21036 8842
rect 21192 8634 21220 9522
rect 21376 9518 21404 9551
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21192 8106 21220 8570
rect 21192 8078 21312 8106
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20812 7472 20864 7478
rect 21100 7426 21128 7822
rect 20812 7414 20864 7420
rect 20732 7002 20760 7414
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20732 6662 20760 6938
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20824 5778 20852 7414
rect 21008 7398 21128 7426
rect 21192 7410 21220 7958
rect 21284 7818 21312 8078
rect 21376 7954 21404 8774
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21180 7404 21232 7410
rect 21008 7342 21036 7398
rect 21180 7346 21232 7352
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 21008 6866 21036 7278
rect 21376 6905 21404 7890
rect 21362 6896 21418 6905
rect 20996 6860 21048 6866
rect 21362 6831 21418 6840
rect 20996 6802 21048 6808
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 21008 5642 21036 6802
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 21100 6225 21128 6666
rect 21086 6216 21142 6225
rect 21086 6151 21088 6160
rect 21140 6151 21142 6160
rect 21088 6122 21140 6128
rect 21548 5840 21600 5846
rect 21548 5782 21600 5788
rect 20996 5636 21048 5642
rect 20996 5578 21048 5584
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 20350 5536 20406 5545
rect 19883 5468 20191 5477
rect 20350 5471 20406 5480
rect 19883 5466 19889 5468
rect 19945 5466 19969 5468
rect 20025 5466 20049 5468
rect 20105 5466 20129 5468
rect 20185 5466 20191 5468
rect 19945 5414 19947 5466
rect 20127 5414 20129 5466
rect 19883 5412 19889 5414
rect 19945 5412 19969 5414
rect 20025 5412 20049 5414
rect 20105 5412 20129 5414
rect 20185 5412 20191 5414
rect 19883 5403 20191 5412
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 4622 19104 5102
rect 19223 4924 19531 4933
rect 19223 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19469 4924
rect 19525 4922 19531 4924
rect 19285 4870 19287 4922
rect 19467 4870 19469 4922
rect 19223 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19469 4870
rect 19525 4868 19531 4870
rect 19223 4859 19531 4868
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19883 4380 20191 4389
rect 19883 4378 19889 4380
rect 19945 4378 19969 4380
rect 20025 4378 20049 4380
rect 20105 4378 20129 4380
rect 20185 4378 20191 4380
rect 19945 4326 19947 4378
rect 20127 4326 20129 4378
rect 19883 4324 19889 4326
rect 19945 4324 19969 4326
rect 20025 4324 20049 4326
rect 20105 4324 20129 4326
rect 20185 4324 20191 4326
rect 19883 4315 20191 4324
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 18984 3738 19012 4218
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 19892 4072 19944 4078
rect 19812 4032 19892 4060
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 18708 2990 18736 3402
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 3126 18920 3334
rect 19076 3126 19104 3878
rect 19223 3836 19531 3845
rect 19223 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19469 3836
rect 19525 3834 19531 3836
rect 19285 3782 19287 3834
rect 19467 3782 19469 3834
rect 19223 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19469 3782
rect 19525 3780 19531 3782
rect 19223 3771 19531 3780
rect 19720 3466 19748 3946
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19812 3194 19840 4032
rect 19892 4014 19944 4020
rect 20640 3738 20668 4150
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20916 3738 20944 3946
rect 21008 3942 21036 5578
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21192 5370 21220 5510
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21376 4622 21404 4966
rect 21468 4842 21496 5578
rect 21560 5234 21588 5782
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21546 4856 21602 4865
rect 21468 4814 21546 4842
rect 21546 4791 21548 4800
rect 21600 4791 21602 4800
rect 21548 4762 21600 4768
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 20640 3398 20668 3674
rect 21008 3534 21036 3878
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 20996 3528 21048 3534
rect 21376 3505 21404 3538
rect 20996 3470 21048 3476
rect 21362 3496 21418 3505
rect 21362 3431 21418 3440
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 19883 3292 20191 3301
rect 19883 3290 19889 3292
rect 19945 3290 19969 3292
rect 20025 3290 20049 3292
rect 20105 3290 20129 3292
rect 20185 3290 20191 3292
rect 19945 3238 19947 3290
rect 20127 3238 20129 3290
rect 19883 3236 19889 3238
rect 19945 3236 19969 3238
rect 20025 3236 20049 3238
rect 20105 3236 20129 3238
rect 20185 3236 20191 3238
rect 19883 3227 20191 3236
rect 21376 3194 21404 3431
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18708 2446 18736 2926
rect 19223 2748 19531 2757
rect 19223 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19469 2748
rect 19525 2746 19531 2748
rect 19285 2694 19287 2746
rect 19467 2694 19469 2746
rect 19223 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19469 2694
rect 19525 2692 19531 2694
rect 19223 2683 19531 2692
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18708 800 18736 2246
rect 19883 2204 20191 2213
rect 19883 2202 19889 2204
rect 19945 2202 19969 2204
rect 20025 2202 20049 2204
rect 20105 2202 20129 2204
rect 20185 2202 20191 2204
rect 19945 2150 19947 2202
rect 20127 2150 20129 2202
rect 19883 2148 19889 2150
rect 19945 2148 19969 2150
rect 20025 2148 20049 2150
rect 20105 2148 20129 2150
rect 20185 2148 20191 2150
rect 19883 2139 20191 2148
rect 16868 734 17080 762
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
<< via2 >>
rect 4226 22874 4282 22876
rect 4306 22874 4362 22876
rect 4386 22874 4442 22876
rect 4466 22874 4522 22876
rect 4226 22822 4272 22874
rect 4272 22822 4282 22874
rect 4306 22822 4336 22874
rect 4336 22822 4348 22874
rect 4348 22822 4362 22874
rect 4386 22822 4400 22874
rect 4400 22822 4412 22874
rect 4412 22822 4442 22874
rect 4466 22822 4476 22874
rect 4476 22822 4522 22874
rect 4226 22820 4282 22822
rect 4306 22820 4362 22822
rect 4386 22820 4442 22822
rect 4466 22820 4522 22822
rect 1306 19080 1362 19136
rect 3566 22330 3622 22332
rect 3646 22330 3702 22332
rect 3726 22330 3782 22332
rect 3806 22330 3862 22332
rect 3566 22278 3612 22330
rect 3612 22278 3622 22330
rect 3646 22278 3676 22330
rect 3676 22278 3688 22330
rect 3688 22278 3702 22330
rect 3726 22278 3740 22330
rect 3740 22278 3752 22330
rect 3752 22278 3782 22330
rect 3806 22278 3816 22330
rect 3816 22278 3862 22330
rect 3566 22276 3622 22278
rect 3646 22276 3702 22278
rect 3726 22276 3782 22278
rect 3806 22276 3862 22278
rect 3054 21800 3110 21856
rect 4226 21786 4282 21788
rect 4306 21786 4362 21788
rect 4386 21786 4442 21788
rect 4466 21786 4522 21788
rect 4226 21734 4272 21786
rect 4272 21734 4282 21786
rect 4306 21734 4336 21786
rect 4336 21734 4348 21786
rect 4348 21734 4362 21786
rect 4386 21734 4400 21786
rect 4400 21734 4412 21786
rect 4412 21734 4442 21786
rect 4466 21734 4476 21786
rect 4476 21734 4522 21786
rect 4226 21732 4282 21734
rect 4306 21732 4362 21734
rect 4386 21732 4442 21734
rect 4466 21732 4522 21734
rect 3566 21242 3622 21244
rect 3646 21242 3702 21244
rect 3726 21242 3782 21244
rect 3806 21242 3862 21244
rect 3566 21190 3612 21242
rect 3612 21190 3622 21242
rect 3646 21190 3676 21242
rect 3676 21190 3688 21242
rect 3688 21190 3702 21242
rect 3726 21190 3740 21242
rect 3740 21190 3752 21242
rect 3752 21190 3782 21242
rect 3806 21190 3816 21242
rect 3816 21190 3862 21242
rect 3566 21188 3622 21190
rect 3646 21188 3702 21190
rect 3726 21188 3782 21190
rect 3806 21188 3862 21190
rect 4226 20698 4282 20700
rect 4306 20698 4362 20700
rect 4386 20698 4442 20700
rect 4466 20698 4522 20700
rect 4226 20646 4272 20698
rect 4272 20646 4282 20698
rect 4306 20646 4336 20698
rect 4336 20646 4348 20698
rect 4348 20646 4362 20698
rect 4386 20646 4400 20698
rect 4400 20646 4412 20698
rect 4412 20646 4442 20698
rect 4466 20646 4476 20698
rect 4476 20646 4522 20698
rect 4226 20644 4282 20646
rect 4306 20644 4362 20646
rect 4386 20644 4442 20646
rect 4466 20644 4522 20646
rect 2686 20440 2742 20496
rect 3566 20154 3622 20156
rect 3646 20154 3702 20156
rect 3726 20154 3782 20156
rect 3806 20154 3862 20156
rect 3566 20102 3612 20154
rect 3612 20102 3622 20154
rect 3646 20102 3676 20154
rect 3676 20102 3688 20154
rect 3688 20102 3702 20154
rect 3726 20102 3740 20154
rect 3740 20102 3752 20154
rect 3752 20102 3782 20154
rect 3806 20102 3816 20154
rect 3816 20102 3862 20154
rect 3566 20100 3622 20102
rect 3646 20100 3702 20102
rect 3726 20100 3782 20102
rect 3806 20100 3862 20102
rect 2778 17720 2834 17776
rect 3566 19066 3622 19068
rect 3646 19066 3702 19068
rect 3726 19066 3782 19068
rect 3806 19066 3862 19068
rect 3566 19014 3612 19066
rect 3612 19014 3622 19066
rect 3646 19014 3676 19066
rect 3676 19014 3688 19066
rect 3688 19014 3702 19066
rect 3726 19014 3740 19066
rect 3740 19014 3752 19066
rect 3752 19014 3782 19066
rect 3806 19014 3816 19066
rect 3816 19014 3862 19066
rect 3566 19012 3622 19014
rect 3646 19012 3702 19014
rect 3726 19012 3782 19014
rect 3806 19012 3862 19014
rect 3566 17978 3622 17980
rect 3646 17978 3702 17980
rect 3726 17978 3782 17980
rect 3806 17978 3862 17980
rect 3566 17926 3612 17978
rect 3612 17926 3622 17978
rect 3646 17926 3676 17978
rect 3676 17926 3688 17978
rect 3688 17926 3702 17978
rect 3726 17926 3740 17978
rect 3740 17926 3752 17978
rect 3752 17926 3782 17978
rect 3806 17926 3816 17978
rect 3816 17926 3862 17978
rect 3566 17924 3622 17926
rect 3646 17924 3702 17926
rect 3726 17924 3782 17926
rect 3806 17924 3862 17926
rect 3054 17212 3056 17232
rect 3056 17212 3108 17232
rect 3108 17212 3110 17232
rect 3054 17176 3110 17212
rect 4226 19610 4282 19612
rect 4306 19610 4362 19612
rect 4386 19610 4442 19612
rect 4466 19610 4522 19612
rect 4226 19558 4272 19610
rect 4272 19558 4282 19610
rect 4306 19558 4336 19610
rect 4336 19558 4348 19610
rect 4348 19558 4362 19610
rect 4386 19558 4400 19610
rect 4400 19558 4412 19610
rect 4412 19558 4442 19610
rect 4466 19558 4476 19610
rect 4476 19558 4522 19610
rect 4226 19556 4282 19558
rect 4306 19556 4362 19558
rect 4386 19556 4442 19558
rect 4466 19556 4522 19558
rect 4802 19760 4858 19816
rect 4226 18522 4282 18524
rect 4306 18522 4362 18524
rect 4386 18522 4442 18524
rect 4466 18522 4522 18524
rect 4226 18470 4272 18522
rect 4272 18470 4282 18522
rect 4306 18470 4336 18522
rect 4336 18470 4348 18522
rect 4348 18470 4362 18522
rect 4386 18470 4400 18522
rect 4400 18470 4412 18522
rect 4412 18470 4442 18522
rect 4466 18470 4476 18522
rect 4476 18470 4522 18522
rect 4226 18468 4282 18470
rect 4306 18468 4362 18470
rect 4386 18468 4442 18470
rect 4466 18468 4522 18470
rect 4342 18264 4398 18320
rect 4226 17434 4282 17436
rect 4306 17434 4362 17436
rect 4386 17434 4442 17436
rect 4466 17434 4522 17436
rect 4226 17382 4272 17434
rect 4272 17382 4282 17434
rect 4306 17382 4336 17434
rect 4336 17382 4348 17434
rect 4348 17382 4362 17434
rect 4386 17382 4400 17434
rect 4400 17382 4412 17434
rect 4412 17382 4442 17434
rect 4466 17382 4476 17434
rect 4476 17382 4522 17434
rect 4226 17380 4282 17382
rect 4306 17380 4362 17382
rect 4386 17380 4442 17382
rect 4466 17380 4522 17382
rect 3566 16890 3622 16892
rect 3646 16890 3702 16892
rect 3726 16890 3782 16892
rect 3806 16890 3862 16892
rect 3566 16838 3612 16890
rect 3612 16838 3622 16890
rect 3646 16838 3676 16890
rect 3676 16838 3688 16890
rect 3688 16838 3702 16890
rect 3726 16838 3740 16890
rect 3740 16838 3752 16890
rect 3752 16838 3782 16890
rect 3806 16838 3816 16890
rect 3816 16838 3862 16890
rect 3566 16836 3622 16838
rect 3646 16836 3702 16838
rect 3726 16836 3782 16838
rect 3806 16836 3862 16838
rect 3566 15802 3622 15804
rect 3646 15802 3702 15804
rect 3726 15802 3782 15804
rect 3806 15802 3862 15804
rect 3566 15750 3612 15802
rect 3612 15750 3622 15802
rect 3646 15750 3676 15802
rect 3676 15750 3688 15802
rect 3688 15750 3702 15802
rect 3726 15750 3740 15802
rect 3740 15750 3752 15802
rect 3752 15750 3782 15802
rect 3806 15750 3816 15802
rect 3816 15750 3862 15802
rect 3566 15748 3622 15750
rect 3646 15748 3702 15750
rect 3726 15748 3782 15750
rect 3806 15748 3862 15750
rect 3146 15680 3202 15736
rect 4226 16346 4282 16348
rect 4306 16346 4362 16348
rect 4386 16346 4442 16348
rect 4466 16346 4522 16348
rect 4226 16294 4272 16346
rect 4272 16294 4282 16346
rect 4306 16294 4336 16346
rect 4336 16294 4348 16346
rect 4348 16294 4362 16346
rect 4386 16294 4400 16346
rect 4400 16294 4412 16346
rect 4412 16294 4442 16346
rect 4466 16294 4476 16346
rect 4476 16294 4522 16346
rect 4226 16292 4282 16294
rect 4306 16292 4362 16294
rect 4386 16292 4442 16294
rect 4466 16292 4522 16294
rect 2870 12960 2926 13016
rect 2778 12280 2834 12336
rect 1306 10240 1362 10296
rect 4226 15258 4282 15260
rect 4306 15258 4362 15260
rect 4386 15258 4442 15260
rect 4466 15258 4522 15260
rect 4226 15206 4272 15258
rect 4272 15206 4282 15258
rect 4306 15206 4336 15258
rect 4336 15206 4348 15258
rect 4348 15206 4362 15258
rect 4386 15206 4400 15258
rect 4400 15206 4412 15258
rect 4412 15206 4442 15258
rect 4466 15206 4476 15258
rect 4476 15206 4522 15258
rect 4226 15204 4282 15206
rect 4306 15204 4362 15206
rect 4386 15204 4442 15206
rect 4466 15204 4522 15206
rect 4894 16496 4950 16552
rect 3566 14714 3622 14716
rect 3646 14714 3702 14716
rect 3726 14714 3782 14716
rect 3806 14714 3862 14716
rect 3566 14662 3612 14714
rect 3612 14662 3622 14714
rect 3646 14662 3676 14714
rect 3676 14662 3688 14714
rect 3688 14662 3702 14714
rect 3726 14662 3740 14714
rect 3740 14662 3752 14714
rect 3752 14662 3782 14714
rect 3806 14662 3816 14714
rect 3816 14662 3862 14714
rect 3566 14660 3622 14662
rect 3646 14660 3702 14662
rect 3726 14660 3782 14662
rect 3806 14660 3862 14662
rect 3566 13626 3622 13628
rect 3646 13626 3702 13628
rect 3726 13626 3782 13628
rect 3806 13626 3862 13628
rect 3566 13574 3612 13626
rect 3612 13574 3622 13626
rect 3646 13574 3676 13626
rect 3676 13574 3688 13626
rect 3688 13574 3702 13626
rect 3726 13574 3740 13626
rect 3740 13574 3752 13626
rect 3752 13574 3782 13626
rect 3806 13574 3816 13626
rect 3816 13574 3862 13626
rect 3566 13572 3622 13574
rect 3646 13572 3702 13574
rect 3726 13572 3782 13574
rect 3806 13572 3862 13574
rect 4226 14170 4282 14172
rect 4306 14170 4362 14172
rect 4386 14170 4442 14172
rect 4466 14170 4522 14172
rect 4226 14118 4272 14170
rect 4272 14118 4282 14170
rect 4306 14118 4336 14170
rect 4336 14118 4348 14170
rect 4348 14118 4362 14170
rect 4386 14118 4400 14170
rect 4400 14118 4412 14170
rect 4412 14118 4442 14170
rect 4466 14118 4476 14170
rect 4476 14118 4522 14170
rect 4226 14116 4282 14118
rect 4306 14116 4362 14118
rect 4386 14116 4442 14118
rect 4466 14116 4522 14118
rect 9447 22874 9503 22876
rect 9527 22874 9583 22876
rect 9607 22874 9663 22876
rect 9687 22874 9743 22876
rect 9447 22822 9493 22874
rect 9493 22822 9503 22874
rect 9527 22822 9557 22874
rect 9557 22822 9569 22874
rect 9569 22822 9583 22874
rect 9607 22822 9621 22874
rect 9621 22822 9633 22874
rect 9633 22822 9663 22874
rect 9687 22822 9697 22874
rect 9697 22822 9743 22874
rect 9447 22820 9503 22822
rect 9527 22820 9583 22822
rect 9607 22820 9663 22822
rect 9687 22820 9743 22822
rect 6182 19488 6238 19544
rect 5354 17040 5410 17096
rect 4226 13082 4282 13084
rect 4306 13082 4362 13084
rect 4386 13082 4442 13084
rect 4466 13082 4522 13084
rect 4226 13030 4272 13082
rect 4272 13030 4282 13082
rect 4306 13030 4336 13082
rect 4336 13030 4348 13082
rect 4348 13030 4362 13082
rect 4386 13030 4400 13082
rect 4400 13030 4412 13082
rect 4412 13030 4442 13082
rect 4466 13030 4476 13082
rect 4476 13030 4522 13082
rect 4226 13028 4282 13030
rect 4306 13028 4362 13030
rect 4386 13028 4442 13030
rect 4466 13028 4522 13030
rect 5446 14320 5502 14376
rect 3566 12538 3622 12540
rect 3646 12538 3702 12540
rect 3726 12538 3782 12540
rect 3806 12538 3862 12540
rect 3566 12486 3612 12538
rect 3612 12486 3622 12538
rect 3646 12486 3676 12538
rect 3676 12486 3688 12538
rect 3688 12486 3702 12538
rect 3726 12486 3740 12538
rect 3740 12486 3752 12538
rect 3752 12486 3782 12538
rect 3806 12486 3816 12538
rect 3816 12486 3862 12538
rect 3566 12484 3622 12486
rect 3646 12484 3702 12486
rect 3726 12484 3782 12486
rect 3806 12484 3862 12486
rect 4226 11994 4282 11996
rect 4306 11994 4362 11996
rect 4386 11994 4442 11996
rect 4466 11994 4522 11996
rect 4226 11942 4272 11994
rect 4272 11942 4282 11994
rect 4306 11942 4336 11994
rect 4336 11942 4348 11994
rect 4348 11942 4362 11994
rect 4386 11942 4400 11994
rect 4400 11942 4412 11994
rect 4412 11942 4442 11994
rect 4466 11942 4476 11994
rect 4476 11942 4522 11994
rect 4226 11940 4282 11942
rect 4306 11940 4362 11942
rect 4386 11940 4442 11942
rect 4466 11940 4522 11942
rect 3238 11600 3294 11656
rect 3566 11450 3622 11452
rect 3646 11450 3702 11452
rect 3726 11450 3782 11452
rect 3806 11450 3862 11452
rect 3566 11398 3612 11450
rect 3612 11398 3622 11450
rect 3646 11398 3676 11450
rect 3676 11398 3688 11450
rect 3688 11398 3702 11450
rect 3726 11398 3740 11450
rect 3740 11398 3752 11450
rect 3752 11398 3782 11450
rect 3806 11398 3816 11450
rect 3816 11398 3862 11450
rect 3566 11396 3622 11398
rect 3646 11396 3702 11398
rect 3726 11396 3782 11398
rect 3806 11396 3862 11398
rect 4066 10920 4122 10976
rect 3566 10362 3622 10364
rect 3646 10362 3702 10364
rect 3726 10362 3782 10364
rect 3806 10362 3862 10364
rect 3566 10310 3612 10362
rect 3612 10310 3622 10362
rect 3646 10310 3676 10362
rect 3676 10310 3688 10362
rect 3688 10310 3702 10362
rect 3726 10310 3740 10362
rect 3740 10310 3752 10362
rect 3752 10310 3782 10362
rect 3806 10310 3816 10362
rect 3816 10310 3862 10362
rect 3566 10308 3622 10310
rect 3646 10308 3702 10310
rect 3726 10308 3782 10310
rect 3806 10308 3862 10310
rect 3882 9596 3884 9616
rect 3884 9596 3936 9616
rect 3936 9596 3938 9616
rect 3882 9560 3938 9596
rect 4226 10906 4282 10908
rect 4306 10906 4362 10908
rect 4386 10906 4442 10908
rect 4466 10906 4522 10908
rect 4226 10854 4272 10906
rect 4272 10854 4282 10906
rect 4306 10854 4336 10906
rect 4336 10854 4348 10906
rect 4348 10854 4362 10906
rect 4386 10854 4400 10906
rect 4400 10854 4412 10906
rect 4412 10854 4442 10906
rect 4466 10854 4476 10906
rect 4476 10854 4522 10906
rect 4226 10852 4282 10854
rect 4306 10852 4362 10854
rect 4386 10852 4442 10854
rect 4466 10852 4522 10854
rect 4226 9818 4282 9820
rect 4306 9818 4362 9820
rect 4386 9818 4442 9820
rect 4466 9818 4522 9820
rect 4226 9766 4272 9818
rect 4272 9766 4282 9818
rect 4306 9766 4336 9818
rect 4336 9766 4348 9818
rect 4348 9766 4362 9818
rect 4386 9766 4400 9818
rect 4400 9766 4412 9818
rect 4412 9766 4442 9818
rect 4466 9766 4476 9818
rect 4476 9766 4522 9818
rect 4226 9764 4282 9766
rect 4306 9764 4362 9766
rect 4386 9764 4442 9766
rect 4466 9764 4522 9766
rect 1306 8880 1362 8936
rect 1122 6840 1178 6896
rect 2778 7404 2834 7440
rect 2778 7384 2780 7404
rect 2780 7384 2832 7404
rect 2832 7384 2834 7404
rect 3566 9274 3622 9276
rect 3646 9274 3702 9276
rect 3726 9274 3782 9276
rect 3806 9274 3862 9276
rect 3566 9222 3612 9274
rect 3612 9222 3622 9274
rect 3646 9222 3676 9274
rect 3676 9222 3688 9274
rect 3688 9222 3702 9274
rect 3726 9222 3740 9274
rect 3740 9222 3752 9274
rect 3752 9222 3782 9274
rect 3806 9222 3816 9274
rect 3816 9222 3862 9274
rect 3566 9220 3622 9222
rect 3646 9220 3702 9222
rect 3726 9220 3782 9222
rect 3806 9220 3862 9222
rect 3566 8186 3622 8188
rect 3646 8186 3702 8188
rect 3726 8186 3782 8188
rect 3806 8186 3862 8188
rect 3566 8134 3612 8186
rect 3612 8134 3622 8186
rect 3646 8134 3676 8186
rect 3676 8134 3688 8186
rect 3688 8134 3702 8186
rect 3726 8134 3740 8186
rect 3740 8134 3752 8186
rect 3752 8134 3782 8186
rect 3806 8134 3816 8186
rect 3816 8134 3862 8186
rect 3566 8132 3622 8134
rect 3646 8132 3702 8134
rect 3726 8132 3782 8134
rect 3806 8132 3862 8134
rect 3790 7520 3846 7576
rect 4226 8730 4282 8732
rect 4306 8730 4362 8732
rect 4386 8730 4442 8732
rect 4466 8730 4522 8732
rect 4226 8678 4272 8730
rect 4272 8678 4282 8730
rect 4306 8678 4336 8730
rect 4336 8678 4348 8730
rect 4348 8678 4362 8730
rect 4386 8678 4400 8730
rect 4400 8678 4412 8730
rect 4412 8678 4442 8730
rect 4466 8678 4476 8730
rect 4476 8678 4522 8730
rect 4226 8676 4282 8678
rect 4306 8676 4362 8678
rect 4386 8676 4442 8678
rect 4466 8676 4522 8678
rect 3882 7384 3938 7440
rect 4226 7642 4282 7644
rect 4306 7642 4362 7644
rect 4386 7642 4442 7644
rect 4466 7642 4522 7644
rect 4226 7590 4272 7642
rect 4272 7590 4282 7642
rect 4306 7590 4336 7642
rect 4336 7590 4348 7642
rect 4348 7590 4362 7642
rect 4386 7590 4400 7642
rect 4400 7590 4412 7642
rect 4412 7590 4442 7642
rect 4466 7590 4476 7642
rect 4476 7590 4522 7642
rect 4226 7588 4282 7590
rect 4306 7588 4362 7590
rect 4386 7588 4442 7590
rect 4466 7588 4522 7590
rect 3566 7098 3622 7100
rect 3646 7098 3702 7100
rect 3726 7098 3782 7100
rect 3806 7098 3862 7100
rect 3566 7046 3612 7098
rect 3612 7046 3622 7098
rect 3646 7046 3676 7098
rect 3676 7046 3688 7098
rect 3688 7046 3702 7098
rect 3726 7046 3740 7098
rect 3740 7046 3752 7098
rect 3752 7046 3782 7098
rect 3806 7046 3816 7098
rect 3816 7046 3862 7098
rect 3566 7044 3622 7046
rect 3646 7044 3702 7046
rect 3726 7044 3782 7046
rect 3806 7044 3862 7046
rect 2962 6160 3018 6216
rect 2778 4140 2834 4176
rect 2778 4120 2780 4140
rect 2780 4120 2832 4140
rect 2832 4120 2834 4140
rect 2778 2760 2834 2816
rect 2962 2080 3018 2136
rect 3566 6010 3622 6012
rect 3646 6010 3702 6012
rect 3726 6010 3782 6012
rect 3806 6010 3862 6012
rect 3566 5958 3612 6010
rect 3612 5958 3622 6010
rect 3646 5958 3676 6010
rect 3676 5958 3688 6010
rect 3688 5958 3702 6010
rect 3726 5958 3740 6010
rect 3740 5958 3752 6010
rect 3752 5958 3782 6010
rect 3806 5958 3816 6010
rect 3816 5958 3862 6010
rect 3566 5956 3622 5958
rect 3646 5956 3702 5958
rect 3726 5956 3782 5958
rect 3806 5956 3862 5958
rect 3566 4922 3622 4924
rect 3646 4922 3702 4924
rect 3726 4922 3782 4924
rect 3806 4922 3862 4924
rect 3566 4870 3612 4922
rect 3612 4870 3622 4922
rect 3646 4870 3676 4922
rect 3676 4870 3688 4922
rect 3688 4870 3702 4922
rect 3726 4870 3740 4922
rect 3740 4870 3752 4922
rect 3752 4870 3782 4922
rect 3806 4870 3816 4922
rect 3816 4870 3862 4922
rect 3566 4868 3622 4870
rect 3646 4868 3702 4870
rect 3726 4868 3782 4870
rect 3806 4868 3862 4870
rect 3422 4800 3478 4856
rect 4226 6554 4282 6556
rect 4306 6554 4362 6556
rect 4386 6554 4442 6556
rect 4466 6554 4522 6556
rect 4226 6502 4272 6554
rect 4272 6502 4282 6554
rect 4306 6502 4336 6554
rect 4336 6502 4348 6554
rect 4348 6502 4362 6554
rect 4386 6502 4400 6554
rect 4400 6502 4412 6554
rect 4412 6502 4442 6554
rect 4466 6502 4476 6554
rect 4476 6502 4522 6554
rect 4226 6500 4282 6502
rect 4306 6500 4362 6502
rect 4386 6500 4442 6502
rect 4466 6500 4522 6502
rect 4894 7928 4950 7984
rect 8787 22330 8843 22332
rect 8867 22330 8923 22332
rect 8947 22330 9003 22332
rect 9027 22330 9083 22332
rect 8787 22278 8833 22330
rect 8833 22278 8843 22330
rect 8867 22278 8897 22330
rect 8897 22278 8909 22330
rect 8909 22278 8923 22330
rect 8947 22278 8961 22330
rect 8961 22278 8973 22330
rect 8973 22278 9003 22330
rect 9027 22278 9037 22330
rect 9037 22278 9083 22330
rect 8787 22276 8843 22278
rect 8867 22276 8923 22278
rect 8947 22276 9003 22278
rect 9027 22276 9083 22278
rect 8022 19508 8078 19544
rect 8022 19488 8024 19508
rect 8024 19488 8076 19508
rect 8076 19488 8078 19508
rect 8787 21242 8843 21244
rect 8867 21242 8923 21244
rect 8947 21242 9003 21244
rect 9027 21242 9083 21244
rect 8787 21190 8833 21242
rect 8833 21190 8843 21242
rect 8867 21190 8897 21242
rect 8897 21190 8909 21242
rect 8909 21190 8923 21242
rect 8947 21190 8961 21242
rect 8961 21190 8973 21242
rect 8973 21190 9003 21242
rect 9027 21190 9037 21242
rect 9037 21190 9083 21242
rect 8787 21188 8843 21190
rect 8867 21188 8923 21190
rect 8947 21188 9003 21190
rect 9027 21188 9083 21190
rect 9447 21786 9503 21788
rect 9527 21786 9583 21788
rect 9607 21786 9663 21788
rect 9687 21786 9743 21788
rect 9447 21734 9493 21786
rect 9493 21734 9503 21786
rect 9527 21734 9557 21786
rect 9557 21734 9569 21786
rect 9569 21734 9583 21786
rect 9607 21734 9621 21786
rect 9621 21734 9633 21786
rect 9633 21734 9663 21786
rect 9687 21734 9697 21786
rect 9697 21734 9743 21786
rect 9447 21732 9503 21734
rect 9527 21732 9583 21734
rect 9607 21732 9663 21734
rect 9687 21732 9743 21734
rect 8787 20154 8843 20156
rect 8867 20154 8923 20156
rect 8947 20154 9003 20156
rect 9027 20154 9083 20156
rect 8787 20102 8833 20154
rect 8833 20102 8843 20154
rect 8867 20102 8897 20154
rect 8897 20102 8909 20154
rect 8909 20102 8923 20154
rect 8947 20102 8961 20154
rect 8961 20102 8973 20154
rect 8973 20102 9003 20154
rect 9027 20102 9037 20154
rect 9037 20102 9083 20154
rect 8787 20100 8843 20102
rect 8867 20100 8923 20102
rect 8947 20100 9003 20102
rect 9027 20100 9083 20102
rect 9447 20698 9503 20700
rect 9527 20698 9583 20700
rect 9607 20698 9663 20700
rect 9687 20698 9743 20700
rect 9447 20646 9493 20698
rect 9493 20646 9503 20698
rect 9527 20646 9557 20698
rect 9557 20646 9569 20698
rect 9569 20646 9583 20698
rect 9607 20646 9621 20698
rect 9621 20646 9633 20698
rect 9633 20646 9663 20698
rect 9687 20646 9697 20698
rect 9697 20646 9743 20698
rect 9447 20644 9503 20646
rect 9527 20644 9583 20646
rect 9607 20644 9663 20646
rect 9687 20644 9743 20646
rect 9447 19610 9503 19612
rect 9527 19610 9583 19612
rect 9607 19610 9663 19612
rect 9687 19610 9743 19612
rect 9447 19558 9493 19610
rect 9493 19558 9503 19610
rect 9527 19558 9557 19610
rect 9557 19558 9569 19610
rect 9569 19558 9583 19610
rect 9607 19558 9621 19610
rect 9621 19558 9633 19610
rect 9633 19558 9663 19610
rect 9687 19558 9697 19610
rect 9697 19558 9743 19610
rect 9447 19556 9503 19558
rect 9527 19556 9583 19558
rect 9607 19556 9663 19558
rect 9687 19556 9743 19558
rect 8574 19372 8630 19408
rect 8574 19352 8576 19372
rect 8576 19352 8628 19372
rect 8628 19352 8630 19372
rect 8787 19066 8843 19068
rect 8867 19066 8923 19068
rect 8947 19066 9003 19068
rect 9027 19066 9083 19068
rect 8787 19014 8833 19066
rect 8833 19014 8843 19066
rect 8867 19014 8897 19066
rect 8897 19014 8909 19066
rect 8909 19014 8923 19066
rect 8947 19014 8961 19066
rect 8961 19014 8973 19066
rect 8973 19014 9003 19066
rect 9027 19014 9037 19066
rect 9037 19014 9083 19066
rect 8787 19012 8843 19014
rect 8867 19012 8923 19014
rect 8947 19012 9003 19014
rect 9027 19012 9083 19014
rect 8022 17212 8024 17232
rect 8024 17212 8076 17232
rect 8076 17212 8078 17232
rect 8022 17176 8078 17212
rect 9447 18522 9503 18524
rect 9527 18522 9583 18524
rect 9607 18522 9663 18524
rect 9687 18522 9743 18524
rect 9447 18470 9493 18522
rect 9493 18470 9503 18522
rect 9527 18470 9557 18522
rect 9557 18470 9569 18522
rect 9569 18470 9583 18522
rect 9607 18470 9621 18522
rect 9621 18470 9633 18522
rect 9633 18470 9663 18522
rect 9687 18470 9697 18522
rect 9697 18470 9743 18522
rect 9447 18468 9503 18470
rect 9527 18468 9583 18470
rect 9607 18468 9663 18470
rect 9687 18468 9743 18470
rect 8787 17978 8843 17980
rect 8867 17978 8923 17980
rect 8947 17978 9003 17980
rect 9027 17978 9083 17980
rect 8787 17926 8833 17978
rect 8833 17926 8843 17978
rect 8867 17926 8897 17978
rect 8897 17926 8909 17978
rect 8909 17926 8923 17978
rect 8947 17926 8961 17978
rect 8961 17926 8973 17978
rect 8973 17926 9003 17978
rect 9027 17926 9037 17978
rect 9037 17926 9083 17978
rect 8787 17924 8843 17926
rect 8867 17924 8923 17926
rect 8947 17924 9003 17926
rect 9027 17924 9083 17926
rect 5906 15000 5962 15056
rect 6458 13368 6514 13424
rect 3974 5480 4030 5536
rect 4226 5466 4282 5468
rect 4306 5466 4362 5468
rect 4386 5466 4442 5468
rect 4466 5466 4522 5468
rect 4226 5414 4272 5466
rect 4272 5414 4282 5466
rect 4306 5414 4336 5466
rect 4336 5414 4348 5466
rect 4348 5414 4362 5466
rect 4386 5414 4400 5466
rect 4400 5414 4412 5466
rect 4412 5414 4442 5466
rect 4466 5414 4476 5466
rect 4476 5414 4522 5466
rect 4226 5412 4282 5414
rect 4306 5412 4362 5414
rect 4386 5412 4442 5414
rect 4466 5412 4522 5414
rect 4226 4378 4282 4380
rect 4306 4378 4362 4380
rect 4386 4378 4442 4380
rect 4466 4378 4522 4380
rect 4226 4326 4272 4378
rect 4272 4326 4282 4378
rect 4306 4326 4336 4378
rect 4336 4326 4348 4378
rect 4348 4326 4362 4378
rect 4386 4326 4400 4378
rect 4400 4326 4412 4378
rect 4412 4326 4442 4378
rect 4466 4326 4476 4378
rect 4476 4326 4522 4378
rect 4226 4324 4282 4326
rect 4306 4324 4362 4326
rect 4386 4324 4442 4326
rect 4466 4324 4522 4326
rect 3566 3834 3622 3836
rect 3646 3834 3702 3836
rect 3726 3834 3782 3836
rect 3806 3834 3862 3836
rect 3566 3782 3612 3834
rect 3612 3782 3622 3834
rect 3646 3782 3676 3834
rect 3676 3782 3688 3834
rect 3688 3782 3702 3834
rect 3726 3782 3740 3834
rect 3740 3782 3752 3834
rect 3752 3782 3782 3834
rect 3806 3782 3816 3834
rect 3816 3782 3862 3834
rect 3566 3780 3622 3782
rect 3646 3780 3702 3782
rect 3726 3780 3782 3782
rect 3806 3780 3862 3782
rect 3566 2746 3622 2748
rect 3646 2746 3702 2748
rect 3726 2746 3782 2748
rect 3806 2746 3862 2748
rect 3566 2694 3612 2746
rect 3612 2694 3622 2746
rect 3646 2694 3676 2746
rect 3676 2694 3688 2746
rect 3688 2694 3702 2746
rect 3726 2694 3740 2746
rect 3740 2694 3752 2746
rect 3752 2694 3782 2746
rect 3806 2694 3816 2746
rect 3816 2694 3862 2746
rect 3566 2692 3622 2694
rect 3646 2692 3702 2694
rect 3726 2692 3782 2694
rect 3806 2692 3862 2694
rect 3422 856 3478 912
rect 4226 3290 4282 3292
rect 4306 3290 4362 3292
rect 4386 3290 4442 3292
rect 4466 3290 4522 3292
rect 4226 3238 4272 3290
rect 4272 3238 4282 3290
rect 4306 3238 4336 3290
rect 4336 3238 4348 3290
rect 4348 3238 4362 3290
rect 4386 3238 4400 3290
rect 4400 3238 4412 3290
rect 4412 3238 4442 3290
rect 4466 3238 4476 3290
rect 4476 3238 4522 3290
rect 4226 3236 4282 3238
rect 4306 3236 4362 3238
rect 4386 3236 4442 3238
rect 4466 3236 4522 3238
rect 4226 2202 4282 2204
rect 4306 2202 4362 2204
rect 4386 2202 4442 2204
rect 4466 2202 4522 2204
rect 4226 2150 4272 2202
rect 4272 2150 4282 2202
rect 4306 2150 4336 2202
rect 4336 2150 4348 2202
rect 4348 2150 4362 2202
rect 4386 2150 4400 2202
rect 4400 2150 4412 2202
rect 4412 2150 4442 2202
rect 4466 2150 4476 2202
rect 4476 2150 4522 2202
rect 4226 2148 4282 2150
rect 4306 2148 4362 2150
rect 4386 2148 4442 2150
rect 4466 2148 4522 2150
rect 4986 3440 5042 3496
rect 9447 17434 9503 17436
rect 9527 17434 9583 17436
rect 9607 17434 9663 17436
rect 9687 17434 9743 17436
rect 9447 17382 9493 17434
rect 9493 17382 9503 17434
rect 9527 17382 9557 17434
rect 9557 17382 9569 17434
rect 9569 17382 9583 17434
rect 9607 17382 9621 17434
rect 9621 17382 9633 17434
rect 9633 17382 9663 17434
rect 9687 17382 9697 17434
rect 9697 17382 9743 17434
rect 9447 17380 9503 17382
rect 9527 17380 9583 17382
rect 9607 17380 9663 17382
rect 9687 17380 9743 17382
rect 8787 16890 8843 16892
rect 8867 16890 8923 16892
rect 8947 16890 9003 16892
rect 9027 16890 9083 16892
rect 8787 16838 8833 16890
rect 8833 16838 8843 16890
rect 8867 16838 8897 16890
rect 8897 16838 8909 16890
rect 8909 16838 8923 16890
rect 8947 16838 8961 16890
rect 8961 16838 8973 16890
rect 8973 16838 9003 16890
rect 9027 16838 9037 16890
rect 9037 16838 9083 16890
rect 8787 16836 8843 16838
rect 8867 16836 8923 16838
rect 8947 16836 9003 16838
rect 9027 16836 9083 16838
rect 9447 16346 9503 16348
rect 9527 16346 9583 16348
rect 9607 16346 9663 16348
rect 9687 16346 9743 16348
rect 9447 16294 9493 16346
rect 9493 16294 9503 16346
rect 9527 16294 9557 16346
rect 9557 16294 9569 16346
rect 9569 16294 9583 16346
rect 9607 16294 9621 16346
rect 9621 16294 9633 16346
rect 9633 16294 9663 16346
rect 9687 16294 9697 16346
rect 9697 16294 9743 16346
rect 9447 16292 9503 16294
rect 9527 16292 9583 16294
rect 9607 16292 9663 16294
rect 9687 16292 9743 16294
rect 8787 15802 8843 15804
rect 8867 15802 8923 15804
rect 8947 15802 9003 15804
rect 9027 15802 9083 15804
rect 8787 15750 8833 15802
rect 8833 15750 8843 15802
rect 8867 15750 8897 15802
rect 8897 15750 8909 15802
rect 8909 15750 8923 15802
rect 8947 15750 8961 15802
rect 8961 15750 8973 15802
rect 8973 15750 9003 15802
rect 9027 15750 9037 15802
rect 9037 15750 9083 15802
rect 8787 15748 8843 15750
rect 8867 15748 8923 15750
rect 8947 15748 9003 15750
rect 9027 15748 9083 15750
rect 9447 15258 9503 15260
rect 9527 15258 9583 15260
rect 9607 15258 9663 15260
rect 9687 15258 9743 15260
rect 9447 15206 9493 15258
rect 9493 15206 9503 15258
rect 9527 15206 9557 15258
rect 9557 15206 9569 15258
rect 9569 15206 9583 15258
rect 9607 15206 9621 15258
rect 9621 15206 9633 15258
rect 9633 15206 9663 15258
rect 9687 15206 9697 15258
rect 9697 15206 9743 15258
rect 9447 15204 9503 15206
rect 9527 15204 9583 15206
rect 9607 15204 9663 15206
rect 9687 15204 9743 15206
rect 8787 14714 8843 14716
rect 8867 14714 8923 14716
rect 8947 14714 9003 14716
rect 9027 14714 9083 14716
rect 8787 14662 8833 14714
rect 8833 14662 8843 14714
rect 8867 14662 8897 14714
rect 8897 14662 8909 14714
rect 8909 14662 8923 14714
rect 8947 14662 8961 14714
rect 8961 14662 8973 14714
rect 8973 14662 9003 14714
rect 9027 14662 9037 14714
rect 9037 14662 9083 14714
rect 8787 14660 8843 14662
rect 8867 14660 8923 14662
rect 8947 14660 9003 14662
rect 9027 14660 9083 14662
rect 8787 13626 8843 13628
rect 8867 13626 8923 13628
rect 8947 13626 9003 13628
rect 9027 13626 9083 13628
rect 8787 13574 8833 13626
rect 8833 13574 8843 13626
rect 8867 13574 8897 13626
rect 8897 13574 8909 13626
rect 8909 13574 8923 13626
rect 8947 13574 8961 13626
rect 8961 13574 8973 13626
rect 8973 13574 9003 13626
rect 9027 13574 9037 13626
rect 9037 13574 9083 13626
rect 8787 13572 8843 13574
rect 8867 13572 8923 13574
rect 8947 13572 9003 13574
rect 9027 13572 9083 13574
rect 9447 14170 9503 14172
rect 9527 14170 9583 14172
rect 9607 14170 9663 14172
rect 9687 14170 9743 14172
rect 9447 14118 9493 14170
rect 9493 14118 9503 14170
rect 9527 14118 9557 14170
rect 9557 14118 9569 14170
rect 9569 14118 9583 14170
rect 9607 14118 9621 14170
rect 9621 14118 9633 14170
rect 9633 14118 9663 14170
rect 9687 14118 9697 14170
rect 9697 14118 9743 14170
rect 9447 14116 9503 14118
rect 9527 14116 9583 14118
rect 9607 14116 9663 14118
rect 9687 14116 9743 14118
rect 9862 13912 9918 13968
rect 9447 13082 9503 13084
rect 9527 13082 9583 13084
rect 9607 13082 9663 13084
rect 9687 13082 9743 13084
rect 9447 13030 9493 13082
rect 9493 13030 9503 13082
rect 9527 13030 9557 13082
rect 9557 13030 9569 13082
rect 9569 13030 9583 13082
rect 9607 13030 9621 13082
rect 9621 13030 9633 13082
rect 9633 13030 9663 13082
rect 9687 13030 9697 13082
rect 9697 13030 9743 13082
rect 9447 13028 9503 13030
rect 9527 13028 9583 13030
rect 9607 13028 9663 13030
rect 9687 13028 9743 13030
rect 8787 12538 8843 12540
rect 8867 12538 8923 12540
rect 8947 12538 9003 12540
rect 9027 12538 9083 12540
rect 8787 12486 8833 12538
rect 8833 12486 8843 12538
rect 8867 12486 8897 12538
rect 8897 12486 8909 12538
rect 8909 12486 8923 12538
rect 8947 12486 8961 12538
rect 8961 12486 8973 12538
rect 8973 12486 9003 12538
rect 9027 12486 9037 12538
rect 9037 12486 9083 12538
rect 8787 12484 8843 12486
rect 8867 12484 8923 12486
rect 8947 12484 9003 12486
rect 9027 12484 9083 12486
rect 8787 11450 8843 11452
rect 8867 11450 8923 11452
rect 8947 11450 9003 11452
rect 9027 11450 9083 11452
rect 8787 11398 8833 11450
rect 8833 11398 8843 11450
rect 8867 11398 8897 11450
rect 8897 11398 8909 11450
rect 8909 11398 8923 11450
rect 8947 11398 8961 11450
rect 8961 11398 8973 11450
rect 8973 11398 9003 11450
rect 9027 11398 9037 11450
rect 9037 11398 9083 11450
rect 8787 11396 8843 11398
rect 8867 11396 8923 11398
rect 8947 11396 9003 11398
rect 9027 11396 9083 11398
rect 9447 11994 9503 11996
rect 9527 11994 9583 11996
rect 9607 11994 9663 11996
rect 9687 11994 9743 11996
rect 9447 11942 9493 11994
rect 9493 11942 9503 11994
rect 9527 11942 9557 11994
rect 9557 11942 9569 11994
rect 9569 11942 9583 11994
rect 9607 11942 9621 11994
rect 9621 11942 9633 11994
rect 9633 11942 9663 11994
rect 9687 11942 9697 11994
rect 9697 11942 9743 11994
rect 9447 11940 9503 11942
rect 9527 11940 9583 11942
rect 9607 11940 9663 11942
rect 9687 11940 9743 11942
rect 9447 10906 9503 10908
rect 9527 10906 9583 10908
rect 9607 10906 9663 10908
rect 9687 10906 9743 10908
rect 9447 10854 9493 10906
rect 9493 10854 9503 10906
rect 9527 10854 9557 10906
rect 9557 10854 9569 10906
rect 9569 10854 9583 10906
rect 9607 10854 9621 10906
rect 9621 10854 9633 10906
rect 9633 10854 9663 10906
rect 9687 10854 9697 10906
rect 9697 10854 9743 10906
rect 9447 10852 9503 10854
rect 9527 10852 9583 10854
rect 9607 10852 9663 10854
rect 9687 10852 9743 10854
rect 8787 10362 8843 10364
rect 8867 10362 8923 10364
rect 8947 10362 9003 10364
rect 9027 10362 9083 10364
rect 8787 10310 8833 10362
rect 8833 10310 8843 10362
rect 8867 10310 8897 10362
rect 8897 10310 8909 10362
rect 8909 10310 8923 10362
rect 8947 10310 8961 10362
rect 8961 10310 8973 10362
rect 8973 10310 9003 10362
rect 9027 10310 9037 10362
rect 9037 10310 9083 10362
rect 8787 10308 8843 10310
rect 8867 10308 8923 10310
rect 8947 10308 9003 10310
rect 9027 10308 9083 10310
rect 9447 9818 9503 9820
rect 9527 9818 9583 9820
rect 9607 9818 9663 9820
rect 9687 9818 9743 9820
rect 9447 9766 9493 9818
rect 9493 9766 9503 9818
rect 9527 9766 9557 9818
rect 9557 9766 9569 9818
rect 9569 9766 9583 9818
rect 9607 9766 9621 9818
rect 9621 9766 9633 9818
rect 9633 9766 9663 9818
rect 9687 9766 9697 9818
rect 9697 9766 9743 9818
rect 9447 9764 9503 9766
rect 9527 9764 9583 9766
rect 9607 9764 9663 9766
rect 9687 9764 9743 9766
rect 8787 9274 8843 9276
rect 8867 9274 8923 9276
rect 8947 9274 9003 9276
rect 9027 9274 9083 9276
rect 8787 9222 8833 9274
rect 8833 9222 8843 9274
rect 8867 9222 8897 9274
rect 8897 9222 8909 9274
rect 8909 9222 8923 9274
rect 8947 9222 8961 9274
rect 8961 9222 8973 9274
rect 8973 9222 9003 9274
rect 9027 9222 9037 9274
rect 9037 9222 9083 9274
rect 8787 9220 8843 9222
rect 8867 9220 8923 9222
rect 8947 9220 9003 9222
rect 9027 9220 9083 9222
rect 8787 8186 8843 8188
rect 8867 8186 8923 8188
rect 8947 8186 9003 8188
rect 9027 8186 9083 8188
rect 8787 8134 8833 8186
rect 8833 8134 8843 8186
rect 8867 8134 8897 8186
rect 8897 8134 8909 8186
rect 8909 8134 8923 8186
rect 8947 8134 8961 8186
rect 8961 8134 8973 8186
rect 8973 8134 9003 8186
rect 9027 8134 9037 8186
rect 9037 8134 9083 8186
rect 8787 8132 8843 8134
rect 8867 8132 8923 8134
rect 8947 8132 9003 8134
rect 9027 8132 9083 8134
rect 8787 7098 8843 7100
rect 8867 7098 8923 7100
rect 8947 7098 9003 7100
rect 9027 7098 9083 7100
rect 8787 7046 8833 7098
rect 8833 7046 8843 7098
rect 8867 7046 8897 7098
rect 8897 7046 8909 7098
rect 8909 7046 8923 7098
rect 8947 7046 8961 7098
rect 8961 7046 8973 7098
rect 8973 7046 9003 7098
rect 9027 7046 9037 7098
rect 9037 7046 9083 7098
rect 8787 7044 8843 7046
rect 8867 7044 8923 7046
rect 8947 7044 9003 7046
rect 9027 7044 9083 7046
rect 9447 8730 9503 8732
rect 9527 8730 9583 8732
rect 9607 8730 9663 8732
rect 9687 8730 9743 8732
rect 9447 8678 9493 8730
rect 9493 8678 9503 8730
rect 9527 8678 9557 8730
rect 9557 8678 9569 8730
rect 9569 8678 9583 8730
rect 9607 8678 9621 8730
rect 9621 8678 9633 8730
rect 9633 8678 9663 8730
rect 9687 8678 9697 8730
rect 9697 8678 9743 8730
rect 9447 8676 9503 8678
rect 9527 8676 9583 8678
rect 9607 8676 9663 8678
rect 9687 8676 9743 8678
rect 9447 7642 9503 7644
rect 9527 7642 9583 7644
rect 9607 7642 9663 7644
rect 9687 7642 9743 7644
rect 9447 7590 9493 7642
rect 9493 7590 9503 7642
rect 9527 7590 9557 7642
rect 9557 7590 9569 7642
rect 9569 7590 9583 7642
rect 9607 7590 9621 7642
rect 9621 7590 9633 7642
rect 9633 7590 9663 7642
rect 9687 7590 9697 7642
rect 9697 7590 9743 7642
rect 9447 7588 9503 7590
rect 9527 7588 9583 7590
rect 9607 7588 9663 7590
rect 9687 7588 9743 7590
rect 9218 7384 9274 7440
rect 9218 6976 9274 7032
rect 9447 6554 9503 6556
rect 9527 6554 9583 6556
rect 9607 6554 9663 6556
rect 9687 6554 9743 6556
rect 9447 6502 9493 6554
rect 9493 6502 9503 6554
rect 9527 6502 9557 6554
rect 9557 6502 9569 6554
rect 9569 6502 9583 6554
rect 9607 6502 9621 6554
rect 9621 6502 9633 6554
rect 9633 6502 9663 6554
rect 9687 6502 9697 6554
rect 9697 6502 9743 6554
rect 9447 6500 9503 6502
rect 9527 6500 9583 6502
rect 9607 6500 9663 6502
rect 9687 6500 9743 6502
rect 8787 6010 8843 6012
rect 8867 6010 8923 6012
rect 8947 6010 9003 6012
rect 9027 6010 9083 6012
rect 8787 5958 8833 6010
rect 8833 5958 8843 6010
rect 8867 5958 8897 6010
rect 8897 5958 8909 6010
rect 8909 5958 8923 6010
rect 8947 5958 8961 6010
rect 8961 5958 8973 6010
rect 8973 5958 9003 6010
rect 9027 5958 9037 6010
rect 9037 5958 9083 6010
rect 8787 5956 8843 5958
rect 8867 5956 8923 5958
rect 8947 5956 9003 5958
rect 9027 5956 9083 5958
rect 5170 1400 5226 1456
rect 8787 4922 8843 4924
rect 8867 4922 8923 4924
rect 8947 4922 9003 4924
rect 9027 4922 9083 4924
rect 8787 4870 8833 4922
rect 8833 4870 8843 4922
rect 8867 4870 8897 4922
rect 8897 4870 8909 4922
rect 8909 4870 8923 4922
rect 8947 4870 8961 4922
rect 8961 4870 8973 4922
rect 8973 4870 9003 4922
rect 9027 4870 9037 4922
rect 9037 4870 9083 4922
rect 8787 4868 8843 4870
rect 8867 4868 8923 4870
rect 8947 4868 9003 4870
rect 9027 4868 9083 4870
rect 9954 6976 10010 7032
rect 11518 12280 11574 12336
rect 9954 6160 10010 6216
rect 9447 5466 9503 5468
rect 9527 5466 9583 5468
rect 9607 5466 9663 5468
rect 9687 5466 9743 5468
rect 9447 5414 9493 5466
rect 9493 5414 9503 5466
rect 9527 5414 9557 5466
rect 9557 5414 9569 5466
rect 9569 5414 9583 5466
rect 9607 5414 9621 5466
rect 9621 5414 9633 5466
rect 9633 5414 9663 5466
rect 9687 5414 9697 5466
rect 9697 5414 9743 5466
rect 9447 5412 9503 5414
rect 9527 5412 9583 5414
rect 9607 5412 9663 5414
rect 9687 5412 9743 5414
rect 9447 4378 9503 4380
rect 9527 4378 9583 4380
rect 9607 4378 9663 4380
rect 9687 4378 9743 4380
rect 9447 4326 9493 4378
rect 9493 4326 9503 4378
rect 9527 4326 9557 4378
rect 9557 4326 9569 4378
rect 9569 4326 9583 4378
rect 9607 4326 9621 4378
rect 9621 4326 9633 4378
rect 9633 4326 9663 4378
rect 9687 4326 9697 4378
rect 9697 4326 9743 4378
rect 9447 4324 9503 4326
rect 9527 4324 9583 4326
rect 9607 4324 9663 4326
rect 9687 4324 9743 4326
rect 8787 3834 8843 3836
rect 8867 3834 8923 3836
rect 8947 3834 9003 3836
rect 9027 3834 9083 3836
rect 8787 3782 8833 3834
rect 8833 3782 8843 3834
rect 8867 3782 8897 3834
rect 8897 3782 8909 3834
rect 8909 3782 8923 3834
rect 8947 3782 8961 3834
rect 8961 3782 8973 3834
rect 8973 3782 9003 3834
rect 9027 3782 9037 3834
rect 9037 3782 9083 3834
rect 8787 3780 8843 3782
rect 8867 3780 8923 3782
rect 8947 3780 9003 3782
rect 9027 3780 9083 3782
rect 9447 3290 9503 3292
rect 9527 3290 9583 3292
rect 9607 3290 9663 3292
rect 9687 3290 9743 3292
rect 9447 3238 9493 3290
rect 9493 3238 9503 3290
rect 9527 3238 9557 3290
rect 9557 3238 9569 3290
rect 9569 3238 9583 3290
rect 9607 3238 9621 3290
rect 9621 3238 9633 3290
rect 9633 3238 9663 3290
rect 9687 3238 9697 3290
rect 9697 3238 9743 3290
rect 9447 3236 9503 3238
rect 9527 3236 9583 3238
rect 9607 3236 9663 3238
rect 9687 3236 9743 3238
rect 8787 2746 8843 2748
rect 8867 2746 8923 2748
rect 8947 2746 9003 2748
rect 9027 2746 9083 2748
rect 8787 2694 8833 2746
rect 8833 2694 8843 2746
rect 8867 2694 8897 2746
rect 8897 2694 8909 2746
rect 8909 2694 8923 2746
rect 8947 2694 8961 2746
rect 8961 2694 8973 2746
rect 8973 2694 9003 2746
rect 9027 2694 9037 2746
rect 9037 2694 9083 2746
rect 8787 2692 8843 2694
rect 8867 2692 8923 2694
rect 8947 2692 9003 2694
rect 9027 2692 9083 2694
rect 9447 2202 9503 2204
rect 9527 2202 9583 2204
rect 9607 2202 9663 2204
rect 9687 2202 9743 2204
rect 9447 2150 9493 2202
rect 9493 2150 9503 2202
rect 9527 2150 9557 2202
rect 9557 2150 9569 2202
rect 9569 2150 9583 2202
rect 9607 2150 9621 2202
rect 9621 2150 9633 2202
rect 9633 2150 9663 2202
rect 9687 2150 9697 2202
rect 9697 2150 9743 2202
rect 9447 2148 9503 2150
rect 9527 2148 9583 2150
rect 9607 2148 9663 2150
rect 9687 2148 9743 2150
rect 10966 6316 11022 6352
rect 10966 6296 10968 6316
rect 10968 6296 11020 6316
rect 11020 6296 11022 6316
rect 14008 22330 14064 22332
rect 14088 22330 14144 22332
rect 14168 22330 14224 22332
rect 14248 22330 14304 22332
rect 14008 22278 14054 22330
rect 14054 22278 14064 22330
rect 14088 22278 14118 22330
rect 14118 22278 14130 22330
rect 14130 22278 14144 22330
rect 14168 22278 14182 22330
rect 14182 22278 14194 22330
rect 14194 22278 14224 22330
rect 14248 22278 14258 22330
rect 14258 22278 14304 22330
rect 14008 22276 14064 22278
rect 14088 22276 14144 22278
rect 14168 22276 14224 22278
rect 14248 22276 14304 22278
rect 14008 21242 14064 21244
rect 14088 21242 14144 21244
rect 14168 21242 14224 21244
rect 14248 21242 14304 21244
rect 14008 21190 14054 21242
rect 14054 21190 14064 21242
rect 14088 21190 14118 21242
rect 14118 21190 14130 21242
rect 14130 21190 14144 21242
rect 14168 21190 14182 21242
rect 14182 21190 14194 21242
rect 14194 21190 14224 21242
rect 14248 21190 14258 21242
rect 14258 21190 14304 21242
rect 14008 21188 14064 21190
rect 14088 21188 14144 21190
rect 14168 21188 14224 21190
rect 14248 21188 14304 21190
rect 14008 20154 14064 20156
rect 14088 20154 14144 20156
rect 14168 20154 14224 20156
rect 14248 20154 14304 20156
rect 14008 20102 14054 20154
rect 14054 20102 14064 20154
rect 14088 20102 14118 20154
rect 14118 20102 14130 20154
rect 14130 20102 14144 20154
rect 14168 20102 14182 20154
rect 14182 20102 14194 20154
rect 14194 20102 14224 20154
rect 14248 20102 14258 20154
rect 14258 20102 14304 20154
rect 14008 20100 14064 20102
rect 14088 20100 14144 20102
rect 14168 20100 14224 20102
rect 14248 20100 14304 20102
rect 14668 22874 14724 22876
rect 14748 22874 14804 22876
rect 14828 22874 14884 22876
rect 14908 22874 14964 22876
rect 14668 22822 14714 22874
rect 14714 22822 14724 22874
rect 14748 22822 14778 22874
rect 14778 22822 14790 22874
rect 14790 22822 14804 22874
rect 14828 22822 14842 22874
rect 14842 22822 14854 22874
rect 14854 22822 14884 22874
rect 14908 22822 14918 22874
rect 14918 22822 14964 22874
rect 14668 22820 14724 22822
rect 14748 22820 14804 22822
rect 14828 22820 14884 22822
rect 14908 22820 14964 22822
rect 14668 21786 14724 21788
rect 14748 21786 14804 21788
rect 14828 21786 14884 21788
rect 14908 21786 14964 21788
rect 14668 21734 14714 21786
rect 14714 21734 14724 21786
rect 14748 21734 14778 21786
rect 14778 21734 14790 21786
rect 14790 21734 14804 21786
rect 14828 21734 14842 21786
rect 14842 21734 14854 21786
rect 14854 21734 14884 21786
rect 14908 21734 14918 21786
rect 14918 21734 14964 21786
rect 14668 21732 14724 21734
rect 14748 21732 14804 21734
rect 14828 21732 14884 21734
rect 14908 21732 14964 21734
rect 14668 20698 14724 20700
rect 14748 20698 14804 20700
rect 14828 20698 14884 20700
rect 14908 20698 14964 20700
rect 14668 20646 14714 20698
rect 14714 20646 14724 20698
rect 14748 20646 14778 20698
rect 14778 20646 14790 20698
rect 14790 20646 14804 20698
rect 14828 20646 14842 20698
rect 14842 20646 14854 20698
rect 14854 20646 14884 20698
rect 14908 20646 14918 20698
rect 14918 20646 14964 20698
rect 14668 20644 14724 20646
rect 14748 20644 14804 20646
rect 14828 20644 14884 20646
rect 14908 20644 14964 20646
rect 14008 19066 14064 19068
rect 14088 19066 14144 19068
rect 14168 19066 14224 19068
rect 14248 19066 14304 19068
rect 14008 19014 14054 19066
rect 14054 19014 14064 19066
rect 14088 19014 14118 19066
rect 14118 19014 14130 19066
rect 14130 19014 14144 19066
rect 14168 19014 14182 19066
rect 14182 19014 14194 19066
rect 14194 19014 14224 19066
rect 14248 19014 14258 19066
rect 14258 19014 14304 19066
rect 14008 19012 14064 19014
rect 14088 19012 14144 19014
rect 14168 19012 14224 19014
rect 14248 19012 14304 19014
rect 14738 19780 14794 19816
rect 14738 19760 14740 19780
rect 14740 19760 14792 19780
rect 14792 19760 14794 19780
rect 14668 19610 14724 19612
rect 14748 19610 14804 19612
rect 14828 19610 14884 19612
rect 14908 19610 14964 19612
rect 14668 19558 14714 19610
rect 14714 19558 14724 19610
rect 14748 19558 14778 19610
rect 14778 19558 14790 19610
rect 14790 19558 14804 19610
rect 14828 19558 14842 19610
rect 14842 19558 14854 19610
rect 14854 19558 14884 19610
rect 14908 19558 14918 19610
rect 14918 19558 14964 19610
rect 14668 19556 14724 19558
rect 14748 19556 14804 19558
rect 14828 19556 14884 19558
rect 14908 19556 14964 19558
rect 14738 19352 14794 19408
rect 14668 18522 14724 18524
rect 14748 18522 14804 18524
rect 14828 18522 14884 18524
rect 14908 18522 14964 18524
rect 14668 18470 14714 18522
rect 14714 18470 14724 18522
rect 14748 18470 14778 18522
rect 14778 18470 14790 18522
rect 14790 18470 14804 18522
rect 14828 18470 14842 18522
rect 14842 18470 14854 18522
rect 14854 18470 14884 18522
rect 14908 18470 14918 18522
rect 14918 18470 14964 18522
rect 14668 18468 14724 18470
rect 14748 18468 14804 18470
rect 14828 18468 14884 18470
rect 14908 18468 14964 18470
rect 15014 18264 15070 18320
rect 14008 17978 14064 17980
rect 14088 17978 14144 17980
rect 14168 17978 14224 17980
rect 14248 17978 14304 17980
rect 14008 17926 14054 17978
rect 14054 17926 14064 17978
rect 14088 17926 14118 17978
rect 14118 17926 14130 17978
rect 14130 17926 14144 17978
rect 14168 17926 14182 17978
rect 14182 17926 14194 17978
rect 14194 17926 14224 17978
rect 14248 17926 14258 17978
rect 14258 17926 14304 17978
rect 14008 17924 14064 17926
rect 14088 17924 14144 17926
rect 14168 17924 14224 17926
rect 14248 17924 14304 17926
rect 14008 16890 14064 16892
rect 14088 16890 14144 16892
rect 14168 16890 14224 16892
rect 14248 16890 14304 16892
rect 14008 16838 14054 16890
rect 14054 16838 14064 16890
rect 14088 16838 14118 16890
rect 14118 16838 14130 16890
rect 14130 16838 14144 16890
rect 14168 16838 14182 16890
rect 14182 16838 14194 16890
rect 14194 16838 14224 16890
rect 14248 16838 14258 16890
rect 14258 16838 14304 16890
rect 14008 16836 14064 16838
rect 14088 16836 14144 16838
rect 14168 16836 14224 16838
rect 14248 16836 14304 16838
rect 14668 17434 14724 17436
rect 14748 17434 14804 17436
rect 14828 17434 14884 17436
rect 14908 17434 14964 17436
rect 14668 17382 14714 17434
rect 14714 17382 14724 17434
rect 14748 17382 14778 17434
rect 14778 17382 14790 17434
rect 14790 17382 14804 17434
rect 14828 17382 14842 17434
rect 14842 17382 14854 17434
rect 14854 17382 14884 17434
rect 14908 17382 14918 17434
rect 14918 17382 14964 17434
rect 14668 17380 14724 17382
rect 14748 17380 14804 17382
rect 14828 17380 14884 17382
rect 14908 17380 14964 17382
rect 15014 17176 15070 17232
rect 14462 16088 14518 16144
rect 14008 15802 14064 15804
rect 14088 15802 14144 15804
rect 14168 15802 14224 15804
rect 14248 15802 14304 15804
rect 14008 15750 14054 15802
rect 14054 15750 14064 15802
rect 14088 15750 14118 15802
rect 14118 15750 14130 15802
rect 14130 15750 14144 15802
rect 14168 15750 14182 15802
rect 14182 15750 14194 15802
rect 14194 15750 14224 15802
rect 14248 15750 14258 15802
rect 14258 15750 14304 15802
rect 14008 15748 14064 15750
rect 14088 15748 14144 15750
rect 14168 15748 14224 15750
rect 14248 15748 14304 15750
rect 14008 14714 14064 14716
rect 14088 14714 14144 14716
rect 14168 14714 14224 14716
rect 14248 14714 14304 14716
rect 14008 14662 14054 14714
rect 14054 14662 14064 14714
rect 14088 14662 14118 14714
rect 14118 14662 14130 14714
rect 14130 14662 14144 14714
rect 14168 14662 14182 14714
rect 14182 14662 14194 14714
rect 14194 14662 14224 14714
rect 14248 14662 14258 14714
rect 14258 14662 14304 14714
rect 14008 14660 14064 14662
rect 14088 14660 14144 14662
rect 14168 14660 14224 14662
rect 14248 14660 14304 14662
rect 13542 13912 13598 13968
rect 13266 12300 13322 12336
rect 13266 12280 13268 12300
rect 13268 12280 13320 12300
rect 13320 12280 13322 12300
rect 14008 13626 14064 13628
rect 14088 13626 14144 13628
rect 14168 13626 14224 13628
rect 14248 13626 14304 13628
rect 14008 13574 14054 13626
rect 14054 13574 14064 13626
rect 14088 13574 14118 13626
rect 14118 13574 14130 13626
rect 14130 13574 14144 13626
rect 14168 13574 14182 13626
rect 14182 13574 14194 13626
rect 14194 13574 14224 13626
rect 14248 13574 14258 13626
rect 14258 13574 14304 13626
rect 14008 13572 14064 13574
rect 14088 13572 14144 13574
rect 14168 13572 14224 13574
rect 14248 13572 14304 13574
rect 14668 16346 14724 16348
rect 14748 16346 14804 16348
rect 14828 16346 14884 16348
rect 14908 16346 14964 16348
rect 14668 16294 14714 16346
rect 14714 16294 14724 16346
rect 14748 16294 14778 16346
rect 14778 16294 14790 16346
rect 14790 16294 14804 16346
rect 14828 16294 14842 16346
rect 14842 16294 14854 16346
rect 14854 16294 14884 16346
rect 14908 16294 14918 16346
rect 14918 16294 14964 16346
rect 14668 16292 14724 16294
rect 14748 16292 14804 16294
rect 14828 16292 14884 16294
rect 14908 16292 14964 16294
rect 14668 15258 14724 15260
rect 14748 15258 14804 15260
rect 14828 15258 14884 15260
rect 14908 15258 14964 15260
rect 14668 15206 14714 15258
rect 14714 15206 14724 15258
rect 14748 15206 14778 15258
rect 14778 15206 14790 15258
rect 14790 15206 14804 15258
rect 14828 15206 14842 15258
rect 14842 15206 14854 15258
rect 14854 15206 14884 15258
rect 14908 15206 14918 15258
rect 14918 15206 14964 15258
rect 14668 15204 14724 15206
rect 14748 15204 14804 15206
rect 14828 15204 14884 15206
rect 14908 15204 14964 15206
rect 14668 14170 14724 14172
rect 14748 14170 14804 14172
rect 14828 14170 14884 14172
rect 14908 14170 14964 14172
rect 14668 14118 14714 14170
rect 14714 14118 14724 14170
rect 14748 14118 14778 14170
rect 14778 14118 14790 14170
rect 14790 14118 14804 14170
rect 14828 14118 14842 14170
rect 14842 14118 14854 14170
rect 14854 14118 14884 14170
rect 14908 14118 14918 14170
rect 14918 14118 14964 14170
rect 14668 14116 14724 14118
rect 14748 14116 14804 14118
rect 14828 14116 14884 14118
rect 14908 14116 14964 14118
rect 14830 13948 14832 13968
rect 14832 13948 14884 13968
rect 14884 13948 14886 13968
rect 14830 13912 14886 13948
rect 14008 12538 14064 12540
rect 14088 12538 14144 12540
rect 14168 12538 14224 12540
rect 14248 12538 14304 12540
rect 14008 12486 14054 12538
rect 14054 12486 14064 12538
rect 14088 12486 14118 12538
rect 14118 12486 14130 12538
rect 14130 12486 14144 12538
rect 14168 12486 14182 12538
rect 14182 12486 14194 12538
rect 14194 12486 14224 12538
rect 14248 12486 14258 12538
rect 14258 12486 14304 12538
rect 14008 12484 14064 12486
rect 14088 12484 14144 12486
rect 14168 12484 14224 12486
rect 14248 12484 14304 12486
rect 14008 11450 14064 11452
rect 14088 11450 14144 11452
rect 14168 11450 14224 11452
rect 14248 11450 14304 11452
rect 14008 11398 14054 11450
rect 14054 11398 14064 11450
rect 14088 11398 14118 11450
rect 14118 11398 14130 11450
rect 14130 11398 14144 11450
rect 14168 11398 14182 11450
rect 14182 11398 14194 11450
rect 14194 11398 14224 11450
rect 14248 11398 14258 11450
rect 14258 11398 14304 11450
rect 14008 11396 14064 11398
rect 14088 11396 14144 11398
rect 14168 11396 14224 11398
rect 14248 11396 14304 11398
rect 14668 13082 14724 13084
rect 14748 13082 14804 13084
rect 14828 13082 14884 13084
rect 14908 13082 14964 13084
rect 14668 13030 14714 13082
rect 14714 13030 14724 13082
rect 14748 13030 14778 13082
rect 14778 13030 14790 13082
rect 14790 13030 14804 13082
rect 14828 13030 14842 13082
rect 14842 13030 14854 13082
rect 14854 13030 14884 13082
rect 14908 13030 14918 13082
rect 14918 13030 14964 13082
rect 14668 13028 14724 13030
rect 14748 13028 14804 13030
rect 14828 13028 14884 13030
rect 14908 13028 14964 13030
rect 14668 11994 14724 11996
rect 14748 11994 14804 11996
rect 14828 11994 14884 11996
rect 14908 11994 14964 11996
rect 14668 11942 14714 11994
rect 14714 11942 14724 11994
rect 14748 11942 14778 11994
rect 14778 11942 14790 11994
rect 14790 11942 14804 11994
rect 14828 11942 14842 11994
rect 14842 11942 14854 11994
rect 14854 11942 14884 11994
rect 14908 11942 14918 11994
rect 14918 11942 14964 11994
rect 14668 11940 14724 11942
rect 14748 11940 14804 11942
rect 14828 11940 14884 11942
rect 14908 11940 14964 11942
rect 14668 10906 14724 10908
rect 14748 10906 14804 10908
rect 14828 10906 14884 10908
rect 14908 10906 14964 10908
rect 14668 10854 14714 10906
rect 14714 10854 14724 10906
rect 14748 10854 14778 10906
rect 14778 10854 14790 10906
rect 14790 10854 14804 10906
rect 14828 10854 14842 10906
rect 14842 10854 14854 10906
rect 14854 10854 14884 10906
rect 14908 10854 14918 10906
rect 14918 10854 14964 10906
rect 14668 10852 14724 10854
rect 14748 10852 14804 10854
rect 14828 10852 14884 10854
rect 14908 10852 14964 10854
rect 14008 10362 14064 10364
rect 14088 10362 14144 10364
rect 14168 10362 14224 10364
rect 14248 10362 14304 10364
rect 14008 10310 14054 10362
rect 14054 10310 14064 10362
rect 14088 10310 14118 10362
rect 14118 10310 14130 10362
rect 14130 10310 14144 10362
rect 14168 10310 14182 10362
rect 14182 10310 14194 10362
rect 14194 10310 14224 10362
rect 14248 10310 14258 10362
rect 14258 10310 14304 10362
rect 14008 10308 14064 10310
rect 14088 10308 14144 10310
rect 14168 10308 14224 10310
rect 14248 10308 14304 10310
rect 14668 9818 14724 9820
rect 14748 9818 14804 9820
rect 14828 9818 14884 9820
rect 14908 9818 14964 9820
rect 14668 9766 14714 9818
rect 14714 9766 14724 9818
rect 14748 9766 14778 9818
rect 14778 9766 14790 9818
rect 14790 9766 14804 9818
rect 14828 9766 14842 9818
rect 14842 9766 14854 9818
rect 14854 9766 14884 9818
rect 14908 9766 14918 9818
rect 14918 9766 14964 9818
rect 14668 9764 14724 9766
rect 14748 9764 14804 9766
rect 14828 9764 14884 9766
rect 14908 9764 14964 9766
rect 14008 9274 14064 9276
rect 14088 9274 14144 9276
rect 14168 9274 14224 9276
rect 14248 9274 14304 9276
rect 14008 9222 14054 9274
rect 14054 9222 14064 9274
rect 14088 9222 14118 9274
rect 14118 9222 14130 9274
rect 14130 9222 14144 9274
rect 14168 9222 14182 9274
rect 14182 9222 14194 9274
rect 14194 9222 14224 9274
rect 14248 9222 14258 9274
rect 14258 9222 14304 9274
rect 14008 9220 14064 9222
rect 14088 9220 14144 9222
rect 14168 9220 14224 9222
rect 14248 9220 14304 9222
rect 14668 8730 14724 8732
rect 14748 8730 14804 8732
rect 14828 8730 14884 8732
rect 14908 8730 14964 8732
rect 14668 8678 14714 8730
rect 14714 8678 14724 8730
rect 14748 8678 14778 8730
rect 14778 8678 14790 8730
rect 14790 8678 14804 8730
rect 14828 8678 14842 8730
rect 14842 8678 14854 8730
rect 14854 8678 14884 8730
rect 14908 8678 14918 8730
rect 14918 8678 14964 8730
rect 14668 8676 14724 8678
rect 14748 8676 14804 8678
rect 14828 8676 14884 8678
rect 14908 8676 14964 8678
rect 14008 8186 14064 8188
rect 14088 8186 14144 8188
rect 14168 8186 14224 8188
rect 14248 8186 14304 8188
rect 14008 8134 14054 8186
rect 14054 8134 14064 8186
rect 14088 8134 14118 8186
rect 14118 8134 14130 8186
rect 14130 8134 14144 8186
rect 14168 8134 14182 8186
rect 14182 8134 14194 8186
rect 14194 8134 14224 8186
rect 14248 8134 14258 8186
rect 14258 8134 14304 8186
rect 14008 8132 14064 8134
rect 14088 8132 14144 8134
rect 14168 8132 14224 8134
rect 14248 8132 14304 8134
rect 14462 8492 14518 8528
rect 14462 8472 14464 8492
rect 14464 8472 14516 8492
rect 14516 8472 14518 8492
rect 14008 7098 14064 7100
rect 14088 7098 14144 7100
rect 14168 7098 14224 7100
rect 14248 7098 14304 7100
rect 14008 7046 14054 7098
rect 14054 7046 14064 7098
rect 14088 7046 14118 7098
rect 14118 7046 14130 7098
rect 14130 7046 14144 7098
rect 14168 7046 14182 7098
rect 14182 7046 14194 7098
rect 14194 7046 14224 7098
rect 14248 7046 14258 7098
rect 14258 7046 14304 7098
rect 14008 7044 14064 7046
rect 14088 7044 14144 7046
rect 14168 7044 14224 7046
rect 14248 7044 14304 7046
rect 13450 6432 13506 6488
rect 13450 6160 13506 6216
rect 14008 6010 14064 6012
rect 14088 6010 14144 6012
rect 14168 6010 14224 6012
rect 14248 6010 14304 6012
rect 14008 5958 14054 6010
rect 14054 5958 14064 6010
rect 14088 5958 14118 6010
rect 14118 5958 14130 6010
rect 14130 5958 14144 6010
rect 14168 5958 14182 6010
rect 14182 5958 14194 6010
rect 14194 5958 14224 6010
rect 14248 5958 14258 6010
rect 14258 5958 14304 6010
rect 14008 5956 14064 5958
rect 14088 5956 14144 5958
rect 14168 5956 14224 5958
rect 14248 5956 14304 5958
rect 14008 4922 14064 4924
rect 14088 4922 14144 4924
rect 14168 4922 14224 4924
rect 14248 4922 14304 4924
rect 14008 4870 14054 4922
rect 14054 4870 14064 4922
rect 14088 4870 14118 4922
rect 14118 4870 14130 4922
rect 14130 4870 14144 4922
rect 14168 4870 14182 4922
rect 14182 4870 14194 4922
rect 14194 4870 14224 4922
rect 14248 4870 14258 4922
rect 14258 4870 14304 4922
rect 14008 4868 14064 4870
rect 14088 4868 14144 4870
rect 14168 4868 14224 4870
rect 14248 4868 14304 4870
rect 14008 3834 14064 3836
rect 14088 3834 14144 3836
rect 14168 3834 14224 3836
rect 14248 3834 14304 3836
rect 14008 3782 14054 3834
rect 14054 3782 14064 3834
rect 14088 3782 14118 3834
rect 14118 3782 14130 3834
rect 14130 3782 14144 3834
rect 14168 3782 14182 3834
rect 14182 3782 14194 3834
rect 14194 3782 14224 3834
rect 14248 3782 14258 3834
rect 14258 3782 14304 3834
rect 14008 3780 14064 3782
rect 14088 3780 14144 3782
rect 14168 3780 14224 3782
rect 14248 3780 14304 3782
rect 14008 2746 14064 2748
rect 14088 2746 14144 2748
rect 14168 2746 14224 2748
rect 14248 2746 14304 2748
rect 14008 2694 14054 2746
rect 14054 2694 14064 2746
rect 14088 2694 14118 2746
rect 14118 2694 14130 2746
rect 14130 2694 14144 2746
rect 14168 2694 14182 2746
rect 14182 2694 14194 2746
rect 14194 2694 14224 2746
rect 14248 2694 14258 2746
rect 14258 2694 14304 2746
rect 14008 2692 14064 2694
rect 14088 2692 14144 2694
rect 14168 2692 14224 2694
rect 14248 2692 14304 2694
rect 19889 22874 19945 22876
rect 19969 22874 20025 22876
rect 20049 22874 20105 22876
rect 20129 22874 20185 22876
rect 19889 22822 19935 22874
rect 19935 22822 19945 22874
rect 19969 22822 19999 22874
rect 19999 22822 20011 22874
rect 20011 22822 20025 22874
rect 20049 22822 20063 22874
rect 20063 22822 20075 22874
rect 20075 22822 20105 22874
rect 20129 22822 20139 22874
rect 20139 22822 20185 22874
rect 19889 22820 19945 22822
rect 19969 22820 20025 22822
rect 20049 22820 20105 22822
rect 20129 22820 20185 22822
rect 19229 22330 19285 22332
rect 19309 22330 19365 22332
rect 19389 22330 19445 22332
rect 19469 22330 19525 22332
rect 19229 22278 19275 22330
rect 19275 22278 19285 22330
rect 19309 22278 19339 22330
rect 19339 22278 19351 22330
rect 19351 22278 19365 22330
rect 19389 22278 19403 22330
rect 19403 22278 19415 22330
rect 19415 22278 19445 22330
rect 19469 22278 19479 22330
rect 19479 22278 19525 22330
rect 19229 22276 19285 22278
rect 19309 22276 19365 22278
rect 19389 22276 19445 22278
rect 19469 22276 19525 22278
rect 18602 20984 18658 21040
rect 17866 18572 17868 18592
rect 17868 18572 17920 18592
rect 17920 18572 17922 18592
rect 17866 18536 17922 18572
rect 17958 17720 18014 17776
rect 17222 16496 17278 16552
rect 17958 15544 18014 15600
rect 16486 12824 16542 12880
rect 19229 21242 19285 21244
rect 19309 21242 19365 21244
rect 19389 21242 19445 21244
rect 19469 21242 19525 21244
rect 19229 21190 19275 21242
rect 19275 21190 19285 21242
rect 19309 21190 19339 21242
rect 19339 21190 19351 21242
rect 19351 21190 19365 21242
rect 19389 21190 19403 21242
rect 19403 21190 19415 21242
rect 19415 21190 19445 21242
rect 19469 21190 19479 21242
rect 19479 21190 19525 21242
rect 19229 21188 19285 21190
rect 19309 21188 19365 21190
rect 19389 21188 19445 21190
rect 19469 21188 19525 21190
rect 19889 21786 19945 21788
rect 19969 21786 20025 21788
rect 20049 21786 20105 21788
rect 20129 21786 20185 21788
rect 19889 21734 19935 21786
rect 19935 21734 19945 21786
rect 19969 21734 19999 21786
rect 19999 21734 20011 21786
rect 20011 21734 20025 21786
rect 20049 21734 20063 21786
rect 20063 21734 20075 21786
rect 20075 21734 20105 21786
rect 20129 21734 20139 21786
rect 20139 21734 20185 21786
rect 19889 21732 19945 21734
rect 19969 21732 20025 21734
rect 20049 21732 20105 21734
rect 20129 21732 20185 21734
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19469 20154 19525 20156
rect 19229 20102 19275 20154
rect 19275 20102 19285 20154
rect 19309 20102 19339 20154
rect 19339 20102 19351 20154
rect 19351 20102 19365 20154
rect 19389 20102 19403 20154
rect 19403 20102 19415 20154
rect 19415 20102 19445 20154
rect 19469 20102 19479 20154
rect 19479 20102 19525 20154
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19469 20100 19525 20102
rect 19889 20698 19945 20700
rect 19969 20698 20025 20700
rect 20049 20698 20105 20700
rect 20129 20698 20185 20700
rect 19889 20646 19935 20698
rect 19935 20646 19945 20698
rect 19969 20646 19999 20698
rect 19999 20646 20011 20698
rect 20011 20646 20025 20698
rect 20049 20646 20063 20698
rect 20063 20646 20075 20698
rect 20075 20646 20105 20698
rect 20129 20646 20139 20698
rect 20139 20646 20185 20698
rect 19889 20644 19945 20646
rect 19969 20644 20025 20646
rect 20049 20644 20105 20646
rect 20129 20644 20185 20646
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19469 19066 19525 19068
rect 19229 19014 19275 19066
rect 19275 19014 19285 19066
rect 19309 19014 19339 19066
rect 19339 19014 19351 19066
rect 19351 19014 19365 19066
rect 19389 19014 19403 19066
rect 19403 19014 19415 19066
rect 19415 19014 19445 19066
rect 19469 19014 19479 19066
rect 19479 19014 19525 19066
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19469 19012 19525 19014
rect 18970 18808 19026 18864
rect 18694 18284 18750 18320
rect 18694 18264 18696 18284
rect 18696 18264 18748 18284
rect 18748 18264 18750 18284
rect 19889 19610 19945 19612
rect 19969 19610 20025 19612
rect 20049 19610 20105 19612
rect 20129 19610 20185 19612
rect 19889 19558 19935 19610
rect 19935 19558 19945 19610
rect 19969 19558 19999 19610
rect 19999 19558 20011 19610
rect 20011 19558 20025 19610
rect 20049 19558 20063 19610
rect 20063 19558 20075 19610
rect 20075 19558 20105 19610
rect 20129 19558 20139 19610
rect 20139 19558 20185 19610
rect 19889 19556 19945 19558
rect 19969 19556 20025 19558
rect 20049 19556 20105 19558
rect 20129 19556 20185 19558
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19469 17978 19525 17980
rect 19229 17926 19275 17978
rect 19275 17926 19285 17978
rect 19309 17926 19339 17978
rect 19339 17926 19351 17978
rect 19351 17926 19365 17978
rect 19389 17926 19403 17978
rect 19403 17926 19415 17978
rect 19415 17926 19445 17978
rect 19469 17926 19479 17978
rect 19479 17926 19525 17978
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19469 17924 19525 17926
rect 21086 21836 21088 21856
rect 21088 21836 21140 21856
rect 21140 21836 21142 21856
rect 21086 21800 21142 21836
rect 21178 21120 21234 21176
rect 21086 20984 21142 21040
rect 21178 20460 21234 20496
rect 21178 20440 21180 20460
rect 21180 20440 21232 20460
rect 21232 20440 21234 20460
rect 20626 19760 20682 19816
rect 19889 18522 19945 18524
rect 19969 18522 20025 18524
rect 20049 18522 20105 18524
rect 20129 18522 20185 18524
rect 19889 18470 19935 18522
rect 19935 18470 19945 18522
rect 19969 18470 19999 18522
rect 19999 18470 20011 18522
rect 20011 18470 20025 18522
rect 20049 18470 20063 18522
rect 20063 18470 20075 18522
rect 20075 18470 20105 18522
rect 20129 18470 20139 18522
rect 20139 18470 20185 18522
rect 19889 18468 19945 18470
rect 19969 18468 20025 18470
rect 20049 18468 20105 18470
rect 20129 18468 20185 18470
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19469 16890 19525 16892
rect 19229 16838 19275 16890
rect 19275 16838 19285 16890
rect 19309 16838 19339 16890
rect 19339 16838 19351 16890
rect 19351 16838 19365 16890
rect 19389 16838 19403 16890
rect 19403 16838 19415 16890
rect 19415 16838 19445 16890
rect 19469 16838 19479 16890
rect 19479 16838 19525 16890
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19469 16836 19525 16838
rect 19889 17434 19945 17436
rect 19969 17434 20025 17436
rect 20049 17434 20105 17436
rect 20129 17434 20185 17436
rect 19889 17382 19935 17434
rect 19935 17382 19945 17434
rect 19969 17382 19999 17434
rect 19999 17382 20011 17434
rect 20011 17382 20025 17434
rect 20049 17382 20063 17434
rect 20063 17382 20075 17434
rect 20075 17382 20105 17434
rect 20129 17382 20139 17434
rect 20139 17382 20185 17434
rect 19889 17380 19945 17382
rect 19969 17380 20025 17382
rect 20049 17380 20105 17382
rect 20129 17380 20185 17382
rect 19889 16346 19945 16348
rect 19969 16346 20025 16348
rect 20049 16346 20105 16348
rect 20129 16346 20185 16348
rect 19889 16294 19935 16346
rect 19935 16294 19945 16346
rect 19969 16294 19999 16346
rect 19999 16294 20011 16346
rect 20011 16294 20025 16346
rect 20049 16294 20063 16346
rect 20063 16294 20075 16346
rect 20075 16294 20105 16346
rect 20129 16294 20139 16346
rect 20139 16294 20185 16346
rect 19889 16292 19945 16294
rect 19969 16292 20025 16294
rect 20049 16292 20105 16294
rect 20129 16292 20185 16294
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19469 15802 19525 15804
rect 19229 15750 19275 15802
rect 19275 15750 19285 15802
rect 19309 15750 19339 15802
rect 19339 15750 19351 15802
rect 19351 15750 19365 15802
rect 19389 15750 19403 15802
rect 19403 15750 19415 15802
rect 19415 15750 19445 15802
rect 19469 15750 19479 15802
rect 19479 15750 19525 15802
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19469 15748 19525 15750
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19469 14714 19525 14716
rect 19229 14662 19275 14714
rect 19275 14662 19285 14714
rect 19309 14662 19339 14714
rect 19339 14662 19351 14714
rect 19351 14662 19365 14714
rect 19389 14662 19403 14714
rect 19403 14662 19415 14714
rect 19415 14662 19445 14714
rect 19469 14662 19479 14714
rect 19479 14662 19525 14714
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19469 14660 19525 14662
rect 19522 14456 19578 14512
rect 18786 13912 18842 13968
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19469 13626 19525 13628
rect 19229 13574 19275 13626
rect 19275 13574 19285 13626
rect 19309 13574 19339 13626
rect 19339 13574 19351 13626
rect 19351 13574 19365 13626
rect 19389 13574 19403 13626
rect 19403 13574 19415 13626
rect 19415 13574 19445 13626
rect 19469 13574 19479 13626
rect 19479 13574 19525 13626
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19469 13572 19525 13574
rect 14668 7642 14724 7644
rect 14748 7642 14804 7644
rect 14828 7642 14884 7644
rect 14908 7642 14964 7644
rect 14668 7590 14714 7642
rect 14714 7590 14724 7642
rect 14748 7590 14778 7642
rect 14778 7590 14790 7642
rect 14790 7590 14804 7642
rect 14828 7590 14842 7642
rect 14842 7590 14854 7642
rect 14854 7590 14884 7642
rect 14908 7590 14918 7642
rect 14918 7590 14964 7642
rect 14668 7588 14724 7590
rect 14748 7588 14804 7590
rect 14828 7588 14884 7590
rect 14908 7588 14964 7590
rect 17222 10648 17278 10704
rect 14668 6554 14724 6556
rect 14748 6554 14804 6556
rect 14828 6554 14884 6556
rect 14908 6554 14964 6556
rect 14668 6502 14714 6554
rect 14714 6502 14724 6554
rect 14748 6502 14778 6554
rect 14778 6502 14790 6554
rect 14790 6502 14804 6554
rect 14828 6502 14842 6554
rect 14842 6502 14854 6554
rect 14854 6502 14884 6554
rect 14908 6502 14918 6554
rect 14918 6502 14964 6554
rect 14668 6500 14724 6502
rect 14748 6500 14804 6502
rect 14828 6500 14884 6502
rect 14908 6500 14964 6502
rect 14668 5466 14724 5468
rect 14748 5466 14804 5468
rect 14828 5466 14884 5468
rect 14908 5466 14964 5468
rect 14668 5414 14714 5466
rect 14714 5414 14724 5466
rect 14748 5414 14778 5466
rect 14778 5414 14790 5466
rect 14790 5414 14804 5466
rect 14828 5414 14842 5466
rect 14842 5414 14854 5466
rect 14854 5414 14884 5466
rect 14908 5414 14918 5466
rect 14918 5414 14964 5466
rect 14668 5412 14724 5414
rect 14748 5412 14804 5414
rect 14828 5412 14884 5414
rect 14908 5412 14964 5414
rect 14668 4378 14724 4380
rect 14748 4378 14804 4380
rect 14828 4378 14884 4380
rect 14908 4378 14964 4380
rect 14668 4326 14714 4378
rect 14714 4326 14724 4378
rect 14748 4326 14778 4378
rect 14778 4326 14790 4378
rect 14790 4326 14804 4378
rect 14828 4326 14842 4378
rect 14842 4326 14854 4378
rect 14854 4326 14884 4378
rect 14908 4326 14918 4378
rect 14918 4326 14964 4378
rect 14668 4324 14724 4326
rect 14748 4324 14804 4326
rect 14828 4324 14884 4326
rect 14908 4324 14964 4326
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19469 12538 19525 12540
rect 19229 12486 19275 12538
rect 19275 12486 19285 12538
rect 19309 12486 19339 12538
rect 19339 12486 19351 12538
rect 19351 12486 19365 12538
rect 19389 12486 19403 12538
rect 19403 12486 19415 12538
rect 19415 12486 19445 12538
rect 19469 12486 19479 12538
rect 19479 12486 19525 12538
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19469 12484 19525 12486
rect 18602 12316 18604 12336
rect 18604 12316 18656 12336
rect 18656 12316 18658 12336
rect 18602 12280 18658 12316
rect 19889 15258 19945 15260
rect 19969 15258 20025 15260
rect 20049 15258 20105 15260
rect 20129 15258 20185 15260
rect 19889 15206 19935 15258
rect 19935 15206 19945 15258
rect 19969 15206 19999 15258
rect 19999 15206 20011 15258
rect 20011 15206 20025 15258
rect 20049 15206 20063 15258
rect 20063 15206 20075 15258
rect 20075 15206 20105 15258
rect 20129 15206 20139 15258
rect 20139 15206 20185 15258
rect 19889 15204 19945 15206
rect 19969 15204 20025 15206
rect 20049 15204 20105 15206
rect 20129 15204 20185 15206
rect 19889 14170 19945 14172
rect 19969 14170 20025 14172
rect 20049 14170 20105 14172
rect 20129 14170 20185 14172
rect 19889 14118 19935 14170
rect 19935 14118 19945 14170
rect 19969 14118 19999 14170
rect 19999 14118 20011 14170
rect 20011 14118 20025 14170
rect 20049 14118 20063 14170
rect 20063 14118 20075 14170
rect 20075 14118 20105 14170
rect 20129 14118 20139 14170
rect 20139 14118 20185 14170
rect 19889 14116 19945 14118
rect 19969 14116 20025 14118
rect 20049 14116 20105 14118
rect 20129 14116 20185 14118
rect 19889 13082 19945 13084
rect 19969 13082 20025 13084
rect 20049 13082 20105 13084
rect 20129 13082 20185 13084
rect 19889 13030 19935 13082
rect 19935 13030 19945 13082
rect 19969 13030 19999 13082
rect 19999 13030 20011 13082
rect 20011 13030 20025 13082
rect 20049 13030 20063 13082
rect 20063 13030 20075 13082
rect 20075 13030 20105 13082
rect 20129 13030 20139 13082
rect 20139 13030 20185 13082
rect 19889 13028 19945 13030
rect 19969 13028 20025 13030
rect 20049 13028 20105 13030
rect 20129 13028 20185 13030
rect 20718 15000 20774 15056
rect 19889 11994 19945 11996
rect 19969 11994 20025 11996
rect 20049 11994 20105 11996
rect 20129 11994 20185 11996
rect 19889 11942 19935 11994
rect 19935 11942 19945 11994
rect 19969 11942 19999 11994
rect 19999 11942 20011 11994
rect 20011 11942 20025 11994
rect 20049 11942 20063 11994
rect 20063 11942 20075 11994
rect 20075 11942 20105 11994
rect 20129 11942 20139 11994
rect 20139 11942 20185 11994
rect 19889 11940 19945 11942
rect 19969 11940 20025 11942
rect 20049 11940 20105 11942
rect 20129 11940 20185 11942
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19469 11450 19525 11452
rect 19229 11398 19275 11450
rect 19275 11398 19285 11450
rect 19309 11398 19339 11450
rect 19339 11398 19351 11450
rect 19351 11398 19365 11450
rect 19389 11398 19403 11450
rect 19403 11398 19415 11450
rect 19415 11398 19445 11450
rect 19469 11398 19479 11450
rect 19479 11398 19525 11450
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19469 11396 19525 11398
rect 18050 10104 18106 10160
rect 17038 7384 17094 7440
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19469 10362 19525 10364
rect 19229 10310 19275 10362
rect 19275 10310 19285 10362
rect 19309 10310 19339 10362
rect 19339 10310 19351 10362
rect 19351 10310 19365 10362
rect 19389 10310 19403 10362
rect 19403 10310 19415 10362
rect 19415 10310 19445 10362
rect 19469 10310 19479 10362
rect 19479 10310 19525 10362
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19469 10308 19525 10310
rect 19889 10906 19945 10908
rect 19969 10906 20025 10908
rect 20049 10906 20105 10908
rect 20129 10906 20185 10908
rect 19889 10854 19935 10906
rect 19935 10854 19945 10906
rect 19969 10854 19999 10906
rect 19999 10854 20011 10906
rect 20011 10854 20025 10906
rect 20049 10854 20063 10906
rect 20063 10854 20075 10906
rect 20075 10854 20105 10906
rect 20129 10854 20139 10906
rect 20139 10854 20185 10906
rect 19889 10852 19945 10854
rect 19969 10852 20025 10854
rect 20049 10852 20105 10854
rect 20129 10852 20185 10854
rect 19889 9818 19945 9820
rect 19969 9818 20025 9820
rect 20049 9818 20105 9820
rect 20129 9818 20185 9820
rect 19889 9766 19935 9818
rect 19935 9766 19945 9818
rect 19969 9766 19999 9818
rect 19999 9766 20011 9818
rect 20011 9766 20025 9818
rect 20049 9766 20063 9818
rect 20063 9766 20075 9818
rect 20075 9766 20105 9818
rect 20129 9766 20139 9818
rect 20139 9766 20185 9818
rect 19889 9764 19945 9766
rect 19969 9764 20025 9766
rect 20049 9764 20105 9766
rect 20129 9764 20185 9766
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19469 9274 19525 9276
rect 19229 9222 19275 9274
rect 19275 9222 19285 9274
rect 19309 9222 19339 9274
rect 19339 9222 19351 9274
rect 19351 9222 19365 9274
rect 19389 9222 19403 9274
rect 19403 9222 19415 9274
rect 19415 9222 19445 9274
rect 19469 9222 19479 9274
rect 19479 9222 19525 9274
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19469 9220 19525 9222
rect 18142 8472 18198 8528
rect 14668 3290 14724 3292
rect 14748 3290 14804 3292
rect 14828 3290 14884 3292
rect 14908 3290 14964 3292
rect 14668 3238 14714 3290
rect 14714 3238 14724 3290
rect 14748 3238 14778 3290
rect 14778 3238 14790 3290
rect 14790 3238 14804 3290
rect 14828 3238 14842 3290
rect 14842 3238 14854 3290
rect 14854 3238 14884 3290
rect 14908 3238 14918 3290
rect 14918 3238 14964 3290
rect 14668 3236 14724 3238
rect 14748 3236 14804 3238
rect 14828 3236 14884 3238
rect 14908 3236 14964 3238
rect 14668 2202 14724 2204
rect 14748 2202 14804 2204
rect 14828 2202 14884 2204
rect 14908 2202 14964 2204
rect 14668 2150 14714 2202
rect 14714 2150 14724 2202
rect 14748 2150 14778 2202
rect 14778 2150 14790 2202
rect 14790 2150 14804 2202
rect 14828 2150 14842 2202
rect 14842 2150 14854 2202
rect 14854 2150 14884 2202
rect 14908 2150 14918 2202
rect 14918 2150 14964 2202
rect 14668 2148 14724 2150
rect 14748 2148 14804 2150
rect 14828 2148 14884 2150
rect 14908 2148 14964 2150
rect 18050 6296 18106 6352
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19469 8186 19525 8188
rect 19229 8134 19275 8186
rect 19275 8134 19285 8186
rect 19309 8134 19339 8186
rect 19339 8134 19351 8186
rect 19351 8134 19365 8186
rect 19389 8134 19403 8186
rect 19403 8134 19415 8186
rect 19415 8134 19445 8186
rect 19469 8134 19479 8186
rect 19479 8134 19525 8186
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19469 8132 19525 8134
rect 19889 8730 19945 8732
rect 19969 8730 20025 8732
rect 20049 8730 20105 8732
rect 20129 8730 20185 8732
rect 19889 8678 19935 8730
rect 19935 8678 19945 8730
rect 19969 8678 19999 8730
rect 19999 8678 20011 8730
rect 20011 8678 20025 8730
rect 20049 8678 20063 8730
rect 20063 8678 20075 8730
rect 20075 8678 20105 8730
rect 20129 8678 20139 8730
rect 20139 8678 20185 8730
rect 19889 8676 19945 8678
rect 19969 8676 20025 8678
rect 20049 8676 20105 8678
rect 20129 8676 20185 8678
rect 21270 17040 21326 17096
rect 21546 18400 21602 18456
rect 21454 14476 21510 14512
rect 21454 14456 21456 14476
rect 21456 14456 21508 14476
rect 21508 14456 21510 14476
rect 21362 14320 21418 14376
rect 21546 13640 21602 13696
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19469 7098 19525 7100
rect 19229 7046 19275 7098
rect 19275 7046 19285 7098
rect 19309 7046 19339 7098
rect 19339 7046 19351 7098
rect 19351 7046 19365 7098
rect 19389 7046 19403 7098
rect 19403 7046 19415 7098
rect 19415 7046 19445 7098
rect 19469 7046 19479 7098
rect 19479 7046 19525 7098
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19469 7044 19525 7046
rect 18418 4120 18474 4176
rect 19889 7642 19945 7644
rect 19969 7642 20025 7644
rect 20049 7642 20105 7644
rect 20129 7642 20185 7644
rect 19889 7590 19935 7642
rect 19935 7590 19945 7642
rect 19969 7590 19999 7642
rect 19999 7590 20011 7642
rect 20011 7590 20025 7642
rect 20049 7590 20063 7642
rect 20063 7590 20075 7642
rect 20075 7590 20105 7642
rect 20129 7590 20139 7642
rect 20139 7590 20185 7642
rect 19889 7588 19945 7590
rect 19969 7588 20025 7590
rect 20049 7588 20105 7590
rect 20129 7588 20185 7590
rect 19889 6554 19945 6556
rect 19969 6554 20025 6556
rect 20049 6554 20105 6556
rect 20129 6554 20185 6556
rect 19889 6502 19935 6554
rect 19935 6502 19945 6554
rect 19969 6502 19999 6554
rect 19999 6502 20011 6554
rect 20011 6502 20025 6554
rect 20049 6502 20063 6554
rect 20063 6502 20075 6554
rect 20075 6502 20105 6554
rect 20129 6502 20139 6554
rect 20139 6502 20185 6554
rect 19889 6500 19945 6502
rect 19969 6500 20025 6502
rect 20049 6500 20105 6502
rect 20129 6500 20185 6502
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19469 6010 19525 6012
rect 19229 5958 19275 6010
rect 19275 5958 19285 6010
rect 19309 5958 19339 6010
rect 19339 5958 19351 6010
rect 19351 5958 19365 6010
rect 19389 5958 19403 6010
rect 19403 5958 19415 6010
rect 19415 5958 19445 6010
rect 19469 5958 19479 6010
rect 19479 5958 19525 6010
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19469 5956 19525 5958
rect 21362 11600 21418 11656
rect 21362 9560 21418 9616
rect 20810 8880 20866 8936
rect 20626 8200 20682 8256
rect 21362 6840 21418 6896
rect 21086 6180 21142 6216
rect 21086 6160 21088 6180
rect 21088 6160 21140 6180
rect 21140 6160 21142 6180
rect 20350 5480 20406 5536
rect 19889 5466 19945 5468
rect 19969 5466 20025 5468
rect 20049 5466 20105 5468
rect 20129 5466 20185 5468
rect 19889 5414 19935 5466
rect 19935 5414 19945 5466
rect 19969 5414 19999 5466
rect 19999 5414 20011 5466
rect 20011 5414 20025 5466
rect 20049 5414 20063 5466
rect 20063 5414 20075 5466
rect 20075 5414 20105 5466
rect 20129 5414 20139 5466
rect 20139 5414 20185 5466
rect 19889 5412 19945 5414
rect 19969 5412 20025 5414
rect 20049 5412 20105 5414
rect 20129 5412 20185 5414
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19469 4922 19525 4924
rect 19229 4870 19275 4922
rect 19275 4870 19285 4922
rect 19309 4870 19339 4922
rect 19339 4870 19351 4922
rect 19351 4870 19365 4922
rect 19389 4870 19403 4922
rect 19403 4870 19415 4922
rect 19415 4870 19445 4922
rect 19469 4870 19479 4922
rect 19479 4870 19525 4922
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19469 4868 19525 4870
rect 19889 4378 19945 4380
rect 19969 4378 20025 4380
rect 20049 4378 20105 4380
rect 20129 4378 20185 4380
rect 19889 4326 19935 4378
rect 19935 4326 19945 4378
rect 19969 4326 19999 4378
rect 19999 4326 20011 4378
rect 20011 4326 20025 4378
rect 20049 4326 20063 4378
rect 20063 4326 20075 4378
rect 20075 4326 20105 4378
rect 20129 4326 20139 4378
rect 20139 4326 20185 4378
rect 19889 4324 19945 4326
rect 19969 4324 20025 4326
rect 20049 4324 20105 4326
rect 20129 4324 20185 4326
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19469 3834 19525 3836
rect 19229 3782 19275 3834
rect 19275 3782 19285 3834
rect 19309 3782 19339 3834
rect 19339 3782 19351 3834
rect 19351 3782 19365 3834
rect 19389 3782 19403 3834
rect 19403 3782 19415 3834
rect 19415 3782 19445 3834
rect 19469 3782 19479 3834
rect 19479 3782 19525 3834
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19469 3780 19525 3782
rect 21546 4820 21602 4856
rect 21546 4800 21548 4820
rect 21548 4800 21600 4820
rect 21600 4800 21602 4820
rect 21362 3440 21418 3496
rect 19889 3290 19945 3292
rect 19969 3290 20025 3292
rect 20049 3290 20105 3292
rect 20129 3290 20185 3292
rect 19889 3238 19935 3290
rect 19935 3238 19945 3290
rect 19969 3238 19999 3290
rect 19999 3238 20011 3290
rect 20011 3238 20025 3290
rect 20049 3238 20063 3290
rect 20063 3238 20075 3290
rect 20075 3238 20105 3290
rect 20129 3238 20139 3290
rect 20139 3238 20185 3290
rect 19889 3236 19945 3238
rect 19969 3236 20025 3238
rect 20049 3236 20105 3238
rect 20129 3236 20185 3238
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19469 2746 19525 2748
rect 19229 2694 19275 2746
rect 19275 2694 19285 2746
rect 19309 2694 19339 2746
rect 19339 2694 19351 2746
rect 19351 2694 19365 2746
rect 19389 2694 19403 2746
rect 19403 2694 19415 2746
rect 19415 2694 19445 2746
rect 19469 2694 19479 2746
rect 19479 2694 19525 2746
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19469 2692 19525 2694
rect 19889 2202 19945 2204
rect 19969 2202 20025 2204
rect 20049 2202 20105 2204
rect 20129 2202 20185 2204
rect 19889 2150 19935 2202
rect 19935 2150 19945 2202
rect 19969 2150 19999 2202
rect 19999 2150 20011 2202
rect 20011 2150 20025 2202
rect 20049 2150 20063 2202
rect 20063 2150 20075 2202
rect 20075 2150 20105 2202
rect 20129 2150 20139 2202
rect 20139 2150 20185 2202
rect 19889 2148 19945 2150
rect 19969 2148 20025 2150
rect 20049 2148 20105 2150
rect 20129 2148 20185 2150
<< metal3 >>
rect 4216 22880 4532 22881
rect 4216 22816 4222 22880
rect 4286 22816 4302 22880
rect 4366 22816 4382 22880
rect 4446 22816 4462 22880
rect 4526 22816 4532 22880
rect 4216 22815 4532 22816
rect 9437 22880 9753 22881
rect 9437 22816 9443 22880
rect 9507 22816 9523 22880
rect 9587 22816 9603 22880
rect 9667 22816 9683 22880
rect 9747 22816 9753 22880
rect 9437 22815 9753 22816
rect 14658 22880 14974 22881
rect 14658 22816 14664 22880
rect 14728 22816 14744 22880
rect 14808 22816 14824 22880
rect 14888 22816 14904 22880
rect 14968 22816 14974 22880
rect 14658 22815 14974 22816
rect 19879 22880 20195 22881
rect 19879 22816 19885 22880
rect 19949 22816 19965 22880
rect 20029 22816 20045 22880
rect 20109 22816 20125 22880
rect 20189 22816 20195 22880
rect 19879 22815 20195 22816
rect 3556 22336 3872 22337
rect 3556 22272 3562 22336
rect 3626 22272 3642 22336
rect 3706 22272 3722 22336
rect 3786 22272 3802 22336
rect 3866 22272 3872 22336
rect 3556 22271 3872 22272
rect 8777 22336 9093 22337
rect 8777 22272 8783 22336
rect 8847 22272 8863 22336
rect 8927 22272 8943 22336
rect 9007 22272 9023 22336
rect 9087 22272 9093 22336
rect 8777 22271 9093 22272
rect 13998 22336 14314 22337
rect 13998 22272 14004 22336
rect 14068 22272 14084 22336
rect 14148 22272 14164 22336
rect 14228 22272 14244 22336
rect 14308 22272 14314 22336
rect 13998 22271 14314 22272
rect 19219 22336 19535 22337
rect 19219 22272 19225 22336
rect 19289 22272 19305 22336
rect 19369 22272 19385 22336
rect 19449 22272 19465 22336
rect 19529 22272 19535 22336
rect 19219 22271 19535 22272
rect 0 21858 800 21888
rect 3049 21858 3115 21861
rect 0 21856 3115 21858
rect 0 21800 3054 21856
rect 3110 21800 3115 21856
rect 0 21798 3115 21800
rect 0 21768 800 21798
rect 3049 21795 3115 21798
rect 21081 21858 21147 21861
rect 22331 21858 23131 21888
rect 21081 21856 23131 21858
rect 21081 21800 21086 21856
rect 21142 21800 23131 21856
rect 21081 21798 23131 21800
rect 21081 21795 21147 21798
rect 4216 21792 4532 21793
rect 4216 21728 4222 21792
rect 4286 21728 4302 21792
rect 4366 21728 4382 21792
rect 4446 21728 4462 21792
rect 4526 21728 4532 21792
rect 4216 21727 4532 21728
rect 9437 21792 9753 21793
rect 9437 21728 9443 21792
rect 9507 21728 9523 21792
rect 9587 21728 9603 21792
rect 9667 21728 9683 21792
rect 9747 21728 9753 21792
rect 9437 21727 9753 21728
rect 14658 21792 14974 21793
rect 14658 21728 14664 21792
rect 14728 21728 14744 21792
rect 14808 21728 14824 21792
rect 14888 21728 14904 21792
rect 14968 21728 14974 21792
rect 14658 21727 14974 21728
rect 19879 21792 20195 21793
rect 19879 21728 19885 21792
rect 19949 21728 19965 21792
rect 20029 21728 20045 21792
rect 20109 21728 20125 21792
rect 20189 21728 20195 21792
rect 22331 21768 23131 21798
rect 19879 21727 20195 21728
rect 3556 21248 3872 21249
rect 0 21178 800 21208
rect 3556 21184 3562 21248
rect 3626 21184 3642 21248
rect 3706 21184 3722 21248
rect 3786 21184 3802 21248
rect 3866 21184 3872 21248
rect 3556 21183 3872 21184
rect 8777 21248 9093 21249
rect 8777 21184 8783 21248
rect 8847 21184 8863 21248
rect 8927 21184 8943 21248
rect 9007 21184 9023 21248
rect 9087 21184 9093 21248
rect 8777 21183 9093 21184
rect 13998 21248 14314 21249
rect 13998 21184 14004 21248
rect 14068 21184 14084 21248
rect 14148 21184 14164 21248
rect 14228 21184 14244 21248
rect 14308 21184 14314 21248
rect 13998 21183 14314 21184
rect 19219 21248 19535 21249
rect 19219 21184 19225 21248
rect 19289 21184 19305 21248
rect 19369 21184 19385 21248
rect 19449 21184 19465 21248
rect 19529 21184 19535 21248
rect 19219 21183 19535 21184
rect 2998 21178 3004 21180
rect 0 21118 3004 21178
rect 0 21088 800 21118
rect 2998 21116 3004 21118
rect 3068 21116 3074 21180
rect 21173 21178 21239 21181
rect 22331 21178 23131 21208
rect 21173 21176 23131 21178
rect 21173 21120 21178 21176
rect 21234 21120 23131 21176
rect 21173 21118 23131 21120
rect 21173 21115 21239 21118
rect 22331 21088 23131 21118
rect 18597 21042 18663 21045
rect 21081 21042 21147 21045
rect 18597 21040 21147 21042
rect 18597 20984 18602 21040
rect 18658 20984 21086 21040
rect 21142 20984 21147 21040
rect 18597 20982 21147 20984
rect 18597 20979 18663 20982
rect 21081 20979 21147 20982
rect 4216 20704 4532 20705
rect 4216 20640 4222 20704
rect 4286 20640 4302 20704
rect 4366 20640 4382 20704
rect 4446 20640 4462 20704
rect 4526 20640 4532 20704
rect 4216 20639 4532 20640
rect 9437 20704 9753 20705
rect 9437 20640 9443 20704
rect 9507 20640 9523 20704
rect 9587 20640 9603 20704
rect 9667 20640 9683 20704
rect 9747 20640 9753 20704
rect 9437 20639 9753 20640
rect 14658 20704 14974 20705
rect 14658 20640 14664 20704
rect 14728 20640 14744 20704
rect 14808 20640 14824 20704
rect 14888 20640 14904 20704
rect 14968 20640 14974 20704
rect 14658 20639 14974 20640
rect 19879 20704 20195 20705
rect 19879 20640 19885 20704
rect 19949 20640 19965 20704
rect 20029 20640 20045 20704
rect 20109 20640 20125 20704
rect 20189 20640 20195 20704
rect 19879 20639 20195 20640
rect 0 20498 800 20528
rect 2681 20498 2747 20501
rect 0 20496 2747 20498
rect 0 20440 2686 20496
rect 2742 20440 2747 20496
rect 0 20438 2747 20440
rect 0 20408 800 20438
rect 2681 20435 2747 20438
rect 21173 20498 21239 20501
rect 22331 20498 23131 20528
rect 21173 20496 23131 20498
rect 21173 20440 21178 20496
rect 21234 20440 23131 20496
rect 21173 20438 23131 20440
rect 21173 20435 21239 20438
rect 22331 20408 23131 20438
rect 3556 20160 3872 20161
rect 3556 20096 3562 20160
rect 3626 20096 3642 20160
rect 3706 20096 3722 20160
rect 3786 20096 3802 20160
rect 3866 20096 3872 20160
rect 3556 20095 3872 20096
rect 8777 20160 9093 20161
rect 8777 20096 8783 20160
rect 8847 20096 8863 20160
rect 8927 20096 8943 20160
rect 9007 20096 9023 20160
rect 9087 20096 9093 20160
rect 8777 20095 9093 20096
rect 13998 20160 14314 20161
rect 13998 20096 14004 20160
rect 14068 20096 14084 20160
rect 14148 20096 14164 20160
rect 14228 20096 14244 20160
rect 14308 20096 14314 20160
rect 13998 20095 14314 20096
rect 19219 20160 19535 20161
rect 19219 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19465 20160
rect 19529 20096 19535 20160
rect 19219 20095 19535 20096
rect 0 19818 800 19848
rect 4797 19818 4863 19821
rect 14733 19818 14799 19821
rect 0 19816 4863 19818
rect 0 19760 4802 19816
rect 4858 19760 4863 19816
rect 0 19758 4863 19760
rect 0 19728 800 19758
rect 4797 19755 4863 19758
rect 14414 19816 14799 19818
rect 14414 19760 14738 19816
rect 14794 19760 14799 19816
rect 14414 19758 14799 19760
rect 4216 19616 4532 19617
rect 4216 19552 4222 19616
rect 4286 19552 4302 19616
rect 4366 19552 4382 19616
rect 4446 19552 4462 19616
rect 4526 19552 4532 19616
rect 4216 19551 4532 19552
rect 9437 19616 9753 19617
rect 9437 19552 9443 19616
rect 9507 19552 9523 19616
rect 9587 19552 9603 19616
rect 9667 19552 9683 19616
rect 9747 19552 9753 19616
rect 9437 19551 9753 19552
rect 6177 19546 6243 19549
rect 8017 19546 8083 19549
rect 6177 19544 8083 19546
rect 6177 19488 6182 19544
rect 6238 19488 8022 19544
rect 8078 19488 8083 19544
rect 6177 19486 8083 19488
rect 6177 19483 6243 19486
rect 8017 19483 8083 19486
rect 8569 19412 8635 19413
rect 8518 19348 8524 19412
rect 8588 19410 8635 19412
rect 14414 19410 14474 19758
rect 14733 19755 14799 19758
rect 20621 19818 20687 19821
rect 22331 19818 23131 19848
rect 20621 19816 23131 19818
rect 20621 19760 20626 19816
rect 20682 19760 23131 19816
rect 20621 19758 23131 19760
rect 20621 19755 20687 19758
rect 22331 19728 23131 19758
rect 14658 19616 14974 19617
rect 14658 19552 14664 19616
rect 14728 19552 14744 19616
rect 14808 19552 14824 19616
rect 14888 19552 14904 19616
rect 14968 19552 14974 19616
rect 14658 19551 14974 19552
rect 19879 19616 20195 19617
rect 19879 19552 19885 19616
rect 19949 19552 19965 19616
rect 20029 19552 20045 19616
rect 20109 19552 20125 19616
rect 20189 19552 20195 19616
rect 19879 19551 20195 19552
rect 14733 19410 14799 19413
rect 8588 19408 8680 19410
rect 8630 19352 8680 19408
rect 8588 19350 8680 19352
rect 14414 19408 14799 19410
rect 14414 19352 14738 19408
rect 14794 19352 14799 19408
rect 14414 19350 14799 19352
rect 8588 19348 8635 19350
rect 8569 19347 8635 19348
rect 14733 19347 14799 19350
rect 0 19138 800 19168
rect 1301 19138 1367 19141
rect 22331 19138 23131 19168
rect 0 19136 1367 19138
rect 0 19080 1306 19136
rect 1362 19080 1367 19136
rect 0 19078 1367 19080
rect 0 19048 800 19078
rect 1301 19075 1367 19078
rect 19934 19078 23131 19138
rect 3556 19072 3872 19073
rect 3556 19008 3562 19072
rect 3626 19008 3642 19072
rect 3706 19008 3722 19072
rect 3786 19008 3802 19072
rect 3866 19008 3872 19072
rect 3556 19007 3872 19008
rect 8777 19072 9093 19073
rect 8777 19008 8783 19072
rect 8847 19008 8863 19072
rect 8927 19008 8943 19072
rect 9007 19008 9023 19072
rect 9087 19008 9093 19072
rect 8777 19007 9093 19008
rect 13998 19072 14314 19073
rect 13998 19008 14004 19072
rect 14068 19008 14084 19072
rect 14148 19008 14164 19072
rect 14228 19008 14244 19072
rect 14308 19008 14314 19072
rect 13998 19007 14314 19008
rect 19219 19072 19535 19073
rect 19219 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19465 19072
rect 19529 19008 19535 19072
rect 19219 19007 19535 19008
rect 18965 18866 19031 18869
rect 19934 18866 19994 19078
rect 22331 19048 23131 19078
rect 18965 18864 19994 18866
rect 18965 18808 18970 18864
rect 19026 18808 19994 18864
rect 18965 18806 19994 18808
rect 18965 18803 19031 18806
rect 17718 18532 17724 18596
rect 17788 18594 17794 18596
rect 17861 18594 17927 18597
rect 17788 18592 17927 18594
rect 17788 18536 17866 18592
rect 17922 18536 17927 18592
rect 17788 18534 17927 18536
rect 17788 18532 17794 18534
rect 17861 18531 17927 18534
rect 4216 18528 4532 18529
rect 0 18458 800 18488
rect 4216 18464 4222 18528
rect 4286 18464 4302 18528
rect 4366 18464 4382 18528
rect 4446 18464 4462 18528
rect 4526 18464 4532 18528
rect 4216 18463 4532 18464
rect 9437 18528 9753 18529
rect 9437 18464 9443 18528
rect 9507 18464 9523 18528
rect 9587 18464 9603 18528
rect 9667 18464 9683 18528
rect 9747 18464 9753 18528
rect 9437 18463 9753 18464
rect 14658 18528 14974 18529
rect 14658 18464 14664 18528
rect 14728 18464 14744 18528
rect 14808 18464 14824 18528
rect 14888 18464 14904 18528
rect 14968 18464 14974 18528
rect 14658 18463 14974 18464
rect 19879 18528 20195 18529
rect 19879 18464 19885 18528
rect 19949 18464 19965 18528
rect 20029 18464 20045 18528
rect 20109 18464 20125 18528
rect 20189 18464 20195 18528
rect 19879 18463 20195 18464
rect 21541 18458 21607 18461
rect 22331 18458 23131 18488
rect 0 18398 2790 18458
rect 0 18368 800 18398
rect 2730 18322 2790 18398
rect 21541 18456 23131 18458
rect 21541 18400 21546 18456
rect 21602 18400 23131 18456
rect 21541 18398 23131 18400
rect 21541 18395 21607 18398
rect 22331 18368 23131 18398
rect 4337 18322 4403 18325
rect 2730 18320 4403 18322
rect 2730 18264 4342 18320
rect 4398 18264 4403 18320
rect 2730 18262 4403 18264
rect 4337 18259 4403 18262
rect 15009 18322 15075 18325
rect 18689 18322 18755 18325
rect 15009 18320 18755 18322
rect 15009 18264 15014 18320
rect 15070 18264 18694 18320
rect 18750 18264 18755 18320
rect 15009 18262 18755 18264
rect 15009 18259 15075 18262
rect 18689 18259 18755 18262
rect 3556 17984 3872 17985
rect 3556 17920 3562 17984
rect 3626 17920 3642 17984
rect 3706 17920 3722 17984
rect 3786 17920 3802 17984
rect 3866 17920 3872 17984
rect 3556 17919 3872 17920
rect 8777 17984 9093 17985
rect 8777 17920 8783 17984
rect 8847 17920 8863 17984
rect 8927 17920 8943 17984
rect 9007 17920 9023 17984
rect 9087 17920 9093 17984
rect 8777 17919 9093 17920
rect 13998 17984 14314 17985
rect 13998 17920 14004 17984
rect 14068 17920 14084 17984
rect 14148 17920 14164 17984
rect 14228 17920 14244 17984
rect 14308 17920 14314 17984
rect 13998 17919 14314 17920
rect 19219 17984 19535 17985
rect 19219 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19465 17984
rect 19529 17920 19535 17984
rect 19219 17919 19535 17920
rect 0 17778 800 17808
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17688 800 17718
rect 2773 17715 2839 17718
rect 17953 17778 18019 17781
rect 22331 17778 23131 17808
rect 17953 17776 23131 17778
rect 17953 17720 17958 17776
rect 18014 17720 23131 17776
rect 17953 17718 23131 17720
rect 17953 17715 18019 17718
rect 22331 17688 23131 17718
rect 4216 17440 4532 17441
rect 4216 17376 4222 17440
rect 4286 17376 4302 17440
rect 4366 17376 4382 17440
rect 4446 17376 4462 17440
rect 4526 17376 4532 17440
rect 4216 17375 4532 17376
rect 9437 17440 9753 17441
rect 9437 17376 9443 17440
rect 9507 17376 9523 17440
rect 9587 17376 9603 17440
rect 9667 17376 9683 17440
rect 9747 17376 9753 17440
rect 9437 17375 9753 17376
rect 14658 17440 14974 17441
rect 14658 17376 14664 17440
rect 14728 17376 14744 17440
rect 14808 17376 14824 17440
rect 14888 17376 14904 17440
rect 14968 17376 14974 17440
rect 14658 17375 14974 17376
rect 19879 17440 20195 17441
rect 19879 17376 19885 17440
rect 19949 17376 19965 17440
rect 20029 17376 20045 17440
rect 20109 17376 20125 17440
rect 20189 17376 20195 17440
rect 19879 17375 20195 17376
rect 3049 17234 3115 17237
rect 8017 17234 8083 17237
rect 8518 17234 8524 17236
rect 3049 17232 8524 17234
rect 3049 17176 3054 17232
rect 3110 17176 8022 17232
rect 8078 17176 8524 17232
rect 3049 17174 8524 17176
rect 3049 17171 3115 17174
rect 8017 17171 8083 17174
rect 8518 17172 8524 17174
rect 8588 17234 8594 17236
rect 14406 17234 14412 17236
rect 8588 17174 14412 17234
rect 8588 17172 8594 17174
rect 14406 17172 14412 17174
rect 14476 17234 14482 17236
rect 15009 17234 15075 17237
rect 14476 17232 15075 17234
rect 14476 17176 15014 17232
rect 15070 17176 15075 17232
rect 14476 17174 15075 17176
rect 14476 17172 14482 17174
rect 15009 17171 15075 17174
rect 0 17098 800 17128
rect 5349 17098 5415 17101
rect 0 17096 5415 17098
rect 0 17040 5354 17096
rect 5410 17040 5415 17096
rect 0 17038 5415 17040
rect 0 17008 800 17038
rect 5349 17035 5415 17038
rect 21265 17098 21331 17101
rect 22331 17098 23131 17128
rect 21265 17096 23131 17098
rect 21265 17040 21270 17096
rect 21326 17040 23131 17096
rect 21265 17038 23131 17040
rect 21265 17035 21331 17038
rect 22331 17008 23131 17038
rect 3556 16896 3872 16897
rect 3556 16832 3562 16896
rect 3626 16832 3642 16896
rect 3706 16832 3722 16896
rect 3786 16832 3802 16896
rect 3866 16832 3872 16896
rect 3556 16831 3872 16832
rect 8777 16896 9093 16897
rect 8777 16832 8783 16896
rect 8847 16832 8863 16896
rect 8927 16832 8943 16896
rect 9007 16832 9023 16896
rect 9087 16832 9093 16896
rect 8777 16831 9093 16832
rect 13998 16896 14314 16897
rect 13998 16832 14004 16896
rect 14068 16832 14084 16896
rect 14148 16832 14164 16896
rect 14228 16832 14244 16896
rect 14308 16832 14314 16896
rect 13998 16831 14314 16832
rect 19219 16896 19535 16897
rect 19219 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19465 16896
rect 19529 16832 19535 16896
rect 19219 16831 19535 16832
rect 4889 16554 4955 16557
rect 2730 16552 4955 16554
rect 2730 16496 4894 16552
rect 4950 16496 4955 16552
rect 2730 16494 4955 16496
rect 0 16418 800 16448
rect 2730 16418 2790 16494
rect 4889 16491 4955 16494
rect 17217 16554 17283 16557
rect 17217 16552 20362 16554
rect 17217 16496 17222 16552
rect 17278 16496 20362 16552
rect 17217 16494 20362 16496
rect 17217 16491 17283 16494
rect 0 16358 2790 16418
rect 20302 16418 20362 16494
rect 22331 16418 23131 16448
rect 20302 16358 23131 16418
rect 0 16328 800 16358
rect 4216 16352 4532 16353
rect 4216 16288 4222 16352
rect 4286 16288 4302 16352
rect 4366 16288 4382 16352
rect 4446 16288 4462 16352
rect 4526 16288 4532 16352
rect 4216 16287 4532 16288
rect 9437 16352 9753 16353
rect 9437 16288 9443 16352
rect 9507 16288 9523 16352
rect 9587 16288 9603 16352
rect 9667 16288 9683 16352
rect 9747 16288 9753 16352
rect 9437 16287 9753 16288
rect 14658 16352 14974 16353
rect 14658 16288 14664 16352
rect 14728 16288 14744 16352
rect 14808 16288 14824 16352
rect 14888 16288 14904 16352
rect 14968 16288 14974 16352
rect 14658 16287 14974 16288
rect 19879 16352 20195 16353
rect 19879 16288 19885 16352
rect 19949 16288 19965 16352
rect 20029 16288 20045 16352
rect 20109 16288 20125 16352
rect 20189 16288 20195 16352
rect 22331 16328 23131 16358
rect 19879 16287 20195 16288
rect 14457 16146 14523 16149
rect 17718 16146 17724 16148
rect 14457 16144 17724 16146
rect 14457 16088 14462 16144
rect 14518 16088 17724 16144
rect 14457 16086 17724 16088
rect 14457 16083 14523 16086
rect 17718 16084 17724 16086
rect 17788 16084 17794 16148
rect 3556 15808 3872 15809
rect 0 15738 800 15768
rect 3556 15744 3562 15808
rect 3626 15744 3642 15808
rect 3706 15744 3722 15808
rect 3786 15744 3802 15808
rect 3866 15744 3872 15808
rect 3556 15743 3872 15744
rect 8777 15808 9093 15809
rect 8777 15744 8783 15808
rect 8847 15744 8863 15808
rect 8927 15744 8943 15808
rect 9007 15744 9023 15808
rect 9087 15744 9093 15808
rect 8777 15743 9093 15744
rect 13998 15808 14314 15809
rect 13998 15744 14004 15808
rect 14068 15744 14084 15808
rect 14148 15744 14164 15808
rect 14228 15744 14244 15808
rect 14308 15744 14314 15808
rect 13998 15743 14314 15744
rect 19219 15808 19535 15809
rect 19219 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19465 15808
rect 19529 15744 19535 15808
rect 19219 15743 19535 15744
rect 3141 15738 3207 15741
rect 22331 15738 23131 15768
rect 0 15736 3207 15738
rect 0 15680 3146 15736
rect 3202 15680 3207 15736
rect 0 15678 3207 15680
rect 0 15648 800 15678
rect 3141 15675 3207 15678
rect 19750 15678 23131 15738
rect 17953 15602 18019 15605
rect 19750 15602 19810 15678
rect 22331 15648 23131 15678
rect 17953 15600 19810 15602
rect 17953 15544 17958 15600
rect 18014 15544 19810 15600
rect 17953 15542 19810 15544
rect 17953 15539 18019 15542
rect 4216 15264 4532 15265
rect 4216 15200 4222 15264
rect 4286 15200 4302 15264
rect 4366 15200 4382 15264
rect 4446 15200 4462 15264
rect 4526 15200 4532 15264
rect 4216 15199 4532 15200
rect 9437 15264 9753 15265
rect 9437 15200 9443 15264
rect 9507 15200 9523 15264
rect 9587 15200 9603 15264
rect 9667 15200 9683 15264
rect 9747 15200 9753 15264
rect 9437 15199 9753 15200
rect 14658 15264 14974 15265
rect 14658 15200 14664 15264
rect 14728 15200 14744 15264
rect 14808 15200 14824 15264
rect 14888 15200 14904 15264
rect 14968 15200 14974 15264
rect 14658 15199 14974 15200
rect 19879 15264 20195 15265
rect 19879 15200 19885 15264
rect 19949 15200 19965 15264
rect 20029 15200 20045 15264
rect 20109 15200 20125 15264
rect 20189 15200 20195 15264
rect 19879 15199 20195 15200
rect 0 15058 800 15088
rect 5901 15058 5967 15061
rect 0 15056 5967 15058
rect 0 15000 5906 15056
rect 5962 15000 5967 15056
rect 0 14998 5967 15000
rect 0 14968 800 14998
rect 5901 14995 5967 14998
rect 20713 15058 20779 15061
rect 22331 15058 23131 15088
rect 20713 15056 23131 15058
rect 20713 15000 20718 15056
rect 20774 15000 23131 15056
rect 20713 14998 23131 15000
rect 20713 14995 20779 14998
rect 22331 14968 23131 14998
rect 3556 14720 3872 14721
rect 3556 14656 3562 14720
rect 3626 14656 3642 14720
rect 3706 14656 3722 14720
rect 3786 14656 3802 14720
rect 3866 14656 3872 14720
rect 3556 14655 3872 14656
rect 8777 14720 9093 14721
rect 8777 14656 8783 14720
rect 8847 14656 8863 14720
rect 8927 14656 8943 14720
rect 9007 14656 9023 14720
rect 9087 14656 9093 14720
rect 8777 14655 9093 14656
rect 13998 14720 14314 14721
rect 13998 14656 14004 14720
rect 14068 14656 14084 14720
rect 14148 14656 14164 14720
rect 14228 14656 14244 14720
rect 14308 14656 14314 14720
rect 13998 14655 14314 14656
rect 19219 14720 19535 14721
rect 19219 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19465 14720
rect 19529 14656 19535 14720
rect 19219 14655 19535 14656
rect 19517 14514 19583 14517
rect 21449 14514 21515 14517
rect 19517 14512 21515 14514
rect 19517 14456 19522 14512
rect 19578 14456 21454 14512
rect 21510 14456 21515 14512
rect 19517 14454 21515 14456
rect 19517 14451 19583 14454
rect 21449 14451 21515 14454
rect 0 14378 800 14408
rect 5441 14378 5507 14381
rect 0 14376 5507 14378
rect 0 14320 5446 14376
rect 5502 14320 5507 14376
rect 0 14318 5507 14320
rect 0 14288 800 14318
rect 5441 14315 5507 14318
rect 21357 14378 21423 14381
rect 22331 14378 23131 14408
rect 21357 14376 23131 14378
rect 21357 14320 21362 14376
rect 21418 14320 23131 14376
rect 21357 14318 23131 14320
rect 21357 14315 21423 14318
rect 22331 14288 23131 14318
rect 4216 14176 4532 14177
rect 4216 14112 4222 14176
rect 4286 14112 4302 14176
rect 4366 14112 4382 14176
rect 4446 14112 4462 14176
rect 4526 14112 4532 14176
rect 4216 14111 4532 14112
rect 9437 14176 9753 14177
rect 9437 14112 9443 14176
rect 9507 14112 9523 14176
rect 9587 14112 9603 14176
rect 9667 14112 9683 14176
rect 9747 14112 9753 14176
rect 9437 14111 9753 14112
rect 14658 14176 14974 14177
rect 14658 14112 14664 14176
rect 14728 14112 14744 14176
rect 14808 14112 14824 14176
rect 14888 14112 14904 14176
rect 14968 14112 14974 14176
rect 14658 14111 14974 14112
rect 19879 14176 20195 14177
rect 19879 14112 19885 14176
rect 19949 14112 19965 14176
rect 20029 14112 20045 14176
rect 20109 14112 20125 14176
rect 20189 14112 20195 14176
rect 19879 14111 20195 14112
rect 9857 13970 9923 13973
rect 13537 13970 13603 13973
rect 14825 13970 14891 13973
rect 18781 13970 18847 13973
rect 9857 13968 18847 13970
rect 9857 13912 9862 13968
rect 9918 13912 13542 13968
rect 13598 13912 14830 13968
rect 14886 13912 18786 13968
rect 18842 13912 18847 13968
rect 9857 13910 18847 13912
rect 9857 13907 9923 13910
rect 13537 13907 13603 13910
rect 14825 13907 14891 13910
rect 18781 13907 18847 13910
rect 0 13698 800 13728
rect 21541 13698 21607 13701
rect 22331 13698 23131 13728
rect 0 13638 2790 13698
rect 0 13608 800 13638
rect 2730 13426 2790 13638
rect 21541 13696 23131 13698
rect 21541 13640 21546 13696
rect 21602 13640 23131 13696
rect 21541 13638 23131 13640
rect 21541 13635 21607 13638
rect 3556 13632 3872 13633
rect 3556 13568 3562 13632
rect 3626 13568 3642 13632
rect 3706 13568 3722 13632
rect 3786 13568 3802 13632
rect 3866 13568 3872 13632
rect 3556 13567 3872 13568
rect 8777 13632 9093 13633
rect 8777 13568 8783 13632
rect 8847 13568 8863 13632
rect 8927 13568 8943 13632
rect 9007 13568 9023 13632
rect 9087 13568 9093 13632
rect 8777 13567 9093 13568
rect 13998 13632 14314 13633
rect 13998 13568 14004 13632
rect 14068 13568 14084 13632
rect 14148 13568 14164 13632
rect 14228 13568 14244 13632
rect 14308 13568 14314 13632
rect 13998 13567 14314 13568
rect 19219 13632 19535 13633
rect 19219 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19465 13632
rect 19529 13568 19535 13632
rect 22331 13608 23131 13638
rect 19219 13567 19535 13568
rect 6453 13426 6519 13429
rect 2730 13424 6519 13426
rect 2730 13368 6458 13424
rect 6514 13368 6519 13424
rect 2730 13366 6519 13368
rect 6453 13363 6519 13366
rect 4216 13088 4532 13089
rect 0 13018 800 13048
rect 4216 13024 4222 13088
rect 4286 13024 4302 13088
rect 4366 13024 4382 13088
rect 4446 13024 4462 13088
rect 4526 13024 4532 13088
rect 4216 13023 4532 13024
rect 9437 13088 9753 13089
rect 9437 13024 9443 13088
rect 9507 13024 9523 13088
rect 9587 13024 9603 13088
rect 9667 13024 9683 13088
rect 9747 13024 9753 13088
rect 9437 13023 9753 13024
rect 14658 13088 14974 13089
rect 14658 13024 14664 13088
rect 14728 13024 14744 13088
rect 14808 13024 14824 13088
rect 14888 13024 14904 13088
rect 14968 13024 14974 13088
rect 14658 13023 14974 13024
rect 19879 13088 20195 13089
rect 19879 13024 19885 13088
rect 19949 13024 19965 13088
rect 20029 13024 20045 13088
rect 20109 13024 20125 13088
rect 20189 13024 20195 13088
rect 19879 13023 20195 13024
rect 2865 13018 2931 13021
rect 22331 13018 23131 13048
rect 0 13016 2931 13018
rect 0 12960 2870 13016
rect 2926 12960 2931 13016
rect 0 12958 2931 12960
rect 0 12928 800 12958
rect 2865 12955 2931 12958
rect 20302 12958 23131 13018
rect 16481 12882 16547 12885
rect 20302 12882 20362 12958
rect 22331 12928 23131 12958
rect 16481 12880 20362 12882
rect 16481 12824 16486 12880
rect 16542 12824 20362 12880
rect 16481 12822 20362 12824
rect 16481 12819 16547 12822
rect 3556 12544 3872 12545
rect 3556 12480 3562 12544
rect 3626 12480 3642 12544
rect 3706 12480 3722 12544
rect 3786 12480 3802 12544
rect 3866 12480 3872 12544
rect 3556 12479 3872 12480
rect 8777 12544 9093 12545
rect 8777 12480 8783 12544
rect 8847 12480 8863 12544
rect 8927 12480 8943 12544
rect 9007 12480 9023 12544
rect 9087 12480 9093 12544
rect 8777 12479 9093 12480
rect 13998 12544 14314 12545
rect 13998 12480 14004 12544
rect 14068 12480 14084 12544
rect 14148 12480 14164 12544
rect 14228 12480 14244 12544
rect 14308 12480 14314 12544
rect 13998 12479 14314 12480
rect 19219 12544 19535 12545
rect 19219 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19465 12544
rect 19529 12480 19535 12544
rect 19219 12479 19535 12480
rect 0 12338 800 12368
rect 2773 12338 2839 12341
rect 0 12336 2839 12338
rect 0 12280 2778 12336
rect 2834 12280 2839 12336
rect 0 12278 2839 12280
rect 0 12248 800 12278
rect 2773 12275 2839 12278
rect 2998 12276 3004 12340
rect 3068 12338 3074 12340
rect 11513 12338 11579 12341
rect 3068 12336 11579 12338
rect 3068 12280 11518 12336
rect 11574 12280 11579 12336
rect 3068 12278 11579 12280
rect 3068 12276 3074 12278
rect 11513 12275 11579 12278
rect 13261 12338 13327 12341
rect 14406 12338 14412 12340
rect 13261 12336 14412 12338
rect 13261 12280 13266 12336
rect 13322 12280 14412 12336
rect 13261 12278 14412 12280
rect 13261 12275 13327 12278
rect 14406 12276 14412 12278
rect 14476 12276 14482 12340
rect 18597 12338 18663 12341
rect 22331 12338 23131 12368
rect 18597 12336 23131 12338
rect 18597 12280 18602 12336
rect 18658 12280 23131 12336
rect 18597 12278 23131 12280
rect 18597 12275 18663 12278
rect 22331 12248 23131 12278
rect 4216 12000 4532 12001
rect 4216 11936 4222 12000
rect 4286 11936 4302 12000
rect 4366 11936 4382 12000
rect 4446 11936 4462 12000
rect 4526 11936 4532 12000
rect 4216 11935 4532 11936
rect 9437 12000 9753 12001
rect 9437 11936 9443 12000
rect 9507 11936 9523 12000
rect 9587 11936 9603 12000
rect 9667 11936 9683 12000
rect 9747 11936 9753 12000
rect 9437 11935 9753 11936
rect 14658 12000 14974 12001
rect 14658 11936 14664 12000
rect 14728 11936 14744 12000
rect 14808 11936 14824 12000
rect 14888 11936 14904 12000
rect 14968 11936 14974 12000
rect 14658 11935 14974 11936
rect 19879 12000 20195 12001
rect 19879 11936 19885 12000
rect 19949 11936 19965 12000
rect 20029 11936 20045 12000
rect 20109 11936 20125 12000
rect 20189 11936 20195 12000
rect 19879 11935 20195 11936
rect 0 11658 800 11688
rect 3233 11658 3299 11661
rect 0 11656 3299 11658
rect 0 11600 3238 11656
rect 3294 11600 3299 11656
rect 0 11598 3299 11600
rect 0 11568 800 11598
rect 3233 11595 3299 11598
rect 21357 11658 21423 11661
rect 22331 11658 23131 11688
rect 21357 11656 23131 11658
rect 21357 11600 21362 11656
rect 21418 11600 23131 11656
rect 21357 11598 23131 11600
rect 21357 11595 21423 11598
rect 22331 11568 23131 11598
rect 3556 11456 3872 11457
rect 3556 11392 3562 11456
rect 3626 11392 3642 11456
rect 3706 11392 3722 11456
rect 3786 11392 3802 11456
rect 3866 11392 3872 11456
rect 3556 11391 3872 11392
rect 8777 11456 9093 11457
rect 8777 11392 8783 11456
rect 8847 11392 8863 11456
rect 8927 11392 8943 11456
rect 9007 11392 9023 11456
rect 9087 11392 9093 11456
rect 8777 11391 9093 11392
rect 13998 11456 14314 11457
rect 13998 11392 14004 11456
rect 14068 11392 14084 11456
rect 14148 11392 14164 11456
rect 14228 11392 14244 11456
rect 14308 11392 14314 11456
rect 13998 11391 14314 11392
rect 19219 11456 19535 11457
rect 19219 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19465 11456
rect 19529 11392 19535 11456
rect 19219 11391 19535 11392
rect 0 10978 800 11008
rect 4061 10978 4127 10981
rect 22331 10978 23131 11008
rect 0 10976 4127 10978
rect 0 10920 4066 10976
rect 4122 10920 4127 10976
rect 0 10918 4127 10920
rect 0 10888 800 10918
rect 4061 10915 4127 10918
rect 20302 10918 23131 10978
rect 4216 10912 4532 10913
rect 4216 10848 4222 10912
rect 4286 10848 4302 10912
rect 4366 10848 4382 10912
rect 4446 10848 4462 10912
rect 4526 10848 4532 10912
rect 4216 10847 4532 10848
rect 9437 10912 9753 10913
rect 9437 10848 9443 10912
rect 9507 10848 9523 10912
rect 9587 10848 9603 10912
rect 9667 10848 9683 10912
rect 9747 10848 9753 10912
rect 9437 10847 9753 10848
rect 14658 10912 14974 10913
rect 14658 10848 14664 10912
rect 14728 10848 14744 10912
rect 14808 10848 14824 10912
rect 14888 10848 14904 10912
rect 14968 10848 14974 10912
rect 14658 10847 14974 10848
rect 19879 10912 20195 10913
rect 19879 10848 19885 10912
rect 19949 10848 19965 10912
rect 20029 10848 20045 10912
rect 20109 10848 20125 10912
rect 20189 10848 20195 10912
rect 19879 10847 20195 10848
rect 17217 10706 17283 10709
rect 20302 10706 20362 10918
rect 22331 10888 23131 10918
rect 17217 10704 20362 10706
rect 17217 10648 17222 10704
rect 17278 10648 20362 10704
rect 17217 10646 20362 10648
rect 17217 10643 17283 10646
rect 3556 10368 3872 10369
rect 0 10298 800 10328
rect 3556 10304 3562 10368
rect 3626 10304 3642 10368
rect 3706 10304 3722 10368
rect 3786 10304 3802 10368
rect 3866 10304 3872 10368
rect 3556 10303 3872 10304
rect 8777 10368 9093 10369
rect 8777 10304 8783 10368
rect 8847 10304 8863 10368
rect 8927 10304 8943 10368
rect 9007 10304 9023 10368
rect 9087 10304 9093 10368
rect 8777 10303 9093 10304
rect 13998 10368 14314 10369
rect 13998 10304 14004 10368
rect 14068 10304 14084 10368
rect 14148 10304 14164 10368
rect 14228 10304 14244 10368
rect 14308 10304 14314 10368
rect 13998 10303 14314 10304
rect 19219 10368 19535 10369
rect 19219 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19465 10368
rect 19529 10304 19535 10368
rect 19219 10303 19535 10304
rect 1301 10298 1367 10301
rect 22331 10298 23131 10328
rect 0 10296 1367 10298
rect 0 10240 1306 10296
rect 1362 10240 1367 10296
rect 0 10238 1367 10240
rect 0 10208 800 10238
rect 1301 10235 1367 10238
rect 19750 10238 23131 10298
rect 18045 10162 18111 10165
rect 19750 10162 19810 10238
rect 22331 10208 23131 10238
rect 18045 10160 19810 10162
rect 18045 10104 18050 10160
rect 18106 10104 19810 10160
rect 18045 10102 19810 10104
rect 18045 10099 18111 10102
rect 4216 9824 4532 9825
rect 4216 9760 4222 9824
rect 4286 9760 4302 9824
rect 4366 9760 4382 9824
rect 4446 9760 4462 9824
rect 4526 9760 4532 9824
rect 4216 9759 4532 9760
rect 9437 9824 9753 9825
rect 9437 9760 9443 9824
rect 9507 9760 9523 9824
rect 9587 9760 9603 9824
rect 9667 9760 9683 9824
rect 9747 9760 9753 9824
rect 9437 9759 9753 9760
rect 14658 9824 14974 9825
rect 14658 9760 14664 9824
rect 14728 9760 14744 9824
rect 14808 9760 14824 9824
rect 14888 9760 14904 9824
rect 14968 9760 14974 9824
rect 14658 9759 14974 9760
rect 19879 9824 20195 9825
rect 19879 9760 19885 9824
rect 19949 9760 19965 9824
rect 20029 9760 20045 9824
rect 20109 9760 20125 9824
rect 20189 9760 20195 9824
rect 19879 9759 20195 9760
rect 0 9618 800 9648
rect 3877 9618 3943 9621
rect 0 9616 3943 9618
rect 0 9560 3882 9616
rect 3938 9560 3943 9616
rect 0 9558 3943 9560
rect 0 9528 800 9558
rect 3877 9555 3943 9558
rect 21357 9618 21423 9621
rect 22331 9618 23131 9648
rect 21357 9616 23131 9618
rect 21357 9560 21362 9616
rect 21418 9560 23131 9616
rect 21357 9558 23131 9560
rect 21357 9555 21423 9558
rect 22331 9528 23131 9558
rect 3556 9280 3872 9281
rect 3556 9216 3562 9280
rect 3626 9216 3642 9280
rect 3706 9216 3722 9280
rect 3786 9216 3802 9280
rect 3866 9216 3872 9280
rect 3556 9215 3872 9216
rect 8777 9280 9093 9281
rect 8777 9216 8783 9280
rect 8847 9216 8863 9280
rect 8927 9216 8943 9280
rect 9007 9216 9023 9280
rect 9087 9216 9093 9280
rect 8777 9215 9093 9216
rect 13998 9280 14314 9281
rect 13998 9216 14004 9280
rect 14068 9216 14084 9280
rect 14148 9216 14164 9280
rect 14228 9216 14244 9280
rect 14308 9216 14314 9280
rect 13998 9215 14314 9216
rect 19219 9280 19535 9281
rect 19219 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19465 9280
rect 19529 9216 19535 9280
rect 19219 9215 19535 9216
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 20805 8938 20871 8941
rect 22331 8938 23131 8968
rect 20805 8936 23131 8938
rect 20805 8880 20810 8936
rect 20866 8880 23131 8936
rect 20805 8878 23131 8880
rect 20805 8875 20871 8878
rect 22331 8848 23131 8878
rect 4216 8736 4532 8737
rect 4216 8672 4222 8736
rect 4286 8672 4302 8736
rect 4366 8672 4382 8736
rect 4446 8672 4462 8736
rect 4526 8672 4532 8736
rect 4216 8671 4532 8672
rect 9437 8736 9753 8737
rect 9437 8672 9443 8736
rect 9507 8672 9523 8736
rect 9587 8672 9603 8736
rect 9667 8672 9683 8736
rect 9747 8672 9753 8736
rect 9437 8671 9753 8672
rect 14658 8736 14974 8737
rect 14658 8672 14664 8736
rect 14728 8672 14744 8736
rect 14808 8672 14824 8736
rect 14888 8672 14904 8736
rect 14968 8672 14974 8736
rect 14658 8671 14974 8672
rect 19879 8736 20195 8737
rect 19879 8672 19885 8736
rect 19949 8672 19965 8736
rect 20029 8672 20045 8736
rect 20109 8672 20125 8736
rect 20189 8672 20195 8736
rect 19879 8671 20195 8672
rect 14457 8532 14523 8533
rect 14406 8468 14412 8532
rect 14476 8530 14523 8532
rect 18137 8530 18203 8533
rect 14476 8528 18203 8530
rect 14518 8472 18142 8528
rect 18198 8472 18203 8528
rect 14476 8470 18203 8472
rect 14476 8468 14523 8470
rect 14457 8467 14523 8468
rect 18137 8467 18203 8470
rect 0 8258 800 8288
rect 20621 8258 20687 8261
rect 22331 8258 23131 8288
rect 0 8198 2514 8258
rect 0 8168 800 8198
rect 2454 7986 2514 8198
rect 20621 8256 23131 8258
rect 20621 8200 20626 8256
rect 20682 8200 23131 8256
rect 20621 8198 23131 8200
rect 20621 8195 20687 8198
rect 3556 8192 3872 8193
rect 3556 8128 3562 8192
rect 3626 8128 3642 8192
rect 3706 8128 3722 8192
rect 3786 8128 3802 8192
rect 3866 8128 3872 8192
rect 3556 8127 3872 8128
rect 8777 8192 9093 8193
rect 8777 8128 8783 8192
rect 8847 8128 8863 8192
rect 8927 8128 8943 8192
rect 9007 8128 9023 8192
rect 9087 8128 9093 8192
rect 8777 8127 9093 8128
rect 13998 8192 14314 8193
rect 13998 8128 14004 8192
rect 14068 8128 14084 8192
rect 14148 8128 14164 8192
rect 14228 8128 14244 8192
rect 14308 8128 14314 8192
rect 13998 8127 14314 8128
rect 19219 8192 19535 8193
rect 19219 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19465 8192
rect 19529 8128 19535 8192
rect 22331 8168 23131 8198
rect 19219 8127 19535 8128
rect 4889 7986 4955 7989
rect 2454 7984 4955 7986
rect 2454 7928 4894 7984
rect 4950 7928 4955 7984
rect 2454 7926 4955 7928
rect 4889 7923 4955 7926
rect 4216 7648 4532 7649
rect 0 7578 800 7608
rect 4216 7584 4222 7648
rect 4286 7584 4302 7648
rect 4366 7584 4382 7648
rect 4446 7584 4462 7648
rect 4526 7584 4532 7648
rect 4216 7583 4532 7584
rect 9437 7648 9753 7649
rect 9437 7584 9443 7648
rect 9507 7584 9523 7648
rect 9587 7584 9603 7648
rect 9667 7584 9683 7648
rect 9747 7584 9753 7648
rect 9437 7583 9753 7584
rect 14658 7648 14974 7649
rect 14658 7584 14664 7648
rect 14728 7584 14744 7648
rect 14808 7584 14824 7648
rect 14888 7584 14904 7648
rect 14968 7584 14974 7648
rect 14658 7583 14974 7584
rect 19879 7648 20195 7649
rect 19879 7584 19885 7648
rect 19949 7584 19965 7648
rect 20029 7584 20045 7648
rect 20109 7584 20125 7648
rect 20189 7584 20195 7648
rect 19879 7583 20195 7584
rect 3785 7578 3851 7581
rect 22331 7578 23131 7608
rect 0 7576 3851 7578
rect 0 7520 3790 7576
rect 3846 7520 3851 7576
rect 0 7518 3851 7520
rect 0 7488 800 7518
rect 3785 7515 3851 7518
rect 20302 7518 23131 7578
rect 2773 7442 2839 7445
rect 3877 7442 3943 7445
rect 9213 7442 9279 7445
rect 2773 7440 9279 7442
rect 2773 7384 2778 7440
rect 2834 7384 3882 7440
rect 3938 7384 9218 7440
rect 9274 7384 9279 7440
rect 2773 7382 9279 7384
rect 2773 7379 2839 7382
rect 3877 7379 3943 7382
rect 9213 7379 9279 7382
rect 17033 7442 17099 7445
rect 20302 7442 20362 7518
rect 22331 7488 23131 7518
rect 17033 7440 20362 7442
rect 17033 7384 17038 7440
rect 17094 7384 20362 7440
rect 17033 7382 20362 7384
rect 17033 7379 17099 7382
rect 3556 7104 3872 7105
rect 3556 7040 3562 7104
rect 3626 7040 3642 7104
rect 3706 7040 3722 7104
rect 3786 7040 3802 7104
rect 3866 7040 3872 7104
rect 3556 7039 3872 7040
rect 8777 7104 9093 7105
rect 8777 7040 8783 7104
rect 8847 7040 8863 7104
rect 8927 7040 8943 7104
rect 9007 7040 9023 7104
rect 9087 7040 9093 7104
rect 8777 7039 9093 7040
rect 13998 7104 14314 7105
rect 13998 7040 14004 7104
rect 14068 7040 14084 7104
rect 14148 7040 14164 7104
rect 14228 7040 14244 7104
rect 14308 7040 14314 7104
rect 13998 7039 14314 7040
rect 19219 7104 19535 7105
rect 19219 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19465 7104
rect 19529 7040 19535 7104
rect 19219 7039 19535 7040
rect 9213 7034 9279 7037
rect 9949 7034 10015 7037
rect 9213 7032 10015 7034
rect 9213 6976 9218 7032
rect 9274 6976 9954 7032
rect 10010 6976 10015 7032
rect 9213 6974 10015 6976
rect 9213 6971 9279 6974
rect 9949 6971 10015 6974
rect 0 6898 800 6928
rect 1117 6898 1183 6901
rect 0 6896 1183 6898
rect 0 6840 1122 6896
rect 1178 6840 1183 6896
rect 0 6838 1183 6840
rect 0 6808 800 6838
rect 1117 6835 1183 6838
rect 21357 6898 21423 6901
rect 22331 6898 23131 6928
rect 21357 6896 23131 6898
rect 21357 6840 21362 6896
rect 21418 6840 23131 6896
rect 21357 6838 23131 6840
rect 21357 6835 21423 6838
rect 22331 6808 23131 6838
rect 4216 6560 4532 6561
rect 4216 6496 4222 6560
rect 4286 6496 4302 6560
rect 4366 6496 4382 6560
rect 4446 6496 4462 6560
rect 4526 6496 4532 6560
rect 4216 6495 4532 6496
rect 9437 6560 9753 6561
rect 9437 6496 9443 6560
rect 9507 6496 9523 6560
rect 9587 6496 9603 6560
rect 9667 6496 9683 6560
rect 9747 6496 9753 6560
rect 9437 6495 9753 6496
rect 14658 6560 14974 6561
rect 14658 6496 14664 6560
rect 14728 6496 14744 6560
rect 14808 6496 14824 6560
rect 14888 6496 14904 6560
rect 14968 6496 14974 6560
rect 14658 6495 14974 6496
rect 19879 6560 20195 6561
rect 19879 6496 19885 6560
rect 19949 6496 19965 6560
rect 20029 6496 20045 6560
rect 20109 6496 20125 6560
rect 20189 6496 20195 6560
rect 19879 6495 20195 6496
rect 13445 6490 13511 6493
rect 14406 6490 14412 6492
rect 13445 6488 14412 6490
rect 13445 6432 13450 6488
rect 13506 6432 14412 6488
rect 13445 6430 14412 6432
rect 13445 6427 13511 6430
rect 14406 6428 14412 6430
rect 14476 6428 14482 6492
rect 10961 6354 11027 6357
rect 18045 6354 18111 6357
rect 10961 6352 18111 6354
rect 10961 6296 10966 6352
rect 11022 6296 18050 6352
rect 18106 6296 18111 6352
rect 10961 6294 18111 6296
rect 10961 6291 11027 6294
rect 18045 6291 18111 6294
rect 0 6218 800 6248
rect 2957 6218 3023 6221
rect 0 6216 3023 6218
rect 0 6160 2962 6216
rect 3018 6160 3023 6216
rect 0 6158 3023 6160
rect 0 6128 800 6158
rect 2957 6155 3023 6158
rect 9949 6218 10015 6221
rect 13445 6218 13511 6221
rect 9949 6216 13511 6218
rect 9949 6160 9954 6216
rect 10010 6160 13450 6216
rect 13506 6160 13511 6216
rect 9949 6158 13511 6160
rect 9949 6155 10015 6158
rect 13445 6155 13511 6158
rect 21081 6218 21147 6221
rect 22331 6218 23131 6248
rect 21081 6216 23131 6218
rect 21081 6160 21086 6216
rect 21142 6160 23131 6216
rect 21081 6158 23131 6160
rect 21081 6155 21147 6158
rect 22331 6128 23131 6158
rect 3556 6016 3872 6017
rect 3556 5952 3562 6016
rect 3626 5952 3642 6016
rect 3706 5952 3722 6016
rect 3786 5952 3802 6016
rect 3866 5952 3872 6016
rect 3556 5951 3872 5952
rect 8777 6016 9093 6017
rect 8777 5952 8783 6016
rect 8847 5952 8863 6016
rect 8927 5952 8943 6016
rect 9007 5952 9023 6016
rect 9087 5952 9093 6016
rect 8777 5951 9093 5952
rect 13998 6016 14314 6017
rect 13998 5952 14004 6016
rect 14068 5952 14084 6016
rect 14148 5952 14164 6016
rect 14228 5952 14244 6016
rect 14308 5952 14314 6016
rect 13998 5951 14314 5952
rect 19219 6016 19535 6017
rect 19219 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19465 6016
rect 19529 5952 19535 6016
rect 19219 5951 19535 5952
rect 0 5538 800 5568
rect 3969 5538 4035 5541
rect 0 5536 4035 5538
rect 0 5480 3974 5536
rect 4030 5480 4035 5536
rect 0 5478 4035 5480
rect 0 5448 800 5478
rect 3969 5475 4035 5478
rect 20345 5538 20411 5541
rect 22331 5538 23131 5568
rect 20345 5536 23131 5538
rect 20345 5480 20350 5536
rect 20406 5480 23131 5536
rect 20345 5478 23131 5480
rect 20345 5475 20411 5478
rect 4216 5472 4532 5473
rect 4216 5408 4222 5472
rect 4286 5408 4302 5472
rect 4366 5408 4382 5472
rect 4446 5408 4462 5472
rect 4526 5408 4532 5472
rect 4216 5407 4532 5408
rect 9437 5472 9753 5473
rect 9437 5408 9443 5472
rect 9507 5408 9523 5472
rect 9587 5408 9603 5472
rect 9667 5408 9683 5472
rect 9747 5408 9753 5472
rect 9437 5407 9753 5408
rect 14658 5472 14974 5473
rect 14658 5408 14664 5472
rect 14728 5408 14744 5472
rect 14808 5408 14824 5472
rect 14888 5408 14904 5472
rect 14968 5408 14974 5472
rect 14658 5407 14974 5408
rect 19879 5472 20195 5473
rect 19879 5408 19885 5472
rect 19949 5408 19965 5472
rect 20029 5408 20045 5472
rect 20109 5408 20125 5472
rect 20189 5408 20195 5472
rect 22331 5448 23131 5478
rect 19879 5407 20195 5408
rect 3556 4928 3872 4929
rect 0 4858 800 4888
rect 3556 4864 3562 4928
rect 3626 4864 3642 4928
rect 3706 4864 3722 4928
rect 3786 4864 3802 4928
rect 3866 4864 3872 4928
rect 3556 4863 3872 4864
rect 8777 4928 9093 4929
rect 8777 4864 8783 4928
rect 8847 4864 8863 4928
rect 8927 4864 8943 4928
rect 9007 4864 9023 4928
rect 9087 4864 9093 4928
rect 8777 4863 9093 4864
rect 13998 4928 14314 4929
rect 13998 4864 14004 4928
rect 14068 4864 14084 4928
rect 14148 4864 14164 4928
rect 14228 4864 14244 4928
rect 14308 4864 14314 4928
rect 13998 4863 14314 4864
rect 19219 4928 19535 4929
rect 19219 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19465 4928
rect 19529 4864 19535 4928
rect 19219 4863 19535 4864
rect 3417 4858 3483 4861
rect 0 4856 3483 4858
rect 0 4800 3422 4856
rect 3478 4800 3483 4856
rect 0 4798 3483 4800
rect 0 4768 800 4798
rect 3417 4795 3483 4798
rect 21541 4858 21607 4861
rect 22331 4858 23131 4888
rect 21541 4856 23131 4858
rect 21541 4800 21546 4856
rect 21602 4800 23131 4856
rect 21541 4798 23131 4800
rect 21541 4795 21607 4798
rect 22331 4768 23131 4798
rect 4216 4384 4532 4385
rect 4216 4320 4222 4384
rect 4286 4320 4302 4384
rect 4366 4320 4382 4384
rect 4446 4320 4462 4384
rect 4526 4320 4532 4384
rect 4216 4319 4532 4320
rect 9437 4384 9753 4385
rect 9437 4320 9443 4384
rect 9507 4320 9523 4384
rect 9587 4320 9603 4384
rect 9667 4320 9683 4384
rect 9747 4320 9753 4384
rect 9437 4319 9753 4320
rect 14658 4384 14974 4385
rect 14658 4320 14664 4384
rect 14728 4320 14744 4384
rect 14808 4320 14824 4384
rect 14888 4320 14904 4384
rect 14968 4320 14974 4384
rect 14658 4319 14974 4320
rect 19879 4384 20195 4385
rect 19879 4320 19885 4384
rect 19949 4320 19965 4384
rect 20029 4320 20045 4384
rect 20109 4320 20125 4384
rect 20189 4320 20195 4384
rect 19879 4319 20195 4320
rect 0 4178 800 4208
rect 2773 4178 2839 4181
rect 0 4176 2839 4178
rect 0 4120 2778 4176
rect 2834 4120 2839 4176
rect 0 4118 2839 4120
rect 0 4088 800 4118
rect 2773 4115 2839 4118
rect 18413 4178 18479 4181
rect 22331 4178 23131 4208
rect 18413 4176 23131 4178
rect 18413 4120 18418 4176
rect 18474 4120 23131 4176
rect 18413 4118 23131 4120
rect 18413 4115 18479 4118
rect 22331 4088 23131 4118
rect 3556 3840 3872 3841
rect 3556 3776 3562 3840
rect 3626 3776 3642 3840
rect 3706 3776 3722 3840
rect 3786 3776 3802 3840
rect 3866 3776 3872 3840
rect 3556 3775 3872 3776
rect 8777 3840 9093 3841
rect 8777 3776 8783 3840
rect 8847 3776 8863 3840
rect 8927 3776 8943 3840
rect 9007 3776 9023 3840
rect 9087 3776 9093 3840
rect 8777 3775 9093 3776
rect 13998 3840 14314 3841
rect 13998 3776 14004 3840
rect 14068 3776 14084 3840
rect 14148 3776 14164 3840
rect 14228 3776 14244 3840
rect 14308 3776 14314 3840
rect 13998 3775 14314 3776
rect 19219 3840 19535 3841
rect 19219 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19465 3840
rect 19529 3776 19535 3840
rect 19219 3775 19535 3776
rect 0 3498 800 3528
rect 4981 3498 5047 3501
rect 0 3496 5047 3498
rect 0 3440 4986 3496
rect 5042 3440 5047 3496
rect 0 3438 5047 3440
rect 0 3408 800 3438
rect 4981 3435 5047 3438
rect 21357 3498 21423 3501
rect 22331 3498 23131 3528
rect 21357 3496 23131 3498
rect 21357 3440 21362 3496
rect 21418 3440 23131 3496
rect 21357 3438 23131 3440
rect 21357 3435 21423 3438
rect 22331 3408 23131 3438
rect 4216 3296 4532 3297
rect 4216 3232 4222 3296
rect 4286 3232 4302 3296
rect 4366 3232 4382 3296
rect 4446 3232 4462 3296
rect 4526 3232 4532 3296
rect 4216 3231 4532 3232
rect 9437 3296 9753 3297
rect 9437 3232 9443 3296
rect 9507 3232 9523 3296
rect 9587 3232 9603 3296
rect 9667 3232 9683 3296
rect 9747 3232 9753 3296
rect 9437 3231 9753 3232
rect 14658 3296 14974 3297
rect 14658 3232 14664 3296
rect 14728 3232 14744 3296
rect 14808 3232 14824 3296
rect 14888 3232 14904 3296
rect 14968 3232 14974 3296
rect 14658 3231 14974 3232
rect 19879 3296 20195 3297
rect 19879 3232 19885 3296
rect 19949 3232 19965 3296
rect 20029 3232 20045 3296
rect 20109 3232 20125 3296
rect 20189 3232 20195 3296
rect 19879 3231 20195 3232
rect 0 2818 800 2848
rect 2773 2818 2839 2821
rect 0 2816 2839 2818
rect 0 2760 2778 2816
rect 2834 2760 2839 2816
rect 0 2758 2839 2760
rect 0 2728 800 2758
rect 2773 2755 2839 2758
rect 3556 2752 3872 2753
rect 3556 2688 3562 2752
rect 3626 2688 3642 2752
rect 3706 2688 3722 2752
rect 3786 2688 3802 2752
rect 3866 2688 3872 2752
rect 3556 2687 3872 2688
rect 8777 2752 9093 2753
rect 8777 2688 8783 2752
rect 8847 2688 8863 2752
rect 8927 2688 8943 2752
rect 9007 2688 9023 2752
rect 9087 2688 9093 2752
rect 8777 2687 9093 2688
rect 13998 2752 14314 2753
rect 13998 2688 14004 2752
rect 14068 2688 14084 2752
rect 14148 2688 14164 2752
rect 14228 2688 14244 2752
rect 14308 2688 14314 2752
rect 13998 2687 14314 2688
rect 19219 2752 19535 2753
rect 19219 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19465 2752
rect 19529 2688 19535 2752
rect 19219 2687 19535 2688
rect 4216 2208 4532 2209
rect 0 2138 800 2168
rect 4216 2144 4222 2208
rect 4286 2144 4302 2208
rect 4366 2144 4382 2208
rect 4446 2144 4462 2208
rect 4526 2144 4532 2208
rect 4216 2143 4532 2144
rect 9437 2208 9753 2209
rect 9437 2144 9443 2208
rect 9507 2144 9523 2208
rect 9587 2144 9603 2208
rect 9667 2144 9683 2208
rect 9747 2144 9753 2208
rect 9437 2143 9753 2144
rect 14658 2208 14974 2209
rect 14658 2144 14664 2208
rect 14728 2144 14744 2208
rect 14808 2144 14824 2208
rect 14888 2144 14904 2208
rect 14968 2144 14974 2208
rect 14658 2143 14974 2144
rect 19879 2208 20195 2209
rect 19879 2144 19885 2208
rect 19949 2144 19965 2208
rect 20029 2144 20045 2208
rect 20109 2144 20125 2208
rect 20189 2144 20195 2208
rect 19879 2143 20195 2144
rect 2957 2138 3023 2141
rect 0 2136 3023 2138
rect 0 2080 2962 2136
rect 3018 2080 3023 2136
rect 0 2078 3023 2080
rect 0 2048 800 2078
rect 2957 2075 3023 2078
rect 0 1458 800 1488
rect 5165 1458 5231 1461
rect 0 1456 5231 1458
rect 0 1400 5170 1456
rect 5226 1400 5231 1456
rect 0 1398 5231 1400
rect 0 1368 800 1398
rect 5165 1395 5231 1398
rect 3417 914 3483 917
rect 1166 912 3483 914
rect 1166 856 3422 912
rect 3478 856 3483 912
rect 1166 854 3483 856
rect 0 778 800 808
rect 1166 778 1226 854
rect 3417 851 3483 854
rect 0 718 1226 778
rect 0 688 800 718
<< via3 >>
rect 4222 22876 4286 22880
rect 4222 22820 4226 22876
rect 4226 22820 4282 22876
rect 4282 22820 4286 22876
rect 4222 22816 4286 22820
rect 4302 22876 4366 22880
rect 4302 22820 4306 22876
rect 4306 22820 4362 22876
rect 4362 22820 4366 22876
rect 4302 22816 4366 22820
rect 4382 22876 4446 22880
rect 4382 22820 4386 22876
rect 4386 22820 4442 22876
rect 4442 22820 4446 22876
rect 4382 22816 4446 22820
rect 4462 22876 4526 22880
rect 4462 22820 4466 22876
rect 4466 22820 4522 22876
rect 4522 22820 4526 22876
rect 4462 22816 4526 22820
rect 9443 22876 9507 22880
rect 9443 22820 9447 22876
rect 9447 22820 9503 22876
rect 9503 22820 9507 22876
rect 9443 22816 9507 22820
rect 9523 22876 9587 22880
rect 9523 22820 9527 22876
rect 9527 22820 9583 22876
rect 9583 22820 9587 22876
rect 9523 22816 9587 22820
rect 9603 22876 9667 22880
rect 9603 22820 9607 22876
rect 9607 22820 9663 22876
rect 9663 22820 9667 22876
rect 9603 22816 9667 22820
rect 9683 22876 9747 22880
rect 9683 22820 9687 22876
rect 9687 22820 9743 22876
rect 9743 22820 9747 22876
rect 9683 22816 9747 22820
rect 14664 22876 14728 22880
rect 14664 22820 14668 22876
rect 14668 22820 14724 22876
rect 14724 22820 14728 22876
rect 14664 22816 14728 22820
rect 14744 22876 14808 22880
rect 14744 22820 14748 22876
rect 14748 22820 14804 22876
rect 14804 22820 14808 22876
rect 14744 22816 14808 22820
rect 14824 22876 14888 22880
rect 14824 22820 14828 22876
rect 14828 22820 14884 22876
rect 14884 22820 14888 22876
rect 14824 22816 14888 22820
rect 14904 22876 14968 22880
rect 14904 22820 14908 22876
rect 14908 22820 14964 22876
rect 14964 22820 14968 22876
rect 14904 22816 14968 22820
rect 19885 22876 19949 22880
rect 19885 22820 19889 22876
rect 19889 22820 19945 22876
rect 19945 22820 19949 22876
rect 19885 22816 19949 22820
rect 19965 22876 20029 22880
rect 19965 22820 19969 22876
rect 19969 22820 20025 22876
rect 20025 22820 20029 22876
rect 19965 22816 20029 22820
rect 20045 22876 20109 22880
rect 20045 22820 20049 22876
rect 20049 22820 20105 22876
rect 20105 22820 20109 22876
rect 20045 22816 20109 22820
rect 20125 22876 20189 22880
rect 20125 22820 20129 22876
rect 20129 22820 20185 22876
rect 20185 22820 20189 22876
rect 20125 22816 20189 22820
rect 3562 22332 3626 22336
rect 3562 22276 3566 22332
rect 3566 22276 3622 22332
rect 3622 22276 3626 22332
rect 3562 22272 3626 22276
rect 3642 22332 3706 22336
rect 3642 22276 3646 22332
rect 3646 22276 3702 22332
rect 3702 22276 3706 22332
rect 3642 22272 3706 22276
rect 3722 22332 3786 22336
rect 3722 22276 3726 22332
rect 3726 22276 3782 22332
rect 3782 22276 3786 22332
rect 3722 22272 3786 22276
rect 3802 22332 3866 22336
rect 3802 22276 3806 22332
rect 3806 22276 3862 22332
rect 3862 22276 3866 22332
rect 3802 22272 3866 22276
rect 8783 22332 8847 22336
rect 8783 22276 8787 22332
rect 8787 22276 8843 22332
rect 8843 22276 8847 22332
rect 8783 22272 8847 22276
rect 8863 22332 8927 22336
rect 8863 22276 8867 22332
rect 8867 22276 8923 22332
rect 8923 22276 8927 22332
rect 8863 22272 8927 22276
rect 8943 22332 9007 22336
rect 8943 22276 8947 22332
rect 8947 22276 9003 22332
rect 9003 22276 9007 22332
rect 8943 22272 9007 22276
rect 9023 22332 9087 22336
rect 9023 22276 9027 22332
rect 9027 22276 9083 22332
rect 9083 22276 9087 22332
rect 9023 22272 9087 22276
rect 14004 22332 14068 22336
rect 14004 22276 14008 22332
rect 14008 22276 14064 22332
rect 14064 22276 14068 22332
rect 14004 22272 14068 22276
rect 14084 22332 14148 22336
rect 14084 22276 14088 22332
rect 14088 22276 14144 22332
rect 14144 22276 14148 22332
rect 14084 22272 14148 22276
rect 14164 22332 14228 22336
rect 14164 22276 14168 22332
rect 14168 22276 14224 22332
rect 14224 22276 14228 22332
rect 14164 22272 14228 22276
rect 14244 22332 14308 22336
rect 14244 22276 14248 22332
rect 14248 22276 14304 22332
rect 14304 22276 14308 22332
rect 14244 22272 14308 22276
rect 19225 22332 19289 22336
rect 19225 22276 19229 22332
rect 19229 22276 19285 22332
rect 19285 22276 19289 22332
rect 19225 22272 19289 22276
rect 19305 22332 19369 22336
rect 19305 22276 19309 22332
rect 19309 22276 19365 22332
rect 19365 22276 19369 22332
rect 19305 22272 19369 22276
rect 19385 22332 19449 22336
rect 19385 22276 19389 22332
rect 19389 22276 19445 22332
rect 19445 22276 19449 22332
rect 19385 22272 19449 22276
rect 19465 22332 19529 22336
rect 19465 22276 19469 22332
rect 19469 22276 19525 22332
rect 19525 22276 19529 22332
rect 19465 22272 19529 22276
rect 4222 21788 4286 21792
rect 4222 21732 4226 21788
rect 4226 21732 4282 21788
rect 4282 21732 4286 21788
rect 4222 21728 4286 21732
rect 4302 21788 4366 21792
rect 4302 21732 4306 21788
rect 4306 21732 4362 21788
rect 4362 21732 4366 21788
rect 4302 21728 4366 21732
rect 4382 21788 4446 21792
rect 4382 21732 4386 21788
rect 4386 21732 4442 21788
rect 4442 21732 4446 21788
rect 4382 21728 4446 21732
rect 4462 21788 4526 21792
rect 4462 21732 4466 21788
rect 4466 21732 4522 21788
rect 4522 21732 4526 21788
rect 4462 21728 4526 21732
rect 9443 21788 9507 21792
rect 9443 21732 9447 21788
rect 9447 21732 9503 21788
rect 9503 21732 9507 21788
rect 9443 21728 9507 21732
rect 9523 21788 9587 21792
rect 9523 21732 9527 21788
rect 9527 21732 9583 21788
rect 9583 21732 9587 21788
rect 9523 21728 9587 21732
rect 9603 21788 9667 21792
rect 9603 21732 9607 21788
rect 9607 21732 9663 21788
rect 9663 21732 9667 21788
rect 9603 21728 9667 21732
rect 9683 21788 9747 21792
rect 9683 21732 9687 21788
rect 9687 21732 9743 21788
rect 9743 21732 9747 21788
rect 9683 21728 9747 21732
rect 14664 21788 14728 21792
rect 14664 21732 14668 21788
rect 14668 21732 14724 21788
rect 14724 21732 14728 21788
rect 14664 21728 14728 21732
rect 14744 21788 14808 21792
rect 14744 21732 14748 21788
rect 14748 21732 14804 21788
rect 14804 21732 14808 21788
rect 14744 21728 14808 21732
rect 14824 21788 14888 21792
rect 14824 21732 14828 21788
rect 14828 21732 14884 21788
rect 14884 21732 14888 21788
rect 14824 21728 14888 21732
rect 14904 21788 14968 21792
rect 14904 21732 14908 21788
rect 14908 21732 14964 21788
rect 14964 21732 14968 21788
rect 14904 21728 14968 21732
rect 19885 21788 19949 21792
rect 19885 21732 19889 21788
rect 19889 21732 19945 21788
rect 19945 21732 19949 21788
rect 19885 21728 19949 21732
rect 19965 21788 20029 21792
rect 19965 21732 19969 21788
rect 19969 21732 20025 21788
rect 20025 21732 20029 21788
rect 19965 21728 20029 21732
rect 20045 21788 20109 21792
rect 20045 21732 20049 21788
rect 20049 21732 20105 21788
rect 20105 21732 20109 21788
rect 20045 21728 20109 21732
rect 20125 21788 20189 21792
rect 20125 21732 20129 21788
rect 20129 21732 20185 21788
rect 20185 21732 20189 21788
rect 20125 21728 20189 21732
rect 3562 21244 3626 21248
rect 3562 21188 3566 21244
rect 3566 21188 3622 21244
rect 3622 21188 3626 21244
rect 3562 21184 3626 21188
rect 3642 21244 3706 21248
rect 3642 21188 3646 21244
rect 3646 21188 3702 21244
rect 3702 21188 3706 21244
rect 3642 21184 3706 21188
rect 3722 21244 3786 21248
rect 3722 21188 3726 21244
rect 3726 21188 3782 21244
rect 3782 21188 3786 21244
rect 3722 21184 3786 21188
rect 3802 21244 3866 21248
rect 3802 21188 3806 21244
rect 3806 21188 3862 21244
rect 3862 21188 3866 21244
rect 3802 21184 3866 21188
rect 8783 21244 8847 21248
rect 8783 21188 8787 21244
rect 8787 21188 8843 21244
rect 8843 21188 8847 21244
rect 8783 21184 8847 21188
rect 8863 21244 8927 21248
rect 8863 21188 8867 21244
rect 8867 21188 8923 21244
rect 8923 21188 8927 21244
rect 8863 21184 8927 21188
rect 8943 21244 9007 21248
rect 8943 21188 8947 21244
rect 8947 21188 9003 21244
rect 9003 21188 9007 21244
rect 8943 21184 9007 21188
rect 9023 21244 9087 21248
rect 9023 21188 9027 21244
rect 9027 21188 9083 21244
rect 9083 21188 9087 21244
rect 9023 21184 9087 21188
rect 14004 21244 14068 21248
rect 14004 21188 14008 21244
rect 14008 21188 14064 21244
rect 14064 21188 14068 21244
rect 14004 21184 14068 21188
rect 14084 21244 14148 21248
rect 14084 21188 14088 21244
rect 14088 21188 14144 21244
rect 14144 21188 14148 21244
rect 14084 21184 14148 21188
rect 14164 21244 14228 21248
rect 14164 21188 14168 21244
rect 14168 21188 14224 21244
rect 14224 21188 14228 21244
rect 14164 21184 14228 21188
rect 14244 21244 14308 21248
rect 14244 21188 14248 21244
rect 14248 21188 14304 21244
rect 14304 21188 14308 21244
rect 14244 21184 14308 21188
rect 19225 21244 19289 21248
rect 19225 21188 19229 21244
rect 19229 21188 19285 21244
rect 19285 21188 19289 21244
rect 19225 21184 19289 21188
rect 19305 21244 19369 21248
rect 19305 21188 19309 21244
rect 19309 21188 19365 21244
rect 19365 21188 19369 21244
rect 19305 21184 19369 21188
rect 19385 21244 19449 21248
rect 19385 21188 19389 21244
rect 19389 21188 19445 21244
rect 19445 21188 19449 21244
rect 19385 21184 19449 21188
rect 19465 21244 19529 21248
rect 19465 21188 19469 21244
rect 19469 21188 19525 21244
rect 19525 21188 19529 21244
rect 19465 21184 19529 21188
rect 3004 21116 3068 21180
rect 4222 20700 4286 20704
rect 4222 20644 4226 20700
rect 4226 20644 4282 20700
rect 4282 20644 4286 20700
rect 4222 20640 4286 20644
rect 4302 20700 4366 20704
rect 4302 20644 4306 20700
rect 4306 20644 4362 20700
rect 4362 20644 4366 20700
rect 4302 20640 4366 20644
rect 4382 20700 4446 20704
rect 4382 20644 4386 20700
rect 4386 20644 4442 20700
rect 4442 20644 4446 20700
rect 4382 20640 4446 20644
rect 4462 20700 4526 20704
rect 4462 20644 4466 20700
rect 4466 20644 4522 20700
rect 4522 20644 4526 20700
rect 4462 20640 4526 20644
rect 9443 20700 9507 20704
rect 9443 20644 9447 20700
rect 9447 20644 9503 20700
rect 9503 20644 9507 20700
rect 9443 20640 9507 20644
rect 9523 20700 9587 20704
rect 9523 20644 9527 20700
rect 9527 20644 9583 20700
rect 9583 20644 9587 20700
rect 9523 20640 9587 20644
rect 9603 20700 9667 20704
rect 9603 20644 9607 20700
rect 9607 20644 9663 20700
rect 9663 20644 9667 20700
rect 9603 20640 9667 20644
rect 9683 20700 9747 20704
rect 9683 20644 9687 20700
rect 9687 20644 9743 20700
rect 9743 20644 9747 20700
rect 9683 20640 9747 20644
rect 14664 20700 14728 20704
rect 14664 20644 14668 20700
rect 14668 20644 14724 20700
rect 14724 20644 14728 20700
rect 14664 20640 14728 20644
rect 14744 20700 14808 20704
rect 14744 20644 14748 20700
rect 14748 20644 14804 20700
rect 14804 20644 14808 20700
rect 14744 20640 14808 20644
rect 14824 20700 14888 20704
rect 14824 20644 14828 20700
rect 14828 20644 14884 20700
rect 14884 20644 14888 20700
rect 14824 20640 14888 20644
rect 14904 20700 14968 20704
rect 14904 20644 14908 20700
rect 14908 20644 14964 20700
rect 14964 20644 14968 20700
rect 14904 20640 14968 20644
rect 19885 20700 19949 20704
rect 19885 20644 19889 20700
rect 19889 20644 19945 20700
rect 19945 20644 19949 20700
rect 19885 20640 19949 20644
rect 19965 20700 20029 20704
rect 19965 20644 19969 20700
rect 19969 20644 20025 20700
rect 20025 20644 20029 20700
rect 19965 20640 20029 20644
rect 20045 20700 20109 20704
rect 20045 20644 20049 20700
rect 20049 20644 20105 20700
rect 20105 20644 20109 20700
rect 20045 20640 20109 20644
rect 20125 20700 20189 20704
rect 20125 20644 20129 20700
rect 20129 20644 20185 20700
rect 20185 20644 20189 20700
rect 20125 20640 20189 20644
rect 3562 20156 3626 20160
rect 3562 20100 3566 20156
rect 3566 20100 3622 20156
rect 3622 20100 3626 20156
rect 3562 20096 3626 20100
rect 3642 20156 3706 20160
rect 3642 20100 3646 20156
rect 3646 20100 3702 20156
rect 3702 20100 3706 20156
rect 3642 20096 3706 20100
rect 3722 20156 3786 20160
rect 3722 20100 3726 20156
rect 3726 20100 3782 20156
rect 3782 20100 3786 20156
rect 3722 20096 3786 20100
rect 3802 20156 3866 20160
rect 3802 20100 3806 20156
rect 3806 20100 3862 20156
rect 3862 20100 3866 20156
rect 3802 20096 3866 20100
rect 8783 20156 8847 20160
rect 8783 20100 8787 20156
rect 8787 20100 8843 20156
rect 8843 20100 8847 20156
rect 8783 20096 8847 20100
rect 8863 20156 8927 20160
rect 8863 20100 8867 20156
rect 8867 20100 8923 20156
rect 8923 20100 8927 20156
rect 8863 20096 8927 20100
rect 8943 20156 9007 20160
rect 8943 20100 8947 20156
rect 8947 20100 9003 20156
rect 9003 20100 9007 20156
rect 8943 20096 9007 20100
rect 9023 20156 9087 20160
rect 9023 20100 9027 20156
rect 9027 20100 9083 20156
rect 9083 20100 9087 20156
rect 9023 20096 9087 20100
rect 14004 20156 14068 20160
rect 14004 20100 14008 20156
rect 14008 20100 14064 20156
rect 14064 20100 14068 20156
rect 14004 20096 14068 20100
rect 14084 20156 14148 20160
rect 14084 20100 14088 20156
rect 14088 20100 14144 20156
rect 14144 20100 14148 20156
rect 14084 20096 14148 20100
rect 14164 20156 14228 20160
rect 14164 20100 14168 20156
rect 14168 20100 14224 20156
rect 14224 20100 14228 20156
rect 14164 20096 14228 20100
rect 14244 20156 14308 20160
rect 14244 20100 14248 20156
rect 14248 20100 14304 20156
rect 14304 20100 14308 20156
rect 14244 20096 14308 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 19465 20156 19529 20160
rect 19465 20100 19469 20156
rect 19469 20100 19525 20156
rect 19525 20100 19529 20156
rect 19465 20096 19529 20100
rect 4222 19612 4286 19616
rect 4222 19556 4226 19612
rect 4226 19556 4282 19612
rect 4282 19556 4286 19612
rect 4222 19552 4286 19556
rect 4302 19612 4366 19616
rect 4302 19556 4306 19612
rect 4306 19556 4362 19612
rect 4362 19556 4366 19612
rect 4302 19552 4366 19556
rect 4382 19612 4446 19616
rect 4382 19556 4386 19612
rect 4386 19556 4442 19612
rect 4442 19556 4446 19612
rect 4382 19552 4446 19556
rect 4462 19612 4526 19616
rect 4462 19556 4466 19612
rect 4466 19556 4522 19612
rect 4522 19556 4526 19612
rect 4462 19552 4526 19556
rect 9443 19612 9507 19616
rect 9443 19556 9447 19612
rect 9447 19556 9503 19612
rect 9503 19556 9507 19612
rect 9443 19552 9507 19556
rect 9523 19612 9587 19616
rect 9523 19556 9527 19612
rect 9527 19556 9583 19612
rect 9583 19556 9587 19612
rect 9523 19552 9587 19556
rect 9603 19612 9667 19616
rect 9603 19556 9607 19612
rect 9607 19556 9663 19612
rect 9663 19556 9667 19612
rect 9603 19552 9667 19556
rect 9683 19612 9747 19616
rect 9683 19556 9687 19612
rect 9687 19556 9743 19612
rect 9743 19556 9747 19612
rect 9683 19552 9747 19556
rect 8524 19408 8588 19412
rect 14664 19612 14728 19616
rect 14664 19556 14668 19612
rect 14668 19556 14724 19612
rect 14724 19556 14728 19612
rect 14664 19552 14728 19556
rect 14744 19612 14808 19616
rect 14744 19556 14748 19612
rect 14748 19556 14804 19612
rect 14804 19556 14808 19612
rect 14744 19552 14808 19556
rect 14824 19612 14888 19616
rect 14824 19556 14828 19612
rect 14828 19556 14884 19612
rect 14884 19556 14888 19612
rect 14824 19552 14888 19556
rect 14904 19612 14968 19616
rect 14904 19556 14908 19612
rect 14908 19556 14964 19612
rect 14964 19556 14968 19612
rect 14904 19552 14968 19556
rect 19885 19612 19949 19616
rect 19885 19556 19889 19612
rect 19889 19556 19945 19612
rect 19945 19556 19949 19612
rect 19885 19552 19949 19556
rect 19965 19612 20029 19616
rect 19965 19556 19969 19612
rect 19969 19556 20025 19612
rect 20025 19556 20029 19612
rect 19965 19552 20029 19556
rect 20045 19612 20109 19616
rect 20045 19556 20049 19612
rect 20049 19556 20105 19612
rect 20105 19556 20109 19612
rect 20045 19552 20109 19556
rect 20125 19612 20189 19616
rect 20125 19556 20129 19612
rect 20129 19556 20185 19612
rect 20185 19556 20189 19612
rect 20125 19552 20189 19556
rect 8524 19352 8574 19408
rect 8574 19352 8588 19408
rect 8524 19348 8588 19352
rect 3562 19068 3626 19072
rect 3562 19012 3566 19068
rect 3566 19012 3622 19068
rect 3622 19012 3626 19068
rect 3562 19008 3626 19012
rect 3642 19068 3706 19072
rect 3642 19012 3646 19068
rect 3646 19012 3702 19068
rect 3702 19012 3706 19068
rect 3642 19008 3706 19012
rect 3722 19068 3786 19072
rect 3722 19012 3726 19068
rect 3726 19012 3782 19068
rect 3782 19012 3786 19068
rect 3722 19008 3786 19012
rect 3802 19068 3866 19072
rect 3802 19012 3806 19068
rect 3806 19012 3862 19068
rect 3862 19012 3866 19068
rect 3802 19008 3866 19012
rect 8783 19068 8847 19072
rect 8783 19012 8787 19068
rect 8787 19012 8843 19068
rect 8843 19012 8847 19068
rect 8783 19008 8847 19012
rect 8863 19068 8927 19072
rect 8863 19012 8867 19068
rect 8867 19012 8923 19068
rect 8923 19012 8927 19068
rect 8863 19008 8927 19012
rect 8943 19068 9007 19072
rect 8943 19012 8947 19068
rect 8947 19012 9003 19068
rect 9003 19012 9007 19068
rect 8943 19008 9007 19012
rect 9023 19068 9087 19072
rect 9023 19012 9027 19068
rect 9027 19012 9083 19068
rect 9083 19012 9087 19068
rect 9023 19008 9087 19012
rect 14004 19068 14068 19072
rect 14004 19012 14008 19068
rect 14008 19012 14064 19068
rect 14064 19012 14068 19068
rect 14004 19008 14068 19012
rect 14084 19068 14148 19072
rect 14084 19012 14088 19068
rect 14088 19012 14144 19068
rect 14144 19012 14148 19068
rect 14084 19008 14148 19012
rect 14164 19068 14228 19072
rect 14164 19012 14168 19068
rect 14168 19012 14224 19068
rect 14224 19012 14228 19068
rect 14164 19008 14228 19012
rect 14244 19068 14308 19072
rect 14244 19012 14248 19068
rect 14248 19012 14304 19068
rect 14304 19012 14308 19068
rect 14244 19008 14308 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 19465 19068 19529 19072
rect 19465 19012 19469 19068
rect 19469 19012 19525 19068
rect 19525 19012 19529 19068
rect 19465 19008 19529 19012
rect 17724 18532 17788 18596
rect 4222 18524 4286 18528
rect 4222 18468 4226 18524
rect 4226 18468 4282 18524
rect 4282 18468 4286 18524
rect 4222 18464 4286 18468
rect 4302 18524 4366 18528
rect 4302 18468 4306 18524
rect 4306 18468 4362 18524
rect 4362 18468 4366 18524
rect 4302 18464 4366 18468
rect 4382 18524 4446 18528
rect 4382 18468 4386 18524
rect 4386 18468 4442 18524
rect 4442 18468 4446 18524
rect 4382 18464 4446 18468
rect 4462 18524 4526 18528
rect 4462 18468 4466 18524
rect 4466 18468 4522 18524
rect 4522 18468 4526 18524
rect 4462 18464 4526 18468
rect 9443 18524 9507 18528
rect 9443 18468 9447 18524
rect 9447 18468 9503 18524
rect 9503 18468 9507 18524
rect 9443 18464 9507 18468
rect 9523 18524 9587 18528
rect 9523 18468 9527 18524
rect 9527 18468 9583 18524
rect 9583 18468 9587 18524
rect 9523 18464 9587 18468
rect 9603 18524 9667 18528
rect 9603 18468 9607 18524
rect 9607 18468 9663 18524
rect 9663 18468 9667 18524
rect 9603 18464 9667 18468
rect 9683 18524 9747 18528
rect 9683 18468 9687 18524
rect 9687 18468 9743 18524
rect 9743 18468 9747 18524
rect 9683 18464 9747 18468
rect 14664 18524 14728 18528
rect 14664 18468 14668 18524
rect 14668 18468 14724 18524
rect 14724 18468 14728 18524
rect 14664 18464 14728 18468
rect 14744 18524 14808 18528
rect 14744 18468 14748 18524
rect 14748 18468 14804 18524
rect 14804 18468 14808 18524
rect 14744 18464 14808 18468
rect 14824 18524 14888 18528
rect 14824 18468 14828 18524
rect 14828 18468 14884 18524
rect 14884 18468 14888 18524
rect 14824 18464 14888 18468
rect 14904 18524 14968 18528
rect 14904 18468 14908 18524
rect 14908 18468 14964 18524
rect 14964 18468 14968 18524
rect 14904 18464 14968 18468
rect 19885 18524 19949 18528
rect 19885 18468 19889 18524
rect 19889 18468 19945 18524
rect 19945 18468 19949 18524
rect 19885 18464 19949 18468
rect 19965 18524 20029 18528
rect 19965 18468 19969 18524
rect 19969 18468 20025 18524
rect 20025 18468 20029 18524
rect 19965 18464 20029 18468
rect 20045 18524 20109 18528
rect 20045 18468 20049 18524
rect 20049 18468 20105 18524
rect 20105 18468 20109 18524
rect 20045 18464 20109 18468
rect 20125 18524 20189 18528
rect 20125 18468 20129 18524
rect 20129 18468 20185 18524
rect 20185 18468 20189 18524
rect 20125 18464 20189 18468
rect 3562 17980 3626 17984
rect 3562 17924 3566 17980
rect 3566 17924 3622 17980
rect 3622 17924 3626 17980
rect 3562 17920 3626 17924
rect 3642 17980 3706 17984
rect 3642 17924 3646 17980
rect 3646 17924 3702 17980
rect 3702 17924 3706 17980
rect 3642 17920 3706 17924
rect 3722 17980 3786 17984
rect 3722 17924 3726 17980
rect 3726 17924 3782 17980
rect 3782 17924 3786 17980
rect 3722 17920 3786 17924
rect 3802 17980 3866 17984
rect 3802 17924 3806 17980
rect 3806 17924 3862 17980
rect 3862 17924 3866 17980
rect 3802 17920 3866 17924
rect 8783 17980 8847 17984
rect 8783 17924 8787 17980
rect 8787 17924 8843 17980
rect 8843 17924 8847 17980
rect 8783 17920 8847 17924
rect 8863 17980 8927 17984
rect 8863 17924 8867 17980
rect 8867 17924 8923 17980
rect 8923 17924 8927 17980
rect 8863 17920 8927 17924
rect 8943 17980 9007 17984
rect 8943 17924 8947 17980
rect 8947 17924 9003 17980
rect 9003 17924 9007 17980
rect 8943 17920 9007 17924
rect 9023 17980 9087 17984
rect 9023 17924 9027 17980
rect 9027 17924 9083 17980
rect 9083 17924 9087 17980
rect 9023 17920 9087 17924
rect 14004 17980 14068 17984
rect 14004 17924 14008 17980
rect 14008 17924 14064 17980
rect 14064 17924 14068 17980
rect 14004 17920 14068 17924
rect 14084 17980 14148 17984
rect 14084 17924 14088 17980
rect 14088 17924 14144 17980
rect 14144 17924 14148 17980
rect 14084 17920 14148 17924
rect 14164 17980 14228 17984
rect 14164 17924 14168 17980
rect 14168 17924 14224 17980
rect 14224 17924 14228 17980
rect 14164 17920 14228 17924
rect 14244 17980 14308 17984
rect 14244 17924 14248 17980
rect 14248 17924 14304 17980
rect 14304 17924 14308 17980
rect 14244 17920 14308 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 19465 17980 19529 17984
rect 19465 17924 19469 17980
rect 19469 17924 19525 17980
rect 19525 17924 19529 17980
rect 19465 17920 19529 17924
rect 4222 17436 4286 17440
rect 4222 17380 4226 17436
rect 4226 17380 4282 17436
rect 4282 17380 4286 17436
rect 4222 17376 4286 17380
rect 4302 17436 4366 17440
rect 4302 17380 4306 17436
rect 4306 17380 4362 17436
rect 4362 17380 4366 17436
rect 4302 17376 4366 17380
rect 4382 17436 4446 17440
rect 4382 17380 4386 17436
rect 4386 17380 4442 17436
rect 4442 17380 4446 17436
rect 4382 17376 4446 17380
rect 4462 17436 4526 17440
rect 4462 17380 4466 17436
rect 4466 17380 4522 17436
rect 4522 17380 4526 17436
rect 4462 17376 4526 17380
rect 9443 17436 9507 17440
rect 9443 17380 9447 17436
rect 9447 17380 9503 17436
rect 9503 17380 9507 17436
rect 9443 17376 9507 17380
rect 9523 17436 9587 17440
rect 9523 17380 9527 17436
rect 9527 17380 9583 17436
rect 9583 17380 9587 17436
rect 9523 17376 9587 17380
rect 9603 17436 9667 17440
rect 9603 17380 9607 17436
rect 9607 17380 9663 17436
rect 9663 17380 9667 17436
rect 9603 17376 9667 17380
rect 9683 17436 9747 17440
rect 9683 17380 9687 17436
rect 9687 17380 9743 17436
rect 9743 17380 9747 17436
rect 9683 17376 9747 17380
rect 14664 17436 14728 17440
rect 14664 17380 14668 17436
rect 14668 17380 14724 17436
rect 14724 17380 14728 17436
rect 14664 17376 14728 17380
rect 14744 17436 14808 17440
rect 14744 17380 14748 17436
rect 14748 17380 14804 17436
rect 14804 17380 14808 17436
rect 14744 17376 14808 17380
rect 14824 17436 14888 17440
rect 14824 17380 14828 17436
rect 14828 17380 14884 17436
rect 14884 17380 14888 17436
rect 14824 17376 14888 17380
rect 14904 17436 14968 17440
rect 14904 17380 14908 17436
rect 14908 17380 14964 17436
rect 14964 17380 14968 17436
rect 14904 17376 14968 17380
rect 19885 17436 19949 17440
rect 19885 17380 19889 17436
rect 19889 17380 19945 17436
rect 19945 17380 19949 17436
rect 19885 17376 19949 17380
rect 19965 17436 20029 17440
rect 19965 17380 19969 17436
rect 19969 17380 20025 17436
rect 20025 17380 20029 17436
rect 19965 17376 20029 17380
rect 20045 17436 20109 17440
rect 20045 17380 20049 17436
rect 20049 17380 20105 17436
rect 20105 17380 20109 17436
rect 20045 17376 20109 17380
rect 20125 17436 20189 17440
rect 20125 17380 20129 17436
rect 20129 17380 20185 17436
rect 20185 17380 20189 17436
rect 20125 17376 20189 17380
rect 8524 17172 8588 17236
rect 14412 17172 14476 17236
rect 3562 16892 3626 16896
rect 3562 16836 3566 16892
rect 3566 16836 3622 16892
rect 3622 16836 3626 16892
rect 3562 16832 3626 16836
rect 3642 16892 3706 16896
rect 3642 16836 3646 16892
rect 3646 16836 3702 16892
rect 3702 16836 3706 16892
rect 3642 16832 3706 16836
rect 3722 16892 3786 16896
rect 3722 16836 3726 16892
rect 3726 16836 3782 16892
rect 3782 16836 3786 16892
rect 3722 16832 3786 16836
rect 3802 16892 3866 16896
rect 3802 16836 3806 16892
rect 3806 16836 3862 16892
rect 3862 16836 3866 16892
rect 3802 16832 3866 16836
rect 8783 16892 8847 16896
rect 8783 16836 8787 16892
rect 8787 16836 8843 16892
rect 8843 16836 8847 16892
rect 8783 16832 8847 16836
rect 8863 16892 8927 16896
rect 8863 16836 8867 16892
rect 8867 16836 8923 16892
rect 8923 16836 8927 16892
rect 8863 16832 8927 16836
rect 8943 16892 9007 16896
rect 8943 16836 8947 16892
rect 8947 16836 9003 16892
rect 9003 16836 9007 16892
rect 8943 16832 9007 16836
rect 9023 16892 9087 16896
rect 9023 16836 9027 16892
rect 9027 16836 9083 16892
rect 9083 16836 9087 16892
rect 9023 16832 9087 16836
rect 14004 16892 14068 16896
rect 14004 16836 14008 16892
rect 14008 16836 14064 16892
rect 14064 16836 14068 16892
rect 14004 16832 14068 16836
rect 14084 16892 14148 16896
rect 14084 16836 14088 16892
rect 14088 16836 14144 16892
rect 14144 16836 14148 16892
rect 14084 16832 14148 16836
rect 14164 16892 14228 16896
rect 14164 16836 14168 16892
rect 14168 16836 14224 16892
rect 14224 16836 14228 16892
rect 14164 16832 14228 16836
rect 14244 16892 14308 16896
rect 14244 16836 14248 16892
rect 14248 16836 14304 16892
rect 14304 16836 14308 16892
rect 14244 16832 14308 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 19465 16892 19529 16896
rect 19465 16836 19469 16892
rect 19469 16836 19525 16892
rect 19525 16836 19529 16892
rect 19465 16832 19529 16836
rect 4222 16348 4286 16352
rect 4222 16292 4226 16348
rect 4226 16292 4282 16348
rect 4282 16292 4286 16348
rect 4222 16288 4286 16292
rect 4302 16348 4366 16352
rect 4302 16292 4306 16348
rect 4306 16292 4362 16348
rect 4362 16292 4366 16348
rect 4302 16288 4366 16292
rect 4382 16348 4446 16352
rect 4382 16292 4386 16348
rect 4386 16292 4442 16348
rect 4442 16292 4446 16348
rect 4382 16288 4446 16292
rect 4462 16348 4526 16352
rect 4462 16292 4466 16348
rect 4466 16292 4522 16348
rect 4522 16292 4526 16348
rect 4462 16288 4526 16292
rect 9443 16348 9507 16352
rect 9443 16292 9447 16348
rect 9447 16292 9503 16348
rect 9503 16292 9507 16348
rect 9443 16288 9507 16292
rect 9523 16348 9587 16352
rect 9523 16292 9527 16348
rect 9527 16292 9583 16348
rect 9583 16292 9587 16348
rect 9523 16288 9587 16292
rect 9603 16348 9667 16352
rect 9603 16292 9607 16348
rect 9607 16292 9663 16348
rect 9663 16292 9667 16348
rect 9603 16288 9667 16292
rect 9683 16348 9747 16352
rect 9683 16292 9687 16348
rect 9687 16292 9743 16348
rect 9743 16292 9747 16348
rect 9683 16288 9747 16292
rect 14664 16348 14728 16352
rect 14664 16292 14668 16348
rect 14668 16292 14724 16348
rect 14724 16292 14728 16348
rect 14664 16288 14728 16292
rect 14744 16348 14808 16352
rect 14744 16292 14748 16348
rect 14748 16292 14804 16348
rect 14804 16292 14808 16348
rect 14744 16288 14808 16292
rect 14824 16348 14888 16352
rect 14824 16292 14828 16348
rect 14828 16292 14884 16348
rect 14884 16292 14888 16348
rect 14824 16288 14888 16292
rect 14904 16348 14968 16352
rect 14904 16292 14908 16348
rect 14908 16292 14964 16348
rect 14964 16292 14968 16348
rect 14904 16288 14968 16292
rect 19885 16348 19949 16352
rect 19885 16292 19889 16348
rect 19889 16292 19945 16348
rect 19945 16292 19949 16348
rect 19885 16288 19949 16292
rect 19965 16348 20029 16352
rect 19965 16292 19969 16348
rect 19969 16292 20025 16348
rect 20025 16292 20029 16348
rect 19965 16288 20029 16292
rect 20045 16348 20109 16352
rect 20045 16292 20049 16348
rect 20049 16292 20105 16348
rect 20105 16292 20109 16348
rect 20045 16288 20109 16292
rect 20125 16348 20189 16352
rect 20125 16292 20129 16348
rect 20129 16292 20185 16348
rect 20185 16292 20189 16348
rect 20125 16288 20189 16292
rect 17724 16084 17788 16148
rect 3562 15804 3626 15808
rect 3562 15748 3566 15804
rect 3566 15748 3622 15804
rect 3622 15748 3626 15804
rect 3562 15744 3626 15748
rect 3642 15804 3706 15808
rect 3642 15748 3646 15804
rect 3646 15748 3702 15804
rect 3702 15748 3706 15804
rect 3642 15744 3706 15748
rect 3722 15804 3786 15808
rect 3722 15748 3726 15804
rect 3726 15748 3782 15804
rect 3782 15748 3786 15804
rect 3722 15744 3786 15748
rect 3802 15804 3866 15808
rect 3802 15748 3806 15804
rect 3806 15748 3862 15804
rect 3862 15748 3866 15804
rect 3802 15744 3866 15748
rect 8783 15804 8847 15808
rect 8783 15748 8787 15804
rect 8787 15748 8843 15804
rect 8843 15748 8847 15804
rect 8783 15744 8847 15748
rect 8863 15804 8927 15808
rect 8863 15748 8867 15804
rect 8867 15748 8923 15804
rect 8923 15748 8927 15804
rect 8863 15744 8927 15748
rect 8943 15804 9007 15808
rect 8943 15748 8947 15804
rect 8947 15748 9003 15804
rect 9003 15748 9007 15804
rect 8943 15744 9007 15748
rect 9023 15804 9087 15808
rect 9023 15748 9027 15804
rect 9027 15748 9083 15804
rect 9083 15748 9087 15804
rect 9023 15744 9087 15748
rect 14004 15804 14068 15808
rect 14004 15748 14008 15804
rect 14008 15748 14064 15804
rect 14064 15748 14068 15804
rect 14004 15744 14068 15748
rect 14084 15804 14148 15808
rect 14084 15748 14088 15804
rect 14088 15748 14144 15804
rect 14144 15748 14148 15804
rect 14084 15744 14148 15748
rect 14164 15804 14228 15808
rect 14164 15748 14168 15804
rect 14168 15748 14224 15804
rect 14224 15748 14228 15804
rect 14164 15744 14228 15748
rect 14244 15804 14308 15808
rect 14244 15748 14248 15804
rect 14248 15748 14304 15804
rect 14304 15748 14308 15804
rect 14244 15744 14308 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 19465 15804 19529 15808
rect 19465 15748 19469 15804
rect 19469 15748 19525 15804
rect 19525 15748 19529 15804
rect 19465 15744 19529 15748
rect 4222 15260 4286 15264
rect 4222 15204 4226 15260
rect 4226 15204 4282 15260
rect 4282 15204 4286 15260
rect 4222 15200 4286 15204
rect 4302 15260 4366 15264
rect 4302 15204 4306 15260
rect 4306 15204 4362 15260
rect 4362 15204 4366 15260
rect 4302 15200 4366 15204
rect 4382 15260 4446 15264
rect 4382 15204 4386 15260
rect 4386 15204 4442 15260
rect 4442 15204 4446 15260
rect 4382 15200 4446 15204
rect 4462 15260 4526 15264
rect 4462 15204 4466 15260
rect 4466 15204 4522 15260
rect 4522 15204 4526 15260
rect 4462 15200 4526 15204
rect 9443 15260 9507 15264
rect 9443 15204 9447 15260
rect 9447 15204 9503 15260
rect 9503 15204 9507 15260
rect 9443 15200 9507 15204
rect 9523 15260 9587 15264
rect 9523 15204 9527 15260
rect 9527 15204 9583 15260
rect 9583 15204 9587 15260
rect 9523 15200 9587 15204
rect 9603 15260 9667 15264
rect 9603 15204 9607 15260
rect 9607 15204 9663 15260
rect 9663 15204 9667 15260
rect 9603 15200 9667 15204
rect 9683 15260 9747 15264
rect 9683 15204 9687 15260
rect 9687 15204 9743 15260
rect 9743 15204 9747 15260
rect 9683 15200 9747 15204
rect 14664 15260 14728 15264
rect 14664 15204 14668 15260
rect 14668 15204 14724 15260
rect 14724 15204 14728 15260
rect 14664 15200 14728 15204
rect 14744 15260 14808 15264
rect 14744 15204 14748 15260
rect 14748 15204 14804 15260
rect 14804 15204 14808 15260
rect 14744 15200 14808 15204
rect 14824 15260 14888 15264
rect 14824 15204 14828 15260
rect 14828 15204 14884 15260
rect 14884 15204 14888 15260
rect 14824 15200 14888 15204
rect 14904 15260 14968 15264
rect 14904 15204 14908 15260
rect 14908 15204 14964 15260
rect 14964 15204 14968 15260
rect 14904 15200 14968 15204
rect 19885 15260 19949 15264
rect 19885 15204 19889 15260
rect 19889 15204 19945 15260
rect 19945 15204 19949 15260
rect 19885 15200 19949 15204
rect 19965 15260 20029 15264
rect 19965 15204 19969 15260
rect 19969 15204 20025 15260
rect 20025 15204 20029 15260
rect 19965 15200 20029 15204
rect 20045 15260 20109 15264
rect 20045 15204 20049 15260
rect 20049 15204 20105 15260
rect 20105 15204 20109 15260
rect 20045 15200 20109 15204
rect 20125 15260 20189 15264
rect 20125 15204 20129 15260
rect 20129 15204 20185 15260
rect 20185 15204 20189 15260
rect 20125 15200 20189 15204
rect 3562 14716 3626 14720
rect 3562 14660 3566 14716
rect 3566 14660 3622 14716
rect 3622 14660 3626 14716
rect 3562 14656 3626 14660
rect 3642 14716 3706 14720
rect 3642 14660 3646 14716
rect 3646 14660 3702 14716
rect 3702 14660 3706 14716
rect 3642 14656 3706 14660
rect 3722 14716 3786 14720
rect 3722 14660 3726 14716
rect 3726 14660 3782 14716
rect 3782 14660 3786 14716
rect 3722 14656 3786 14660
rect 3802 14716 3866 14720
rect 3802 14660 3806 14716
rect 3806 14660 3862 14716
rect 3862 14660 3866 14716
rect 3802 14656 3866 14660
rect 8783 14716 8847 14720
rect 8783 14660 8787 14716
rect 8787 14660 8843 14716
rect 8843 14660 8847 14716
rect 8783 14656 8847 14660
rect 8863 14716 8927 14720
rect 8863 14660 8867 14716
rect 8867 14660 8923 14716
rect 8923 14660 8927 14716
rect 8863 14656 8927 14660
rect 8943 14716 9007 14720
rect 8943 14660 8947 14716
rect 8947 14660 9003 14716
rect 9003 14660 9007 14716
rect 8943 14656 9007 14660
rect 9023 14716 9087 14720
rect 9023 14660 9027 14716
rect 9027 14660 9083 14716
rect 9083 14660 9087 14716
rect 9023 14656 9087 14660
rect 14004 14716 14068 14720
rect 14004 14660 14008 14716
rect 14008 14660 14064 14716
rect 14064 14660 14068 14716
rect 14004 14656 14068 14660
rect 14084 14716 14148 14720
rect 14084 14660 14088 14716
rect 14088 14660 14144 14716
rect 14144 14660 14148 14716
rect 14084 14656 14148 14660
rect 14164 14716 14228 14720
rect 14164 14660 14168 14716
rect 14168 14660 14224 14716
rect 14224 14660 14228 14716
rect 14164 14656 14228 14660
rect 14244 14716 14308 14720
rect 14244 14660 14248 14716
rect 14248 14660 14304 14716
rect 14304 14660 14308 14716
rect 14244 14656 14308 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 19465 14716 19529 14720
rect 19465 14660 19469 14716
rect 19469 14660 19525 14716
rect 19525 14660 19529 14716
rect 19465 14656 19529 14660
rect 4222 14172 4286 14176
rect 4222 14116 4226 14172
rect 4226 14116 4282 14172
rect 4282 14116 4286 14172
rect 4222 14112 4286 14116
rect 4302 14172 4366 14176
rect 4302 14116 4306 14172
rect 4306 14116 4362 14172
rect 4362 14116 4366 14172
rect 4302 14112 4366 14116
rect 4382 14172 4446 14176
rect 4382 14116 4386 14172
rect 4386 14116 4442 14172
rect 4442 14116 4446 14172
rect 4382 14112 4446 14116
rect 4462 14172 4526 14176
rect 4462 14116 4466 14172
rect 4466 14116 4522 14172
rect 4522 14116 4526 14172
rect 4462 14112 4526 14116
rect 9443 14172 9507 14176
rect 9443 14116 9447 14172
rect 9447 14116 9503 14172
rect 9503 14116 9507 14172
rect 9443 14112 9507 14116
rect 9523 14172 9587 14176
rect 9523 14116 9527 14172
rect 9527 14116 9583 14172
rect 9583 14116 9587 14172
rect 9523 14112 9587 14116
rect 9603 14172 9667 14176
rect 9603 14116 9607 14172
rect 9607 14116 9663 14172
rect 9663 14116 9667 14172
rect 9603 14112 9667 14116
rect 9683 14172 9747 14176
rect 9683 14116 9687 14172
rect 9687 14116 9743 14172
rect 9743 14116 9747 14172
rect 9683 14112 9747 14116
rect 14664 14172 14728 14176
rect 14664 14116 14668 14172
rect 14668 14116 14724 14172
rect 14724 14116 14728 14172
rect 14664 14112 14728 14116
rect 14744 14172 14808 14176
rect 14744 14116 14748 14172
rect 14748 14116 14804 14172
rect 14804 14116 14808 14172
rect 14744 14112 14808 14116
rect 14824 14172 14888 14176
rect 14824 14116 14828 14172
rect 14828 14116 14884 14172
rect 14884 14116 14888 14172
rect 14824 14112 14888 14116
rect 14904 14172 14968 14176
rect 14904 14116 14908 14172
rect 14908 14116 14964 14172
rect 14964 14116 14968 14172
rect 14904 14112 14968 14116
rect 19885 14172 19949 14176
rect 19885 14116 19889 14172
rect 19889 14116 19945 14172
rect 19945 14116 19949 14172
rect 19885 14112 19949 14116
rect 19965 14172 20029 14176
rect 19965 14116 19969 14172
rect 19969 14116 20025 14172
rect 20025 14116 20029 14172
rect 19965 14112 20029 14116
rect 20045 14172 20109 14176
rect 20045 14116 20049 14172
rect 20049 14116 20105 14172
rect 20105 14116 20109 14172
rect 20045 14112 20109 14116
rect 20125 14172 20189 14176
rect 20125 14116 20129 14172
rect 20129 14116 20185 14172
rect 20185 14116 20189 14172
rect 20125 14112 20189 14116
rect 3562 13628 3626 13632
rect 3562 13572 3566 13628
rect 3566 13572 3622 13628
rect 3622 13572 3626 13628
rect 3562 13568 3626 13572
rect 3642 13628 3706 13632
rect 3642 13572 3646 13628
rect 3646 13572 3702 13628
rect 3702 13572 3706 13628
rect 3642 13568 3706 13572
rect 3722 13628 3786 13632
rect 3722 13572 3726 13628
rect 3726 13572 3782 13628
rect 3782 13572 3786 13628
rect 3722 13568 3786 13572
rect 3802 13628 3866 13632
rect 3802 13572 3806 13628
rect 3806 13572 3862 13628
rect 3862 13572 3866 13628
rect 3802 13568 3866 13572
rect 8783 13628 8847 13632
rect 8783 13572 8787 13628
rect 8787 13572 8843 13628
rect 8843 13572 8847 13628
rect 8783 13568 8847 13572
rect 8863 13628 8927 13632
rect 8863 13572 8867 13628
rect 8867 13572 8923 13628
rect 8923 13572 8927 13628
rect 8863 13568 8927 13572
rect 8943 13628 9007 13632
rect 8943 13572 8947 13628
rect 8947 13572 9003 13628
rect 9003 13572 9007 13628
rect 8943 13568 9007 13572
rect 9023 13628 9087 13632
rect 9023 13572 9027 13628
rect 9027 13572 9083 13628
rect 9083 13572 9087 13628
rect 9023 13568 9087 13572
rect 14004 13628 14068 13632
rect 14004 13572 14008 13628
rect 14008 13572 14064 13628
rect 14064 13572 14068 13628
rect 14004 13568 14068 13572
rect 14084 13628 14148 13632
rect 14084 13572 14088 13628
rect 14088 13572 14144 13628
rect 14144 13572 14148 13628
rect 14084 13568 14148 13572
rect 14164 13628 14228 13632
rect 14164 13572 14168 13628
rect 14168 13572 14224 13628
rect 14224 13572 14228 13628
rect 14164 13568 14228 13572
rect 14244 13628 14308 13632
rect 14244 13572 14248 13628
rect 14248 13572 14304 13628
rect 14304 13572 14308 13628
rect 14244 13568 14308 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 19465 13628 19529 13632
rect 19465 13572 19469 13628
rect 19469 13572 19525 13628
rect 19525 13572 19529 13628
rect 19465 13568 19529 13572
rect 4222 13084 4286 13088
rect 4222 13028 4226 13084
rect 4226 13028 4282 13084
rect 4282 13028 4286 13084
rect 4222 13024 4286 13028
rect 4302 13084 4366 13088
rect 4302 13028 4306 13084
rect 4306 13028 4362 13084
rect 4362 13028 4366 13084
rect 4302 13024 4366 13028
rect 4382 13084 4446 13088
rect 4382 13028 4386 13084
rect 4386 13028 4442 13084
rect 4442 13028 4446 13084
rect 4382 13024 4446 13028
rect 4462 13084 4526 13088
rect 4462 13028 4466 13084
rect 4466 13028 4522 13084
rect 4522 13028 4526 13084
rect 4462 13024 4526 13028
rect 9443 13084 9507 13088
rect 9443 13028 9447 13084
rect 9447 13028 9503 13084
rect 9503 13028 9507 13084
rect 9443 13024 9507 13028
rect 9523 13084 9587 13088
rect 9523 13028 9527 13084
rect 9527 13028 9583 13084
rect 9583 13028 9587 13084
rect 9523 13024 9587 13028
rect 9603 13084 9667 13088
rect 9603 13028 9607 13084
rect 9607 13028 9663 13084
rect 9663 13028 9667 13084
rect 9603 13024 9667 13028
rect 9683 13084 9747 13088
rect 9683 13028 9687 13084
rect 9687 13028 9743 13084
rect 9743 13028 9747 13084
rect 9683 13024 9747 13028
rect 14664 13084 14728 13088
rect 14664 13028 14668 13084
rect 14668 13028 14724 13084
rect 14724 13028 14728 13084
rect 14664 13024 14728 13028
rect 14744 13084 14808 13088
rect 14744 13028 14748 13084
rect 14748 13028 14804 13084
rect 14804 13028 14808 13084
rect 14744 13024 14808 13028
rect 14824 13084 14888 13088
rect 14824 13028 14828 13084
rect 14828 13028 14884 13084
rect 14884 13028 14888 13084
rect 14824 13024 14888 13028
rect 14904 13084 14968 13088
rect 14904 13028 14908 13084
rect 14908 13028 14964 13084
rect 14964 13028 14968 13084
rect 14904 13024 14968 13028
rect 19885 13084 19949 13088
rect 19885 13028 19889 13084
rect 19889 13028 19945 13084
rect 19945 13028 19949 13084
rect 19885 13024 19949 13028
rect 19965 13084 20029 13088
rect 19965 13028 19969 13084
rect 19969 13028 20025 13084
rect 20025 13028 20029 13084
rect 19965 13024 20029 13028
rect 20045 13084 20109 13088
rect 20045 13028 20049 13084
rect 20049 13028 20105 13084
rect 20105 13028 20109 13084
rect 20045 13024 20109 13028
rect 20125 13084 20189 13088
rect 20125 13028 20129 13084
rect 20129 13028 20185 13084
rect 20185 13028 20189 13084
rect 20125 13024 20189 13028
rect 3562 12540 3626 12544
rect 3562 12484 3566 12540
rect 3566 12484 3622 12540
rect 3622 12484 3626 12540
rect 3562 12480 3626 12484
rect 3642 12540 3706 12544
rect 3642 12484 3646 12540
rect 3646 12484 3702 12540
rect 3702 12484 3706 12540
rect 3642 12480 3706 12484
rect 3722 12540 3786 12544
rect 3722 12484 3726 12540
rect 3726 12484 3782 12540
rect 3782 12484 3786 12540
rect 3722 12480 3786 12484
rect 3802 12540 3866 12544
rect 3802 12484 3806 12540
rect 3806 12484 3862 12540
rect 3862 12484 3866 12540
rect 3802 12480 3866 12484
rect 8783 12540 8847 12544
rect 8783 12484 8787 12540
rect 8787 12484 8843 12540
rect 8843 12484 8847 12540
rect 8783 12480 8847 12484
rect 8863 12540 8927 12544
rect 8863 12484 8867 12540
rect 8867 12484 8923 12540
rect 8923 12484 8927 12540
rect 8863 12480 8927 12484
rect 8943 12540 9007 12544
rect 8943 12484 8947 12540
rect 8947 12484 9003 12540
rect 9003 12484 9007 12540
rect 8943 12480 9007 12484
rect 9023 12540 9087 12544
rect 9023 12484 9027 12540
rect 9027 12484 9083 12540
rect 9083 12484 9087 12540
rect 9023 12480 9087 12484
rect 14004 12540 14068 12544
rect 14004 12484 14008 12540
rect 14008 12484 14064 12540
rect 14064 12484 14068 12540
rect 14004 12480 14068 12484
rect 14084 12540 14148 12544
rect 14084 12484 14088 12540
rect 14088 12484 14144 12540
rect 14144 12484 14148 12540
rect 14084 12480 14148 12484
rect 14164 12540 14228 12544
rect 14164 12484 14168 12540
rect 14168 12484 14224 12540
rect 14224 12484 14228 12540
rect 14164 12480 14228 12484
rect 14244 12540 14308 12544
rect 14244 12484 14248 12540
rect 14248 12484 14304 12540
rect 14304 12484 14308 12540
rect 14244 12480 14308 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 19465 12540 19529 12544
rect 19465 12484 19469 12540
rect 19469 12484 19525 12540
rect 19525 12484 19529 12540
rect 19465 12480 19529 12484
rect 3004 12276 3068 12340
rect 14412 12276 14476 12340
rect 4222 11996 4286 12000
rect 4222 11940 4226 11996
rect 4226 11940 4282 11996
rect 4282 11940 4286 11996
rect 4222 11936 4286 11940
rect 4302 11996 4366 12000
rect 4302 11940 4306 11996
rect 4306 11940 4362 11996
rect 4362 11940 4366 11996
rect 4302 11936 4366 11940
rect 4382 11996 4446 12000
rect 4382 11940 4386 11996
rect 4386 11940 4442 11996
rect 4442 11940 4446 11996
rect 4382 11936 4446 11940
rect 4462 11996 4526 12000
rect 4462 11940 4466 11996
rect 4466 11940 4522 11996
rect 4522 11940 4526 11996
rect 4462 11936 4526 11940
rect 9443 11996 9507 12000
rect 9443 11940 9447 11996
rect 9447 11940 9503 11996
rect 9503 11940 9507 11996
rect 9443 11936 9507 11940
rect 9523 11996 9587 12000
rect 9523 11940 9527 11996
rect 9527 11940 9583 11996
rect 9583 11940 9587 11996
rect 9523 11936 9587 11940
rect 9603 11996 9667 12000
rect 9603 11940 9607 11996
rect 9607 11940 9663 11996
rect 9663 11940 9667 11996
rect 9603 11936 9667 11940
rect 9683 11996 9747 12000
rect 9683 11940 9687 11996
rect 9687 11940 9743 11996
rect 9743 11940 9747 11996
rect 9683 11936 9747 11940
rect 14664 11996 14728 12000
rect 14664 11940 14668 11996
rect 14668 11940 14724 11996
rect 14724 11940 14728 11996
rect 14664 11936 14728 11940
rect 14744 11996 14808 12000
rect 14744 11940 14748 11996
rect 14748 11940 14804 11996
rect 14804 11940 14808 11996
rect 14744 11936 14808 11940
rect 14824 11996 14888 12000
rect 14824 11940 14828 11996
rect 14828 11940 14884 11996
rect 14884 11940 14888 11996
rect 14824 11936 14888 11940
rect 14904 11996 14968 12000
rect 14904 11940 14908 11996
rect 14908 11940 14964 11996
rect 14964 11940 14968 11996
rect 14904 11936 14968 11940
rect 19885 11996 19949 12000
rect 19885 11940 19889 11996
rect 19889 11940 19945 11996
rect 19945 11940 19949 11996
rect 19885 11936 19949 11940
rect 19965 11996 20029 12000
rect 19965 11940 19969 11996
rect 19969 11940 20025 11996
rect 20025 11940 20029 11996
rect 19965 11936 20029 11940
rect 20045 11996 20109 12000
rect 20045 11940 20049 11996
rect 20049 11940 20105 11996
rect 20105 11940 20109 11996
rect 20045 11936 20109 11940
rect 20125 11996 20189 12000
rect 20125 11940 20129 11996
rect 20129 11940 20185 11996
rect 20185 11940 20189 11996
rect 20125 11936 20189 11940
rect 3562 11452 3626 11456
rect 3562 11396 3566 11452
rect 3566 11396 3622 11452
rect 3622 11396 3626 11452
rect 3562 11392 3626 11396
rect 3642 11452 3706 11456
rect 3642 11396 3646 11452
rect 3646 11396 3702 11452
rect 3702 11396 3706 11452
rect 3642 11392 3706 11396
rect 3722 11452 3786 11456
rect 3722 11396 3726 11452
rect 3726 11396 3782 11452
rect 3782 11396 3786 11452
rect 3722 11392 3786 11396
rect 3802 11452 3866 11456
rect 3802 11396 3806 11452
rect 3806 11396 3862 11452
rect 3862 11396 3866 11452
rect 3802 11392 3866 11396
rect 8783 11452 8847 11456
rect 8783 11396 8787 11452
rect 8787 11396 8843 11452
rect 8843 11396 8847 11452
rect 8783 11392 8847 11396
rect 8863 11452 8927 11456
rect 8863 11396 8867 11452
rect 8867 11396 8923 11452
rect 8923 11396 8927 11452
rect 8863 11392 8927 11396
rect 8943 11452 9007 11456
rect 8943 11396 8947 11452
rect 8947 11396 9003 11452
rect 9003 11396 9007 11452
rect 8943 11392 9007 11396
rect 9023 11452 9087 11456
rect 9023 11396 9027 11452
rect 9027 11396 9083 11452
rect 9083 11396 9087 11452
rect 9023 11392 9087 11396
rect 14004 11452 14068 11456
rect 14004 11396 14008 11452
rect 14008 11396 14064 11452
rect 14064 11396 14068 11452
rect 14004 11392 14068 11396
rect 14084 11452 14148 11456
rect 14084 11396 14088 11452
rect 14088 11396 14144 11452
rect 14144 11396 14148 11452
rect 14084 11392 14148 11396
rect 14164 11452 14228 11456
rect 14164 11396 14168 11452
rect 14168 11396 14224 11452
rect 14224 11396 14228 11452
rect 14164 11392 14228 11396
rect 14244 11452 14308 11456
rect 14244 11396 14248 11452
rect 14248 11396 14304 11452
rect 14304 11396 14308 11452
rect 14244 11392 14308 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 19465 11452 19529 11456
rect 19465 11396 19469 11452
rect 19469 11396 19525 11452
rect 19525 11396 19529 11452
rect 19465 11392 19529 11396
rect 4222 10908 4286 10912
rect 4222 10852 4226 10908
rect 4226 10852 4282 10908
rect 4282 10852 4286 10908
rect 4222 10848 4286 10852
rect 4302 10908 4366 10912
rect 4302 10852 4306 10908
rect 4306 10852 4362 10908
rect 4362 10852 4366 10908
rect 4302 10848 4366 10852
rect 4382 10908 4446 10912
rect 4382 10852 4386 10908
rect 4386 10852 4442 10908
rect 4442 10852 4446 10908
rect 4382 10848 4446 10852
rect 4462 10908 4526 10912
rect 4462 10852 4466 10908
rect 4466 10852 4522 10908
rect 4522 10852 4526 10908
rect 4462 10848 4526 10852
rect 9443 10908 9507 10912
rect 9443 10852 9447 10908
rect 9447 10852 9503 10908
rect 9503 10852 9507 10908
rect 9443 10848 9507 10852
rect 9523 10908 9587 10912
rect 9523 10852 9527 10908
rect 9527 10852 9583 10908
rect 9583 10852 9587 10908
rect 9523 10848 9587 10852
rect 9603 10908 9667 10912
rect 9603 10852 9607 10908
rect 9607 10852 9663 10908
rect 9663 10852 9667 10908
rect 9603 10848 9667 10852
rect 9683 10908 9747 10912
rect 9683 10852 9687 10908
rect 9687 10852 9743 10908
rect 9743 10852 9747 10908
rect 9683 10848 9747 10852
rect 14664 10908 14728 10912
rect 14664 10852 14668 10908
rect 14668 10852 14724 10908
rect 14724 10852 14728 10908
rect 14664 10848 14728 10852
rect 14744 10908 14808 10912
rect 14744 10852 14748 10908
rect 14748 10852 14804 10908
rect 14804 10852 14808 10908
rect 14744 10848 14808 10852
rect 14824 10908 14888 10912
rect 14824 10852 14828 10908
rect 14828 10852 14884 10908
rect 14884 10852 14888 10908
rect 14824 10848 14888 10852
rect 14904 10908 14968 10912
rect 14904 10852 14908 10908
rect 14908 10852 14964 10908
rect 14964 10852 14968 10908
rect 14904 10848 14968 10852
rect 19885 10908 19949 10912
rect 19885 10852 19889 10908
rect 19889 10852 19945 10908
rect 19945 10852 19949 10908
rect 19885 10848 19949 10852
rect 19965 10908 20029 10912
rect 19965 10852 19969 10908
rect 19969 10852 20025 10908
rect 20025 10852 20029 10908
rect 19965 10848 20029 10852
rect 20045 10908 20109 10912
rect 20045 10852 20049 10908
rect 20049 10852 20105 10908
rect 20105 10852 20109 10908
rect 20045 10848 20109 10852
rect 20125 10908 20189 10912
rect 20125 10852 20129 10908
rect 20129 10852 20185 10908
rect 20185 10852 20189 10908
rect 20125 10848 20189 10852
rect 3562 10364 3626 10368
rect 3562 10308 3566 10364
rect 3566 10308 3622 10364
rect 3622 10308 3626 10364
rect 3562 10304 3626 10308
rect 3642 10364 3706 10368
rect 3642 10308 3646 10364
rect 3646 10308 3702 10364
rect 3702 10308 3706 10364
rect 3642 10304 3706 10308
rect 3722 10364 3786 10368
rect 3722 10308 3726 10364
rect 3726 10308 3782 10364
rect 3782 10308 3786 10364
rect 3722 10304 3786 10308
rect 3802 10364 3866 10368
rect 3802 10308 3806 10364
rect 3806 10308 3862 10364
rect 3862 10308 3866 10364
rect 3802 10304 3866 10308
rect 8783 10364 8847 10368
rect 8783 10308 8787 10364
rect 8787 10308 8843 10364
rect 8843 10308 8847 10364
rect 8783 10304 8847 10308
rect 8863 10364 8927 10368
rect 8863 10308 8867 10364
rect 8867 10308 8923 10364
rect 8923 10308 8927 10364
rect 8863 10304 8927 10308
rect 8943 10364 9007 10368
rect 8943 10308 8947 10364
rect 8947 10308 9003 10364
rect 9003 10308 9007 10364
rect 8943 10304 9007 10308
rect 9023 10364 9087 10368
rect 9023 10308 9027 10364
rect 9027 10308 9083 10364
rect 9083 10308 9087 10364
rect 9023 10304 9087 10308
rect 14004 10364 14068 10368
rect 14004 10308 14008 10364
rect 14008 10308 14064 10364
rect 14064 10308 14068 10364
rect 14004 10304 14068 10308
rect 14084 10364 14148 10368
rect 14084 10308 14088 10364
rect 14088 10308 14144 10364
rect 14144 10308 14148 10364
rect 14084 10304 14148 10308
rect 14164 10364 14228 10368
rect 14164 10308 14168 10364
rect 14168 10308 14224 10364
rect 14224 10308 14228 10364
rect 14164 10304 14228 10308
rect 14244 10364 14308 10368
rect 14244 10308 14248 10364
rect 14248 10308 14304 10364
rect 14304 10308 14308 10364
rect 14244 10304 14308 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 19465 10364 19529 10368
rect 19465 10308 19469 10364
rect 19469 10308 19525 10364
rect 19525 10308 19529 10364
rect 19465 10304 19529 10308
rect 4222 9820 4286 9824
rect 4222 9764 4226 9820
rect 4226 9764 4282 9820
rect 4282 9764 4286 9820
rect 4222 9760 4286 9764
rect 4302 9820 4366 9824
rect 4302 9764 4306 9820
rect 4306 9764 4362 9820
rect 4362 9764 4366 9820
rect 4302 9760 4366 9764
rect 4382 9820 4446 9824
rect 4382 9764 4386 9820
rect 4386 9764 4442 9820
rect 4442 9764 4446 9820
rect 4382 9760 4446 9764
rect 4462 9820 4526 9824
rect 4462 9764 4466 9820
rect 4466 9764 4522 9820
rect 4522 9764 4526 9820
rect 4462 9760 4526 9764
rect 9443 9820 9507 9824
rect 9443 9764 9447 9820
rect 9447 9764 9503 9820
rect 9503 9764 9507 9820
rect 9443 9760 9507 9764
rect 9523 9820 9587 9824
rect 9523 9764 9527 9820
rect 9527 9764 9583 9820
rect 9583 9764 9587 9820
rect 9523 9760 9587 9764
rect 9603 9820 9667 9824
rect 9603 9764 9607 9820
rect 9607 9764 9663 9820
rect 9663 9764 9667 9820
rect 9603 9760 9667 9764
rect 9683 9820 9747 9824
rect 9683 9764 9687 9820
rect 9687 9764 9743 9820
rect 9743 9764 9747 9820
rect 9683 9760 9747 9764
rect 14664 9820 14728 9824
rect 14664 9764 14668 9820
rect 14668 9764 14724 9820
rect 14724 9764 14728 9820
rect 14664 9760 14728 9764
rect 14744 9820 14808 9824
rect 14744 9764 14748 9820
rect 14748 9764 14804 9820
rect 14804 9764 14808 9820
rect 14744 9760 14808 9764
rect 14824 9820 14888 9824
rect 14824 9764 14828 9820
rect 14828 9764 14884 9820
rect 14884 9764 14888 9820
rect 14824 9760 14888 9764
rect 14904 9820 14968 9824
rect 14904 9764 14908 9820
rect 14908 9764 14964 9820
rect 14964 9764 14968 9820
rect 14904 9760 14968 9764
rect 19885 9820 19949 9824
rect 19885 9764 19889 9820
rect 19889 9764 19945 9820
rect 19945 9764 19949 9820
rect 19885 9760 19949 9764
rect 19965 9820 20029 9824
rect 19965 9764 19969 9820
rect 19969 9764 20025 9820
rect 20025 9764 20029 9820
rect 19965 9760 20029 9764
rect 20045 9820 20109 9824
rect 20045 9764 20049 9820
rect 20049 9764 20105 9820
rect 20105 9764 20109 9820
rect 20045 9760 20109 9764
rect 20125 9820 20189 9824
rect 20125 9764 20129 9820
rect 20129 9764 20185 9820
rect 20185 9764 20189 9820
rect 20125 9760 20189 9764
rect 3562 9276 3626 9280
rect 3562 9220 3566 9276
rect 3566 9220 3622 9276
rect 3622 9220 3626 9276
rect 3562 9216 3626 9220
rect 3642 9276 3706 9280
rect 3642 9220 3646 9276
rect 3646 9220 3702 9276
rect 3702 9220 3706 9276
rect 3642 9216 3706 9220
rect 3722 9276 3786 9280
rect 3722 9220 3726 9276
rect 3726 9220 3782 9276
rect 3782 9220 3786 9276
rect 3722 9216 3786 9220
rect 3802 9276 3866 9280
rect 3802 9220 3806 9276
rect 3806 9220 3862 9276
rect 3862 9220 3866 9276
rect 3802 9216 3866 9220
rect 8783 9276 8847 9280
rect 8783 9220 8787 9276
rect 8787 9220 8843 9276
rect 8843 9220 8847 9276
rect 8783 9216 8847 9220
rect 8863 9276 8927 9280
rect 8863 9220 8867 9276
rect 8867 9220 8923 9276
rect 8923 9220 8927 9276
rect 8863 9216 8927 9220
rect 8943 9276 9007 9280
rect 8943 9220 8947 9276
rect 8947 9220 9003 9276
rect 9003 9220 9007 9276
rect 8943 9216 9007 9220
rect 9023 9276 9087 9280
rect 9023 9220 9027 9276
rect 9027 9220 9083 9276
rect 9083 9220 9087 9276
rect 9023 9216 9087 9220
rect 14004 9276 14068 9280
rect 14004 9220 14008 9276
rect 14008 9220 14064 9276
rect 14064 9220 14068 9276
rect 14004 9216 14068 9220
rect 14084 9276 14148 9280
rect 14084 9220 14088 9276
rect 14088 9220 14144 9276
rect 14144 9220 14148 9276
rect 14084 9216 14148 9220
rect 14164 9276 14228 9280
rect 14164 9220 14168 9276
rect 14168 9220 14224 9276
rect 14224 9220 14228 9276
rect 14164 9216 14228 9220
rect 14244 9276 14308 9280
rect 14244 9220 14248 9276
rect 14248 9220 14304 9276
rect 14304 9220 14308 9276
rect 14244 9216 14308 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 19465 9276 19529 9280
rect 19465 9220 19469 9276
rect 19469 9220 19525 9276
rect 19525 9220 19529 9276
rect 19465 9216 19529 9220
rect 4222 8732 4286 8736
rect 4222 8676 4226 8732
rect 4226 8676 4282 8732
rect 4282 8676 4286 8732
rect 4222 8672 4286 8676
rect 4302 8732 4366 8736
rect 4302 8676 4306 8732
rect 4306 8676 4362 8732
rect 4362 8676 4366 8732
rect 4302 8672 4366 8676
rect 4382 8732 4446 8736
rect 4382 8676 4386 8732
rect 4386 8676 4442 8732
rect 4442 8676 4446 8732
rect 4382 8672 4446 8676
rect 4462 8732 4526 8736
rect 4462 8676 4466 8732
rect 4466 8676 4522 8732
rect 4522 8676 4526 8732
rect 4462 8672 4526 8676
rect 9443 8732 9507 8736
rect 9443 8676 9447 8732
rect 9447 8676 9503 8732
rect 9503 8676 9507 8732
rect 9443 8672 9507 8676
rect 9523 8732 9587 8736
rect 9523 8676 9527 8732
rect 9527 8676 9583 8732
rect 9583 8676 9587 8732
rect 9523 8672 9587 8676
rect 9603 8732 9667 8736
rect 9603 8676 9607 8732
rect 9607 8676 9663 8732
rect 9663 8676 9667 8732
rect 9603 8672 9667 8676
rect 9683 8732 9747 8736
rect 9683 8676 9687 8732
rect 9687 8676 9743 8732
rect 9743 8676 9747 8732
rect 9683 8672 9747 8676
rect 14664 8732 14728 8736
rect 14664 8676 14668 8732
rect 14668 8676 14724 8732
rect 14724 8676 14728 8732
rect 14664 8672 14728 8676
rect 14744 8732 14808 8736
rect 14744 8676 14748 8732
rect 14748 8676 14804 8732
rect 14804 8676 14808 8732
rect 14744 8672 14808 8676
rect 14824 8732 14888 8736
rect 14824 8676 14828 8732
rect 14828 8676 14884 8732
rect 14884 8676 14888 8732
rect 14824 8672 14888 8676
rect 14904 8732 14968 8736
rect 14904 8676 14908 8732
rect 14908 8676 14964 8732
rect 14964 8676 14968 8732
rect 14904 8672 14968 8676
rect 19885 8732 19949 8736
rect 19885 8676 19889 8732
rect 19889 8676 19945 8732
rect 19945 8676 19949 8732
rect 19885 8672 19949 8676
rect 19965 8732 20029 8736
rect 19965 8676 19969 8732
rect 19969 8676 20025 8732
rect 20025 8676 20029 8732
rect 19965 8672 20029 8676
rect 20045 8732 20109 8736
rect 20045 8676 20049 8732
rect 20049 8676 20105 8732
rect 20105 8676 20109 8732
rect 20045 8672 20109 8676
rect 20125 8732 20189 8736
rect 20125 8676 20129 8732
rect 20129 8676 20185 8732
rect 20185 8676 20189 8732
rect 20125 8672 20189 8676
rect 14412 8528 14476 8532
rect 14412 8472 14462 8528
rect 14462 8472 14476 8528
rect 14412 8468 14476 8472
rect 3562 8188 3626 8192
rect 3562 8132 3566 8188
rect 3566 8132 3622 8188
rect 3622 8132 3626 8188
rect 3562 8128 3626 8132
rect 3642 8188 3706 8192
rect 3642 8132 3646 8188
rect 3646 8132 3702 8188
rect 3702 8132 3706 8188
rect 3642 8128 3706 8132
rect 3722 8188 3786 8192
rect 3722 8132 3726 8188
rect 3726 8132 3782 8188
rect 3782 8132 3786 8188
rect 3722 8128 3786 8132
rect 3802 8188 3866 8192
rect 3802 8132 3806 8188
rect 3806 8132 3862 8188
rect 3862 8132 3866 8188
rect 3802 8128 3866 8132
rect 8783 8188 8847 8192
rect 8783 8132 8787 8188
rect 8787 8132 8843 8188
rect 8843 8132 8847 8188
rect 8783 8128 8847 8132
rect 8863 8188 8927 8192
rect 8863 8132 8867 8188
rect 8867 8132 8923 8188
rect 8923 8132 8927 8188
rect 8863 8128 8927 8132
rect 8943 8188 9007 8192
rect 8943 8132 8947 8188
rect 8947 8132 9003 8188
rect 9003 8132 9007 8188
rect 8943 8128 9007 8132
rect 9023 8188 9087 8192
rect 9023 8132 9027 8188
rect 9027 8132 9083 8188
rect 9083 8132 9087 8188
rect 9023 8128 9087 8132
rect 14004 8188 14068 8192
rect 14004 8132 14008 8188
rect 14008 8132 14064 8188
rect 14064 8132 14068 8188
rect 14004 8128 14068 8132
rect 14084 8188 14148 8192
rect 14084 8132 14088 8188
rect 14088 8132 14144 8188
rect 14144 8132 14148 8188
rect 14084 8128 14148 8132
rect 14164 8188 14228 8192
rect 14164 8132 14168 8188
rect 14168 8132 14224 8188
rect 14224 8132 14228 8188
rect 14164 8128 14228 8132
rect 14244 8188 14308 8192
rect 14244 8132 14248 8188
rect 14248 8132 14304 8188
rect 14304 8132 14308 8188
rect 14244 8128 14308 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 19465 8188 19529 8192
rect 19465 8132 19469 8188
rect 19469 8132 19525 8188
rect 19525 8132 19529 8188
rect 19465 8128 19529 8132
rect 4222 7644 4286 7648
rect 4222 7588 4226 7644
rect 4226 7588 4282 7644
rect 4282 7588 4286 7644
rect 4222 7584 4286 7588
rect 4302 7644 4366 7648
rect 4302 7588 4306 7644
rect 4306 7588 4362 7644
rect 4362 7588 4366 7644
rect 4302 7584 4366 7588
rect 4382 7644 4446 7648
rect 4382 7588 4386 7644
rect 4386 7588 4442 7644
rect 4442 7588 4446 7644
rect 4382 7584 4446 7588
rect 4462 7644 4526 7648
rect 4462 7588 4466 7644
rect 4466 7588 4522 7644
rect 4522 7588 4526 7644
rect 4462 7584 4526 7588
rect 9443 7644 9507 7648
rect 9443 7588 9447 7644
rect 9447 7588 9503 7644
rect 9503 7588 9507 7644
rect 9443 7584 9507 7588
rect 9523 7644 9587 7648
rect 9523 7588 9527 7644
rect 9527 7588 9583 7644
rect 9583 7588 9587 7644
rect 9523 7584 9587 7588
rect 9603 7644 9667 7648
rect 9603 7588 9607 7644
rect 9607 7588 9663 7644
rect 9663 7588 9667 7644
rect 9603 7584 9667 7588
rect 9683 7644 9747 7648
rect 9683 7588 9687 7644
rect 9687 7588 9743 7644
rect 9743 7588 9747 7644
rect 9683 7584 9747 7588
rect 14664 7644 14728 7648
rect 14664 7588 14668 7644
rect 14668 7588 14724 7644
rect 14724 7588 14728 7644
rect 14664 7584 14728 7588
rect 14744 7644 14808 7648
rect 14744 7588 14748 7644
rect 14748 7588 14804 7644
rect 14804 7588 14808 7644
rect 14744 7584 14808 7588
rect 14824 7644 14888 7648
rect 14824 7588 14828 7644
rect 14828 7588 14884 7644
rect 14884 7588 14888 7644
rect 14824 7584 14888 7588
rect 14904 7644 14968 7648
rect 14904 7588 14908 7644
rect 14908 7588 14964 7644
rect 14964 7588 14968 7644
rect 14904 7584 14968 7588
rect 19885 7644 19949 7648
rect 19885 7588 19889 7644
rect 19889 7588 19945 7644
rect 19945 7588 19949 7644
rect 19885 7584 19949 7588
rect 19965 7644 20029 7648
rect 19965 7588 19969 7644
rect 19969 7588 20025 7644
rect 20025 7588 20029 7644
rect 19965 7584 20029 7588
rect 20045 7644 20109 7648
rect 20045 7588 20049 7644
rect 20049 7588 20105 7644
rect 20105 7588 20109 7644
rect 20045 7584 20109 7588
rect 20125 7644 20189 7648
rect 20125 7588 20129 7644
rect 20129 7588 20185 7644
rect 20185 7588 20189 7644
rect 20125 7584 20189 7588
rect 3562 7100 3626 7104
rect 3562 7044 3566 7100
rect 3566 7044 3622 7100
rect 3622 7044 3626 7100
rect 3562 7040 3626 7044
rect 3642 7100 3706 7104
rect 3642 7044 3646 7100
rect 3646 7044 3702 7100
rect 3702 7044 3706 7100
rect 3642 7040 3706 7044
rect 3722 7100 3786 7104
rect 3722 7044 3726 7100
rect 3726 7044 3782 7100
rect 3782 7044 3786 7100
rect 3722 7040 3786 7044
rect 3802 7100 3866 7104
rect 3802 7044 3806 7100
rect 3806 7044 3862 7100
rect 3862 7044 3866 7100
rect 3802 7040 3866 7044
rect 8783 7100 8847 7104
rect 8783 7044 8787 7100
rect 8787 7044 8843 7100
rect 8843 7044 8847 7100
rect 8783 7040 8847 7044
rect 8863 7100 8927 7104
rect 8863 7044 8867 7100
rect 8867 7044 8923 7100
rect 8923 7044 8927 7100
rect 8863 7040 8927 7044
rect 8943 7100 9007 7104
rect 8943 7044 8947 7100
rect 8947 7044 9003 7100
rect 9003 7044 9007 7100
rect 8943 7040 9007 7044
rect 9023 7100 9087 7104
rect 9023 7044 9027 7100
rect 9027 7044 9083 7100
rect 9083 7044 9087 7100
rect 9023 7040 9087 7044
rect 14004 7100 14068 7104
rect 14004 7044 14008 7100
rect 14008 7044 14064 7100
rect 14064 7044 14068 7100
rect 14004 7040 14068 7044
rect 14084 7100 14148 7104
rect 14084 7044 14088 7100
rect 14088 7044 14144 7100
rect 14144 7044 14148 7100
rect 14084 7040 14148 7044
rect 14164 7100 14228 7104
rect 14164 7044 14168 7100
rect 14168 7044 14224 7100
rect 14224 7044 14228 7100
rect 14164 7040 14228 7044
rect 14244 7100 14308 7104
rect 14244 7044 14248 7100
rect 14248 7044 14304 7100
rect 14304 7044 14308 7100
rect 14244 7040 14308 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 19465 7100 19529 7104
rect 19465 7044 19469 7100
rect 19469 7044 19525 7100
rect 19525 7044 19529 7100
rect 19465 7040 19529 7044
rect 4222 6556 4286 6560
rect 4222 6500 4226 6556
rect 4226 6500 4282 6556
rect 4282 6500 4286 6556
rect 4222 6496 4286 6500
rect 4302 6556 4366 6560
rect 4302 6500 4306 6556
rect 4306 6500 4362 6556
rect 4362 6500 4366 6556
rect 4302 6496 4366 6500
rect 4382 6556 4446 6560
rect 4382 6500 4386 6556
rect 4386 6500 4442 6556
rect 4442 6500 4446 6556
rect 4382 6496 4446 6500
rect 4462 6556 4526 6560
rect 4462 6500 4466 6556
rect 4466 6500 4522 6556
rect 4522 6500 4526 6556
rect 4462 6496 4526 6500
rect 9443 6556 9507 6560
rect 9443 6500 9447 6556
rect 9447 6500 9503 6556
rect 9503 6500 9507 6556
rect 9443 6496 9507 6500
rect 9523 6556 9587 6560
rect 9523 6500 9527 6556
rect 9527 6500 9583 6556
rect 9583 6500 9587 6556
rect 9523 6496 9587 6500
rect 9603 6556 9667 6560
rect 9603 6500 9607 6556
rect 9607 6500 9663 6556
rect 9663 6500 9667 6556
rect 9603 6496 9667 6500
rect 9683 6556 9747 6560
rect 9683 6500 9687 6556
rect 9687 6500 9743 6556
rect 9743 6500 9747 6556
rect 9683 6496 9747 6500
rect 14664 6556 14728 6560
rect 14664 6500 14668 6556
rect 14668 6500 14724 6556
rect 14724 6500 14728 6556
rect 14664 6496 14728 6500
rect 14744 6556 14808 6560
rect 14744 6500 14748 6556
rect 14748 6500 14804 6556
rect 14804 6500 14808 6556
rect 14744 6496 14808 6500
rect 14824 6556 14888 6560
rect 14824 6500 14828 6556
rect 14828 6500 14884 6556
rect 14884 6500 14888 6556
rect 14824 6496 14888 6500
rect 14904 6556 14968 6560
rect 14904 6500 14908 6556
rect 14908 6500 14964 6556
rect 14964 6500 14968 6556
rect 14904 6496 14968 6500
rect 19885 6556 19949 6560
rect 19885 6500 19889 6556
rect 19889 6500 19945 6556
rect 19945 6500 19949 6556
rect 19885 6496 19949 6500
rect 19965 6556 20029 6560
rect 19965 6500 19969 6556
rect 19969 6500 20025 6556
rect 20025 6500 20029 6556
rect 19965 6496 20029 6500
rect 20045 6556 20109 6560
rect 20045 6500 20049 6556
rect 20049 6500 20105 6556
rect 20105 6500 20109 6556
rect 20045 6496 20109 6500
rect 20125 6556 20189 6560
rect 20125 6500 20129 6556
rect 20129 6500 20185 6556
rect 20185 6500 20189 6556
rect 20125 6496 20189 6500
rect 14412 6428 14476 6492
rect 3562 6012 3626 6016
rect 3562 5956 3566 6012
rect 3566 5956 3622 6012
rect 3622 5956 3626 6012
rect 3562 5952 3626 5956
rect 3642 6012 3706 6016
rect 3642 5956 3646 6012
rect 3646 5956 3702 6012
rect 3702 5956 3706 6012
rect 3642 5952 3706 5956
rect 3722 6012 3786 6016
rect 3722 5956 3726 6012
rect 3726 5956 3782 6012
rect 3782 5956 3786 6012
rect 3722 5952 3786 5956
rect 3802 6012 3866 6016
rect 3802 5956 3806 6012
rect 3806 5956 3862 6012
rect 3862 5956 3866 6012
rect 3802 5952 3866 5956
rect 8783 6012 8847 6016
rect 8783 5956 8787 6012
rect 8787 5956 8843 6012
rect 8843 5956 8847 6012
rect 8783 5952 8847 5956
rect 8863 6012 8927 6016
rect 8863 5956 8867 6012
rect 8867 5956 8923 6012
rect 8923 5956 8927 6012
rect 8863 5952 8927 5956
rect 8943 6012 9007 6016
rect 8943 5956 8947 6012
rect 8947 5956 9003 6012
rect 9003 5956 9007 6012
rect 8943 5952 9007 5956
rect 9023 6012 9087 6016
rect 9023 5956 9027 6012
rect 9027 5956 9083 6012
rect 9083 5956 9087 6012
rect 9023 5952 9087 5956
rect 14004 6012 14068 6016
rect 14004 5956 14008 6012
rect 14008 5956 14064 6012
rect 14064 5956 14068 6012
rect 14004 5952 14068 5956
rect 14084 6012 14148 6016
rect 14084 5956 14088 6012
rect 14088 5956 14144 6012
rect 14144 5956 14148 6012
rect 14084 5952 14148 5956
rect 14164 6012 14228 6016
rect 14164 5956 14168 6012
rect 14168 5956 14224 6012
rect 14224 5956 14228 6012
rect 14164 5952 14228 5956
rect 14244 6012 14308 6016
rect 14244 5956 14248 6012
rect 14248 5956 14304 6012
rect 14304 5956 14308 6012
rect 14244 5952 14308 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 19465 6012 19529 6016
rect 19465 5956 19469 6012
rect 19469 5956 19525 6012
rect 19525 5956 19529 6012
rect 19465 5952 19529 5956
rect 4222 5468 4286 5472
rect 4222 5412 4226 5468
rect 4226 5412 4282 5468
rect 4282 5412 4286 5468
rect 4222 5408 4286 5412
rect 4302 5468 4366 5472
rect 4302 5412 4306 5468
rect 4306 5412 4362 5468
rect 4362 5412 4366 5468
rect 4302 5408 4366 5412
rect 4382 5468 4446 5472
rect 4382 5412 4386 5468
rect 4386 5412 4442 5468
rect 4442 5412 4446 5468
rect 4382 5408 4446 5412
rect 4462 5468 4526 5472
rect 4462 5412 4466 5468
rect 4466 5412 4522 5468
rect 4522 5412 4526 5468
rect 4462 5408 4526 5412
rect 9443 5468 9507 5472
rect 9443 5412 9447 5468
rect 9447 5412 9503 5468
rect 9503 5412 9507 5468
rect 9443 5408 9507 5412
rect 9523 5468 9587 5472
rect 9523 5412 9527 5468
rect 9527 5412 9583 5468
rect 9583 5412 9587 5468
rect 9523 5408 9587 5412
rect 9603 5468 9667 5472
rect 9603 5412 9607 5468
rect 9607 5412 9663 5468
rect 9663 5412 9667 5468
rect 9603 5408 9667 5412
rect 9683 5468 9747 5472
rect 9683 5412 9687 5468
rect 9687 5412 9743 5468
rect 9743 5412 9747 5468
rect 9683 5408 9747 5412
rect 14664 5468 14728 5472
rect 14664 5412 14668 5468
rect 14668 5412 14724 5468
rect 14724 5412 14728 5468
rect 14664 5408 14728 5412
rect 14744 5468 14808 5472
rect 14744 5412 14748 5468
rect 14748 5412 14804 5468
rect 14804 5412 14808 5468
rect 14744 5408 14808 5412
rect 14824 5468 14888 5472
rect 14824 5412 14828 5468
rect 14828 5412 14884 5468
rect 14884 5412 14888 5468
rect 14824 5408 14888 5412
rect 14904 5468 14968 5472
rect 14904 5412 14908 5468
rect 14908 5412 14964 5468
rect 14964 5412 14968 5468
rect 14904 5408 14968 5412
rect 19885 5468 19949 5472
rect 19885 5412 19889 5468
rect 19889 5412 19945 5468
rect 19945 5412 19949 5468
rect 19885 5408 19949 5412
rect 19965 5468 20029 5472
rect 19965 5412 19969 5468
rect 19969 5412 20025 5468
rect 20025 5412 20029 5468
rect 19965 5408 20029 5412
rect 20045 5468 20109 5472
rect 20045 5412 20049 5468
rect 20049 5412 20105 5468
rect 20105 5412 20109 5468
rect 20045 5408 20109 5412
rect 20125 5468 20189 5472
rect 20125 5412 20129 5468
rect 20129 5412 20185 5468
rect 20185 5412 20189 5468
rect 20125 5408 20189 5412
rect 3562 4924 3626 4928
rect 3562 4868 3566 4924
rect 3566 4868 3622 4924
rect 3622 4868 3626 4924
rect 3562 4864 3626 4868
rect 3642 4924 3706 4928
rect 3642 4868 3646 4924
rect 3646 4868 3702 4924
rect 3702 4868 3706 4924
rect 3642 4864 3706 4868
rect 3722 4924 3786 4928
rect 3722 4868 3726 4924
rect 3726 4868 3782 4924
rect 3782 4868 3786 4924
rect 3722 4864 3786 4868
rect 3802 4924 3866 4928
rect 3802 4868 3806 4924
rect 3806 4868 3862 4924
rect 3862 4868 3866 4924
rect 3802 4864 3866 4868
rect 8783 4924 8847 4928
rect 8783 4868 8787 4924
rect 8787 4868 8843 4924
rect 8843 4868 8847 4924
rect 8783 4864 8847 4868
rect 8863 4924 8927 4928
rect 8863 4868 8867 4924
rect 8867 4868 8923 4924
rect 8923 4868 8927 4924
rect 8863 4864 8927 4868
rect 8943 4924 9007 4928
rect 8943 4868 8947 4924
rect 8947 4868 9003 4924
rect 9003 4868 9007 4924
rect 8943 4864 9007 4868
rect 9023 4924 9087 4928
rect 9023 4868 9027 4924
rect 9027 4868 9083 4924
rect 9083 4868 9087 4924
rect 9023 4864 9087 4868
rect 14004 4924 14068 4928
rect 14004 4868 14008 4924
rect 14008 4868 14064 4924
rect 14064 4868 14068 4924
rect 14004 4864 14068 4868
rect 14084 4924 14148 4928
rect 14084 4868 14088 4924
rect 14088 4868 14144 4924
rect 14144 4868 14148 4924
rect 14084 4864 14148 4868
rect 14164 4924 14228 4928
rect 14164 4868 14168 4924
rect 14168 4868 14224 4924
rect 14224 4868 14228 4924
rect 14164 4864 14228 4868
rect 14244 4924 14308 4928
rect 14244 4868 14248 4924
rect 14248 4868 14304 4924
rect 14304 4868 14308 4924
rect 14244 4864 14308 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 19465 4924 19529 4928
rect 19465 4868 19469 4924
rect 19469 4868 19525 4924
rect 19525 4868 19529 4924
rect 19465 4864 19529 4868
rect 4222 4380 4286 4384
rect 4222 4324 4226 4380
rect 4226 4324 4282 4380
rect 4282 4324 4286 4380
rect 4222 4320 4286 4324
rect 4302 4380 4366 4384
rect 4302 4324 4306 4380
rect 4306 4324 4362 4380
rect 4362 4324 4366 4380
rect 4302 4320 4366 4324
rect 4382 4380 4446 4384
rect 4382 4324 4386 4380
rect 4386 4324 4442 4380
rect 4442 4324 4446 4380
rect 4382 4320 4446 4324
rect 4462 4380 4526 4384
rect 4462 4324 4466 4380
rect 4466 4324 4522 4380
rect 4522 4324 4526 4380
rect 4462 4320 4526 4324
rect 9443 4380 9507 4384
rect 9443 4324 9447 4380
rect 9447 4324 9503 4380
rect 9503 4324 9507 4380
rect 9443 4320 9507 4324
rect 9523 4380 9587 4384
rect 9523 4324 9527 4380
rect 9527 4324 9583 4380
rect 9583 4324 9587 4380
rect 9523 4320 9587 4324
rect 9603 4380 9667 4384
rect 9603 4324 9607 4380
rect 9607 4324 9663 4380
rect 9663 4324 9667 4380
rect 9603 4320 9667 4324
rect 9683 4380 9747 4384
rect 9683 4324 9687 4380
rect 9687 4324 9743 4380
rect 9743 4324 9747 4380
rect 9683 4320 9747 4324
rect 14664 4380 14728 4384
rect 14664 4324 14668 4380
rect 14668 4324 14724 4380
rect 14724 4324 14728 4380
rect 14664 4320 14728 4324
rect 14744 4380 14808 4384
rect 14744 4324 14748 4380
rect 14748 4324 14804 4380
rect 14804 4324 14808 4380
rect 14744 4320 14808 4324
rect 14824 4380 14888 4384
rect 14824 4324 14828 4380
rect 14828 4324 14884 4380
rect 14884 4324 14888 4380
rect 14824 4320 14888 4324
rect 14904 4380 14968 4384
rect 14904 4324 14908 4380
rect 14908 4324 14964 4380
rect 14964 4324 14968 4380
rect 14904 4320 14968 4324
rect 19885 4380 19949 4384
rect 19885 4324 19889 4380
rect 19889 4324 19945 4380
rect 19945 4324 19949 4380
rect 19885 4320 19949 4324
rect 19965 4380 20029 4384
rect 19965 4324 19969 4380
rect 19969 4324 20025 4380
rect 20025 4324 20029 4380
rect 19965 4320 20029 4324
rect 20045 4380 20109 4384
rect 20045 4324 20049 4380
rect 20049 4324 20105 4380
rect 20105 4324 20109 4380
rect 20045 4320 20109 4324
rect 20125 4380 20189 4384
rect 20125 4324 20129 4380
rect 20129 4324 20185 4380
rect 20185 4324 20189 4380
rect 20125 4320 20189 4324
rect 3562 3836 3626 3840
rect 3562 3780 3566 3836
rect 3566 3780 3622 3836
rect 3622 3780 3626 3836
rect 3562 3776 3626 3780
rect 3642 3836 3706 3840
rect 3642 3780 3646 3836
rect 3646 3780 3702 3836
rect 3702 3780 3706 3836
rect 3642 3776 3706 3780
rect 3722 3836 3786 3840
rect 3722 3780 3726 3836
rect 3726 3780 3782 3836
rect 3782 3780 3786 3836
rect 3722 3776 3786 3780
rect 3802 3836 3866 3840
rect 3802 3780 3806 3836
rect 3806 3780 3862 3836
rect 3862 3780 3866 3836
rect 3802 3776 3866 3780
rect 8783 3836 8847 3840
rect 8783 3780 8787 3836
rect 8787 3780 8843 3836
rect 8843 3780 8847 3836
rect 8783 3776 8847 3780
rect 8863 3836 8927 3840
rect 8863 3780 8867 3836
rect 8867 3780 8923 3836
rect 8923 3780 8927 3836
rect 8863 3776 8927 3780
rect 8943 3836 9007 3840
rect 8943 3780 8947 3836
rect 8947 3780 9003 3836
rect 9003 3780 9007 3836
rect 8943 3776 9007 3780
rect 9023 3836 9087 3840
rect 9023 3780 9027 3836
rect 9027 3780 9083 3836
rect 9083 3780 9087 3836
rect 9023 3776 9087 3780
rect 14004 3836 14068 3840
rect 14004 3780 14008 3836
rect 14008 3780 14064 3836
rect 14064 3780 14068 3836
rect 14004 3776 14068 3780
rect 14084 3836 14148 3840
rect 14084 3780 14088 3836
rect 14088 3780 14144 3836
rect 14144 3780 14148 3836
rect 14084 3776 14148 3780
rect 14164 3836 14228 3840
rect 14164 3780 14168 3836
rect 14168 3780 14224 3836
rect 14224 3780 14228 3836
rect 14164 3776 14228 3780
rect 14244 3836 14308 3840
rect 14244 3780 14248 3836
rect 14248 3780 14304 3836
rect 14304 3780 14308 3836
rect 14244 3776 14308 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 19465 3836 19529 3840
rect 19465 3780 19469 3836
rect 19469 3780 19525 3836
rect 19525 3780 19529 3836
rect 19465 3776 19529 3780
rect 4222 3292 4286 3296
rect 4222 3236 4226 3292
rect 4226 3236 4282 3292
rect 4282 3236 4286 3292
rect 4222 3232 4286 3236
rect 4302 3292 4366 3296
rect 4302 3236 4306 3292
rect 4306 3236 4362 3292
rect 4362 3236 4366 3292
rect 4302 3232 4366 3236
rect 4382 3292 4446 3296
rect 4382 3236 4386 3292
rect 4386 3236 4442 3292
rect 4442 3236 4446 3292
rect 4382 3232 4446 3236
rect 4462 3292 4526 3296
rect 4462 3236 4466 3292
rect 4466 3236 4522 3292
rect 4522 3236 4526 3292
rect 4462 3232 4526 3236
rect 9443 3292 9507 3296
rect 9443 3236 9447 3292
rect 9447 3236 9503 3292
rect 9503 3236 9507 3292
rect 9443 3232 9507 3236
rect 9523 3292 9587 3296
rect 9523 3236 9527 3292
rect 9527 3236 9583 3292
rect 9583 3236 9587 3292
rect 9523 3232 9587 3236
rect 9603 3292 9667 3296
rect 9603 3236 9607 3292
rect 9607 3236 9663 3292
rect 9663 3236 9667 3292
rect 9603 3232 9667 3236
rect 9683 3292 9747 3296
rect 9683 3236 9687 3292
rect 9687 3236 9743 3292
rect 9743 3236 9747 3292
rect 9683 3232 9747 3236
rect 14664 3292 14728 3296
rect 14664 3236 14668 3292
rect 14668 3236 14724 3292
rect 14724 3236 14728 3292
rect 14664 3232 14728 3236
rect 14744 3292 14808 3296
rect 14744 3236 14748 3292
rect 14748 3236 14804 3292
rect 14804 3236 14808 3292
rect 14744 3232 14808 3236
rect 14824 3292 14888 3296
rect 14824 3236 14828 3292
rect 14828 3236 14884 3292
rect 14884 3236 14888 3292
rect 14824 3232 14888 3236
rect 14904 3292 14968 3296
rect 14904 3236 14908 3292
rect 14908 3236 14964 3292
rect 14964 3236 14968 3292
rect 14904 3232 14968 3236
rect 19885 3292 19949 3296
rect 19885 3236 19889 3292
rect 19889 3236 19945 3292
rect 19945 3236 19949 3292
rect 19885 3232 19949 3236
rect 19965 3292 20029 3296
rect 19965 3236 19969 3292
rect 19969 3236 20025 3292
rect 20025 3236 20029 3292
rect 19965 3232 20029 3236
rect 20045 3292 20109 3296
rect 20045 3236 20049 3292
rect 20049 3236 20105 3292
rect 20105 3236 20109 3292
rect 20045 3232 20109 3236
rect 20125 3292 20189 3296
rect 20125 3236 20129 3292
rect 20129 3236 20185 3292
rect 20185 3236 20189 3292
rect 20125 3232 20189 3236
rect 3562 2748 3626 2752
rect 3562 2692 3566 2748
rect 3566 2692 3622 2748
rect 3622 2692 3626 2748
rect 3562 2688 3626 2692
rect 3642 2748 3706 2752
rect 3642 2692 3646 2748
rect 3646 2692 3702 2748
rect 3702 2692 3706 2748
rect 3642 2688 3706 2692
rect 3722 2748 3786 2752
rect 3722 2692 3726 2748
rect 3726 2692 3782 2748
rect 3782 2692 3786 2748
rect 3722 2688 3786 2692
rect 3802 2748 3866 2752
rect 3802 2692 3806 2748
rect 3806 2692 3862 2748
rect 3862 2692 3866 2748
rect 3802 2688 3866 2692
rect 8783 2748 8847 2752
rect 8783 2692 8787 2748
rect 8787 2692 8843 2748
rect 8843 2692 8847 2748
rect 8783 2688 8847 2692
rect 8863 2748 8927 2752
rect 8863 2692 8867 2748
rect 8867 2692 8923 2748
rect 8923 2692 8927 2748
rect 8863 2688 8927 2692
rect 8943 2748 9007 2752
rect 8943 2692 8947 2748
rect 8947 2692 9003 2748
rect 9003 2692 9007 2748
rect 8943 2688 9007 2692
rect 9023 2748 9087 2752
rect 9023 2692 9027 2748
rect 9027 2692 9083 2748
rect 9083 2692 9087 2748
rect 9023 2688 9087 2692
rect 14004 2748 14068 2752
rect 14004 2692 14008 2748
rect 14008 2692 14064 2748
rect 14064 2692 14068 2748
rect 14004 2688 14068 2692
rect 14084 2748 14148 2752
rect 14084 2692 14088 2748
rect 14088 2692 14144 2748
rect 14144 2692 14148 2748
rect 14084 2688 14148 2692
rect 14164 2748 14228 2752
rect 14164 2692 14168 2748
rect 14168 2692 14224 2748
rect 14224 2692 14228 2748
rect 14164 2688 14228 2692
rect 14244 2748 14308 2752
rect 14244 2692 14248 2748
rect 14248 2692 14304 2748
rect 14304 2692 14308 2748
rect 14244 2688 14308 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 19465 2748 19529 2752
rect 19465 2692 19469 2748
rect 19469 2692 19525 2748
rect 19525 2692 19529 2748
rect 19465 2688 19529 2692
rect 4222 2204 4286 2208
rect 4222 2148 4226 2204
rect 4226 2148 4282 2204
rect 4282 2148 4286 2204
rect 4222 2144 4286 2148
rect 4302 2204 4366 2208
rect 4302 2148 4306 2204
rect 4306 2148 4362 2204
rect 4362 2148 4366 2204
rect 4302 2144 4366 2148
rect 4382 2204 4446 2208
rect 4382 2148 4386 2204
rect 4386 2148 4442 2204
rect 4442 2148 4446 2204
rect 4382 2144 4446 2148
rect 4462 2204 4526 2208
rect 4462 2148 4466 2204
rect 4466 2148 4522 2204
rect 4522 2148 4526 2204
rect 4462 2144 4526 2148
rect 9443 2204 9507 2208
rect 9443 2148 9447 2204
rect 9447 2148 9503 2204
rect 9503 2148 9507 2204
rect 9443 2144 9507 2148
rect 9523 2204 9587 2208
rect 9523 2148 9527 2204
rect 9527 2148 9583 2204
rect 9583 2148 9587 2204
rect 9523 2144 9587 2148
rect 9603 2204 9667 2208
rect 9603 2148 9607 2204
rect 9607 2148 9663 2204
rect 9663 2148 9667 2204
rect 9603 2144 9667 2148
rect 9683 2204 9747 2208
rect 9683 2148 9687 2204
rect 9687 2148 9743 2204
rect 9743 2148 9747 2204
rect 9683 2144 9747 2148
rect 14664 2204 14728 2208
rect 14664 2148 14668 2204
rect 14668 2148 14724 2204
rect 14724 2148 14728 2204
rect 14664 2144 14728 2148
rect 14744 2204 14808 2208
rect 14744 2148 14748 2204
rect 14748 2148 14804 2204
rect 14804 2148 14808 2204
rect 14744 2144 14808 2148
rect 14824 2204 14888 2208
rect 14824 2148 14828 2204
rect 14828 2148 14884 2204
rect 14884 2148 14888 2204
rect 14824 2144 14888 2148
rect 14904 2204 14968 2208
rect 14904 2148 14908 2204
rect 14908 2148 14964 2204
rect 14964 2148 14968 2204
rect 14904 2144 14968 2148
rect 19885 2204 19949 2208
rect 19885 2148 19889 2204
rect 19889 2148 19945 2204
rect 19945 2148 19949 2204
rect 19885 2144 19949 2148
rect 19965 2204 20029 2208
rect 19965 2148 19969 2204
rect 19969 2148 20025 2204
rect 20025 2148 20029 2204
rect 19965 2144 20029 2148
rect 20045 2204 20109 2208
rect 20045 2148 20049 2204
rect 20049 2148 20105 2204
rect 20105 2148 20109 2204
rect 20045 2144 20109 2148
rect 20125 2204 20189 2208
rect 20125 2148 20129 2204
rect 20129 2148 20185 2204
rect 20185 2148 20189 2204
rect 20125 2144 20189 2148
<< metal4 >>
rect 3554 22336 3874 22896
rect 3554 22272 3562 22336
rect 3626 22272 3642 22336
rect 3706 22272 3722 22336
rect 3786 22272 3802 22336
rect 3866 22272 3874 22336
rect 3554 21248 3874 22272
rect 3554 21184 3562 21248
rect 3626 21184 3642 21248
rect 3706 21184 3722 21248
rect 3786 21184 3802 21248
rect 3866 21184 3874 21248
rect 3003 21180 3069 21181
rect 3003 21116 3004 21180
rect 3068 21116 3069 21180
rect 3003 21115 3069 21116
rect 3006 12341 3066 21115
rect 3554 20382 3874 21184
rect 3554 20160 3596 20382
rect 3832 20160 3874 20382
rect 3554 20096 3562 20160
rect 3626 20096 3642 20146
rect 3706 20096 3722 20146
rect 3786 20096 3802 20146
rect 3866 20096 3874 20160
rect 3554 19072 3874 20096
rect 3554 19008 3562 19072
rect 3626 19008 3642 19072
rect 3706 19008 3722 19072
rect 3786 19008 3802 19072
rect 3866 19008 3874 19072
rect 3554 17984 3874 19008
rect 3554 17920 3562 17984
rect 3626 17920 3642 17984
rect 3706 17920 3722 17984
rect 3786 17920 3802 17984
rect 3866 17920 3874 17984
rect 3554 16896 3874 17920
rect 3554 16832 3562 16896
rect 3626 16832 3642 16896
rect 3706 16832 3722 16896
rect 3786 16832 3802 16896
rect 3866 16832 3874 16896
rect 3554 15808 3874 16832
rect 3554 15744 3562 15808
rect 3626 15744 3642 15808
rect 3706 15744 3722 15808
rect 3786 15744 3802 15808
rect 3866 15744 3874 15808
rect 3554 15214 3874 15744
rect 3554 14978 3596 15214
rect 3832 14978 3874 15214
rect 3554 14720 3874 14978
rect 3554 14656 3562 14720
rect 3626 14656 3642 14720
rect 3706 14656 3722 14720
rect 3786 14656 3802 14720
rect 3866 14656 3874 14720
rect 3554 13632 3874 14656
rect 3554 13568 3562 13632
rect 3626 13568 3642 13632
rect 3706 13568 3722 13632
rect 3786 13568 3802 13632
rect 3866 13568 3874 13632
rect 3554 12544 3874 13568
rect 3554 12480 3562 12544
rect 3626 12480 3642 12544
rect 3706 12480 3722 12544
rect 3786 12480 3802 12544
rect 3866 12480 3874 12544
rect 3003 12340 3069 12341
rect 3003 12276 3004 12340
rect 3068 12276 3069 12340
rect 3003 12275 3069 12276
rect 3554 11456 3874 12480
rect 3554 11392 3562 11456
rect 3626 11392 3642 11456
rect 3706 11392 3722 11456
rect 3786 11392 3802 11456
rect 3866 11392 3874 11456
rect 3554 10368 3874 11392
rect 3554 10304 3562 10368
rect 3626 10304 3642 10368
rect 3706 10304 3722 10368
rect 3786 10304 3802 10368
rect 3866 10304 3874 10368
rect 3554 10046 3874 10304
rect 3554 9810 3596 10046
rect 3832 9810 3874 10046
rect 3554 9280 3874 9810
rect 3554 9216 3562 9280
rect 3626 9216 3642 9280
rect 3706 9216 3722 9280
rect 3786 9216 3802 9280
rect 3866 9216 3874 9280
rect 3554 8192 3874 9216
rect 3554 8128 3562 8192
rect 3626 8128 3642 8192
rect 3706 8128 3722 8192
rect 3786 8128 3802 8192
rect 3866 8128 3874 8192
rect 3554 7104 3874 8128
rect 3554 7040 3562 7104
rect 3626 7040 3642 7104
rect 3706 7040 3722 7104
rect 3786 7040 3802 7104
rect 3866 7040 3874 7104
rect 3554 6016 3874 7040
rect 3554 5952 3562 6016
rect 3626 5952 3642 6016
rect 3706 5952 3722 6016
rect 3786 5952 3802 6016
rect 3866 5952 3874 6016
rect 3554 4928 3874 5952
rect 3554 4864 3562 4928
rect 3626 4878 3642 4928
rect 3706 4878 3722 4928
rect 3786 4878 3802 4928
rect 3866 4864 3874 4928
rect 3554 4642 3596 4864
rect 3832 4642 3874 4864
rect 3554 3840 3874 4642
rect 3554 3776 3562 3840
rect 3626 3776 3642 3840
rect 3706 3776 3722 3840
rect 3786 3776 3802 3840
rect 3866 3776 3874 3840
rect 3554 2752 3874 3776
rect 3554 2688 3562 2752
rect 3626 2688 3642 2752
rect 3706 2688 3722 2752
rect 3786 2688 3802 2752
rect 3866 2688 3874 2752
rect 3554 2128 3874 2688
rect 4214 22880 4534 22896
rect 4214 22816 4222 22880
rect 4286 22816 4302 22880
rect 4366 22816 4382 22880
rect 4446 22816 4462 22880
rect 4526 22816 4534 22880
rect 4214 21792 4534 22816
rect 4214 21728 4222 21792
rect 4286 21728 4302 21792
rect 4366 21728 4382 21792
rect 4446 21728 4462 21792
rect 4526 21728 4534 21792
rect 4214 21042 4534 21728
rect 4214 20806 4256 21042
rect 4492 20806 4534 21042
rect 4214 20704 4534 20806
rect 4214 20640 4222 20704
rect 4286 20640 4302 20704
rect 4366 20640 4382 20704
rect 4446 20640 4462 20704
rect 4526 20640 4534 20704
rect 4214 19616 4534 20640
rect 4214 19552 4222 19616
rect 4286 19552 4302 19616
rect 4366 19552 4382 19616
rect 4446 19552 4462 19616
rect 4526 19552 4534 19616
rect 4214 18528 4534 19552
rect 8775 22336 9095 22896
rect 8775 22272 8783 22336
rect 8847 22272 8863 22336
rect 8927 22272 8943 22336
rect 9007 22272 9023 22336
rect 9087 22272 9095 22336
rect 8775 21248 9095 22272
rect 8775 21184 8783 21248
rect 8847 21184 8863 21248
rect 8927 21184 8943 21248
rect 9007 21184 9023 21248
rect 9087 21184 9095 21248
rect 8775 20382 9095 21184
rect 8775 20160 8817 20382
rect 9053 20160 9095 20382
rect 8775 20096 8783 20160
rect 8847 20096 8863 20146
rect 8927 20096 8943 20146
rect 9007 20096 9023 20146
rect 9087 20096 9095 20160
rect 8523 19412 8589 19413
rect 8523 19348 8524 19412
rect 8588 19348 8589 19412
rect 8523 19347 8589 19348
rect 4214 18464 4222 18528
rect 4286 18464 4302 18528
rect 4366 18464 4382 18528
rect 4446 18464 4462 18528
rect 4526 18464 4534 18528
rect 4214 17440 4534 18464
rect 4214 17376 4222 17440
rect 4286 17376 4302 17440
rect 4366 17376 4382 17440
rect 4446 17376 4462 17440
rect 4526 17376 4534 17440
rect 4214 16352 4534 17376
rect 8526 17237 8586 19347
rect 8775 19072 9095 20096
rect 8775 19008 8783 19072
rect 8847 19008 8863 19072
rect 8927 19008 8943 19072
rect 9007 19008 9023 19072
rect 9087 19008 9095 19072
rect 8775 17984 9095 19008
rect 8775 17920 8783 17984
rect 8847 17920 8863 17984
rect 8927 17920 8943 17984
rect 9007 17920 9023 17984
rect 9087 17920 9095 17984
rect 8523 17236 8589 17237
rect 8523 17172 8524 17236
rect 8588 17172 8589 17236
rect 8523 17171 8589 17172
rect 4214 16288 4222 16352
rect 4286 16288 4302 16352
rect 4366 16288 4382 16352
rect 4446 16288 4462 16352
rect 4526 16288 4534 16352
rect 4214 15874 4534 16288
rect 4214 15638 4256 15874
rect 4492 15638 4534 15874
rect 4214 15264 4534 15638
rect 4214 15200 4222 15264
rect 4286 15200 4302 15264
rect 4366 15200 4382 15264
rect 4446 15200 4462 15264
rect 4526 15200 4534 15264
rect 4214 14176 4534 15200
rect 4214 14112 4222 14176
rect 4286 14112 4302 14176
rect 4366 14112 4382 14176
rect 4446 14112 4462 14176
rect 4526 14112 4534 14176
rect 4214 13088 4534 14112
rect 4214 13024 4222 13088
rect 4286 13024 4302 13088
rect 4366 13024 4382 13088
rect 4446 13024 4462 13088
rect 4526 13024 4534 13088
rect 4214 12000 4534 13024
rect 4214 11936 4222 12000
rect 4286 11936 4302 12000
rect 4366 11936 4382 12000
rect 4446 11936 4462 12000
rect 4526 11936 4534 12000
rect 4214 10912 4534 11936
rect 4214 10848 4222 10912
rect 4286 10848 4302 10912
rect 4366 10848 4382 10912
rect 4446 10848 4462 10912
rect 4526 10848 4534 10912
rect 4214 10706 4534 10848
rect 4214 10470 4256 10706
rect 4492 10470 4534 10706
rect 4214 9824 4534 10470
rect 4214 9760 4222 9824
rect 4286 9760 4302 9824
rect 4366 9760 4382 9824
rect 4446 9760 4462 9824
rect 4526 9760 4534 9824
rect 4214 8736 4534 9760
rect 4214 8672 4222 8736
rect 4286 8672 4302 8736
rect 4366 8672 4382 8736
rect 4446 8672 4462 8736
rect 4526 8672 4534 8736
rect 4214 7648 4534 8672
rect 4214 7584 4222 7648
rect 4286 7584 4302 7648
rect 4366 7584 4382 7648
rect 4446 7584 4462 7648
rect 4526 7584 4534 7648
rect 4214 6560 4534 7584
rect 4214 6496 4222 6560
rect 4286 6496 4302 6560
rect 4366 6496 4382 6560
rect 4446 6496 4462 6560
rect 4526 6496 4534 6560
rect 4214 5538 4534 6496
rect 4214 5472 4256 5538
rect 4492 5472 4534 5538
rect 4214 5408 4222 5472
rect 4526 5408 4534 5472
rect 4214 5302 4256 5408
rect 4492 5302 4534 5408
rect 4214 4384 4534 5302
rect 4214 4320 4222 4384
rect 4286 4320 4302 4384
rect 4366 4320 4382 4384
rect 4446 4320 4462 4384
rect 4526 4320 4534 4384
rect 4214 3296 4534 4320
rect 4214 3232 4222 3296
rect 4286 3232 4302 3296
rect 4366 3232 4382 3296
rect 4446 3232 4462 3296
rect 4526 3232 4534 3296
rect 4214 2208 4534 3232
rect 4214 2144 4222 2208
rect 4286 2144 4302 2208
rect 4366 2144 4382 2208
rect 4446 2144 4462 2208
rect 4526 2144 4534 2208
rect 4214 2128 4534 2144
rect 8775 16896 9095 17920
rect 8775 16832 8783 16896
rect 8847 16832 8863 16896
rect 8927 16832 8943 16896
rect 9007 16832 9023 16896
rect 9087 16832 9095 16896
rect 8775 15808 9095 16832
rect 8775 15744 8783 15808
rect 8847 15744 8863 15808
rect 8927 15744 8943 15808
rect 9007 15744 9023 15808
rect 9087 15744 9095 15808
rect 8775 15214 9095 15744
rect 8775 14978 8817 15214
rect 9053 14978 9095 15214
rect 8775 14720 9095 14978
rect 8775 14656 8783 14720
rect 8847 14656 8863 14720
rect 8927 14656 8943 14720
rect 9007 14656 9023 14720
rect 9087 14656 9095 14720
rect 8775 13632 9095 14656
rect 8775 13568 8783 13632
rect 8847 13568 8863 13632
rect 8927 13568 8943 13632
rect 9007 13568 9023 13632
rect 9087 13568 9095 13632
rect 8775 12544 9095 13568
rect 8775 12480 8783 12544
rect 8847 12480 8863 12544
rect 8927 12480 8943 12544
rect 9007 12480 9023 12544
rect 9087 12480 9095 12544
rect 8775 11456 9095 12480
rect 8775 11392 8783 11456
rect 8847 11392 8863 11456
rect 8927 11392 8943 11456
rect 9007 11392 9023 11456
rect 9087 11392 9095 11456
rect 8775 10368 9095 11392
rect 8775 10304 8783 10368
rect 8847 10304 8863 10368
rect 8927 10304 8943 10368
rect 9007 10304 9023 10368
rect 9087 10304 9095 10368
rect 8775 10046 9095 10304
rect 8775 9810 8817 10046
rect 9053 9810 9095 10046
rect 8775 9280 9095 9810
rect 8775 9216 8783 9280
rect 8847 9216 8863 9280
rect 8927 9216 8943 9280
rect 9007 9216 9023 9280
rect 9087 9216 9095 9280
rect 8775 8192 9095 9216
rect 8775 8128 8783 8192
rect 8847 8128 8863 8192
rect 8927 8128 8943 8192
rect 9007 8128 9023 8192
rect 9087 8128 9095 8192
rect 8775 7104 9095 8128
rect 8775 7040 8783 7104
rect 8847 7040 8863 7104
rect 8927 7040 8943 7104
rect 9007 7040 9023 7104
rect 9087 7040 9095 7104
rect 8775 6016 9095 7040
rect 8775 5952 8783 6016
rect 8847 5952 8863 6016
rect 8927 5952 8943 6016
rect 9007 5952 9023 6016
rect 9087 5952 9095 6016
rect 8775 4928 9095 5952
rect 8775 4864 8783 4928
rect 8847 4878 8863 4928
rect 8927 4878 8943 4928
rect 9007 4878 9023 4928
rect 9087 4864 9095 4928
rect 8775 4642 8817 4864
rect 9053 4642 9095 4864
rect 8775 3840 9095 4642
rect 8775 3776 8783 3840
rect 8847 3776 8863 3840
rect 8927 3776 8943 3840
rect 9007 3776 9023 3840
rect 9087 3776 9095 3840
rect 8775 2752 9095 3776
rect 8775 2688 8783 2752
rect 8847 2688 8863 2752
rect 8927 2688 8943 2752
rect 9007 2688 9023 2752
rect 9087 2688 9095 2752
rect 8775 2128 9095 2688
rect 9435 22880 9755 22896
rect 9435 22816 9443 22880
rect 9507 22816 9523 22880
rect 9587 22816 9603 22880
rect 9667 22816 9683 22880
rect 9747 22816 9755 22880
rect 9435 21792 9755 22816
rect 9435 21728 9443 21792
rect 9507 21728 9523 21792
rect 9587 21728 9603 21792
rect 9667 21728 9683 21792
rect 9747 21728 9755 21792
rect 9435 21042 9755 21728
rect 9435 20806 9477 21042
rect 9713 20806 9755 21042
rect 9435 20704 9755 20806
rect 9435 20640 9443 20704
rect 9507 20640 9523 20704
rect 9587 20640 9603 20704
rect 9667 20640 9683 20704
rect 9747 20640 9755 20704
rect 9435 19616 9755 20640
rect 9435 19552 9443 19616
rect 9507 19552 9523 19616
rect 9587 19552 9603 19616
rect 9667 19552 9683 19616
rect 9747 19552 9755 19616
rect 9435 18528 9755 19552
rect 9435 18464 9443 18528
rect 9507 18464 9523 18528
rect 9587 18464 9603 18528
rect 9667 18464 9683 18528
rect 9747 18464 9755 18528
rect 9435 17440 9755 18464
rect 9435 17376 9443 17440
rect 9507 17376 9523 17440
rect 9587 17376 9603 17440
rect 9667 17376 9683 17440
rect 9747 17376 9755 17440
rect 9435 16352 9755 17376
rect 9435 16288 9443 16352
rect 9507 16288 9523 16352
rect 9587 16288 9603 16352
rect 9667 16288 9683 16352
rect 9747 16288 9755 16352
rect 9435 15874 9755 16288
rect 9435 15638 9477 15874
rect 9713 15638 9755 15874
rect 9435 15264 9755 15638
rect 9435 15200 9443 15264
rect 9507 15200 9523 15264
rect 9587 15200 9603 15264
rect 9667 15200 9683 15264
rect 9747 15200 9755 15264
rect 9435 14176 9755 15200
rect 9435 14112 9443 14176
rect 9507 14112 9523 14176
rect 9587 14112 9603 14176
rect 9667 14112 9683 14176
rect 9747 14112 9755 14176
rect 9435 13088 9755 14112
rect 9435 13024 9443 13088
rect 9507 13024 9523 13088
rect 9587 13024 9603 13088
rect 9667 13024 9683 13088
rect 9747 13024 9755 13088
rect 9435 12000 9755 13024
rect 9435 11936 9443 12000
rect 9507 11936 9523 12000
rect 9587 11936 9603 12000
rect 9667 11936 9683 12000
rect 9747 11936 9755 12000
rect 9435 10912 9755 11936
rect 9435 10848 9443 10912
rect 9507 10848 9523 10912
rect 9587 10848 9603 10912
rect 9667 10848 9683 10912
rect 9747 10848 9755 10912
rect 9435 10706 9755 10848
rect 9435 10470 9477 10706
rect 9713 10470 9755 10706
rect 9435 9824 9755 10470
rect 9435 9760 9443 9824
rect 9507 9760 9523 9824
rect 9587 9760 9603 9824
rect 9667 9760 9683 9824
rect 9747 9760 9755 9824
rect 9435 8736 9755 9760
rect 9435 8672 9443 8736
rect 9507 8672 9523 8736
rect 9587 8672 9603 8736
rect 9667 8672 9683 8736
rect 9747 8672 9755 8736
rect 9435 7648 9755 8672
rect 9435 7584 9443 7648
rect 9507 7584 9523 7648
rect 9587 7584 9603 7648
rect 9667 7584 9683 7648
rect 9747 7584 9755 7648
rect 9435 6560 9755 7584
rect 9435 6496 9443 6560
rect 9507 6496 9523 6560
rect 9587 6496 9603 6560
rect 9667 6496 9683 6560
rect 9747 6496 9755 6560
rect 9435 5538 9755 6496
rect 9435 5472 9477 5538
rect 9713 5472 9755 5538
rect 9435 5408 9443 5472
rect 9747 5408 9755 5472
rect 9435 5302 9477 5408
rect 9713 5302 9755 5408
rect 9435 4384 9755 5302
rect 9435 4320 9443 4384
rect 9507 4320 9523 4384
rect 9587 4320 9603 4384
rect 9667 4320 9683 4384
rect 9747 4320 9755 4384
rect 9435 3296 9755 4320
rect 9435 3232 9443 3296
rect 9507 3232 9523 3296
rect 9587 3232 9603 3296
rect 9667 3232 9683 3296
rect 9747 3232 9755 3296
rect 9435 2208 9755 3232
rect 9435 2144 9443 2208
rect 9507 2144 9523 2208
rect 9587 2144 9603 2208
rect 9667 2144 9683 2208
rect 9747 2144 9755 2208
rect 9435 2128 9755 2144
rect 13996 22336 14316 22896
rect 13996 22272 14004 22336
rect 14068 22272 14084 22336
rect 14148 22272 14164 22336
rect 14228 22272 14244 22336
rect 14308 22272 14316 22336
rect 13996 21248 14316 22272
rect 13996 21184 14004 21248
rect 14068 21184 14084 21248
rect 14148 21184 14164 21248
rect 14228 21184 14244 21248
rect 14308 21184 14316 21248
rect 13996 20382 14316 21184
rect 13996 20160 14038 20382
rect 14274 20160 14316 20382
rect 13996 20096 14004 20160
rect 14068 20096 14084 20146
rect 14148 20096 14164 20146
rect 14228 20096 14244 20146
rect 14308 20096 14316 20160
rect 13996 19072 14316 20096
rect 13996 19008 14004 19072
rect 14068 19008 14084 19072
rect 14148 19008 14164 19072
rect 14228 19008 14244 19072
rect 14308 19008 14316 19072
rect 13996 17984 14316 19008
rect 13996 17920 14004 17984
rect 14068 17920 14084 17984
rect 14148 17920 14164 17984
rect 14228 17920 14244 17984
rect 14308 17920 14316 17984
rect 13996 16896 14316 17920
rect 14656 22880 14976 22896
rect 14656 22816 14664 22880
rect 14728 22816 14744 22880
rect 14808 22816 14824 22880
rect 14888 22816 14904 22880
rect 14968 22816 14976 22880
rect 14656 21792 14976 22816
rect 14656 21728 14664 21792
rect 14728 21728 14744 21792
rect 14808 21728 14824 21792
rect 14888 21728 14904 21792
rect 14968 21728 14976 21792
rect 14656 21042 14976 21728
rect 14656 20806 14698 21042
rect 14934 20806 14976 21042
rect 14656 20704 14976 20806
rect 14656 20640 14664 20704
rect 14728 20640 14744 20704
rect 14808 20640 14824 20704
rect 14888 20640 14904 20704
rect 14968 20640 14976 20704
rect 14656 19616 14976 20640
rect 14656 19552 14664 19616
rect 14728 19552 14744 19616
rect 14808 19552 14824 19616
rect 14888 19552 14904 19616
rect 14968 19552 14976 19616
rect 14656 18528 14976 19552
rect 19217 22336 19537 22896
rect 19217 22272 19225 22336
rect 19289 22272 19305 22336
rect 19369 22272 19385 22336
rect 19449 22272 19465 22336
rect 19529 22272 19537 22336
rect 19217 21248 19537 22272
rect 19217 21184 19225 21248
rect 19289 21184 19305 21248
rect 19369 21184 19385 21248
rect 19449 21184 19465 21248
rect 19529 21184 19537 21248
rect 19217 20382 19537 21184
rect 19217 20160 19259 20382
rect 19495 20160 19537 20382
rect 19217 20096 19225 20160
rect 19289 20096 19305 20146
rect 19369 20096 19385 20146
rect 19449 20096 19465 20146
rect 19529 20096 19537 20160
rect 19217 19072 19537 20096
rect 19217 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19465 19072
rect 19529 19008 19537 19072
rect 17723 18596 17789 18597
rect 17723 18532 17724 18596
rect 17788 18532 17789 18596
rect 17723 18531 17789 18532
rect 14656 18464 14664 18528
rect 14728 18464 14744 18528
rect 14808 18464 14824 18528
rect 14888 18464 14904 18528
rect 14968 18464 14976 18528
rect 14656 17440 14976 18464
rect 14656 17376 14664 17440
rect 14728 17376 14744 17440
rect 14808 17376 14824 17440
rect 14888 17376 14904 17440
rect 14968 17376 14976 17440
rect 14411 17236 14477 17237
rect 14411 17172 14412 17236
rect 14476 17172 14477 17236
rect 14411 17171 14477 17172
rect 13996 16832 14004 16896
rect 14068 16832 14084 16896
rect 14148 16832 14164 16896
rect 14228 16832 14244 16896
rect 14308 16832 14316 16896
rect 13996 15808 14316 16832
rect 13996 15744 14004 15808
rect 14068 15744 14084 15808
rect 14148 15744 14164 15808
rect 14228 15744 14244 15808
rect 14308 15744 14316 15808
rect 13996 15214 14316 15744
rect 13996 14978 14038 15214
rect 14274 14978 14316 15214
rect 13996 14720 14316 14978
rect 13996 14656 14004 14720
rect 14068 14656 14084 14720
rect 14148 14656 14164 14720
rect 14228 14656 14244 14720
rect 14308 14656 14316 14720
rect 13996 13632 14316 14656
rect 13996 13568 14004 13632
rect 14068 13568 14084 13632
rect 14148 13568 14164 13632
rect 14228 13568 14244 13632
rect 14308 13568 14316 13632
rect 13996 12544 14316 13568
rect 13996 12480 14004 12544
rect 14068 12480 14084 12544
rect 14148 12480 14164 12544
rect 14228 12480 14244 12544
rect 14308 12480 14316 12544
rect 13996 11456 14316 12480
rect 14414 12341 14474 17171
rect 14656 16352 14976 17376
rect 14656 16288 14664 16352
rect 14728 16288 14744 16352
rect 14808 16288 14824 16352
rect 14888 16288 14904 16352
rect 14968 16288 14976 16352
rect 14656 15874 14976 16288
rect 17726 16149 17786 18531
rect 19217 17984 19537 19008
rect 19217 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19465 17984
rect 19529 17920 19537 17984
rect 19217 16896 19537 17920
rect 19217 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19465 16896
rect 19529 16832 19537 16896
rect 17723 16148 17789 16149
rect 17723 16084 17724 16148
rect 17788 16084 17789 16148
rect 17723 16083 17789 16084
rect 14656 15638 14698 15874
rect 14934 15638 14976 15874
rect 14656 15264 14976 15638
rect 14656 15200 14664 15264
rect 14728 15200 14744 15264
rect 14808 15200 14824 15264
rect 14888 15200 14904 15264
rect 14968 15200 14976 15264
rect 14656 14176 14976 15200
rect 14656 14112 14664 14176
rect 14728 14112 14744 14176
rect 14808 14112 14824 14176
rect 14888 14112 14904 14176
rect 14968 14112 14976 14176
rect 14656 13088 14976 14112
rect 14656 13024 14664 13088
rect 14728 13024 14744 13088
rect 14808 13024 14824 13088
rect 14888 13024 14904 13088
rect 14968 13024 14976 13088
rect 14411 12340 14477 12341
rect 14411 12276 14412 12340
rect 14476 12276 14477 12340
rect 14411 12275 14477 12276
rect 13996 11392 14004 11456
rect 14068 11392 14084 11456
rect 14148 11392 14164 11456
rect 14228 11392 14244 11456
rect 14308 11392 14316 11456
rect 13996 10368 14316 11392
rect 13996 10304 14004 10368
rect 14068 10304 14084 10368
rect 14148 10304 14164 10368
rect 14228 10304 14244 10368
rect 14308 10304 14316 10368
rect 13996 10046 14316 10304
rect 13996 9810 14038 10046
rect 14274 9810 14316 10046
rect 13996 9280 14316 9810
rect 13996 9216 14004 9280
rect 14068 9216 14084 9280
rect 14148 9216 14164 9280
rect 14228 9216 14244 9280
rect 14308 9216 14316 9280
rect 13996 8192 14316 9216
rect 14414 8533 14474 12275
rect 14656 12000 14976 13024
rect 14656 11936 14664 12000
rect 14728 11936 14744 12000
rect 14808 11936 14824 12000
rect 14888 11936 14904 12000
rect 14968 11936 14976 12000
rect 14656 10912 14976 11936
rect 14656 10848 14664 10912
rect 14728 10848 14744 10912
rect 14808 10848 14824 10912
rect 14888 10848 14904 10912
rect 14968 10848 14976 10912
rect 14656 10706 14976 10848
rect 14656 10470 14698 10706
rect 14934 10470 14976 10706
rect 14656 9824 14976 10470
rect 14656 9760 14664 9824
rect 14728 9760 14744 9824
rect 14808 9760 14824 9824
rect 14888 9760 14904 9824
rect 14968 9760 14976 9824
rect 14656 8736 14976 9760
rect 14656 8672 14664 8736
rect 14728 8672 14744 8736
rect 14808 8672 14824 8736
rect 14888 8672 14904 8736
rect 14968 8672 14976 8736
rect 14411 8532 14477 8533
rect 14411 8468 14412 8532
rect 14476 8468 14477 8532
rect 14411 8467 14477 8468
rect 13996 8128 14004 8192
rect 14068 8128 14084 8192
rect 14148 8128 14164 8192
rect 14228 8128 14244 8192
rect 14308 8128 14316 8192
rect 13996 7104 14316 8128
rect 13996 7040 14004 7104
rect 14068 7040 14084 7104
rect 14148 7040 14164 7104
rect 14228 7040 14244 7104
rect 14308 7040 14316 7104
rect 13996 6016 14316 7040
rect 14414 6493 14474 8467
rect 14656 7648 14976 8672
rect 14656 7584 14664 7648
rect 14728 7584 14744 7648
rect 14808 7584 14824 7648
rect 14888 7584 14904 7648
rect 14968 7584 14976 7648
rect 14656 6560 14976 7584
rect 14656 6496 14664 6560
rect 14728 6496 14744 6560
rect 14808 6496 14824 6560
rect 14888 6496 14904 6560
rect 14968 6496 14976 6560
rect 14411 6492 14477 6493
rect 14411 6428 14412 6492
rect 14476 6428 14477 6492
rect 14411 6427 14477 6428
rect 13996 5952 14004 6016
rect 14068 5952 14084 6016
rect 14148 5952 14164 6016
rect 14228 5952 14244 6016
rect 14308 5952 14316 6016
rect 13996 4928 14316 5952
rect 13996 4864 14004 4928
rect 14068 4878 14084 4928
rect 14148 4878 14164 4928
rect 14228 4878 14244 4928
rect 14308 4864 14316 4928
rect 13996 4642 14038 4864
rect 14274 4642 14316 4864
rect 13996 3840 14316 4642
rect 13996 3776 14004 3840
rect 14068 3776 14084 3840
rect 14148 3776 14164 3840
rect 14228 3776 14244 3840
rect 14308 3776 14316 3840
rect 13996 2752 14316 3776
rect 13996 2688 14004 2752
rect 14068 2688 14084 2752
rect 14148 2688 14164 2752
rect 14228 2688 14244 2752
rect 14308 2688 14316 2752
rect 13996 2128 14316 2688
rect 14656 5538 14976 6496
rect 14656 5472 14698 5538
rect 14934 5472 14976 5538
rect 14656 5408 14664 5472
rect 14968 5408 14976 5472
rect 14656 5302 14698 5408
rect 14934 5302 14976 5408
rect 14656 4384 14976 5302
rect 14656 4320 14664 4384
rect 14728 4320 14744 4384
rect 14808 4320 14824 4384
rect 14888 4320 14904 4384
rect 14968 4320 14976 4384
rect 14656 3296 14976 4320
rect 14656 3232 14664 3296
rect 14728 3232 14744 3296
rect 14808 3232 14824 3296
rect 14888 3232 14904 3296
rect 14968 3232 14976 3296
rect 14656 2208 14976 3232
rect 14656 2144 14664 2208
rect 14728 2144 14744 2208
rect 14808 2144 14824 2208
rect 14888 2144 14904 2208
rect 14968 2144 14976 2208
rect 14656 2128 14976 2144
rect 19217 15808 19537 16832
rect 19217 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19465 15808
rect 19529 15744 19537 15808
rect 19217 15214 19537 15744
rect 19217 14978 19259 15214
rect 19495 14978 19537 15214
rect 19217 14720 19537 14978
rect 19217 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19465 14720
rect 19529 14656 19537 14720
rect 19217 13632 19537 14656
rect 19217 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19465 13632
rect 19529 13568 19537 13632
rect 19217 12544 19537 13568
rect 19217 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19465 12544
rect 19529 12480 19537 12544
rect 19217 11456 19537 12480
rect 19217 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19465 11456
rect 19529 11392 19537 11456
rect 19217 10368 19537 11392
rect 19217 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19465 10368
rect 19529 10304 19537 10368
rect 19217 10046 19537 10304
rect 19217 9810 19259 10046
rect 19495 9810 19537 10046
rect 19217 9280 19537 9810
rect 19217 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19465 9280
rect 19529 9216 19537 9280
rect 19217 8192 19537 9216
rect 19217 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19465 8192
rect 19529 8128 19537 8192
rect 19217 7104 19537 8128
rect 19217 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19465 7104
rect 19529 7040 19537 7104
rect 19217 6016 19537 7040
rect 19217 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19465 6016
rect 19529 5952 19537 6016
rect 19217 4928 19537 5952
rect 19217 4864 19225 4928
rect 19289 4878 19305 4928
rect 19369 4878 19385 4928
rect 19449 4878 19465 4928
rect 19529 4864 19537 4928
rect 19217 4642 19259 4864
rect 19495 4642 19537 4864
rect 19217 3840 19537 4642
rect 19217 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19465 3840
rect 19529 3776 19537 3840
rect 19217 2752 19537 3776
rect 19217 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19465 2752
rect 19529 2688 19537 2752
rect 19217 2128 19537 2688
rect 19877 22880 20197 22896
rect 19877 22816 19885 22880
rect 19949 22816 19965 22880
rect 20029 22816 20045 22880
rect 20109 22816 20125 22880
rect 20189 22816 20197 22880
rect 19877 21792 20197 22816
rect 19877 21728 19885 21792
rect 19949 21728 19965 21792
rect 20029 21728 20045 21792
rect 20109 21728 20125 21792
rect 20189 21728 20197 21792
rect 19877 21042 20197 21728
rect 19877 20806 19919 21042
rect 20155 20806 20197 21042
rect 19877 20704 20197 20806
rect 19877 20640 19885 20704
rect 19949 20640 19965 20704
rect 20029 20640 20045 20704
rect 20109 20640 20125 20704
rect 20189 20640 20197 20704
rect 19877 19616 20197 20640
rect 19877 19552 19885 19616
rect 19949 19552 19965 19616
rect 20029 19552 20045 19616
rect 20109 19552 20125 19616
rect 20189 19552 20197 19616
rect 19877 18528 20197 19552
rect 19877 18464 19885 18528
rect 19949 18464 19965 18528
rect 20029 18464 20045 18528
rect 20109 18464 20125 18528
rect 20189 18464 20197 18528
rect 19877 17440 20197 18464
rect 19877 17376 19885 17440
rect 19949 17376 19965 17440
rect 20029 17376 20045 17440
rect 20109 17376 20125 17440
rect 20189 17376 20197 17440
rect 19877 16352 20197 17376
rect 19877 16288 19885 16352
rect 19949 16288 19965 16352
rect 20029 16288 20045 16352
rect 20109 16288 20125 16352
rect 20189 16288 20197 16352
rect 19877 15874 20197 16288
rect 19877 15638 19919 15874
rect 20155 15638 20197 15874
rect 19877 15264 20197 15638
rect 19877 15200 19885 15264
rect 19949 15200 19965 15264
rect 20029 15200 20045 15264
rect 20109 15200 20125 15264
rect 20189 15200 20197 15264
rect 19877 14176 20197 15200
rect 19877 14112 19885 14176
rect 19949 14112 19965 14176
rect 20029 14112 20045 14176
rect 20109 14112 20125 14176
rect 20189 14112 20197 14176
rect 19877 13088 20197 14112
rect 19877 13024 19885 13088
rect 19949 13024 19965 13088
rect 20029 13024 20045 13088
rect 20109 13024 20125 13088
rect 20189 13024 20197 13088
rect 19877 12000 20197 13024
rect 19877 11936 19885 12000
rect 19949 11936 19965 12000
rect 20029 11936 20045 12000
rect 20109 11936 20125 12000
rect 20189 11936 20197 12000
rect 19877 10912 20197 11936
rect 19877 10848 19885 10912
rect 19949 10848 19965 10912
rect 20029 10848 20045 10912
rect 20109 10848 20125 10912
rect 20189 10848 20197 10912
rect 19877 10706 20197 10848
rect 19877 10470 19919 10706
rect 20155 10470 20197 10706
rect 19877 9824 20197 10470
rect 19877 9760 19885 9824
rect 19949 9760 19965 9824
rect 20029 9760 20045 9824
rect 20109 9760 20125 9824
rect 20189 9760 20197 9824
rect 19877 8736 20197 9760
rect 19877 8672 19885 8736
rect 19949 8672 19965 8736
rect 20029 8672 20045 8736
rect 20109 8672 20125 8736
rect 20189 8672 20197 8736
rect 19877 7648 20197 8672
rect 19877 7584 19885 7648
rect 19949 7584 19965 7648
rect 20029 7584 20045 7648
rect 20109 7584 20125 7648
rect 20189 7584 20197 7648
rect 19877 6560 20197 7584
rect 19877 6496 19885 6560
rect 19949 6496 19965 6560
rect 20029 6496 20045 6560
rect 20109 6496 20125 6560
rect 20189 6496 20197 6560
rect 19877 5538 20197 6496
rect 19877 5472 19919 5538
rect 20155 5472 20197 5538
rect 19877 5408 19885 5472
rect 20189 5408 20197 5472
rect 19877 5302 19919 5408
rect 20155 5302 20197 5408
rect 19877 4384 20197 5302
rect 19877 4320 19885 4384
rect 19949 4320 19965 4384
rect 20029 4320 20045 4384
rect 20109 4320 20125 4384
rect 20189 4320 20197 4384
rect 19877 3296 20197 4320
rect 19877 3232 19885 3296
rect 19949 3232 19965 3296
rect 20029 3232 20045 3296
rect 20109 3232 20125 3296
rect 20189 3232 20197 3296
rect 19877 2208 20197 3232
rect 19877 2144 19885 2208
rect 19949 2144 19965 2208
rect 20029 2144 20045 2208
rect 20109 2144 20125 2208
rect 20189 2144 20197 2208
rect 19877 2128 20197 2144
<< via4 >>
rect 3596 20160 3832 20382
rect 3596 20146 3626 20160
rect 3626 20146 3642 20160
rect 3642 20146 3706 20160
rect 3706 20146 3722 20160
rect 3722 20146 3786 20160
rect 3786 20146 3802 20160
rect 3802 20146 3832 20160
rect 3596 14978 3832 15214
rect 3596 9810 3832 10046
rect 3596 4864 3626 4878
rect 3626 4864 3642 4878
rect 3642 4864 3706 4878
rect 3706 4864 3722 4878
rect 3722 4864 3786 4878
rect 3786 4864 3802 4878
rect 3802 4864 3832 4878
rect 3596 4642 3832 4864
rect 4256 20806 4492 21042
rect 8817 20160 9053 20382
rect 8817 20146 8847 20160
rect 8847 20146 8863 20160
rect 8863 20146 8927 20160
rect 8927 20146 8943 20160
rect 8943 20146 9007 20160
rect 9007 20146 9023 20160
rect 9023 20146 9053 20160
rect 4256 15638 4492 15874
rect 4256 10470 4492 10706
rect 4256 5472 4492 5538
rect 4256 5408 4286 5472
rect 4286 5408 4302 5472
rect 4302 5408 4366 5472
rect 4366 5408 4382 5472
rect 4382 5408 4446 5472
rect 4446 5408 4462 5472
rect 4462 5408 4492 5472
rect 4256 5302 4492 5408
rect 8817 14978 9053 15214
rect 8817 9810 9053 10046
rect 8817 4864 8847 4878
rect 8847 4864 8863 4878
rect 8863 4864 8927 4878
rect 8927 4864 8943 4878
rect 8943 4864 9007 4878
rect 9007 4864 9023 4878
rect 9023 4864 9053 4878
rect 8817 4642 9053 4864
rect 9477 20806 9713 21042
rect 9477 15638 9713 15874
rect 9477 10470 9713 10706
rect 9477 5472 9713 5538
rect 9477 5408 9507 5472
rect 9507 5408 9523 5472
rect 9523 5408 9587 5472
rect 9587 5408 9603 5472
rect 9603 5408 9667 5472
rect 9667 5408 9683 5472
rect 9683 5408 9713 5472
rect 9477 5302 9713 5408
rect 14038 20160 14274 20382
rect 14038 20146 14068 20160
rect 14068 20146 14084 20160
rect 14084 20146 14148 20160
rect 14148 20146 14164 20160
rect 14164 20146 14228 20160
rect 14228 20146 14244 20160
rect 14244 20146 14274 20160
rect 14698 20806 14934 21042
rect 19259 20160 19495 20382
rect 19259 20146 19289 20160
rect 19289 20146 19305 20160
rect 19305 20146 19369 20160
rect 19369 20146 19385 20160
rect 19385 20146 19449 20160
rect 19449 20146 19465 20160
rect 19465 20146 19495 20160
rect 14038 14978 14274 15214
rect 14698 15638 14934 15874
rect 14038 9810 14274 10046
rect 14698 10470 14934 10706
rect 14038 4864 14068 4878
rect 14068 4864 14084 4878
rect 14084 4864 14148 4878
rect 14148 4864 14164 4878
rect 14164 4864 14228 4878
rect 14228 4864 14244 4878
rect 14244 4864 14274 4878
rect 14038 4642 14274 4864
rect 14698 5472 14934 5538
rect 14698 5408 14728 5472
rect 14728 5408 14744 5472
rect 14744 5408 14808 5472
rect 14808 5408 14824 5472
rect 14824 5408 14888 5472
rect 14888 5408 14904 5472
rect 14904 5408 14934 5472
rect 14698 5302 14934 5408
rect 19259 14978 19495 15214
rect 19259 9810 19495 10046
rect 19259 4864 19289 4878
rect 19289 4864 19305 4878
rect 19305 4864 19369 4878
rect 19369 4864 19385 4878
rect 19385 4864 19449 4878
rect 19449 4864 19465 4878
rect 19465 4864 19495 4878
rect 19259 4642 19495 4864
rect 19919 20806 20155 21042
rect 19919 15638 20155 15874
rect 19919 10470 20155 10706
rect 19919 5472 20155 5538
rect 19919 5408 19949 5472
rect 19949 5408 19965 5472
rect 19965 5408 20029 5472
rect 20029 5408 20045 5472
rect 20045 5408 20109 5472
rect 20109 5408 20125 5472
rect 20125 5408 20155 5472
rect 19919 5302 20155 5408
<< metal5 >>
rect 1056 21042 22036 21084
rect 1056 20806 4256 21042
rect 4492 20806 9477 21042
rect 9713 20806 14698 21042
rect 14934 20806 19919 21042
rect 20155 20806 22036 21042
rect 1056 20764 22036 20806
rect 1056 20382 22036 20424
rect 1056 20146 3596 20382
rect 3832 20146 8817 20382
rect 9053 20146 14038 20382
rect 14274 20146 19259 20382
rect 19495 20146 22036 20382
rect 1056 20104 22036 20146
rect 1056 15874 22036 15916
rect 1056 15638 4256 15874
rect 4492 15638 9477 15874
rect 9713 15638 14698 15874
rect 14934 15638 19919 15874
rect 20155 15638 22036 15874
rect 1056 15596 22036 15638
rect 1056 15214 22036 15256
rect 1056 14978 3596 15214
rect 3832 14978 8817 15214
rect 9053 14978 14038 15214
rect 14274 14978 19259 15214
rect 19495 14978 22036 15214
rect 1056 14936 22036 14978
rect 1056 10706 22036 10748
rect 1056 10470 4256 10706
rect 4492 10470 9477 10706
rect 9713 10470 14698 10706
rect 14934 10470 19919 10706
rect 20155 10470 22036 10706
rect 1056 10428 22036 10470
rect 1056 10046 22036 10088
rect 1056 9810 3596 10046
rect 3832 9810 8817 10046
rect 9053 9810 14038 10046
rect 14274 9810 19259 10046
rect 19495 9810 22036 10046
rect 1056 9768 22036 9810
rect 1056 5538 22036 5580
rect 1056 5302 4256 5538
rect 4492 5302 9477 5538
rect 9713 5302 14698 5538
rect 14934 5302 19919 5538
rect 20155 5302 22036 5538
rect 1056 5260 22036 5302
rect 1056 4878 22036 4920
rect 1056 4642 3596 4878
rect 3832 4642 8817 4878
rect 9053 4642 14038 4878
rect 14274 4642 19259 4878
rect 19495 4642 22036 4878
rect 1056 4600 22036 4642
use sky130_fd_sc_hd__and4b_2  _0478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10120 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9476 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0480_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0481_
timestamp 1704896540
transform 1 0 10948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_1  _0482_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10304 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0483_
timestamp 1704896540
transform -1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6900 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _0485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4968 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7084 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0489_
timestamp 1704896540
transform -1 0 6532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10304 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8832 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _0492_
timestamp 1704896540
transform -1 0 10764 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10396 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13524 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _0495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_2  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10120 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__or3b_2  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9200 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _0498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9016 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _0499_
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0500_
timestamp 1704896540
transform 1 0 7360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0501_
timestamp 1704896540
transform 1 0 7912 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0502_
timestamp 1704896540
transform -1 0 9200 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _0503_
timestamp 1704896540
transform -1 0 4600 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _0504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9476 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _0505_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9844 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1704896540
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0508_
timestamp 1704896540
transform 1 0 13432 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_2  _0509_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11776 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_2  _0510_
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1704896540
transform -1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0513_
timestamp 1704896540
transform -1 0 2944 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _0514_
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0515_
timestamp 1704896540
transform -1 0 4232 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0516_
timestamp 1704896540
transform -1 0 11408 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _0517_
timestamp 1704896540
transform 1 0 4876 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0518_
timestamp 1704896540
transform 1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0519_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10396 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0520_
timestamp 1704896540
transform -1 0 9936 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0521_
timestamp 1704896540
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0522_
timestamp 1704896540
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0523_
timestamp 1704896540
transform -1 0 7544 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0524_
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0525_
timestamp 1704896540
transform -1 0 3680 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0526_
timestamp 1704896540
transform 1 0 17756 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0528_
timestamp 1704896540
transform -1 0 16560 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0529_
timestamp 1704896540
transform -1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0530_
timestamp 1704896540
transform 1 0 15916 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0531_
timestamp 1704896540
transform 1 0 18492 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0532_
timestamp 1704896540
transform 1 0 17020 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0533_
timestamp 1704896540
transform -1 0 14076 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0534_
timestamp 1704896540
transform 1 0 19504 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0535_
timestamp 1704896540
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0536_
timestamp 1704896540
transform 1 0 10488 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0537_
timestamp 1704896540
transform -1 0 18860 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0538_
timestamp 1704896540
transform -1 0 19136 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0539_
timestamp 1704896540
transform 1 0 6164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0540_
timestamp 1704896540
transform 1 0 15732 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0541_
timestamp 1704896540
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0542_
timestamp 1704896540
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0543_
timestamp 1704896540
transform 1 0 18216 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0544_
timestamp 1704896540
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0545_
timestamp 1704896540
transform 1 0 20056 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0546_
timestamp 1704896540
transform 1 0 19504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0547_
timestamp 1704896540
transform 1 0 20148 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0548_
timestamp 1704896540
transform -1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1704896540
transform -1 0 7820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0550_
timestamp 1704896540
transform -1 0 10856 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0551_
timestamp 1704896540
transform -1 0 8832 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _0552_
timestamp 1704896540
transform 1 0 7912 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0553_
timestamp 1704896540
transform -1 0 7636 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_2  _0554_
timestamp 1704896540
transform 1 0 7544 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_2  _0555_
timestamp 1704896540
transform 1 0 6164 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0556_
timestamp 1704896540
transform -1 0 10120 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o41ai_4  _0557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 -1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__a22o_2  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0559_
timestamp 1704896540
transform 1 0 3956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0560_
timestamp 1704896540
transform 1 0 4692 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0561_
timestamp 1704896540
transform 1 0 5060 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0562_
timestamp 1704896540
transform -1 0 7268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0564_
timestamp 1704896540
transform -1 0 7820 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0565_
timestamp 1704896540
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0566_
timestamp 1704896540
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0567_
timestamp 1704896540
transform 1 0 9568 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0568_
timestamp 1704896540
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0569_
timestamp 1704896540
transform -1 0 10120 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0570_
timestamp 1704896540
transform 1 0 8096 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0571_
timestamp 1704896540
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0572_
timestamp 1704896540
transform 1 0 7176 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _0573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _0574_
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0575_
timestamp 1704896540
transform 1 0 8096 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _0577_
timestamp 1704896540
transform 1 0 7268 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0578_
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0579_
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0580_
timestamp 1704896540
transform 1 0 5612 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0581_
timestamp 1704896540
transform -1 0 8004 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0582_
timestamp 1704896540
transform 1 0 6440 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0583_
timestamp 1704896540
transform 1 0 6808 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0584_
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0585_
timestamp 1704896540
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0586_
timestamp 1704896540
transform 1 0 4324 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0587_
timestamp 1704896540
transform -1 0 6900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0588_
timestamp 1704896540
transform 1 0 5612 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0589_
timestamp 1704896540
transform 1 0 8464 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0590_
timestamp 1704896540
transform 1 0 6072 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0591_
timestamp 1704896540
transform 1 0 5796 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0592_
timestamp 1704896540
transform 1 0 6532 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0593_
timestamp 1704896540
transform -1 0 9660 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0594_
timestamp 1704896540
transform 1 0 7544 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0595_
timestamp 1704896540
transform 1 0 8188 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0596_
timestamp 1704896540
transform 1 0 3772 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0597_
timestamp 1704896540
transform 1 0 4600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0598_
timestamp 1704896540
transform 1 0 4876 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0599_
timestamp 1704896540
transform -1 0 9384 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0600_
timestamp 1704896540
transform 1 0 7544 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0601_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6256 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0602_
timestamp 1704896540
transform -1 0 5152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0603_
timestamp 1704896540
transform 1 0 3220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0604_
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0605_
timestamp 1704896540
transform 1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0606_
timestamp 1704896540
transform 1 0 3956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0607_
timestamp 1704896540
transform 1 0 3128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0608_
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0609_
timestamp 1704896540
transform -1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0610_
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0611_
timestamp 1704896540
transform -1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0612_
timestamp 1704896540
transform 1 0 2208 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0613_
timestamp 1704896540
transform -1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0614_
timestamp 1704896540
transform 1 0 2300 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0615_
timestamp 1704896540
transform -1 0 2300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0616_
timestamp 1704896540
transform 1 0 4692 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0617_
timestamp 1704896540
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0618_
timestamp 1704896540
transform 1 0 1656 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0619_
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0620_
timestamp 1704896540
transform 1 0 1656 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0621_
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0622_
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0623_
timestamp 1704896540
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0624_
timestamp 1704896540
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0625_
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0626_
timestamp 1704896540
transform 1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0627_
timestamp 1704896540
transform 1 0 8004 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0628_
timestamp 1704896540
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0629_
timestamp 1704896540
transform 1 0 4508 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0630_
timestamp 1704896540
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0631_
timestamp 1704896540
transform 1 0 3220 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0632_
timestamp 1704896540
transform 1 0 1472 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0633_
timestamp 1704896540
transform 1 0 4968 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0634_
timestamp 1704896540
transform -1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0635_
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0636_
timestamp 1704896540
transform -1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0637_
timestamp 1704896540
transform 1 0 2300 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0638_
timestamp 1704896540
transform -1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0639_
timestamp 1704896540
transform 1 0 4784 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0640_
timestamp 1704896540
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0641_
timestamp 1704896540
transform 1 0 8004 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0642_
timestamp 1704896540
transform 1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0643_
timestamp 1704896540
transform 1 0 6992 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0644_
timestamp 1704896540
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0645_
timestamp 1704896540
transform 1 0 2576 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0646_
timestamp 1704896540
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0647_
timestamp 1704896540
transform 1 0 2300 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0648_
timestamp 1704896540
transform -1 0 2208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0649_
timestamp 1704896540
transform 1 0 3956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0650_
timestamp 1704896540
transform 1 0 3312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0651_
timestamp 1704896540
transform 1 0 1748 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0652_
timestamp 1704896540
transform -1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9844 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_2  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0655_
timestamp 1704896540
transform 1 0 9844 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0656_
timestamp 1704896540
transform 1 0 14076 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0657_
timestamp 1704896540
transform 1 0 12696 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0658_
timestamp 1704896540
transform 1 0 13064 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0659_
timestamp 1704896540
transform 1 0 12144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0660_
timestamp 1704896540
transform 1 0 11500 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0661_
timestamp 1704896540
transform 1 0 11224 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0662_
timestamp 1704896540
transform 1 0 8924 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0663_
timestamp 1704896540
transform -1 0 9200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0664_
timestamp 1704896540
transform 1 0 3404 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0665_
timestamp 1704896540
transform -1 0 3220 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0666_
timestamp 1704896540
transform 1 0 3128 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0667_
timestamp 1704896540
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0668_
timestamp 1704896540
transform 1 0 2208 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0669_
timestamp 1704896540
transform -1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0670_
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0671_
timestamp 1704896540
transform -1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0672_
timestamp 1704896540
transform 1 0 10120 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0673_
timestamp 1704896540
transform -1 0 15272 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0674_
timestamp 1704896540
transform -1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0675_
timestamp 1704896540
transform 1 0 12052 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0676_
timestamp 1704896540
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0677_
timestamp 1704896540
transform 1 0 11960 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0678_
timestamp 1704896540
transform -1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0679_
timestamp 1704896540
transform -1 0 11132 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0680_
timestamp 1704896540
transform -1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0681_
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0682_
timestamp 1704896540
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0683_
timestamp 1704896540
transform -1 0 11224 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0684_
timestamp 1704896540
transform -1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0685_
timestamp 1704896540
transform 1 0 12512 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0686_
timestamp 1704896540
transform 1 0 11776 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0687_
timestamp 1704896540
transform 1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0688_
timestamp 1704896540
transform -1 0 12420 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0689_
timestamp 1704896540
transform 1 0 10304 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0690_
timestamp 1704896540
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0691_
timestamp 1704896540
transform 1 0 17940 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0692_
timestamp 1704896540
transform -1 0 17756 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0693_
timestamp 1704896540
transform 1 0 18216 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0694_
timestamp 1704896540
transform -1 0 17940 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0695_
timestamp 1704896540
transform -1 0 20148 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0696_
timestamp 1704896540
transform -1 0 21620 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0697_
timestamp 1704896540
transform -1 0 19044 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0698_
timestamp 1704896540
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0699_
timestamp 1704896540
transform 1 0 15732 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0700_
timestamp 1704896540
transform -1 0 16008 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0701_
timestamp 1704896540
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0702_
timestamp 1704896540
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0703_
timestamp 1704896540
transform -1 0 20148 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0704_
timestamp 1704896540
transform -1 0 20148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0705_
timestamp 1704896540
transform -1 0 21620 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0706_
timestamp 1704896540
transform -1 0 19872 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0707_
timestamp 1704896540
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0708_
timestamp 1704896540
transform 1 0 16652 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_2  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0710_
timestamp 1704896540
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0711_
timestamp 1704896540
transform 1 0 16376 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0712_
timestamp 1704896540
transform 1 0 16100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0713_
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0714_
timestamp 1704896540
transform -1 0 16560 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0715_
timestamp 1704896540
transform -1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0716_
timestamp 1704896540
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0717_
timestamp 1704896540
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0718_
timestamp 1704896540
transform 1 0 14076 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0719_
timestamp 1704896540
transform 1 0 13248 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0720_
timestamp 1704896540
transform 1 0 9568 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0721_
timestamp 1704896540
transform 1 0 8924 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0722_
timestamp 1704896540
transform 1 0 8280 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0723_
timestamp 1704896540
transform 1 0 6992 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0724_
timestamp 1704896540
transform 1 0 6440 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0725_
timestamp 1704896540
transform 1 0 5520 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0726_
timestamp 1704896540
transform 1 0 6900 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0727_
timestamp 1704896540
transform 1 0 5428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0728_
timestamp 1704896540
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0729_
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0730_
timestamp 1704896540
transform 1 0 10764 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0731_
timestamp 1704896540
transform -1 0 10764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0732_
timestamp 1704896540
transform 1 0 6992 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0733_
timestamp 1704896540
transform 1 0 6532 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0734_
timestamp 1704896540
transform -1 0 6624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0735_
timestamp 1704896540
transform -1 0 14812 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0736_
timestamp 1704896540
transform 1 0 14076 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0737_
timestamp 1704896540
transform -1 0 13248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0738_
timestamp 1704896540
transform 1 0 13984 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0739_
timestamp 1704896540
transform 1 0 13064 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0740_
timestamp 1704896540
transform -1 0 13064 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0741_
timestamp 1704896540
transform 1 0 11592 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0742_
timestamp 1704896540
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0743_
timestamp 1704896540
transform -1 0 11868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0744_
timestamp 1704896540
transform 1 0 9108 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0745_
timestamp 1704896540
transform -1 0 8832 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0746_
timestamp 1704896540
transform -1 0 9200 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0747_
timestamp 1704896540
transform 1 0 2852 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0748_
timestamp 1704896540
transform 1 0 2208 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0749_
timestamp 1704896540
transform -1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0750_
timestamp 1704896540
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0751_
timestamp 1704896540
transform 1 0 2024 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0752_
timestamp 1704896540
transform -1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0753_
timestamp 1704896540
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0754_
timestamp 1704896540
transform 1 0 1748 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0755_
timestamp 1704896540
transform -1 0 1748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0756_
timestamp 1704896540
transform 1 0 3128 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0757_
timestamp 1704896540
transform 1 0 1932 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0758_
timestamp 1704896540
transform -1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0759_
timestamp 1704896540
transform 1 0 10212 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0760_
timestamp 1704896540
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0761_
timestamp 1704896540
transform 1 0 15272 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0762_
timestamp 1704896540
transform 1 0 14536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0763_
timestamp 1704896540
transform 1 0 17480 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0764_
timestamp 1704896540
transform 1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0765_
timestamp 1704896540
transform -1 0 20884 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0766_
timestamp 1704896540
transform -1 0 21528 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0767_
timestamp 1704896540
transform -1 0 21252 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0768_
timestamp 1704896540
transform -1 0 19504 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0769_
timestamp 1704896540
transform 1 0 15456 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0770_
timestamp 1704896540
transform -1 0 15548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0771_
timestamp 1704896540
transform 1 0 17664 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0772_
timestamp 1704896540
transform 1 0 17020 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0773_
timestamp 1704896540
transform -1 0 20792 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0774_
timestamp 1704896540
transform -1 0 21620 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0775_
timestamp 1704896540
transform 1 0 19228 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0776_
timestamp 1704896540
transform -1 0 19044 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0777_
timestamp 1704896540
transform 1 0 17112 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0778_
timestamp 1704896540
transform 1 0 12788 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0779_
timestamp 1704896540
transform 1 0 14260 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0780_
timestamp 1704896540
transform -1 0 16192 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0781_
timestamp 1704896540
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0782_
timestamp 1704896540
transform -1 0 19136 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0783_
timestamp 1704896540
transform -1 0 19136 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0784_
timestamp 1704896540
transform -1 0 21528 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0785_
timestamp 1704896540
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0786_
timestamp 1704896540
transform -1 0 16560 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0787_
timestamp 1704896540
transform 1 0 20792 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0788_
timestamp 1704896540
transform -1 0 21712 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0789_
timestamp 1704896540
transform 1 0 17940 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0790_
timestamp 1704896540
transform -1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0791_
timestamp 1704896540
transform -1 0 15824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0792_
timestamp 1704896540
transform 1 0 12880 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0793_
timestamp 1704896540
transform -1 0 11592 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0794_
timestamp 1704896540
transform 1 0 5428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0795_
timestamp 1704896540
transform -1 0 5704 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0796_
timestamp 1704896540
transform 1 0 5520 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0797_
timestamp 1704896540
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _0798_
timestamp 1704896540
transform 1 0 10672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0799_
timestamp 1704896540
transform -1 0 11408 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0800_
timestamp 1704896540
transform -1 0 18032 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0801_
timestamp 1704896540
transform 1 0 15916 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0802_
timestamp 1704896540
transform 1 0 16468 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0803_
timestamp 1704896540
transform 1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0804_
timestamp 1704896540
transform 1 0 15088 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0805_
timestamp 1704896540
transform -1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0806_
timestamp 1704896540
transform 1 0 10028 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0807_
timestamp 1704896540
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0808_
timestamp 1704896540
transform 1 0 8096 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0809_
timestamp 1704896540
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0810_
timestamp 1704896540
transform 1 0 6900 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0811_
timestamp 1704896540
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0812_
timestamp 1704896540
transform 1 0 11500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0813_
timestamp 1704896540
transform 1 0 9568 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0814_
timestamp 1704896540
transform 1 0 7912 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0815_
timestamp 1704896540
transform 1 0 6716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0816_
timestamp 1704896540
transform 1 0 9844 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0817_
timestamp 1704896540
transform 1 0 15272 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0818_
timestamp 1704896540
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0819_
timestamp 1704896540
transform 1 0 14536 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0820_
timestamp 1704896540
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0821_
timestamp 1704896540
transform 1 0 15640 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0822_
timestamp 1704896540
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0823_
timestamp 1704896540
transform 1 0 14168 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0824_
timestamp 1704896540
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0825_
timestamp 1704896540
transform 1 0 15456 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0826_
timestamp 1704896540
transform -1 0 15640 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0827_
timestamp 1704896540
transform 1 0 17572 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0828_
timestamp 1704896540
transform -1 0 17664 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0829_
timestamp 1704896540
transform 1 0 19688 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0830_
timestamp 1704896540
transform 1 0 19228 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0831_
timestamp 1704896540
transform -1 0 21620 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0832_
timestamp 1704896540
transform 1 0 18952 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0833_
timestamp 1704896540
transform -1 0 10212 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0834_
timestamp 1704896540
transform 1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _0835_
timestamp 1704896540
transform -1 0 19136 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _0836_
timestamp 1704896540
transform 1 0 13800 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0837_
timestamp 1704896540
transform 1 0 13524 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0838_
timestamp 1704896540
transform 1 0 12604 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0839_
timestamp 1704896540
transform -1 0 12604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0840_
timestamp 1704896540
transform 1 0 16100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0841_
timestamp 1704896540
transform -1 0 13616 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0842_
timestamp 1704896540
transform -1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0843_
timestamp 1704896540
transform 1 0 10580 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0844_
timestamp 1704896540
transform -1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0845_
timestamp 1704896540
transform 1 0 10856 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0846_
timestamp 1704896540
transform -1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0847_
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0848_
timestamp 1704896540
transform 1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0849_
timestamp 1704896540
transform 1 0 13340 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0850_
timestamp 1704896540
transform 1 0 11500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0851_
timestamp 1704896540
transform 1 0 12420 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0852_
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0853_
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0854_
timestamp 1704896540
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0855_
timestamp 1704896540
transform 1 0 15640 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0856_
timestamp 1704896540
transform -1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0857_
timestamp 1704896540
transform -1 0 18032 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0858_
timestamp 1704896540
transform -1 0 15640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0859_
timestamp 1704896540
transform 1 0 14444 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0860_
timestamp 1704896540
transform -1 0 14168 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0861_
timestamp 1704896540
transform 1 0 16560 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0862_
timestamp 1704896540
transform 1 0 16652 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0863_
timestamp 1704896540
transform -1 0 16560 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0864_
timestamp 1704896540
transform -1 0 18584 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0865_
timestamp 1704896540
transform -1 0 18952 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0866_
timestamp 1704896540
transform -1 0 21344 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0867_
timestamp 1704896540
transform -1 0 21344 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0868_
timestamp 1704896540
transform 1 0 20792 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0869_
timestamp 1704896540
transform 1 0 19688 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0870_
timestamp 1704896540
transform -1 0 16928 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0871_
timestamp 1704896540
transform -1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0872_
timestamp 1704896540
transform 1 0 18308 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0873_
timestamp 1704896540
transform 1 0 16560 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0874_
timestamp 1704896540
transform 1 0 20608 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0875_
timestamp 1704896540
transform 1 0 19872 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0876_
timestamp 1704896540
transform 1 0 20792 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0877_
timestamp 1704896540
transform -1 0 19688 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0878_
timestamp 1704896540
transform 1 0 15732 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0879_
timestamp 1704896540
transform 1 0 14720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0880_
timestamp 1704896540
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0881_
timestamp 1704896540
transform -1 0 17940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0882_
timestamp 1704896540
transform 1 0 16284 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0883_
timestamp 1704896540
transform 1 0 20792 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0884_
timestamp 1704896540
transform -1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0885_
timestamp 1704896540
transform 1 0 19320 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0886_
timestamp 1704896540
transform 1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0887_
timestamp 1704896540
transform -1 0 18124 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0888_
timestamp 1704896540
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0889_
timestamp 1704896540
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0890_
timestamp 1704896540
transform 1 0 16928 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0891_
timestamp 1704896540
transform 1 0 20792 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0892_
timestamp 1704896540
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0893_
timestamp 1704896540
transform 1 0 17940 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0894_
timestamp 1704896540
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0895_
timestamp 1704896540
transform 1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0896_
timestamp 1704896540
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0897_
timestamp 1704896540
transform 1 0 17112 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0898_
timestamp 1704896540
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0899_
timestamp 1704896540
transform -1 0 21712 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0900_
timestamp 1704896540
transform -1 0 21620 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0901_
timestamp 1704896540
transform 1 0 20884 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0902_
timestamp 1704896540
transform 1 0 19136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0903_
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0904_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3956 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _0905_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1704896540
transform -1 0 3128 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1704896540
transform -1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1704896540
transform -1 0 4692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0909_
timestamp 1704896540
transform 1 0 12880 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0910_
timestamp 1704896540
transform 1 0 12604 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0911_
timestamp 1704896540
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0912_
timestamp 1704896540
transform 1 0 12512 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0913_
timestamp 1704896540
transform 1 0 10856 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0914_
timestamp 1704896540
transform 1 0 10488 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0915_
timestamp 1704896540
transform 1 0 7728 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0916_
timestamp 1704896540
transform -1 0 8004 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0917_
timestamp 1704896540
transform -1 0 5336 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0918_
timestamp 1704896540
transform -1 0 6532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0919_
timestamp 1704896540
transform -1 0 8648 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0920_
timestamp 1704896540
transform 1 0 8464 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0921_
timestamp 1704896540
transform -1 0 6256 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0922_
timestamp 1704896540
transform 1 0 5888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1704896540
transform 1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1704896540
transform 1 0 8464 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1704896540
transform 1 0 6624 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11408 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _0928_
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0929_
timestamp 1704896540
transform 1 0 13800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0930_
timestamp 1704896540
transform -1 0 13432 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0931_
timestamp 1704896540
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0932_
timestamp 1704896540
transform 1 0 11408 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0933_
timestamp 1704896540
transform 1 0 10672 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0934_
timestamp 1704896540
transform 1 0 10580 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0935_
timestamp 1704896540
transform -1 0 11500 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0936_
timestamp 1704896540
transform 1 0 11868 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0937_
timestamp 1704896540
transform 1 0 11592 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0938_
timestamp 1704896540
transform -1 0 13892 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0939_
timestamp 1704896540
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0940_
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1704896540
transform -1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0942_
timestamp 1704896540
transform 1 0 14260 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0943_
timestamp 1704896540
transform 1 0 11960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0944_
timestamp 1704896540
transform 1 0 14904 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0945_
timestamp 1704896540
transform -1 0 15180 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0946_
timestamp 1704896540
transform -1 0 15180 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0947_
timestamp 1704896540
transform -1 0 15180 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0948_
timestamp 1704896540
transform 1 0 13156 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1704896540
transform 1 0 12420 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0950_
timestamp 1704896540
transform 1 0 9660 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0951_
timestamp 1704896540
transform -1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0952_
timestamp 1704896540
transform -1 0 5428 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0953_
timestamp 1704896540
transform -1 0 5704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0954_
timestamp 1704896540
transform 1 0 4140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0955_
timestamp 1704896540
transform -1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _0956_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4140 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0957_
timestamp 1704896540
transform 1 0 2760 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0958_
timestamp 1704896540
transform -1 0 18400 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0959_
timestamp 1704896540
transform 1 0 17204 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0960_
timestamp 1704896540
transform 1 0 19228 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0961_
timestamp 1704896540
transform -1 0 18768 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0962_
timestamp 1704896540
transform 1 0 15640 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0963_
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0964_
timestamp 1704896540
transform 1 0 19780 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0965_
timestamp 1704896540
transform 1 0 19320 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0966_
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0967_
timestamp 1704896540
transform 1 0 8004 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0968_
timestamp 1704896540
transform -1 0 8832 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0969_
timestamp 1704896540
transform 1 0 5888 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0970_
timestamp 1704896540
transform 1 0 5980 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0971_
timestamp 1704896540
transform 1 0 6900 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0972_
timestamp 1704896540
transform 1 0 8188 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0973_
timestamp 1704896540
transform 1 0 2116 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0974_
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0975_
timestamp 1704896540
transform 1 0 5336 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0976_
timestamp 1704896540
transform 1 0 5428 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0977_
timestamp 1704896540
transform 1 0 1656 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0978_
timestamp 1704896540
transform 1 0 1656 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0979_
timestamp 1704896540
transform 1 0 4232 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0980_
timestamp 1704896540
transform -1 0 3036 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0981_
timestamp 1704896540
transform 1 0 1564 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0982_
timestamp 1704896540
transform 1 0 1932 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0983_
timestamp 1704896540
transform 1 0 8004 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0984_
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0985_
timestamp 1704896540
transform 1 0 4048 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0986_
timestamp 1704896540
transform 1 0 1748 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0987_
timestamp 1704896540
transform 1 0 4508 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0988_
timestamp 1704896540
transform 1 0 2760 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0989_
timestamp 1704896540
transform 1 0 1564 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0990_
timestamp 1704896540
transform 1 0 3680 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0991_
timestamp 1704896540
transform 1 0 7268 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0992_
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0993_
timestamp 1704896540
transform 1 0 2024 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0994_
timestamp 1704896540
transform 1 0 1564 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0995_
timestamp 1704896540
transform 1 0 3588 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0996_
timestamp 1704896540
transform 1 0 1840 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0997_
timestamp 1704896540
transform 1 0 12972 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0998_
timestamp 1704896540
transform 1 0 12420 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0999_
timestamp 1704896540
transform 1 0 11500 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1704896540
transform 1 0 8188 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1001_
timestamp 1704896540
transform 1 0 2116 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1002_
timestamp 1704896540
transform 1 0 2024 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1003_
timestamp 1704896540
transform 1 0 1840 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1004_
timestamp 1704896540
transform 1 0 2116 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1005_
timestamp 1704896540
transform 1 0 12880 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1006_
timestamp 1704896540
transform 1 0 11960 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1007_
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1008_
timestamp 1704896540
transform 1 0 9752 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1009_
timestamp 1704896540
transform 1 0 9844 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1010_
timestamp 1704896540
transform 1 0 9844 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1011_
timestamp 1704896540
transform 1 0 12052 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1012_
timestamp 1704896540
transform 1 0 11776 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1013_
timestamp 1704896540
transform 1 0 17204 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1014_
timestamp 1704896540
transform 1 0 17388 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1015_
timestamp 1704896540
transform 1 0 19780 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1016_
timestamp 1704896540
transform 1 0 19228 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1017_
timestamp 1704896540
transform 1 0 15272 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1018_
timestamp 1704896540
transform 1 0 18216 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1019_
timestamp 1704896540
transform 1 0 19412 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1020_
timestamp 1704896540
transform 1 0 19228 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1021_
timestamp 1704896540
transform 1 0 16652 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1022_
timestamp 1704896540
transform 1 0 15824 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1023_
timestamp 1704896540
transform 1 0 13248 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1024_
timestamp 1704896540
transform 1 0 8464 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1025_
timestamp 1704896540
transform 1 0 5704 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1026_
timestamp 1704896540
transform 1 0 6348 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1027_
timestamp 1704896540
transform 1 0 9844 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1028_
timestamp 1704896540
transform -1 0 6808 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1029_
timestamp 1704896540
transform 1 0 12420 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1030_
timestamp 1704896540
transform 1 0 12420 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1031_
timestamp 1704896540
transform 1 0 10488 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1032_
timestamp 1704896540
transform -1 0 8832 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1033_
timestamp 1704896540
transform 1 0 1380 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1034_
timestamp 1704896540
transform 1 0 1380 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1035_
timestamp 1704896540
transform 1 0 1380 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1036_
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1037_
timestamp 1704896540
transform 1 0 14812 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1038_
timestamp 1704896540
transform 1 0 17112 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1039_
timestamp 1704896540
transform 1 0 19964 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1040_
timestamp 1704896540
transform 1 0 18860 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1041_
timestamp 1704896540
transform 1 0 14996 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1042_
timestamp 1704896540
transform 1 0 17204 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1043_
timestamp 1704896540
transform 1 0 19964 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1044_
timestamp 1704896540
transform 1 0 18308 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1045_
timestamp 1704896540
transform 1 0 18216 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1046_
timestamp 1704896540
transform 1 0 18032 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1047_
timestamp 1704896540
transform 1 0 20148 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1048_
timestamp 1704896540
transform 1 0 19780 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1049_
timestamp 1704896540
transform 1 0 16376 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1050_
timestamp 1704896540
transform 1 0 19228 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1051_
timestamp 1704896540
transform 1 0 20148 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1052_
timestamp 1704896540
transform 1 0 20148 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1053_
timestamp 1704896540
transform -1 0 18216 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1054_
timestamp 1704896540
transform 1 0 14904 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1055_
timestamp 1704896540
transform -1 0 13984 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1056_
timestamp 1704896540
transform 1 0 9844 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1057_
timestamp 1704896540
transform 1 0 4324 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1058_
timestamp 1704896540
transform 1 0 4324 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1059_
timestamp 1704896540
transform -1 0 5796 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1060_
timestamp 1704896540
transform -1 0 5888 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1061_
timestamp 1704896540
transform 1 0 16192 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1062_
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1063_
timestamp 1704896540
transform 1 0 14812 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1064_
timestamp 1704896540
transform 1 0 8924 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1065_
timestamp 1704896540
transform 1 0 6440 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1066_
timestamp 1704896540
transform 1 0 6532 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1704896540
transform 1 0 10396 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1068_
timestamp 1704896540
transform 1 0 6808 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1069_
timestamp 1704896540
transform 1 0 14536 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1704896540
transform 1 0 14076 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1071_
timestamp 1704896540
transform 1 0 15640 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1072_
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1073_
timestamp 1704896540
transform 1 0 14996 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1074_
timestamp 1704896540
transform 1 0 17112 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1075_
timestamp 1704896540
transform 1 0 19504 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1076_
timestamp 1704896540
transform 1 0 19228 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1077_
timestamp 1704896540
transform -1 0 10580 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _1079_
timestamp 1704896540
transform 1 0 19780 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1080_
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1081_
timestamp 1704896540
transform 1 0 11868 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1082_
timestamp 1704896540
transform 1 0 11592 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1083_
timestamp 1704896540
transform 1 0 9844 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1084_
timestamp 1704896540
transform 1 0 10212 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1704896540
transform 1 0 10028 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1086_
timestamp 1704896540
transform 1 0 12052 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1087_
timestamp 1704896540
transform 1 0 11868 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1088_
timestamp 1704896540
transform 1 0 14536 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1089_
timestamp 1704896540
transform 1 0 14168 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1090_
timestamp 1704896540
transform 1 0 14996 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1091_
timestamp 1704896540
transform 1 0 13800 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1092_
timestamp 1704896540
transform 1 0 15088 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1093_
timestamp 1704896540
transform -1 0 18676 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1094_
timestamp 1704896540
transform 1 0 19964 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1095_
timestamp 1704896540
transform 1 0 19780 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1096_
timestamp 1704896540
transform 1 0 14904 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1097_
timestamp 1704896540
transform 1 0 17112 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1098_
timestamp 1704896540
transform 1 0 20148 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1099_
timestamp 1704896540
transform 1 0 19228 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1100_
timestamp 1704896540
transform 1 0 16560 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1101_
timestamp 1704896540
transform 1 0 17296 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1102_
timestamp 1704896540
transform 1 0 20148 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1103_
timestamp 1704896540
transform 1 0 19228 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1104_
timestamp 1704896540
transform -1 0 18492 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1105_
timestamp 1704896540
transform 1 0 17296 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1106_
timestamp 1704896540
transform 1 0 18952 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1107_
timestamp 1704896540
transform 1 0 17204 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1108_
timestamp 1704896540
transform 1 0 17204 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1109_
timestamp 1704896540
transform 1 0 16560 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1110_
timestamp 1704896540
transform 1 0 20148 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1111_
timestamp 1704896540
transform 1 0 19688 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1112_
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _1113_
timestamp 1704896540
transform 1 0 1564 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1114_
timestamp 1704896540
transform 1 0 1748 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1115_
timestamp 1704896540
transform 1 0 2944 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _1116_
timestamp 1704896540
transform 1 0 13708 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1117_
timestamp 1704896540
transform 1 0 12328 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1118_
timestamp 1704896540
transform -1 0 11316 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1119_
timestamp 1704896540
transform -1 0 8096 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1120_
timestamp 1704896540
transform -1 0 6164 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1121_
timestamp 1704896540
transform 1 0 8924 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1122_
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _1123_
timestamp 1704896540
transform 1 0 7544 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1124_
timestamp 1704896540
transform 1 0 7544 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1125_
timestamp 1704896540
transform 1 0 8096 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1126_
timestamp 1704896540
transform 1 0 5704 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _1127_
timestamp 1704896540
transform -1 0 14720 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1128_
timestamp 1704896540
transform -1 0 13800 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1129_
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1130_
timestamp 1704896540
transform 1 0 10948 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1131_
timestamp 1704896540
transform 1 0 12236 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1132_
timestamp 1704896540
transform -1 0 14260 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1133_
timestamp 1704896540
transform 1 0 10580 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1134_
timestamp 1704896540
transform 1 0 12144 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1135_
timestamp 1704896540
transform 1 0 14536 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1136_
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1137_
timestamp 1704896540
transform -1 0 13156 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1138_
timestamp 1704896540
transform 1 0 9292 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1139_
timestamp 1704896540
transform -1 0 5428 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1140_
timestamp 1704896540
transform 1 0 3312 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_spi_sck $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_spi_sck $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2760 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_spi_sck
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_spi_sck
timestamp 1704896540
transform -1 0 9936 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_spi_sck
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_spi_sck
timestamp 1704896540
transform 1 0 3036 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_spi_sck
timestamp 1704896540
transform -1 0 3312 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_spi_sck
timestamp 1704896540
transform 1 0 8004 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_spi_sck
timestamp 1704896540
transform 1 0 8556 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_spi_sck
timestamp 1704896540
transform 1 0 13432 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_spi_sck
timestamp 1704896540
transform 1 0 14444 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_spi_sck
timestamp 1704896540
transform 1 0 18124 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_spi_sck
timestamp 1704896540
transform 1 0 18952 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_spi_sck
timestamp 1704896540
transform -1 0 15088 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_spi_sck
timestamp 1704896540
transform -1 0 15088 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_spi_sck
timestamp 1704896540
transform 1 0 18676 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_spi_sck
timestamp 1704896540
transform 1 0 19044 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_22
timestamp 1704896540
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49
timestamp 1704896540
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1704896540
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_63
timestamp 1704896540
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_154
timestamp 1704896540
transform 1 0 15272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_158
timestamp 1704896540
transform 1 0 15640 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1704896540
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_192
timestamp 1704896540
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1704896540
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1704896540
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1704896540
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_22
timestamp 1704896540
transform 1 0 3128 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_45
timestamp 1704896540
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_49
timestamp 1704896540
transform 1 0 5612 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_74
timestamp 1704896540
transform 1 0 7912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_92
timestamp 1704896540
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_134
timestamp 1704896540
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_192
timestamp 1704896540
transform 1 0 18768 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_211
timestamp 1704896540
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1704896540
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_46
timestamp 1704896540
transform 1 0 5336 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_73
timestamp 1704896540
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_94
timestamp 1704896540
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_136
timestamp 1704896540
transform 1 0 13616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_223
timestamp 1704896540
transform 1 0 21620 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_24
timestamp 1704896540
transform 1 0 3312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_30
timestamp 1704896540
transform 1 0 3864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_49
timestamp 1704896540
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_88
timestamp 1704896540
transform 1 0 9200 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_136
timestamp 1704896540
transform 1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_173
timestamp 1704896540
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_192
timestamp 1704896540
transform 1 0 18768 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_209
timestamp 1704896540
transform 1 0 20332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_221
timestamp 1704896540
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_7
timestamp 1704896540
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_63
timestamp 1704896540
transform 1 0 6900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_73
timestamp 1704896540
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_102
timestamp 1704896540
transform 1 0 10488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_110
timestamp 1704896540
transform 1 0 11224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1704896540
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_185
timestamp 1704896540
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1704896540
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_197
timestamp 1704896540
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_205
timestamp 1704896540
transform 1 0 19964 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_26
timestamp 1704896540
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_30
timestamp 1704896540
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_40
timestamp 1704896540
transform 1 0 4784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_48
timestamp 1704896540
transform 1 0 5520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1704896540
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_66
timestamp 1704896540
transform 1 0 7176 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_72
timestamp 1704896540
transform 1 0 7728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_89
timestamp 1704896540
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_122
timestamp 1704896540
transform 1 0 12328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_159
timestamp 1704896540
transform 1 0 15732 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_195
timestamp 1704896540
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_199
timestamp 1704896540
transform 1 0 19412 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1704896540
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_21
timestamp 1704896540
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_62
timestamp 1704896540
transform 1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1704896540
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_96
timestamp 1704896540
transform 1 0 9936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_134
timestamp 1704896540
transform 1 0 13432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_167
timestamp 1704896540
transform 1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_171
timestamp 1704896540
transform 1 0 16836 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_192
timestamp 1704896540
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_35
timestamp 1704896540
transform 1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_74
timestamp 1704896540
transform 1 0 7912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_99
timestamp 1704896540
transform 1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1704896540
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_133
timestamp 1704896540
transform 1 0 13340 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_145
timestamp 1704896540
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_158
timestamp 1704896540
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1704896540
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_219
timestamp 1704896540
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1704896540
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_103
timestamp 1704896540
transform 1 0 10580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_115
timestamp 1704896540
transform 1 0 11684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_119
timestamp 1704896540
transform 1 0 12052 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_132
timestamp 1704896540
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1704896540
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_163
timestamp 1704896540
transform 1 0 16100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_171
timestamp 1704896540
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_175
timestamp 1704896540
transform 1 0 17204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_197
timestamp 1704896540
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_11
timestamp 1704896540
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_37
timestamp 1704896540
transform 1 0 4508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_48
timestamp 1704896540
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_65
timestamp 1704896540
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_74
timestamp 1704896540
transform 1 0 7912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_83
timestamp 1704896540
transform 1 0 8740 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_99
timestamp 1704896540
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_131
timestamp 1704896540
transform 1 0 13156 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_139
timestamp 1704896540
transform 1 0 13892 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1704896540
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_219
timestamp 1704896540
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1704896540
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_7
timestamp 1704896540
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1704896540
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_46
timestamp 1704896540
transform 1 0 5336 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_75
timestamp 1704896540
transform 1 0 8004 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1704896540
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_116
timestamp 1704896540
transform 1 0 11776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_135
timestamp 1704896540
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1704896540
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_169
timestamp 1704896540
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1704896540
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_223
timestamp 1704896540
transform 1 0 21620 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_31
timestamp 1704896540
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_61
timestamp 1704896540
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_69
timestamp 1704896540
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_94
timestamp 1704896540
transform 1 0 9752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_156
timestamp 1704896540
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_204
timestamp 1704896540
transform 1 0 19872 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1704896540
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_23
timestamp 1704896540
transform 1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_40
timestamp 1704896540
transform 1 0 4784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_49
timestamp 1704896540
transform 1 0 5612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_115
timestamp 1704896540
transform 1 0 11684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_137
timestamp 1704896540
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1704896540
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_206
timestamp 1704896540
transform 1 0 20056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_21
timestamp 1704896540
transform 1 0 3036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_37
timestamp 1704896540
transform 1 0 4508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_48
timestamp 1704896540
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_98
timestamp 1704896540
transform 1 0 10120 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1704896540
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1704896540
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_134
timestamp 1704896540
transform 1 0 13432 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_147
timestamp 1704896540
transform 1 0 14628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_180
timestamp 1704896540
transform 1 0 17664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_190
timestamp 1704896540
transform 1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1704896540
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_9
timestamp 1704896540
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_66
timestamp 1704896540
transform 1 0 7176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_80
timestamp 1704896540
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_91
timestamp 1704896540
transform 1 0 9476 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_100
timestamp 1704896540
transform 1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_107
timestamp 1704896540
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_111
timestamp 1704896540
transform 1 0 11316 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_121
timestamp 1704896540
transform 1 0 12236 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_134
timestamp 1704896540
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_148
timestamp 1704896540
transform 1 0 14720 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_154
timestamp 1704896540
transform 1 0 15272 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_164
timestamp 1704896540
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_191
timestamp 1704896540
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1704896540
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 1704896540
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_223
timestamp 1704896540
transform 1 0 21620 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_32
timestamp 1704896540
transform 1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1704896540
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_93
timestamp 1704896540
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_106
timestamp 1704896540
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_130
timestamp 1704896540
transform 1 0 13064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_148
timestamp 1704896540
transform 1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_173
timestamp 1704896540
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1704896540
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_24
timestamp 1704896540
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_62
timestamp 1704896540
transform 1 0 6808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_68
timestamp 1704896540
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_98
timestamp 1704896540
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_105
timestamp 1704896540
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_124
timestamp 1704896540
transform 1 0 12512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_150
timestamp 1704896540
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_178
timestamp 1704896540
transform 1 0 17480 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_188
timestamp 1704896540
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1704896540
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1704896540
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_222
timestamp 1704896540
transform 1 0 21528 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_22
timestamp 1704896540
transform 1 0 3128 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_47
timestamp 1704896540
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_69
timestamp 1704896540
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_101
timestamp 1704896540
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_141
timestamp 1704896540
transform 1 0 14076 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_149
timestamp 1704896540
transform 1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_155
timestamp 1704896540
transform 1 0 15364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_173
timestamp 1704896540
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_191
timestamp 1704896540
transform 1 0 18676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_220
timestamp 1704896540
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_12
timestamp 1704896540
transform 1 0 2208 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_22
timestamp 1704896540
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_40
timestamp 1704896540
transform 1 0 4784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_63
timestamp 1704896540
transform 1 0 6900 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_149
timestamp 1704896540
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_167
timestamp 1704896540
transform 1 0 16468 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_191
timestamp 1704896540
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1704896540
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1704896540
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1704896540
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_220
timestamp 1704896540
transform 1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_15
timestamp 1704896540
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_19
timestamp 1704896540
transform 1 0 2852 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_23
timestamp 1704896540
transform 1 0 3220 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_31
timestamp 1704896540
transform 1 0 3956 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_38
timestamp 1704896540
transform 1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_44
timestamp 1704896540
transform 1 0 5152 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_73
timestamp 1704896540
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_88
timestamp 1704896540
transform 1 0 9200 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_92
timestamp 1704896540
transform 1 0 9568 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1704896540
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_126
timestamp 1704896540
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_139
timestamp 1704896540
transform 1 0 13892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_145
timestamp 1704896540
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1704896540
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_172
timestamp 1704896540
transform 1 0 16928 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_196
timestamp 1704896540
transform 1 0 19136 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_204
timestamp 1704896540
transform 1 0 19872 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_215
timestamp 1704896540
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1704896540
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_39
timestamp 1704896540
transform 1 0 4692 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_78
timestamp 1704896540
transform 1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_107
timestamp 1704896540
transform 1 0 10948 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_115
timestamp 1704896540
transform 1 0 11684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1704896540
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_153
timestamp 1704896540
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_172
timestamp 1704896540
transform 1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1704896540
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1704896540
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_200
timestamp 1704896540
transform 1 0 19504 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_204
timestamp 1704896540
transform 1 0 19872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_222
timestamp 1704896540
transform 1 0 21528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_3
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_64
timestamp 1704896540
transform 1 0 6992 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_91
timestamp 1704896540
transform 1 0 9476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_152
timestamp 1704896540
transform 1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1704896540
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1704896540
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_3
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 1704896540
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_42
timestamp 1704896540
transform 1 0 4968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_52
timestamp 1704896540
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_59
timestamp 1704896540
transform 1 0 6532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_63
timestamp 1704896540
transform 1 0 6900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_67
timestamp 1704896540
transform 1 0 7268 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_100
timestamp 1704896540
transform 1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_147
timestamp 1704896540
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1704896540
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_223
timestamp 1704896540
transform 1 0 21620 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_15
timestamp 1704896540
transform 1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_31
timestamp 1704896540
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_43
timestamp 1704896540
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_69
timestamp 1704896540
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_75
timestamp 1704896540
transform 1 0 8004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_97
timestamp 1704896540
transform 1 0 10028 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_122
timestamp 1704896540
transform 1 0 12328 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_135
timestamp 1704896540
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_147
timestamp 1704896540
transform 1 0 14628 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_153
timestamp 1704896540
transform 1 0 15180 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_157
timestamp 1704896540
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_192
timestamp 1704896540
transform 1 0 18768 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_198
timestamp 1704896540
transform 1 0 19320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_202
timestamp 1704896540
transform 1 0 19688 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_38
timestamp 1704896540
transform 1 0 4600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_46
timestamp 1704896540
transform 1 0 5336 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_56
timestamp 1704896540
transform 1 0 6256 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_64
timestamp 1704896540
transform 1 0 6992 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_70
timestamp 1704896540
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1704896540
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_88
timestamp 1704896540
transform 1 0 9200 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_115
timestamp 1704896540
transform 1 0 11684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_127
timestamp 1704896540
transform 1 0 12788 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1704896540
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_153
timestamp 1704896540
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_164
timestamp 1704896540
transform 1 0 16192 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_176
timestamp 1704896540
transform 1 0 17296 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_183
timestamp 1704896540
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1704896540
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1704896540
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_209
timestamp 1704896540
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_221
timestamp 1704896540
transform 1 0 21436 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_3
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1704896540
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_83
timestamp 1704896540
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_102
timestamp 1704896540
transform 1 0 10488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_122
timestamp 1704896540
transform 1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_154
timestamp 1704896540
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_195
timestamp 1704896540
transform 1 0 19044 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_23
timestamp 1704896540
transform 1 0 3220 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_38
timestamp 1704896540
transform 1 0 4600 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_44
timestamp 1704896540
transform 1 0 5152 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_79
timestamp 1704896540
transform 1 0 8372 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_91
timestamp 1704896540
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_118
timestamp 1704896540
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_158
timestamp 1704896540
transform 1 0 15640 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1704896540
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_223
timestamp 1704896540
transform 1 0 21620 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_3
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_32
timestamp 1704896540
transform 1 0 4048 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_36
timestamp 1704896540
transform 1 0 4416 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1704896540
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_60
timestamp 1704896540
transform 1 0 6624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_73
timestamp 1704896540
transform 1 0 7820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_86
timestamp 1704896540
transform 1 0 9016 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_94
timestamp 1704896540
transform 1 0 9752 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_122
timestamp 1704896540
transform 1 0 12328 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_149
timestamp 1704896540
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1704896540
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_178
timestamp 1704896540
transform 1 0 17480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_183
timestamp 1704896540
transform 1 0 17940 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_3
timestamp 1704896540
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_7
timestamp 1704896540
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_38
timestamp 1704896540
transform 1 0 4600 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_68
timestamp 1704896540
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_72
timestamp 1704896540
transform 1 0 7728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_82
timestamp 1704896540
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_91
timestamp 1704896540
transform 1 0 9476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_101
timestamp 1704896540
transform 1 0 10396 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_114
timestamp 1704896540
transform 1 0 11592 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_120
timestamp 1704896540
transform 1 0 12144 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1704896540
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_177
timestamp 1704896540
transform 1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_197
timestamp 1704896540
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_3
timestamp 1704896540
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_33
timestamp 1704896540
transform 1 0 4140 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_51
timestamp 1704896540
transform 1 0 5796 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_74
timestamp 1704896540
transform 1 0 7912 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_106
timestamp 1704896540
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_122
timestamp 1704896540
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_130
timestamp 1704896540
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_153
timestamp 1704896540
transform 1 0 15180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1704896540
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_178
timestamp 1704896540
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_182
timestamp 1704896540
transform 1 0 17848 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_210
timestamp 1704896540
transform 1 0 20424 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_55
timestamp 1704896540
transform 1 0 6164 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_76
timestamp 1704896540
transform 1 0 8096 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_105
timestamp 1704896540
transform 1 0 10764 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_115
timestamp 1704896540
transform 1 0 11684 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_121
timestamp 1704896540
transform 1 0 12236 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1704896540
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_184
timestamp 1704896540
transform 1 0 18032 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1704896540
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_222
timestamp 1704896540
transform 1 0 21528 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_3
timestamp 1704896540
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_9
timestamp 1704896540
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_41
timestamp 1704896540
transform 1 0 4876 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_92
timestamp 1704896540
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1704896540
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_130
timestamp 1704896540
transform 1 0 13064 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1704896540
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1704896540
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1704896540
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1704896540
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_32
timestamp 1704896540
transform 1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_60
timestamp 1704896540
transform 1 0 6624 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_75
timestamp 1704896540
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1704896540
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_94
timestamp 1704896540
transform 1 0 9752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_108
timestamp 1704896540
transform 1 0 11040 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_113
timestamp 1704896540
transform 1 0 11500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_153
timestamp 1704896540
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_161
timestamp 1704896540
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_187
timestamp 1704896540
transform 1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_197
timestamp 1704896540
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_20
timestamp 1704896540
transform 1 0 2944 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_31
timestamp 1704896540
transform 1 0 3956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1704896540
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_85
timestamp 1704896540
transform 1 0 8924 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_96
timestamp 1704896540
transform 1 0 9936 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1704896540
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_126
timestamp 1704896540
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_136
timestamp 1704896540
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_149
timestamp 1704896540
transform 1 0 14812 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_157
timestamp 1704896540
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_177
timestamp 1704896540
transform 1 0 17388 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_181
timestamp 1704896540
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_185
timestamp 1704896540
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1704896540
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_3
timestamp 1704896540
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_9
timestamp 1704896540
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_75
timestamp 1704896540
transform 1 0 8004 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1704896540
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_88
timestamp 1704896540
transform 1 0 9200 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_119
timestamp 1704896540
transform 1 0 12052 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_153
timestamp 1704896540
transform 1 0 15180 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_171
timestamp 1704896540
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_192
timestamp 1704896540
transform 1 0 18768 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_214
timestamp 1704896540
transform 1 0 20792 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_23
timestamp 1704896540
transform 1 0 3220 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_34
timestamp 1704896540
transform 1 0 4232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_52
timestamp 1704896540
transform 1 0 5888 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_63
timestamp 1704896540
transform 1 0 6900 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_73
timestamp 1704896540
transform 1 0 7820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_94
timestamp 1704896540
transform 1 0 9752 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_122
timestamp 1704896540
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1704896540
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_220
timestamp 1704896540
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_3
timestamp 1704896540
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_7
timestamp 1704896540
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_29
timestamp 1704896540
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_88
timestamp 1704896540
transform 1 0 9200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_122
timestamp 1704896540
transform 1 0 12328 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_162
timestamp 1704896540
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_192
timestamp 1704896540
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_197
timestamp 1704896540
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_220
timestamp 1704896540
transform 1 0 21344 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_3
timestamp 1704896540
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_11
timestamp 1704896540
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_21
timestamp 1704896540
transform 1 0 3036 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_27
timestamp 1704896540
transform 1 0 3588 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_29
timestamp 1704896540
transform 1 0 3772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_37
timestamp 1704896540
transform 1 0 4508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1704896540
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1704896540
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_57
timestamp 1704896540
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_67
timestamp 1704896540
transform 1 0 7268 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_94
timestamp 1704896540
transform 1 0 9752 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_106
timestamp 1704896540
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_113
timestamp 1704896540
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_117
timestamp 1704896540
transform 1 0 11868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_132
timestamp 1704896540
transform 1 0 13248 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_141
timestamp 1704896540
transform 1 0 14076 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_153
timestamp 1704896540
transform 1 0 15180 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_159
timestamp 1704896540
transform 1 0 15732 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_185
timestamp 1704896540
transform 1 0 18124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_205
timestamp 1704896540
transform 1 0 19964 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1704896540
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6624 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 6716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 20424 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 19964 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform 1 0 20056 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform -1 0 21712 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform -1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform 1 0 20056 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform -1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform 1 0 4784 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 16560 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform 1 0 4784 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform -1 0 12328 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  max_cap1
timestamp 1704896540
transform -1 0 10120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_38
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_39
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_40
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_41
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_42
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_43
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 21988 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_44
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_45
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 21988 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_46
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_47
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_48
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_49
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 21988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_50
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 21988 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_51
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_52
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_53
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_54
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 21988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_55
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_56
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 21988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_57
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_58
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_59
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_60
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_61
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_62
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 21988 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_63
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 21988 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_64
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 21988 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_65
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 21988 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_66
timestamp 1704896540
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_67
timestamp 1704896540
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_68
timestamp 1704896540
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 21988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_69
timestamp 1704896540
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_70
timestamp 1704896540
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 21988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_71
timestamp 1704896540
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_72
timestamp 1704896540
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 21988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_73
timestamp 1704896540
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1704896540
transform -1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_74
timestamp 1704896540
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1704896540
transform -1 0 21988 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_75
timestamp 1704896540
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1704896540
transform -1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_84
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_85
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_93
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_94
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_97
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_98
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_99
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_100
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_101
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_102
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_103
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_104
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_105
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_106
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_107
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_108
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_109
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_110
timestamp 1704896540
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_111
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_112
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_113
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_114
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_115
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_116
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp 1704896540
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_121
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_122
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_123
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_124
timestamp 1704896540
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_125
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_126
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_127
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_128
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_129
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_130
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_131
timestamp 1704896540
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_132
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_133
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_134
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_135
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_136
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_137
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_138
timestamp 1704896540
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_139
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_140
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_141
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_142
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_143
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_144
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_145
timestamp 1704896540
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_146
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_147
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_148
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_149
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_150
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_151
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_152
timestamp 1704896540
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_153
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_154
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_155
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_156
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_157
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_158
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_159
timestamp 1704896540
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_160
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_161
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_162
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_163
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_164
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_165
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_166
timestamp 1704896540
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_167
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_168
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_169
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_170
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_171
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_172
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_173
timestamp 1704896540
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_174
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_175
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_176
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_177
timestamp 1704896540
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_178
timestamp 1704896540
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_179
timestamp 1704896540
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_180
timestamp 1704896540
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_181
timestamp 1704896540
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_182
timestamp 1704896540
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_183
timestamp 1704896540
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_184
timestamp 1704896540
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_185
timestamp 1704896540
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_186
timestamp 1704896540
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_187
timestamp 1704896540
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_188
timestamp 1704896540
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_189
timestamp 1704896540
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_190
timestamp 1704896540
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_191
timestamp 1704896540
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_192
timestamp 1704896540
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_193
timestamp 1704896540
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_194
timestamp 1704896540
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_195
timestamp 1704896540
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_196
timestamp 1704896540
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_197
timestamp 1704896540
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_198
timestamp 1704896540
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_199
timestamp 1704896540
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_200
timestamp 1704896540
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_201
timestamp 1704896540
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_202
timestamp 1704896540
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_203
timestamp 1704896540
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_204
timestamp 1704896540
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_205
timestamp 1704896540
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_206
timestamp 1704896540
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_207
timestamp 1704896540
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_208
timestamp 1704896540
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_209
timestamp 1704896540
transform 1 0 3680 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_210
timestamp 1704896540
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_211
timestamp 1704896540
transform 1 0 8832 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_212
timestamp 1704896540
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_213
timestamp 1704896540
transform 1 0 13984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_214
timestamp 1704896540
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_215
timestamp 1704896540
transform 1 0 19136 0 -1 22848
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 spi_cs_n
port 0 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 spi_miso
port 1 nsew signal output
flabel metal2 s 16762 24475 16818 25275 0 FreeSans 224 90 0 0 spi_mosi
port 2 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 spi_sck
port 3 nsew signal input
flabel metal4 s 3554 2128 3874 22896 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 8775 2128 9095 22896 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 13996 2128 14316 22896 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 19217 2128 19537 22896 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal5 s 1056 4600 22036 4920 0 FreeSans 2560 0 0 0 vccd1
port 4 nsew power bidirectional
flabel metal5 s 1056 9768 22036 10088 0 FreeSans 2560 0 0 0 vccd1
port 4 nsew power bidirectional
flabel metal5 s 1056 14936 22036 15256 0 FreeSans 2560 0 0 0 vccd1
port 4 nsew power bidirectional
flabel metal5 s 1056 20104 22036 20424 0 FreeSans 2560 0 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 4214 2128 4534 22896 0 FreeSans 1920 90 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal4 s 9435 2128 9755 22896 0 FreeSans 1920 90 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal4 s 14656 2128 14976 22896 0 FreeSans 1920 90 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal4 s 19877 2128 20197 22896 0 FreeSans 1920 90 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal5 s 1056 5260 22036 5580 0 FreeSans 2560 0 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal5 s 1056 10428 22036 10748 0 FreeSans 2560 0 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal5 s 1056 15596 22036 15916 0 FreeSans 2560 0 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal5 s 1056 20764 22036 21084 0 FreeSans 2560 0 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal2 s 17406 24475 17462 25275 0 FreeSans 224 90 0 0 wbs_adr_o[0]
port 6 nsew signal output
flabel metal2 s 12254 24475 12310 25275 0 FreeSans 224 90 0 0 wbs_adr_o[10]
port 7 nsew signal output
flabel metal2 s 9034 24475 9090 25275 0 FreeSans 224 90 0 0 wbs_adr_o[11]
port 8 nsew signal output
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 wbs_adr_o[12]
port 9 nsew signal output
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 wbs_adr_o[13]
port 10 nsew signal output
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 wbs_adr_o[14]
port 11 nsew signal output
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 wbs_adr_o[15]
port 12 nsew signal output
flabel metal2 s 19338 24475 19394 25275 0 FreeSans 224 90 0 0 wbs_adr_o[16]
port 13 nsew signal output
flabel metal3 s 22331 19048 23131 19168 0 FreeSans 480 0 0 0 wbs_adr_o[17]
port 14 nsew signal output
flabel metal3 s 22331 20408 23131 20528 0 FreeSans 480 0 0 0 wbs_adr_o[18]
port 15 nsew signal output
flabel metal3 s 22331 21088 23131 21208 0 FreeSans 480 0 0 0 wbs_adr_o[19]
port 16 nsew signal output
flabel metal3 s 22331 16328 23131 16448 0 FreeSans 480 0 0 0 wbs_adr_o[1]
port 17 nsew signal output
flabel metal2 s 18050 24475 18106 25275 0 FreeSans 224 90 0 0 wbs_adr_o[20]
port 18 nsew signal output
flabel metal3 s 22331 19728 23131 19848 0 FreeSans 480 0 0 0 wbs_adr_o[21]
port 19 nsew signal output
flabel metal3 s 22331 18368 23131 18488 0 FreeSans 480 0 0 0 wbs_adr_o[22]
port 20 nsew signal output
flabel metal3 s 22331 17008 23131 17128 0 FreeSans 480 0 0 0 wbs_adr_o[23]
port 21 nsew signal output
flabel metal2 s 16118 24475 16174 25275 0 FreeSans 224 90 0 0 wbs_adr_o[24]
port 22 nsew signal output
flabel metal3 s 22331 17688 23131 17808 0 FreeSans 480 0 0 0 wbs_adr_o[25]
port 23 nsew signal output
flabel metal2 s 12898 24475 12954 25275 0 FreeSans 224 90 0 0 wbs_adr_o[26]
port 24 nsew signal output
flabel metal2 s 10966 24475 11022 25275 0 FreeSans 224 90 0 0 wbs_adr_o[27]
port 25 nsew signal output
flabel metal2 s 5814 24475 5870 25275 0 FreeSans 224 90 0 0 wbs_adr_o[28]
port 26 nsew signal output
flabel metal2 s 5170 24475 5226 25275 0 FreeSans 224 90 0 0 wbs_adr_o[29]
port 27 nsew signal output
flabel metal2 s 14830 24475 14886 25275 0 FreeSans 224 90 0 0 wbs_adr_o[2]
port 28 nsew signal output
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 wbs_adr_o[30]
port 29 nsew signal output
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 wbs_adr_o[31]
port 30 nsew signal output
flabel metal2 s 9678 24475 9734 25275 0 FreeSans 224 90 0 0 wbs_adr_o[3]
port 31 nsew signal output
flabel metal2 s 7102 24475 7158 25275 0 FreeSans 224 90 0 0 wbs_adr_o[4]
port 32 nsew signal output
flabel metal2 s 7746 24475 7802 25275 0 FreeSans 224 90 0 0 wbs_adr_o[5]
port 33 nsew signal output
flabel metal2 s 11610 24475 11666 25275 0 FreeSans 224 90 0 0 wbs_adr_o[6]
port 34 nsew signal output
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 wbs_adr_o[7]
port 35 nsew signal output
flabel metal2 s 14186 24475 14242 25275 0 FreeSans 224 90 0 0 wbs_adr_o[8]
port 36 nsew signal output
flabel metal2 s 13542 24475 13598 25275 0 FreeSans 224 90 0 0 wbs_adr_o[9]
port 37 nsew signal output
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 wbs_cyc_o
port 38 nsew signal output
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 39 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 40 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 41 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 wbs_dat_i[12]
port 42 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 wbs_dat_i[13]
port 43 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 wbs_dat_i[14]
port 44 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 wbs_dat_i[15]
port 45 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 wbs_dat_i[16]
port 46 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 wbs_dat_i[17]
port 47 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 48 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 49 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 wbs_dat_i[1]
port 50 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 wbs_dat_i[20]
port 51 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 wbs_dat_i[21]
port 52 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 wbs_dat_i[22]
port 53 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 wbs_dat_i[23]
port 54 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 wbs_dat_i[24]
port 55 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 56 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 57 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 58 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 wbs_dat_i[28]
port 59 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 wbs_dat_i[29]
port 60 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 61 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 wbs_dat_i[30]
port 62 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 wbs_dat_i[31]
port 63 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 64 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 wbs_dat_i[4]
port 65 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 wbs_dat_i[5]
port 66 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 wbs_dat_i[6]
port 67 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 wbs_dat_i[7]
port 68 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 wbs_dat_i[8]
port 69 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 70 nsew signal input
flabel metal3 s 22331 4088 23131 4208 0 FreeSans 480 0 0 0 wbs_dat_o[0]
port 71 nsew signal output
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 72 nsew signal output
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 73 nsew signal output
flabel metal3 s 22331 10888 23131 11008 0 FreeSans 480 0 0 0 wbs_dat_o[12]
port 74 nsew signal output
flabel metal3 s 22331 10208 23131 10328 0 FreeSans 480 0 0 0 wbs_dat_o[13]
port 75 nsew signal output
flabel metal3 s 22331 11568 23131 11688 0 FreeSans 480 0 0 0 wbs_dat_o[14]
port 76 nsew signal output
flabel metal3 s 22331 9528 23131 9648 0 FreeSans 480 0 0 0 wbs_dat_o[15]
port 77 nsew signal output
flabel metal3 s 22331 12928 23131 13048 0 FreeSans 480 0 0 0 wbs_dat_o[16]
port 78 nsew signal output
flabel metal3 s 22331 12248 23131 12368 0 FreeSans 480 0 0 0 wbs_dat_o[17]
port 79 nsew signal output
flabel metal3 s 22331 13608 23131 13728 0 FreeSans 480 0 0 0 wbs_dat_o[18]
port 80 nsew signal output
flabel metal3 s 22331 14288 23131 14408 0 FreeSans 480 0 0 0 wbs_dat_o[19]
port 81 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 82 nsew signal output
flabel metal3 s 22331 15648 23131 15768 0 FreeSans 480 0 0 0 wbs_dat_o[20]
port 83 nsew signal output
flabel metal3 s 22331 14968 23131 15088 0 FreeSans 480 0 0 0 wbs_dat_o[21]
port 84 nsew signal output
flabel metal3 s 22331 6808 23131 6928 0 FreeSans 480 0 0 0 wbs_dat_o[22]
port 85 nsew signal output
flabel metal3 s 22331 8168 23131 8288 0 FreeSans 480 0 0 0 wbs_dat_o[23]
port 86 nsew signal output
flabel metal3 s 22331 7488 23131 7608 0 FreeSans 480 0 0 0 wbs_dat_o[24]
port 87 nsew signal output
flabel metal3 s 22331 5448 23131 5568 0 FreeSans 480 0 0 0 wbs_dat_o[25]
port 88 nsew signal output
flabel metal3 s 22331 3408 23131 3528 0 FreeSans 480 0 0 0 wbs_dat_o[26]
port 89 nsew signal output
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 90 nsew signal output
flabel metal3 s 22331 8848 23131 8968 0 FreeSans 480 0 0 0 wbs_dat_o[28]
port 91 nsew signal output
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 92 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 93 nsew signal output
flabel metal3 s 22331 4768 23131 4888 0 FreeSans 480 0 0 0 wbs_dat_o[30]
port 94 nsew signal output
flabel metal3 s 22331 6128 23131 6248 0 FreeSans 480 0 0 0 wbs_dat_o[31]
port 95 nsew signal output
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 96 nsew signal output
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 97 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 98 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 99 nsew signal output
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 100 nsew signal output
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 101 nsew signal output
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 102 nsew signal output
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 wbs_stb_o
port 103 nsew signal output
flabel metal3 s 22331 21768 23131 21888 0 FreeSans 480 0 0 0 wbs_we_o
port 104 nsew signal output
rlabel metal1 11546 22304 11546 22304 0 vccd1
rlabel metal1 11546 22848 11546 22848 0 vssd1
rlabel metal2 1610 14178 1610 14178 0 _0000_
rlabel metal2 2070 13600 2070 13600 0 _0001_
rlabel metal2 3266 14144 3266 14144 0 _0002_
rlabel metal1 7130 12682 7130 12682 0 _0003_
rlabel metal2 2990 14586 2990 14586 0 _0004_
rlabel metal2 3082 13090 3082 13090 0 _0005_
rlabel metal2 4554 13736 4554 13736 0 _0006_
rlabel metal1 8043 11798 8043 11798 0 _0007_
rlabel metal2 8602 13736 8602 13736 0 _0008_
rlabel metal2 9062 15198 9062 15198 0 _0009_
rlabel metal1 6900 14246 6900 14246 0 _0010_
rlabel metal1 3818 17850 3818 17850 0 _0011_
rlabel metal1 3261 16150 3261 16150 0 _0012_
rlabel metal1 18277 7786 18277 7786 0 _0013_
rlabel metal1 17418 5610 17418 5610 0 _0014_
rlabel metal1 19637 3434 19637 3434 0 _0015_
rlabel metal1 18691 3094 18691 3094 0 _0016_
rlabel metal2 16146 8194 16146 8194 0 _0017_
rlabel metal1 16872 5202 16872 5202 0 _0018_
rlabel metal1 19902 5270 19902 5270 0 _0019_
rlabel metal2 19458 6562 19458 6562 0 _0020_
rlabel metal1 6568 6290 6568 6290 0 _0021_
rlabel via1 8321 6358 8321 6358 0 _0022_
rlabel metal2 7958 6290 7958 6290 0 _0023_
rlabel metal2 6578 7650 6578 7650 0 _0024_
rlabel metal1 5964 8874 5964 8874 0 _0025_
rlabel metal2 7590 9316 7590 9316 0 _0026_
rlabel metal1 8034 8534 8034 8534 0 _0027_
rlabel metal1 2238 4522 2238 4522 0 _0028_
rlabel metal1 3710 3434 3710 3434 0 _0029_
rlabel via1 5653 4590 5653 4590 0 _0030_
rlabel metal2 5750 3298 5750 3298 0 _0031_
rlabel via1 1973 8942 1973 8942 0 _0032_
rlabel metal1 2024 10234 2024 10234 0 _0033_
rlabel metal1 4354 9962 4354 9962 0 _0034_
rlabel via1 2718 5678 2718 5678 0 _0035_
rlabel metal1 1778 3094 1778 3094 0 _0036_
rlabel metal1 2152 5202 2152 5202 0 _0037_
rlabel via1 8321 3094 8321 3094 0 _0038_
rlabel metal1 8602 4250 8602 4250 0 _0039_
rlabel metal1 4268 8466 4268 8466 0 _0040_
rlabel metal1 1968 11118 1968 11118 0 _0041_
rlabel metal1 5009 11118 5009 11118 0 _0042_
rlabel metal1 3261 6290 3261 6290 0 _0043_
rlabel metal2 1978 3026 1978 3026 0 _0044_
rlabel metal1 3802 3094 3802 3094 0 _0045_
rlabel metal1 7390 2346 7390 2346 0 _0046_
rlabel metal1 6568 3026 6568 3026 0 _0047_
rlabel metal1 2244 8466 2244 8466 0 _0048_
rlabel via1 1881 11730 1881 11730 0 _0049_
rlabel metal1 3710 11798 3710 11798 0 _0050_
rlabel metal2 2254 7650 2254 7650 0 _0051_
rlabel metal1 13192 21522 13192 21522 0 _0052_
rlabel metal1 12374 16456 12374 16456 0 _0053_
rlabel metal1 11720 19346 11720 19346 0 _0054_
rlabel metal1 8740 21114 8740 21114 0 _0055_
rlabel metal2 2990 21794 2990 21794 0 _0056_
rlabel metal1 2300 19482 2300 19482 0 _0057_
rlabel metal2 1978 17306 1978 17306 0 _0058_
rlabel metal2 2990 15912 2990 15912 0 _0059_
rlabel metal1 13335 8534 13335 8534 0 _0060_
rlabel metal1 12180 7854 12180 7854 0 _0061_
rlabel via1 11817 2414 11817 2414 0 _0062_
rlabel metal1 10759 3094 10759 3094 0 _0063_
rlabel metal1 10391 8466 10391 8466 0 _0064_
rlabel metal1 10897 5270 10897 5270 0 _0065_
rlabel metal1 12174 4522 12174 4522 0 _0066_
rlabel metal1 12139 6358 12139 6358 0 _0067_
rlabel metal2 17526 20706 17526 20706 0 _0068_
rlabel via1 17705 16558 17705 16558 0 _0069_
rlabel metal1 20741 19414 20741 19414 0 _0070_
rlabel metal1 19442 20842 19442 20842 0 _0071_
rlabel metal2 15778 21352 15778 21352 0 _0072_
rlabel metal1 18436 19346 18436 19346 0 _0073_
rlabel metal1 19637 16082 19637 16082 0 _0074_
rlabel metal1 19591 16490 19591 16490 0 _0075_
rlabel via1 16969 19346 16969 19346 0 _0076_
rlabel metal1 16371 16558 16371 16558 0 _0077_
rlabel metal1 13524 18394 13524 18394 0 _0078_
rlabel metal1 8684 18258 8684 18258 0 _0079_
rlabel metal1 5796 22406 5796 22406 0 _0080_
rlabel metal1 6424 18326 6424 18326 0 _0081_
rlabel metal1 10345 17238 10345 17238 0 _0082_
rlabel via1 6490 16558 6490 16558 0 _0083_
rlabel metal1 12875 21998 12875 21998 0 _0084_
rlabel metal1 12783 17238 12783 17238 0 _0085_
rlabel metal1 11362 22406 11362 22406 0 _0086_
rlabel metal1 8878 21862 8878 21862 0 _0087_
rlabel via1 1697 21522 1697 21522 0 _0088_
rlabel metal1 1748 20026 1748 20026 0 _0089_
rlabel metal2 1518 18530 1518 18530 0 _0090_
rlabel metal2 1702 16354 1702 16354 0 _0091_
rlabel metal1 14934 12886 14934 12886 0 _0092_
rlabel metal1 17234 11798 17234 11798 0 _0093_
rlabel via1 20281 13294 20281 13294 0 _0094_
rlabel metal1 19136 13498 19136 13498 0 _0095_
rlabel via1 15313 14382 15313 14382 0 _0096_
rlabel metal1 17296 14042 17296 14042 0 _0097_
rlabel via1 20281 8534 20281 8534 0 _0098_
rlabel metal1 18763 8466 18763 8466 0 _0099_
rlabel via1 18533 21522 18533 21522 0 _0100_
rlabel metal1 18487 17170 18487 17170 0 _0101_
rlabel metal1 20695 19822 20695 19822 0 _0102_
rlabel metal1 21022 22406 21022 22406 0 _0103_
rlabel metal1 16330 22406 16330 22406 0 _0104_
rlabel metal1 20005 18666 20005 18666 0 _0105_
rlabel metal2 21114 16762 21114 16762 0 _0106_
rlabel via1 20465 17170 20465 17170 0 _0107_
rlabel metal2 16790 20910 16790 20910 0 _0108_
rlabel via1 15221 17238 15221 17238 0 _0109_
rlabel metal2 13478 20570 13478 20570 0 _0110_
rlabel metal1 10483 21590 10483 21590 0 _0111_
rlabel metal1 5239 21522 5239 21522 0 _0112_
rlabel metal1 4871 19754 4871 19754 0 _0113_
rlabel metal1 5576 18258 5576 18258 0 _0114_
rlabel via1 5570 16150 5570 16150 0 _0115_
rlabel metal1 16314 18666 16314 18666 0 _0116_
rlabel via1 16969 16082 16969 16082 0 _0117_
rlabel via1 15129 19414 15129 19414 0 _0118_
rlabel metal1 9000 18666 9000 18666 0 _0119_
rlabel metal1 6660 20910 6660 20910 0 _0120_
rlabel metal1 6654 18666 6654 18666 0 _0121_
rlabel metal1 10294 16558 10294 16558 0 _0122_
rlabel metal1 7028 16558 7028 16558 0 _0123_
rlabel metal1 14658 7446 14658 7446 0 _0124_
rlabel metal1 14152 5610 14152 5610 0 _0125_
rlabel metal2 15594 3298 15594 3298 0 _0126_
rlabel metal1 14152 3434 14152 3434 0 _0127_
rlabel metal1 15364 10234 15364 10234 0 _0128_
rlabel metal2 17434 9826 17434 9826 0 _0129_
rlabel metal1 19626 11798 19626 11798 0 _0130_
rlabel metal1 19350 10710 19350 10710 0 _0131_
rlabel metal2 10166 8466 10166 8466 0 _0132_
rlabel metal1 5520 12274 5520 12274 0 _0133_
rlabel metal1 19688 20026 19688 20026 0 _0134_
rlabel metal1 14066 8942 14066 8942 0 _0135_
rlabel via1 12185 8874 12185 8874 0 _0136_
rlabel metal1 12811 3162 12811 3162 0 _0137_
rlabel via1 10161 3502 10161 3502 0 _0138_
rlabel metal1 11035 7854 11035 7854 0 _0139_
rlabel metal1 9936 5338 9936 5338 0 _0140_
rlabel metal1 12036 4182 12036 4182 0 _0141_
rlabel via1 12185 5678 12185 5678 0 _0142_
rlabel via1 14853 6766 14853 6766 0 _0143_
rlabel metal1 14945 5270 14945 5270 0 _0144_
rlabel metal1 15364 2618 15364 2618 0 _0145_
rlabel metal1 14014 3094 14014 3094 0 _0146_
rlabel metal1 15865 11118 15865 11118 0 _0147_
rlabel metal1 18456 10642 18456 10642 0 _0148_
rlabel metal1 20695 11118 20695 11118 0 _0149_
rlabel metal1 20000 10030 20000 10030 0 _0150_
rlabel metal1 15957 12138 15957 12138 0 _0151_
rlabel metal1 17096 12138 17096 12138 0 _0152_
rlabel metal1 20270 15062 20270 15062 0 _0153_
rlabel metal1 19591 14314 19591 14314 0 _0154_
rlabel metal1 15900 14314 15900 14314 0 _0155_
rlabel metal1 17659 13974 17659 13974 0 _0156_
rlabel metal2 21022 8194 21022 8194 0 _0157_
rlabel metal1 19412 6086 19412 6086 0 _0158_
rlabel metal1 18461 7446 18461 7446 0 _0159_
rlabel metal2 17158 6018 17158 6018 0 _0160_
rlabel metal1 19166 3094 19166 3094 0 _0161_
rlabel metal1 17326 2346 17326 2346 0 _0162_
rlabel metal2 16882 8194 16882 8194 0 _0163_
rlabel metal1 16682 4522 16682 4522 0 _0164_
rlabel metal1 20925 4590 20925 4590 0 _0165_
rlabel metal1 19672 6358 19672 6358 0 _0166_
rlabel metal2 5382 6086 5382 6086 0 _0167_
rlabel metal1 13784 16150 13784 16150 0 _0168_
rlabel metal2 12742 18530 12742 18530 0 _0169_
rlabel metal2 10718 19142 10718 19142 0 _0170_
rlabel metal2 7774 20230 7774 20230 0 _0171_
rlabel metal1 6256 17850 6256 17850 0 _0172_
rlabel metal1 9144 16082 9144 16082 0 _0173_
rlabel metal1 6568 16082 6568 16082 0 _0174_
rlabel metal1 8648 12682 8648 12682 0 _0175_
rlabel metal2 7866 14110 7866 14110 0 _0176_
rlabel metal2 7774 14688 7774 14688 0 _0177_
rlabel metal2 6026 13804 6026 13804 0 _0178_
rlabel via1 14402 10710 14402 10710 0 _0179_
rlabel via1 13482 11730 13482 11730 0 _0180_
rlabel metal1 11086 10234 11086 10234 0 _0181_
rlabel via1 11265 11118 11265 11118 0 _0182_
rlabel metal1 12450 13226 12450 13226 0 _0183_
rlabel via1 13942 13974 13942 13974 0 _0184_
rlabel metal1 11173 14382 11173 14382 0 _0185_
rlabel metal2 12466 13906 12466 13906 0 _0186_
rlabel metal1 14904 21114 14904 21114 0 _0187_
rlabel via1 14393 16558 14393 16558 0 _0188_
rlabel via1 12838 19822 12838 19822 0 _0189_
rlabel metal1 9338 21114 9338 21114 0 _0190_
rlabel metal1 5474 21896 5474 21896 0 _0191_
rlabel metal1 3721 19414 3721 19414 0 _0192_
rlabel metal1 9292 10642 9292 10642 0 _0193_
rlabel metal1 4810 2414 4810 2414 0 _0194_
rlabel metal1 8372 13362 8372 13362 0 _0195_
rlabel metal2 10626 15538 10626 15538 0 _0196_
rlabel metal1 10166 11118 10166 11118 0 _0197_
rlabel metal1 5842 11050 5842 11050 0 _0198_
rlabel metal2 7314 12070 7314 12070 0 _0199_
rlabel metal2 5290 13906 5290 13906 0 _0200_
rlabel metal1 7590 13498 7590 13498 0 _0201_
rlabel metal1 9844 14314 9844 14314 0 _0202_
rlabel metal2 6854 13464 6854 13464 0 _0203_
rlabel metal1 8602 14341 8602 14341 0 _0204_
rlabel metal1 10626 12886 10626 12886 0 _0205_
rlabel metal1 9798 13362 9798 13362 0 _0206_
rlabel metal2 13018 13770 13018 13770 0 _0207_
rlabel metal2 10626 11254 10626 11254 0 _0208_
rlabel metal1 10212 13362 10212 13362 0 _0209_
rlabel via1 9246 13294 9246 13294 0 _0210_
rlabel metal2 9154 13872 9154 13872 0 _0211_
rlabel metal1 7406 14450 7406 14450 0 _0212_
rlabel metal1 8510 12818 8510 12818 0 _0213_
rlabel metal1 6118 12784 6118 12784 0 _0214_
rlabel metal2 9890 11152 9890 11152 0 _0215_
rlabel metal1 12006 12818 12006 12818 0 _0216_
rlabel metal2 5658 13566 5658 13566 0 _0217_
rlabel metal1 13110 12410 13110 12410 0 _0218_
rlabel metal1 13754 11288 13754 11288 0 _0219_
rlabel metal2 6946 13396 6946 13396 0 _0220_
rlabel metal1 6394 12886 6394 12886 0 _0221_
rlabel metal2 4002 13770 4002 13770 0 _0222_
rlabel metal1 18400 17510 18400 17510 0 _0223_
rlabel metal2 5658 14178 5658 14178 0 _0224_
rlabel metal2 10718 14382 10718 14382 0 _0225_
rlabel metal1 10442 13498 10442 13498 0 _0226_
rlabel metal1 14214 19754 14214 19754 0 _0227_
rlabel metal1 3680 17646 3680 17646 0 _0228_
rlabel metal1 20976 16422 20976 16422 0 _0229_
rlabel metal1 3772 16558 3772 16558 0 _0230_
rlabel metal1 15180 13226 15180 13226 0 _0231_
rlabel metal1 14444 10030 14444 10030 0 _0232_
rlabel metal1 18446 7854 18446 7854 0 _0233_
rlabel metal1 13248 15334 13248 15334 0 _0234_
rlabel metal1 17158 6290 17158 6290 0 _0235_
rlabel metal1 19550 19822 19550 19822 0 _0236_
rlabel metal1 19449 4114 19449 4114 0 _0237_
rlabel metal1 10902 2414 10902 2414 0 _0238_
rlabel metal1 18906 3502 18906 3502 0 _0239_
rlabel metal1 16330 20468 16330 20468 0 _0240_
rlabel metal2 16330 8364 16330 8364 0 _0241_
rlabel metal1 18354 13158 18354 13158 0 _0242_
rlabel metal1 16376 5202 16376 5202 0 _0243_
rlabel metal2 19550 5508 19550 5508 0 _0244_
rlabel metal2 19642 6732 19642 6732 0 _0245_
rlabel via1 9706 9690 9706 9690 0 _0246_
rlabel metal2 8510 10812 8510 10812 0 _0247_
rlabel metal2 8142 11356 8142 11356 0 _0248_
rlabel metal2 7406 10302 7406 10302 0 _0249_
rlabel metal1 8970 8942 8970 8942 0 _0250_
rlabel metal1 5980 5882 5980 5882 0 _0251_
rlabel metal2 6854 10336 6854 10336 0 _0252_
rlabel metal2 9798 6358 9798 6358 0 _0253_
rlabel metal2 4830 5270 4830 5270 0 _0254_
rlabel metal1 4646 5678 4646 5678 0 _0255_
rlabel metal2 5198 6290 5198 6290 0 _0256_
rlabel metal1 8602 13294 8602 13294 0 _0257_
rlabel metal1 6394 6698 6394 6698 0 _0258_
rlabel metal1 7866 5814 7866 5814 0 _0259_
rlabel metal1 9614 3978 9614 3978 0 _0260_
rlabel metal1 9430 6290 9430 6290 0 _0261_
rlabel metal1 9982 6426 9982 6426 0 _0262_
rlabel metal1 13018 17578 13018 17578 0 _0263_
rlabel metal2 9706 7004 9706 7004 0 _0264_
rlabel metal1 8268 5168 8268 5168 0 _0265_
rlabel metal2 7774 4556 7774 4556 0 _0266_
rlabel metal1 8464 5270 8464 5270 0 _0267_
rlabel metal1 8372 5814 8372 5814 0 _0268_
rlabel metal1 8464 5678 8464 5678 0 _0269_
rlabel metal1 7084 7310 7084 7310 0 _0270_
rlabel metal1 5666 8806 5666 8806 0 _0271_
rlabel metal2 5658 8262 5658 8262 0 _0272_
rlabel metal1 6394 7446 6394 7446 0 _0273_
rlabel metal1 7222 7446 7222 7446 0 _0274_
rlabel metal1 6532 8534 6532 8534 0 _0275_
rlabel metal1 4600 11322 4600 11322 0 _0276_
rlabel metal1 4554 9418 4554 9418 0 _0277_
rlabel metal2 5842 10030 5842 10030 0 _0278_
rlabel metal1 6348 9554 6348 9554 0 _0279_
rlabel metal1 7981 8942 7981 8942 0 _0280_
rlabel metal2 6670 10676 6670 10676 0 _0281_
rlabel metal1 6486 10030 6486 10030 0 _0282_
rlabel metal1 7406 8942 7406 8942 0 _0283_
rlabel metal1 8280 8874 8280 8874 0 _0284_
rlabel metal2 7866 8840 7866 8840 0 _0285_
rlabel metal1 5014 7276 5014 7276 0 _0286_
rlabel metal2 4922 7174 4922 7174 0 _0287_
rlabel metal1 6578 7242 6578 7242 0 _0288_
rlabel metal1 8648 7446 8648 7446 0 _0289_
rlabel metal1 5106 12852 5106 12852 0 _0290_
rlabel metal1 4784 12138 4784 12138 0 _0291_
rlabel metal2 2346 5134 2346 5134 0 _0292_
rlabel metal1 1886 4692 1886 4692 0 _0293_
rlabel metal2 3174 3706 3174 3706 0 _0294_
rlabel metal1 6164 5202 6164 5202 0 _0295_
rlabel metal2 5934 3468 5934 3468 0 _0296_
rlabel metal1 2254 9554 2254 9554 0 _0297_
rlabel metal1 2346 10030 2346 10030 0 _0298_
rlabel metal2 4830 9656 4830 9656 0 _0299_
rlabel metal1 2530 6222 2530 6222 0 _0300_
rlabel metal1 1610 4114 1610 4114 0 _0301_
rlabel metal1 2254 3910 2254 3910 0 _0302_
rlabel metal1 4002 2550 4002 2550 0 _0303_
rlabel metal2 7958 3910 7958 3910 0 _0304_
rlabel metal2 8234 4420 8234 4420 0 _0305_
rlabel metal1 4094 8942 4094 8942 0 _0306_
rlabel metal1 1518 11084 1518 11084 0 _0307_
rlabel metal2 5106 11118 5106 11118 0 _0308_
rlabel metal1 3763 6766 3763 6766 0 _0309_
rlabel metal1 2300 2414 2300 2414 0 _0310_
rlabel metal1 4186 3502 4186 3502 0 _0311_
rlabel metal1 7590 2414 7590 2414 0 _0312_
rlabel metal2 6026 3230 6026 3230 0 _0313_
rlabel metal1 2254 6834 2254 6834 0 _0314_
rlabel metal1 2300 12206 2300 12206 0 _0315_
rlabel metal2 3358 11900 3358 11900 0 _0316_
rlabel metal1 2162 6970 2162 6970 0 _0317_
rlabel metal1 10810 13940 10810 13940 0 _0318_
rlabel metal2 9982 16082 9982 16082 0 _0319_
rlabel metal1 5543 22202 5543 22202 0 _0320_
rlabel metal2 12742 21318 12742 21318 0 _0321_
rlabel metal2 12190 16116 12190 16116 0 _0322_
rlabel metal1 11454 18122 11454 18122 0 _0323_
rlabel metal1 9108 22406 9108 22406 0 _0324_
rlabel metal1 3358 21522 3358 21522 0 _0325_
rlabel metal2 2070 19788 2070 19788 0 _0326_
rlabel metal1 2254 17170 2254 17170 0 _0327_
rlabel metal1 3358 16558 3358 16558 0 _0328_
rlabel metal1 12098 2618 12098 2618 0 _0329_
rlabel metal1 13662 8908 13662 8908 0 _0330_
rlabel metal1 12006 8466 12006 8466 0 _0331_
rlabel metal1 12006 3502 12006 3502 0 _0332_
rlabel metal1 11178 2618 11178 2618 0 _0333_
rlabel metal2 11638 8092 11638 8092 0 _0334_
rlabel metal1 11454 5678 11454 5678 0 _0335_
rlabel metal2 11822 4794 11822 4794 0 _0336_
rlabel metal2 12466 6970 12466 6970 0 _0337_
rlabel metal2 15502 15606 15502 15606 0 _0338_
rlabel metal2 18906 15810 18906 15810 0 _0339_
rlabel metal1 17894 20434 17894 20434 0 _0340_
rlabel metal1 18170 15946 18170 15946 0 _0341_
rlabel metal1 21528 19346 21528 19346 0 _0342_
rlabel metal2 18906 20604 18906 20604 0 _0343_
rlabel metal2 15962 21148 15962 21148 0 _0344_
rlabel metal2 18078 19380 18078 19380 0 _0345_
rlabel metal1 20194 17170 20194 17170 0 _0346_
rlabel metal1 19826 17204 19826 17204 0 _0347_
rlabel via1 14674 17085 14674 17085 0 _0348_
rlabel metal2 16790 18938 16790 18938 0 _0349_
rlabel metal1 2576 20842 2576 20842 0 _0350_
rlabel metal1 11086 22134 11086 22134 0 _0351_
rlabel metal1 16330 19822 16330 19822 0 _0352_
rlabel metal1 16146 16184 16146 16184 0 _0353_
rlabel metal1 16560 15946 16560 15946 0 _0354_
rlabel metal1 14352 19958 14352 19958 0 _0355_
rlabel metal1 7038 22610 7038 22610 0 _0356_
rlabel metal1 13294 18224 13294 18224 0 _0357_
rlabel metal1 9660 19890 9660 19890 0 _0358_
rlabel metal1 8372 18734 8372 18734 0 _0359_
rlabel metal1 7084 21386 7084 21386 0 _0360_
rlabel metal1 6072 22610 6072 22610 0 _0361_
rlabel metal2 5842 19550 5842 19550 0 _0362_
rlabel metal2 6026 18700 6026 18700 0 _0363_
rlabel metal1 11500 15946 11500 15946 0 _0364_
rlabel metal1 10810 17646 10810 17646 0 _0365_
rlabel metal1 7029 17306 7029 17306 0 _0366_
rlabel metal2 6578 17476 6578 17476 0 _0367_
rlabel metal1 14628 20298 14628 20298 0 _0368_
rlabel metal1 13524 22610 13524 22610 0 _0369_
rlabel metal1 13791 17306 13791 17306 0 _0370_
rlabel metal2 13018 18054 13018 18054 0 _0371_
rlabel metal2 11730 20910 11730 20910 0 _0372_
rlabel metal1 11730 22610 11730 22610 0 _0373_
rlabel metal2 8418 22345 8418 22345 0 _0374_
rlabel metal2 8694 22243 8694 22243 0 _0375_
rlabel metal1 2760 22542 2760 22542 0 _0376_
rlabel metal2 2070 22202 2070 22202 0 _0377_
rlabel metal1 2622 21012 2622 21012 0 _0378_
rlabel metal2 1978 20434 1978 20434 0 _0379_
rlabel metal1 2346 18258 2346 18258 0 _0380_
rlabel metal1 1794 18258 1794 18258 0 _0381_
rlabel metal1 3082 14858 3082 14858 0 _0382_
rlabel metal1 1978 16082 1978 16082 0 _0383_
rlabel metal1 15134 11764 15134 11764 0 _0384_
rlabel via1 20378 12818 20378 12818 0 _0385_
rlabel metal2 14582 12988 14582 12988 0 _0386_
rlabel metal1 17250 12614 17250 12614 0 _0387_
rlabel metal2 20746 13294 20746 13294 0 _0388_
rlabel metal1 19688 13294 19688 13294 0 _0389_
rlabel metal1 15594 13804 15594 13804 0 _0390_
rlabel metal2 17066 13702 17066 13702 0 _0391_
rlabel metal2 20654 9724 20654 9724 0 _0392_
rlabel metal1 19173 8942 19173 8942 0 _0393_
rlabel viali 21208 22610 21208 22610 0 _0394_
rlabel metal1 13800 10030 13800 10030 0 _0395_
rlabel metal1 15364 9962 15364 9962 0 _0396_
rlabel metal2 15594 17068 15594 17068 0 _0397_
rlabel metal1 21206 22678 21206 22678 0 _0398_
rlabel metal2 11270 15266 11270 15266 0 _0399_
rlabel metal1 17250 19754 17250 19754 0 _0400_
rlabel metal1 16514 18734 16514 18734 0 _0401_
rlabel metal2 16882 16660 16882 16660 0 _0402_
rlabel metal1 15180 19822 15180 19822 0 _0403_
rlabel metal2 10166 18428 10166 18428 0 _0404_
rlabel metal1 7820 20230 7820 20230 0 _0405_
rlabel metal1 6716 18734 6716 18734 0 _0406_
rlabel metal1 9660 16558 9660 16558 0 _0407_
rlabel metal1 7958 15946 7958 15946 0 _0408_
rlabel metal1 20884 10574 20884 10574 0 _0409_
rlabel metal2 14306 7684 14306 7684 0 _0410_
rlabel metal2 13754 5882 13754 5882 0 _0411_
rlabel metal1 15594 3026 15594 3026 0 _0412_
rlabel metal2 13754 3774 13754 3774 0 _0413_
rlabel metal2 15594 10778 15594 10778 0 _0414_
rlabel metal2 17618 10404 17618 10404 0 _0415_
rlabel metal2 19274 11900 19274 11900 0 _0416_
rlabel metal1 20240 10642 20240 10642 0 _0417_
rlabel metal2 9982 7548 9982 7548 0 _0418_
rlabel metal1 13754 9554 13754 9554 0 _0419_
rlabel metal1 12650 9554 12650 9554 0 _0420_
rlabel metal1 14490 2414 14490 2414 0 _0421_
rlabel metal2 13386 3332 13386 3332 0 _0422_
rlabel metal1 10626 4114 10626 4114 0 _0423_
rlabel metal2 11730 8772 11730 8772 0 _0424_
rlabel metal1 9614 5236 9614 5236 0 _0425_
rlabel metal2 11730 4828 11730 4828 0 _0426_
rlabel metal2 12282 6528 12282 6528 0 _0427_
rlabel metal2 14030 7650 14030 7650 0 _0428_
rlabel metal2 15594 6086 15594 6086 0 _0429_
rlabel metal1 16192 2414 16192 2414 0 _0430_
rlabel metal1 14352 4114 14352 4114 0 _0431_
rlabel metal1 18860 14450 18860 14450 0 _0432_
rlabel metal2 16514 11526 16514 11526 0 _0433_
rlabel metal1 18676 9418 18676 9418 0 _0434_
rlabel metal2 21298 12036 21298 12036 0 _0435_
rlabel metal2 20930 10234 20930 10234 0 _0436_
rlabel metal2 16882 13124 16882 13124 0 _0437_
rlabel metal1 17526 12410 17526 12410 0 _0438_
rlabel metal1 20102 14994 20102 14994 0 _0439_
rlabel metal1 19688 14994 19688 14994 0 _0440_
rlabel metal2 14766 14620 14766 14620 0 _0441_
rlabel metal1 18078 15470 18078 15470 0 _0442_
rlabel metal2 21022 4556 21022 4556 0 _0443_
rlabel metal2 21206 7684 21206 7684 0 _0444_
rlabel metal1 18952 6290 18952 6290 0 _0445_
rlabel metal2 18906 7412 18906 7412 0 _0446_
rlabel metal1 16974 5780 16974 5780 0 _0447_
rlabel metal1 18998 4080 18998 4080 0 _0448_
rlabel metal2 16974 3468 16974 3468 0 _0449_
rlabel metal1 17158 7378 17158 7378 0 _0450_
rlabel metal1 16928 3978 16928 3978 0 _0451_
rlabel metal2 21574 5508 21574 5508 0 _0452_
rlabel metal2 19182 6460 19182 6460 0 _0453_
rlabel metal1 4002 5168 4002 5168 0 _0454_
rlabel metal1 5382 5066 5382 5066 0 _0455_
rlabel metal1 12834 16082 12834 16082 0 _0456_
rlabel metal2 12558 18054 12558 18054 0 _0457_
rlabel metal1 10764 18734 10764 18734 0 _0458_
rlabel metal2 7958 19652 7958 19652 0 _0459_
rlabel metal1 5851 17306 5851 17306 0 _0460_
rlabel metal2 8510 17170 8510 17170 0 _0461_
rlabel metal2 5934 15878 5934 15878 0 _0462_
rlabel metal1 12604 13838 12604 13838 0 _0463_
rlabel metal2 13846 11526 13846 11526 0 _0464_
rlabel metal2 13386 11764 13386 11764 0 _0465_
rlabel metal1 11132 10030 11132 10030 0 _0466_
rlabel metal1 11270 12206 11270 12206 0 _0467_
rlabel metal1 11813 13906 11813 13906 0 _0468_
rlabel metal2 13754 13532 13754 13532 0 _0469_
rlabel metal2 11638 15164 11638 15164 0 _0470_
rlabel metal2 13846 13498 13846 13498 0 _0471_
rlabel metal1 15088 20910 15088 20910 0 _0472_
rlabel metal2 15134 16966 15134 16966 0 _0473_
rlabel metal2 12466 20230 12466 20230 0 _0474_
rlabel metal1 9697 20910 9697 20910 0 _0475_
rlabel metal2 5658 21556 5658 21556 0 _0476_
rlabel metal2 4002 20026 4002 20026 0 _0477_
rlabel metal2 17618 19346 17618 19346 0 addr\[0\]
rlabel metal2 12098 18836 12098 18836 0 addr\[10\]
rlabel metal1 9108 22134 9108 22134 0 addr\[11\]
rlabel metal2 3910 21182 3910 21182 0 addr\[12\]
rlabel metal1 3542 20536 3542 20536 0 addr\[13\]
rlabel metal2 3266 18224 3266 18224 0 addr\[14\]
rlabel metal1 4094 15606 4094 15606 0 addr\[15\]
rlabel metal1 19780 22542 19780 22542 0 addr\[16\]
rlabel metal1 19596 16422 19596 16422 0 addr\[17\]
rlabel metal1 21252 19482 21252 19482 0 addr\[18\]
rlabel metal1 20378 22542 20378 22542 0 addr\[19\]
rlabel metal1 17572 15878 17572 15878 0 addr\[1\]
rlabel metal1 17434 22542 17434 22542 0 addr\[20\]
rlabel metal2 19642 19958 19642 19958 0 addr\[21\]
rlabel metal2 21022 17204 21022 17204 0 addr\[22\]
rlabel metal1 20608 16762 20608 16762 0 addr\[23\]
rlabel metal1 16376 22542 16376 22542 0 addr\[24\]
rlabel metal1 15594 16694 15594 16694 0 addr\[25\]
rlabel metal1 13570 19720 13570 19720 0 addr\[26\]
rlabel metal1 10718 21896 10718 21896 0 addr\[27\]
rlabel metal2 4830 22311 4830 22311 0 addr\[28\]
rlabel metal1 5106 19482 5106 19482 0 addr\[29\]
rlabel metal2 16238 19618 16238 19618 0 addr\[2\]
rlabel metal2 2714 18598 2714 18598 0 addr\[30\]
rlabel metal1 4508 16218 4508 16218 0 addr\[31\]
rlabel metal1 10396 18326 10396 18326 0 addr\[3\]
rlabel metal1 8142 21046 8142 21046 0 addr\[4\]
rlabel metal2 7498 19108 7498 19108 0 addr\[5\]
rlabel metal1 11868 16762 11868 16762 0 addr\[6\]
rlabel metal1 8096 16694 8096 16694 0 addr\[7\]
rlabel metal2 14490 21114 14490 21114 0 addr\[8\]
rlabel metal2 13846 17000 13846 17000 0 addr\[9\]
rlabel metal1 1925 13906 1925 13906 0 bit_count\[0\]
rlabel metal1 3174 13498 3174 13498 0 bit_count\[1\]
rlabel metal2 4738 14076 4738 14076 0 bit_count\[2\]
rlabel metal2 15042 17391 15042 17391 0 clknet_0_spi_sck
rlabel metal1 1978 5236 1978 5236 0 clknet_4_0_0_spi_sck
rlabel metal1 17986 2414 17986 2414 0 clknet_4_10_0_spi_sck
rlabel metal2 17158 11968 17158 11968 0 clknet_4_11_0_spi_sck
rlabel metal1 14306 13838 14306 13838 0 clknet_4_12_0_spi_sck
rlabel metal1 15226 20978 15226 20978 0 clknet_4_13_0_spi_sck
rlabel metal1 19642 17102 19642 17102 0 clknet_4_14_0_spi_sck
rlabel metal1 19550 18734 19550 18734 0 clknet_4_15_0_spi_sck
rlabel metal1 2070 8500 2070 8500 0 clknet_4_1_0_spi_sck
rlabel metal1 8050 6324 8050 6324 0 clknet_4_2_0_spi_sck
rlabel metal2 10534 10064 10534 10064 0 clknet_4_3_0_spi_sck
rlabel metal2 1886 17476 1886 17476 0 clknet_4_4_0_spi_sck
rlabel metal1 1426 21556 1426 21556 0 clknet_4_5_0_spi_sck
rlabel metal1 9890 16626 9890 16626 0 clknet_4_6_0_spi_sck
rlabel metal2 6118 19312 6118 19312 0 clknet_4_7_0_spi_sck
rlabel metal1 13892 3570 13892 3570 0 clknet_4_8_0_spi_sck
rlabel metal1 13846 9010 13846 9010 0 clknet_4_9_0_spi_sck
rlabel metal1 13800 12206 13800 12206 0 command\[0\]
rlabel metal1 13064 11050 13064 11050 0 command\[1\]
rlabel metal2 12558 10880 12558 10880 0 command\[2\]
rlabel metal1 11684 11526 11684 11526 0 command\[3\]
rlabel metal2 13478 14144 13478 14144 0 command\[4\]
rlabel metal1 13064 13702 13064 13702 0 command\[5\]
rlabel metal1 12926 15028 12926 15028 0 command\[6\]
rlabel metal2 13570 14144 13570 14144 0 command\[7\]
rlabel metal1 14352 8602 14352 8602 0 data_in\[0\]
rlabel metal2 17066 3264 17066 3264 0 data_in\[10\]
rlabel metal1 15134 3706 15134 3706 0 data_in\[11\]
rlabel metal1 16238 10778 16238 10778 0 data_in\[12\]
rlabel metal1 18354 10234 18354 10234 0 data_in\[13\]
rlabel metal1 20516 12070 20516 12070 0 data_in\[14\]
rlabel metal1 21206 10710 21206 10710 0 data_in\[15\]
rlabel metal1 16330 13260 16330 13260 0 data_in\[16\]
rlabel metal1 18676 12886 18676 12886 0 data_in\[17\]
rlabel metal1 21298 13498 21298 13498 0 data_in\[18\]
rlabel metal2 20838 14110 20838 14110 0 data_in\[19\]
rlabel metal2 12650 8296 12650 8296 0 data_in\[1\]
rlabel metal1 16146 14246 16146 14246 0 data_in\[20\]
rlabel metal1 18492 14246 18492 14246 0 data_in\[21\]
rlabel metal1 21298 8602 21298 8602 0 data_in\[22\]
rlabel metal2 19734 7888 19734 7888 0 data_in\[23\]
rlabel metal2 16974 8296 16974 8296 0 data_in\[24\]
rlabel metal1 18722 5814 18722 5814 0 data_in\[25\]
rlabel metal2 20654 3944 20654 3944 0 data_in\[26\]
rlabel metal2 18262 3264 18262 3264 0 data_in\[27\]
rlabel metal2 17066 9384 17066 9384 0 data_in\[28\]
rlabel metal2 18078 4624 18078 4624 0 data_in\[29\]
rlabel metal1 12972 2618 12972 2618 0 data_in\[2\]
rlabel metal1 20884 5542 20884 5542 0 data_in\[30\]
rlabel metal2 20746 7208 20746 7208 0 data_in\[31\]
rlabel metal1 10856 2278 10856 2278 0 data_in\[3\]
rlabel metal1 11592 8330 11592 8330 0 data_in\[4\]
rlabel metal2 11270 5848 11270 5848 0 data_in\[5\]
rlabel metal1 13524 5270 13524 5270 0 data_in\[6\]
rlabel metal1 12972 6698 12972 6698 0 data_in\[7\]
rlabel metal1 15870 7820 15870 7820 0 data_in\[8\]
rlabel metal2 15502 6120 15502 6120 0 data_in\[9\]
rlabel metal2 6762 5032 6762 5032 0 data_out\[10\]
rlabel metal2 6946 3944 6946 3944 0 data_out\[11\]
rlabel metal2 3082 8364 3082 8364 0 data_out\[12\]
rlabel metal2 2898 9758 2898 9758 0 data_out\[13\]
rlabel metal2 5658 9758 5658 9758 0 data_out\[14\]
rlabel metal2 3266 6902 3266 6902 0 data_out\[15\]
rlabel metal1 4094 2448 4094 2448 0 data_out\[16\]
rlabel metal1 4002 5338 4002 5338 0 data_out\[17\]
rlabel metal2 9522 3740 9522 3740 0 data_out\[18\]
rlabel metal1 9476 4454 9476 4454 0 data_out\[19\]
rlabel metal1 5336 8602 5336 8602 0 data_out\[20\]
rlabel metal2 3818 10880 3818 10880 0 data_out\[21\]
rlabel metal1 6210 10982 6210 10982 0 data_out\[22\]
rlabel via1 4646 6630 4646 6630 0 data_out\[23\]
rlabel metal1 3358 2414 3358 2414 0 data_out\[24\]
rlabel metal1 5244 4182 5244 4182 0 data_out\[25\]
rlabel metal1 8648 2618 8648 2618 0 data_out\[26\]
rlabel metal1 7544 3434 7544 3434 0 data_out\[27\]
rlabel metal1 3312 8262 3312 8262 0 data_out\[28\]
rlabel metal2 2990 11322 2990 11322 0 data_out\[29\]
rlabel metal1 5566 11594 5566 11594 0 data_out\[30\]
rlabel metal1 3174 7718 3174 7718 0 data_out\[31\]
rlabel metal1 3956 4454 3956 4454 0 data_out\[8\]
rlabel metal2 5290 4148 5290 4148 0 data_out\[9\]
rlabel metal2 9154 10812 9154 10812 0 net1
rlabel metal2 21482 20604 21482 20604 0 net10
rlabel metal1 16974 22610 16974 22610 0 net11
rlabel metal1 20792 22610 20792 22610 0 net12
rlabel metal1 17848 17850 17848 17850 0 net13
rlabel metal2 5474 21658 5474 21658 0 net14
rlabel metal1 12926 20502 12926 20502 0 net15
rlabel metal1 15824 17646 15824 17646 0 net16
rlabel metal2 5382 17340 5382 17340 0 net17
rlabel metal1 11592 21998 11592 21998 0 net18
rlabel metal1 5796 20026 5796 20026 0 net2
rlabel via1 5833 5746 5833 5746 0 net3
rlabel metal2 5566 18190 5566 18190 0 net4
rlabel metal2 21666 17068 21666 17068 0 net5
rlabel metal1 19366 17646 19366 17646 0 net6
rlabel metal1 19182 22610 19182 22610 0 net7
rlabel metal2 20838 19482 20838 19482 0 net8
rlabel metal2 17342 21420 17342 21420 0 net9
rlabel metal2 15962 16286 15962 16286 0 shift_in\[0\]
rlabel metal1 13754 19788 13754 19788 0 shift_in\[1\]
rlabel metal2 9890 18564 9890 18564 0 shift_in\[2\]
rlabel metal2 6670 21080 6670 21080 0 shift_in\[3\]
rlabel metal2 4738 19720 4738 19720 0 shift_in\[4\]
rlabel metal1 11270 16184 11270 16184 0 shift_in\[5\]
rlabel metal1 7682 16218 7682 16218 0 shift_in\[6\]
rlabel metal1 6348 6426 6348 6426 0 shift_out\[0\]
rlabel metal1 7406 6426 7406 6426 0 shift_out\[1\]
rlabel metal1 9890 6732 9890 6732 0 shift_out\[2\]
rlabel metal1 7636 7378 7636 7378 0 shift_out\[3\]
rlabel metal1 7222 8058 7222 8058 0 shift_out\[4\]
rlabel metal1 7544 9146 7544 9146 0 shift_out\[5\]
rlabel metal1 8326 9656 8326 9656 0 shift_out\[6\]
rlabel metal2 9798 7633 9798 7633 0 shift_out\[7\]
rlabel metal1 4692 17102 4692 17102 0 spi_cs_n
rlabel metal1 9982 7514 9982 7514 0 spi_miso
rlabel metal1 16882 18326 16882 18326 0 spi_mosi
rlabel metal3 1855 21148 1855 21148 0 spi_sck
rlabel metal1 9384 12206 9384 12206 0 state\[0\]
rlabel metal1 9338 13872 9338 13872 0 state\[1\]
rlabel metal2 9890 12954 9890 12954 0 state\[2\]
rlabel metal1 9798 12716 9798 12716 0 state\[3\]
rlabel metal1 16974 19788 16974 19788 0 wbs_adr_o[0]
rlabel metal1 12190 21658 12190 21658 0 wbs_adr_o[10]
rlabel metal1 8648 22746 8648 22746 0 wbs_adr_o[11]
rlabel metal1 2944 22678 2944 22678 0 wbs_adr_o[12]
rlabel metal2 2714 20383 2714 20383 0 wbs_adr_o[13]
rlabel metal2 1334 19023 1334 19023 0 wbs_adr_o[14]
rlabel metal2 2806 17085 2806 17085 0 wbs_adr_o[15]
rlabel metal1 19090 22678 19090 22678 0 wbs_adr_o[16]
rlabel metal1 19228 17306 19228 17306 0 wbs_adr_o[17]
rlabel via2 21206 20451 21206 20451 0 wbs_adr_o[18]
rlabel metal2 21160 22610 21160 22610 0 wbs_adr_o[19]
rlabel metal2 17250 16473 17250 16473 0 wbs_adr_o[1]
rlabel via1 17894 22661 17894 22661 0 wbs_adr_o[20]
rlabel metal2 20654 19363 20654 19363 0 wbs_adr_o[21]
rlabel metal2 21574 18139 21574 18139 0 wbs_adr_o[22]
rlabel metal1 21436 17306 21436 17306 0 wbs_adr_o[23]
rlabel metal1 16468 21658 16468 21658 0 wbs_adr_o[24]
rlabel metal1 17158 17306 17158 17306 0 wbs_adr_o[25]
rlabel metal1 12742 21046 12742 21046 0 wbs_adr_o[26]
rlabel metal1 11132 21658 11132 21658 0 wbs_adr_o[27]
rlabel metal2 5796 22508 5796 22508 0 wbs_adr_o[28]
rlabel metal1 5382 20536 5382 20536 0 wbs_adr_o[29]
rlabel metal2 14582 24548 14582 24548 0 wbs_adr_o[2]
rlabel metal3 1717 18428 1717 18428 0 wbs_adr_o[30]
rlabel metal3 1717 16388 1717 16388 0 wbs_adr_o[31]
rlabel metal2 9752 23052 9752 23052 0 wbs_adr_o[3]
rlabel metal1 7084 22746 7084 22746 0 wbs_adr_o[4]
rlabel metal2 7774 23307 7774 23307 0 wbs_adr_o[5]
rlabel metal2 11454 24548 11454 24548 0 wbs_adr_o[6]
rlabel metal2 5382 16915 5382 16915 0 wbs_adr_o[7]
rlabel metal2 14030 24548 14030 24548 0 wbs_adr_o[8]
rlabel metal2 13570 23307 13570 23307 0 wbs_adr_o[9]
rlabel metal2 5934 13923 5934 13923 0 wbs_cyc_o
rlabel metal1 3818 5270 3818 5270 0 wbs_dat_i[0]
rlabel metal2 5198 823 5198 823 0 wbs_dat_i[10]
rlabel metal1 6302 4114 6302 4114 0 wbs_dat_i[11]
rlabel metal3 1004 8908 1004 8908 0 wbs_dat_i[12]
rlabel metal3 1004 10268 1004 10268 0 wbs_dat_i[13]
rlabel via2 3910 9605 3910 9605 0 wbs_dat_i[14]
rlabel metal3 935 748 935 748 0 wbs_dat_i[15]
rlabel metal3 1832 2108 1832 2108 0 wbs_dat_i[16]
rlabel via2 2806 4131 2806 4131 0 wbs_dat_i[17]
rlabel metal2 9706 1231 9706 1231 0 wbs_dat_i[18]
rlabel metal2 9062 823 9062 823 0 wbs_dat_i[19]
rlabel metal2 4002 5593 4002 5593 0 wbs_dat_i[1]
rlabel metal2 3818 7633 3818 7633 0 wbs_dat_i[20]
rlabel metal2 3266 11169 3266 11169 0 wbs_dat_i[21]
rlabel metal3 3074 14348 3074 14348 0 wbs_dat_i[22]
rlabel metal3 2936 1428 2936 1428 0 wbs_dat_i[23]
rlabel metal3 1740 2788 1740 2788 0 wbs_dat_i[24]
rlabel metal2 4554 1367 4554 1367 0 wbs_dat_i[25]
rlabel metal2 8418 2098 8418 2098 0 wbs_dat_i[26]
rlabel metal1 6946 3502 6946 3502 0 wbs_dat_i[27]
rlabel metal2 2990 6443 2990 6443 0 wbs_dat_i[28]
rlabel metal3 1786 12988 1786 12988 0 wbs_dat_i[29]
rlabel metal1 7268 4454 7268 4454 0 wbs_dat_i[2]
rlabel metal2 2806 12257 2806 12257 0 wbs_dat_i[30]
rlabel metal3 912 6868 912 6868 0 wbs_dat_i[31]
rlabel metal2 7774 1707 7774 1707 0 wbs_dat_i[3]
rlabel metal3 1579 8228 1579 8228 0 wbs_dat_i[4]
rlabel metal2 4094 10251 4094 10251 0 wbs_dat_i[5]
rlabel metal3 1924 15708 1924 15708 0 wbs_dat_i[6]
rlabel metal2 5014 3740 5014 3740 0 wbs_dat_i[7]
rlabel metal2 3450 4709 3450 4709 0 wbs_dat_i[8]
rlabel metal1 4140 4114 4140 4114 0 wbs_dat_i[9]
rlabel metal1 16974 8806 16974 8806 0 wbs_dat_o[0]
rlabel metal1 17158 3570 17158 3570 0 wbs_dat_o[10]
rlabel metal1 15272 2482 15272 2482 0 wbs_dat_o[11]
rlabel metal2 17250 10931 17250 10931 0 wbs_dat_o[12]
rlabel metal2 18078 9809 18078 9809 0 wbs_dat_o[13]
rlabel metal2 21390 11475 21390 11475 0 wbs_dat_o[14]
rlabel metal2 21390 9537 21390 9537 0 wbs_dat_o[15]
rlabel metal3 18423 12852 18423 12852 0 wbs_dat_o[16]
rlabel metal1 18676 12818 18676 12818 0 wbs_dat_o[17]
rlabel metal2 21574 14229 21574 14229 0 wbs_dat_o[18]
rlabel metal2 21390 14399 21390 14399 0 wbs_dat_o[19]
rlabel metal2 14214 823 14214 823 0 wbs_dat_o[1]
rlabel via1 17986 15079 17986 15079 0 wbs_dat_o[20]
rlabel metal1 18860 14382 18860 14382 0 wbs_dat_o[21]
rlabel metal2 21390 7395 21390 7395 0 wbs_dat_o[22]
rlabel metal2 20654 8143 20654 8143 0 wbs_dat_o[23]
rlabel metal2 17066 7463 17066 7463 0 wbs_dat_o[24]
rlabel metal1 20102 5746 20102 5746 0 wbs_dat_o[25]
rlabel metal2 21390 3519 21390 3519 0 wbs_dat_o[26]
rlabel metal1 18676 2278 18676 2278 0 wbs_dat_o[27]
rlabel metal1 19734 9146 19734 9146 0 wbs_dat_o[28]
rlabel metal1 17802 4114 17802 4114 0 wbs_dat_o[29]
rlabel metal1 13110 2890 13110 2890 0 wbs_dat_o[2]
rlabel via2 21574 4811 21574 4811 0 wbs_dat_o[30]
rlabel via2 21114 6171 21114 6171 0 wbs_dat_o[31]
rlabel metal1 11132 3366 11132 3366 0 wbs_dat_o[3]
rlabel metal2 12282 1761 12282 1761 0 wbs_dat_o[4]
rlabel metal2 11822 748 11822 748 0 wbs_dat_o[5]
rlabel metal1 13616 4250 13616 4250 0 wbs_dat_o[6]
rlabel metal2 15042 748 15042 748 0 wbs_dat_o[7]
rlabel metal2 16974 748 16974 748 0 wbs_dat_o[8]
rlabel metal1 15870 4998 15870 4998 0 wbs_dat_o[9]
rlabel metal3 1717 13668 1717 13668 0 wbs_stb_o
rlabel metal1 21160 21862 21160 21862 0 wbs_we_o
<< properties >>
string FIXED_BBOX 0 0 23131 25275
<< end >>
