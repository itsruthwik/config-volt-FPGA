##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 01:36:41 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_RAM_IO
  CLASS BLOCK ;
  SIZE 100.2800 BY 30.2600 ;
  FOREIGN S_term_RAM_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.50455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.123 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.3682 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.804 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 7.8600 29.5400 8.2400 30.2600 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.11735 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.491 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.223 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 6.9400 29.5400 7.3200 30.2600 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.37195 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.967 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.8988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 6.0200 29.5400 6.4000 30.2600 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.17555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.885 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 5.1000 29.5400 5.4800 30.2600 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.046 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 29.5400 16.9800 30.2600 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.368 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 29.5400 15.6000 30.2600 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.308 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 14.3000 29.5400 14.6800 30.2600 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.34895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.5876 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.8605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 13.3800 29.5400 13.7600 30.2600 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.58 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 12.0000 29.5400 12.3800 30.2600 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.34895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.428 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 29.5400 11.4600 30.2600 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.846 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 29.5400 10.5400 30.2600 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.77655 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.443 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 11.024 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.083 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 9.2400 29.5400 9.6200 30.2600 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.407 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.4932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.51 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 29.5400 25.2600 30.2600 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.046 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 23.9600 29.5400 24.3400 30.2600 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.5800 29.5400 22.9600 30.2600 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.98175 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.155 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.51 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.4725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 21.6600 29.5400 22.0400 30.2600 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.764 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 29.5400 21.1200 30.2600 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0546 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 29.5400 19.7400 30.2600 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1684 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.292 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 18.4400 29.5400 18.8200 30.2600 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.696 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 17.5200 29.5400 17.9000 30.2600 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.30855 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.363 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.55 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 41.4400 29.5400 41.8200 30.2600 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.96 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 40.5200 29.5400 40.9000 30.2600 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75055 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.883 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.796 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 29.5400 39.9800 30.2600 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.738 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.6800 29.5400 39.0600 30.2600 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.0908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 37.3000 29.5400 37.6800 30.2600 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.3800 29.5400 36.7600 30.2600 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.512 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 29.5400 35.8400 30.2600 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.106 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 29.5400 34.4600 30.2600 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.522 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 29.5400 33.5400 30.2600 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.238 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 32.2400 29.5400 32.6200 30.2600 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.356 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.3200 29.5400 31.7000 30.2600 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.429 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.9400 29.5400 30.3200 30.2600 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 29.5400 29.4000 30.2600 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6896 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.212 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 28.1000 29.5400 28.4800 30.2600 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.7200 29.5400 27.1000 30.2600 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.52235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.476 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 25.8000 29.5400 26.1800 30.2600 ;
    END
  END N4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.0903 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.003 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 45.5800 29.5400 45.9600 30.2600 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.226 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.0638 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.8711 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 44.6600 29.5400 45.0400 30.2600 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.48648 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.9843 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 29.5400 44.1200 30.2600 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19635 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.231 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.89 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.974 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.5519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.311 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 42.8200 29.5400 43.2000 30.2600 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.2628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.866 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6425 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.7642 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 29.5400 62.9800 30.2600 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4613 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.8585 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 61.6800 29.5400 62.0600 30.2600 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.7788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 33.3248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 177.789 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 60.3000 29.5400 60.6800 30.2600 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.50195 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.767 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.9041 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.047 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 59.3800 29.5400 59.7600 30.2600 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9712 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.9972 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.9623 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 29.5400 58.8400 30.2600 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.49 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.9277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 57.5400 29.5400 57.9200 30.2600 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.4356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 35.3487 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.827 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 29.5400 56.5400 30.2600 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.608 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.1255 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.437 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 55.2400 29.5400 55.6200 30.2600 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4538 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.8208 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 54.3200 29.5400 54.7000 30.2600 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7909 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.7158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 48.028 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 253.377 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 52.9400 29.5400 53.3200 30.2600 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.666 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.7179 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.399 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 29.5400 52.4000 30.2600 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.84 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.211 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.5472 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 51.1000 29.5400 51.4800 30.2600 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4575 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.8396 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 50.1800 29.5400 50.5600 30.2600 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.9848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.628 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.4789 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.9465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 48.8000 29.5400 49.1800 30.2600 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9048 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.668 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0513 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.066 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 29.5400 48.2600 30.2600 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 41.6104 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 224.73 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 46.9600 29.5400 47.3400 30.2600 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8632 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3814 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 302.126 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 29.5400 79.5400 30.2600 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.2864 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.3545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.426 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.8085 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.5943 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 78.2400 29.5400 78.6200 30.2600 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4613 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.8585 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.3200 29.5400 77.7000 30.2600 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.49 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.31 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.3632 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 29.5400 76.7800 30.2600 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4513 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.8082 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 29.5400 75.4000 30.2600 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.25 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.8019 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 74.1000 29.5400 74.4800 30.2600 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 74.3752 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 393.447 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 73.1800 29.5400 73.5600 30.2600 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 39.4016 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 206.519 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 29.5400 72.6400 30.2600 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4992 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.26 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.6462 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 143.465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 29.5400 71.2600 30.2600 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.916 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.3428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 69.9600 29.5400 70.3400 30.2600 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.3632 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.3679 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 69.0400 29.5400 69.4200 30.2600 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.1884 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.0786 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 67.6600 29.5400 68.0400 30.2600 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.59755 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.703 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.244 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1055 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5528 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.528 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.655 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.085 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 29.5400 67.1200 30.2600 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.543 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 67.5877 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 363.645 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 65.8200 29.5400 66.2000 30.2600 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.1871 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.4874 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 64.9000 29.5400 65.2800 30.2600 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.856 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 30.5733 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 148.418 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 63.5200 29.5400 63.9000 30.2600 ;
    END
  END S4END[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.431 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.86 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0184 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.055 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 26.0991 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 127.044 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.6088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.8915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.568 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.19 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.3557 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.3302 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2592 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.2185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.1481 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.2925 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.2864 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.3545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.0601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.8522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.3738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 46.4003 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 243.223 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.3614 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.77 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 28.2563 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 137.83 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1016 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.296 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.5955 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.624 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.884 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.63994 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.0094 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2202 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.612 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.3776 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.8105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8299 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.4906 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.2248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 67.062 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 339.283 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.34 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.7594 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7195 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4802 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.9528 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5552 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.304 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.9154 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.903 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.151 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 6.25629 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 34.7767 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.2084 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.606 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 34.8601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 166.827 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.13265 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.509 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4556 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.241 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 22.5594 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 109.346 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.7945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.856 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8953 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.4528 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 41.4664 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 209.931 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.1425 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.5849 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.522 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.5846 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.5377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.7167 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.456 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.322 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5355 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.5503 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.541 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.82987 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.4465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.424 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.8711 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 46.4443 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.811 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.019 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 47.938 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 252.494 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 34.9022 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 181.39 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.718 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 43.6645 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.855 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9648 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.48 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.78333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.0472 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 25.6921 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 129.78 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3272 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.41 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1619 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.6824 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6394 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.971 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8311 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.0283 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.632 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7494 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.044 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.31 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 28.6600 100.2800 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1255 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 26.6200 100.2800 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.852 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 24.9200 100.2800 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 22.8800 100.2800 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.263 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.83 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.7398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 21.1800 100.2800 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.9298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.096 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 19.1400 100.2800 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6815 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 17.4400 100.2800 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 15.7400 100.2800 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 13.7000 100.2800 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 12.0000 100.2800 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.235 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 10.3000 100.2800 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 8.2600 100.2800 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.914 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.9888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.744 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 6.5600 100.2800 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 4.5200 100.2800 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.3286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.36 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 2.8200 100.2800 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.78 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 1.1200 100.2800 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.402 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.142 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 27.6250 100.2800 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 25.9250 100.2800 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.0896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.3705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 24.2250 100.2800 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.472 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 22.5250 100.2800 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.488 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 20.8250 100.2800 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 19.1250 100.2800 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.337 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2824 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.375 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 17.4250 100.2800 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6026 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9355 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 15.7250 100.2800 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1902 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.8365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 14.0250 100.2800 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8874 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.044 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.3944 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.935 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 12.3250 100.2800 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 10.6250 100.2800 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.751 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 8.9250 100.2800 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.6744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 58.2575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.024 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 7.2250 100.2800 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.431 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.86 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.4928 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.427 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 5.5250 100.2800 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0719 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.282 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 3.8250 100.2800 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5406 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.636 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.3844 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.8445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.379 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 2.1250 100.2800 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 21.6355 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.522 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 97.5600 0.0000 97.9400 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.143 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.8676 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.2107 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 96.6400 0.0000 97.0200 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.381 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.1101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 95.7200 0.0000 96.1000 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.54 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.474 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.206 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.9025 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.8000 0.0000 95.1800 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.859 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.3396 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 93.8800 0.0000 94.2600 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.511 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 78.8814 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 389.28 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.9600 0.0000 93.3400 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.8522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.0400 0.0000 92.4200 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.176 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.723 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.9119 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.1200 0.0000 91.5000 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0642 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.213 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5079 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.1541 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.2000 0.0000 90.5800 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.451 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.5884 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.557 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 89.2800 0.0000 89.6600 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.193 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.4173 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.217 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 88.3600 0.0000 88.7400 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.1104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 110.425 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 87.4400 0.0000 87.8200 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.0418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 106.112 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 579.931 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.5200 0.0000 86.9000 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.511 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 33.1494 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 161.362 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 85.6000 0.0000 85.9800 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 42.9047 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.711 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 84.6800 0.0000 85.0600 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.8774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 83.7600 0.0000 84.1400 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.469 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.5632 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.947 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 82.3800 0.0000 82.7600 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 97.5600 29.5400 97.9400 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.1786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 96.6400 29.5400 97.0200 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 95.7200 29.5400 96.1000 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.642 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.8000 29.5400 95.1800 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 93.8800 29.5400 94.2600 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.041 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.9600 29.5400 93.3400 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.0400 29.5400 92.4200 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.665 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.1200 29.5400 91.5000 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.747 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.2000 29.5400 90.5800 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.879 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.2800 29.5400 89.6600 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.844 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.3600 29.5400 88.7400 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.416 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 87.4400 29.5400 87.8200 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.081 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.5200 29.5400 86.9000 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 85.6000 29.5400 85.9800 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.1014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 84.6800 29.5400 85.0600 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 83.7600 29.5400 84.1400 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 82.3800 29.5400 82.7600 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 94.7200 6.0700 ;
        RECT 5.5600 23.0000 94.7200 25.0000 ;
        RECT 92.7200 15.0600 94.7200 15.5400 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 92.7200 9.6200 94.7200 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 92.7200 20.5000 94.7200 20.9800 ;
      LAYER met4 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
        RECT 92.7200 4.0700 94.7200 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 97.7200 3.0700 ;
        RECT 2.5600 26.0000 97.7200 28.0000 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 95.7200 12.3400 97.7200 12.8200 ;
        RECT 95.7200 6.9000 97.7200 7.3800 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 95.7200 17.7800 97.7200 18.2600 ;
      LAYER met4 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
        RECT 95.7200 1.0700 97.7200 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 79.7100 29.3700 100.2800 30.2600 ;
      RECT 78.7900 29.3700 78.9900 30.2600 ;
      RECT 77.8700 29.3700 78.0700 30.2600 ;
      RECT 76.9500 29.3700 77.1500 30.2600 ;
      RECT 75.5700 29.3700 76.2300 30.2600 ;
      RECT 74.6500 29.3700 74.8500 30.2600 ;
      RECT 73.7300 29.3700 73.9300 30.2600 ;
      RECT 72.8100 29.3700 73.0100 30.2600 ;
      RECT 71.4300 29.3700 72.0900 30.2600 ;
      RECT 70.5100 29.3700 70.7100 30.2600 ;
      RECT 69.5900 29.3700 69.7900 30.2600 ;
      RECT 68.2100 29.3700 68.8700 30.2600 ;
      RECT 67.2900 29.3700 67.4900 30.2600 ;
      RECT 66.3700 29.3700 66.5700 30.2600 ;
      RECT 65.4500 29.3700 65.6500 30.2600 ;
      RECT 64.0700 29.3700 64.7300 30.2600 ;
      RECT 63.1500 29.3700 63.3500 30.2600 ;
      RECT 62.2300 29.3700 62.4300 30.2600 ;
      RECT 60.8500 29.3700 61.5100 30.2600 ;
      RECT 59.9300 29.3700 60.1300 30.2600 ;
      RECT 59.0100 29.3700 59.2100 30.2600 ;
      RECT 58.0900 29.3700 58.2900 30.2600 ;
      RECT 56.7100 29.3700 57.3700 30.2600 ;
      RECT 55.7900 29.3700 55.9900 30.2600 ;
      RECT 54.8700 29.3700 55.0700 30.2600 ;
      RECT 53.4900 29.3700 54.1500 30.2600 ;
      RECT 52.5700 29.3700 52.7700 30.2600 ;
      RECT 51.6500 29.3700 51.8500 30.2600 ;
      RECT 50.7300 29.3700 50.9300 30.2600 ;
      RECT 49.3500 29.3700 50.0100 30.2600 ;
      RECT 48.4300 29.3700 48.6300 30.2600 ;
      RECT 47.5100 29.3700 47.7100 30.2600 ;
      RECT 46.1300 29.3700 46.7900 30.2600 ;
      RECT 45.2100 29.3700 45.4100 30.2600 ;
      RECT 44.2900 29.3700 44.4900 30.2600 ;
      RECT 43.3700 29.3700 43.5700 30.2600 ;
      RECT 41.9900 29.3700 42.6500 30.2600 ;
      RECT 41.0700 29.3700 41.2700 30.2600 ;
      RECT 40.1500 29.3700 40.3500 30.2600 ;
      RECT 39.2300 29.3700 39.4300 30.2600 ;
      RECT 37.8500 29.3700 38.5100 30.2600 ;
      RECT 36.9300 29.3700 37.1300 30.2600 ;
      RECT 36.0100 29.3700 36.2100 30.2600 ;
      RECT 34.6300 29.3700 35.2900 30.2600 ;
      RECT 33.7100 29.3700 33.9100 30.2600 ;
      RECT 32.7900 29.3700 32.9900 30.2600 ;
      RECT 31.8700 29.3700 32.0700 30.2600 ;
      RECT 30.4900 29.3700 31.1500 30.2600 ;
      RECT 29.5700 29.3700 29.7700 30.2600 ;
      RECT 28.6500 29.3700 28.8500 30.2600 ;
      RECT 27.2700 29.3700 27.9300 30.2600 ;
      RECT 26.3500 29.3700 26.5500 30.2600 ;
      RECT 25.4300 29.3700 25.6300 30.2600 ;
      RECT 24.5100 29.3700 24.7100 30.2600 ;
      RECT 23.1300 29.3700 23.7900 30.2600 ;
      RECT 22.2100 29.3700 22.4100 30.2600 ;
      RECT 21.2900 29.3700 21.4900 30.2600 ;
      RECT 19.9100 29.3700 20.5700 30.2600 ;
      RECT 18.9900 29.3700 19.1900 30.2600 ;
      RECT 18.0700 29.3700 18.2700 30.2600 ;
      RECT 17.1500 29.3700 17.3500 30.2600 ;
      RECT 15.7700 29.3700 16.4300 30.2600 ;
      RECT 14.8500 29.3700 15.0500 30.2600 ;
      RECT 13.9300 29.3700 14.1300 30.2600 ;
      RECT 12.5500 29.3700 13.2100 30.2600 ;
      RECT 11.6300 29.3700 11.8300 30.2600 ;
      RECT 10.7100 29.3700 10.9100 30.2600 ;
      RECT 9.7900 29.3700 9.9900 30.2600 ;
      RECT 8.4100 29.3700 9.0700 30.2600 ;
      RECT 7.4900 29.3700 7.6900 30.2600 ;
      RECT 6.5700 29.3700 6.7700 30.2600 ;
      RECT 5.6500 29.3700 5.8500 30.2600 ;
      RECT 0.0000 29.3700 4.9300 30.2600 ;
      RECT 0.0000 28.9850 100.2800 29.3700 ;
      RECT 0.5000 28.4750 100.2800 28.9850 ;
      RECT 0.0000 27.9650 100.2800 28.4750 ;
      RECT 0.0000 27.4550 99.7800 27.9650 ;
      RECT 0.0000 26.9450 100.2800 27.4550 ;
      RECT 0.5000 26.4350 100.2800 26.9450 ;
      RECT 0.0000 26.2650 100.2800 26.4350 ;
      RECT 0.0000 25.7550 99.7800 26.2650 ;
      RECT 0.0000 25.2450 100.2800 25.7550 ;
      RECT 0.5000 24.7350 100.2800 25.2450 ;
      RECT 0.0000 24.5650 100.2800 24.7350 ;
      RECT 0.0000 24.0550 99.7800 24.5650 ;
      RECT 0.0000 23.2050 100.2800 24.0550 ;
      RECT 0.5000 22.8650 100.2800 23.2050 ;
      RECT 0.5000 22.6950 99.7800 22.8650 ;
      RECT 0.0000 22.3550 99.7800 22.6950 ;
      RECT 0.0000 21.5050 100.2800 22.3550 ;
      RECT 0.5000 21.1650 100.2800 21.5050 ;
      RECT 0.5000 20.9950 99.7800 21.1650 ;
      RECT 0.0000 20.6550 99.7800 20.9950 ;
      RECT 0.0000 19.4650 100.2800 20.6550 ;
      RECT 0.5000 18.9550 99.7800 19.4650 ;
      RECT 0.0000 17.7650 100.2800 18.9550 ;
      RECT 0.5000 17.2550 99.7800 17.7650 ;
      RECT 0.0000 16.0650 100.2800 17.2550 ;
      RECT 0.5000 15.5550 99.7800 16.0650 ;
      RECT 0.0000 14.3650 100.2800 15.5550 ;
      RECT 0.0000 14.0250 99.7800 14.3650 ;
      RECT 0.5000 13.8550 99.7800 14.0250 ;
      RECT 0.5000 13.5150 100.2800 13.8550 ;
      RECT 0.0000 12.6650 100.2800 13.5150 ;
      RECT 0.0000 12.3250 99.7800 12.6650 ;
      RECT 0.5000 12.1550 99.7800 12.3250 ;
      RECT 0.5000 11.8150 100.2800 12.1550 ;
      RECT 0.0000 10.9650 100.2800 11.8150 ;
      RECT 0.0000 10.6250 99.7800 10.9650 ;
      RECT 0.5000 10.4550 99.7800 10.6250 ;
      RECT 0.5000 10.1150 100.2800 10.4550 ;
      RECT 0.0000 9.2650 100.2800 10.1150 ;
      RECT 0.0000 8.7550 99.7800 9.2650 ;
      RECT 0.0000 8.5850 100.2800 8.7550 ;
      RECT 0.5000 8.0750 100.2800 8.5850 ;
      RECT 0.0000 7.5650 100.2800 8.0750 ;
      RECT 0.0000 7.0550 99.7800 7.5650 ;
      RECT 0.0000 6.8850 100.2800 7.0550 ;
      RECT 0.5000 6.3750 100.2800 6.8850 ;
      RECT 0.0000 5.8650 100.2800 6.3750 ;
      RECT 0.0000 5.3550 99.7800 5.8650 ;
      RECT 0.0000 4.8450 100.2800 5.3550 ;
      RECT 0.5000 4.3350 100.2800 4.8450 ;
      RECT 0.0000 4.1650 100.2800 4.3350 ;
      RECT 0.0000 3.6550 99.7800 4.1650 ;
      RECT 0.0000 3.1450 100.2800 3.6550 ;
      RECT 0.5000 2.6350 100.2800 3.1450 ;
      RECT 0.0000 2.4650 100.2800 2.6350 ;
      RECT 0.0000 1.9550 99.7800 2.4650 ;
      RECT 0.0000 1.4450 100.2800 1.9550 ;
      RECT 0.5000 0.9350 100.2800 1.4450 ;
      RECT 0.0000 0.0000 100.2800 0.9350 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 100.2800 30.2600 ;
    LAYER met2 ;
      RECT 98.0800 29.4000 100.2800 30.2600 ;
      RECT 97.1600 29.4000 97.4200 30.2600 ;
      RECT 96.2400 29.4000 96.5000 30.2600 ;
      RECT 95.3200 29.4000 95.5800 30.2600 ;
      RECT 94.4000 29.4000 94.6600 30.2600 ;
      RECT 93.4800 29.4000 93.7400 30.2600 ;
      RECT 92.5600 29.4000 92.8200 30.2600 ;
      RECT 91.6400 29.4000 91.9000 30.2600 ;
      RECT 90.7200 29.4000 90.9800 30.2600 ;
      RECT 89.8000 29.4000 90.0600 30.2600 ;
      RECT 88.8800 29.4000 89.1400 30.2600 ;
      RECT 87.9600 29.4000 88.2200 30.2600 ;
      RECT 87.0400 29.4000 87.3000 30.2600 ;
      RECT 86.1200 29.4000 86.3800 30.2600 ;
      RECT 85.2000 29.4000 85.4600 30.2600 ;
      RECT 84.2800 29.4000 84.5400 30.2600 ;
      RECT 82.9000 29.4000 83.6200 30.2600 ;
      RECT 0.0000 29.4000 82.2400 30.2600 ;
      RECT 0.0000 28.9400 100.2800 29.4000 ;
      RECT 0.0000 28.5200 99.6550 28.9400 ;
      RECT 0.0000 27.9200 100.2800 28.5200 ;
      RECT 0.6250 27.5000 100.2800 27.9200 ;
      RECT 0.0000 26.9000 100.2800 27.5000 ;
      RECT 0.0000 26.4800 99.6550 26.9000 ;
      RECT 0.0000 26.2200 100.2800 26.4800 ;
      RECT 0.6250 25.8000 100.2800 26.2200 ;
      RECT 0.0000 25.2000 100.2800 25.8000 ;
      RECT 0.0000 24.7800 99.6550 25.2000 ;
      RECT 0.0000 24.5200 100.2800 24.7800 ;
      RECT 0.6250 24.1000 100.2800 24.5200 ;
      RECT 0.0000 23.1600 100.2800 24.1000 ;
      RECT 0.0000 22.8200 99.6550 23.1600 ;
      RECT 0.6250 22.7400 99.6550 22.8200 ;
      RECT 0.6250 22.4000 100.2800 22.7400 ;
      RECT 0.0000 21.4600 100.2800 22.4000 ;
      RECT 0.0000 21.1200 99.6550 21.4600 ;
      RECT 0.6250 21.0400 99.6550 21.1200 ;
      RECT 0.6250 20.7000 100.2800 21.0400 ;
      RECT 0.0000 19.4200 100.2800 20.7000 ;
      RECT 0.6250 19.0000 99.6550 19.4200 ;
      RECT 0.0000 17.7200 100.2800 19.0000 ;
      RECT 0.6250 17.3000 99.6550 17.7200 ;
      RECT 0.0000 16.0200 100.2800 17.3000 ;
      RECT 0.6250 15.6000 99.6550 16.0200 ;
      RECT 0.0000 14.3200 100.2800 15.6000 ;
      RECT 0.6250 13.9800 100.2800 14.3200 ;
      RECT 0.6250 13.9000 99.6550 13.9800 ;
      RECT 0.0000 13.5600 99.6550 13.9000 ;
      RECT 0.0000 12.6200 100.2800 13.5600 ;
      RECT 0.6250 12.2800 100.2800 12.6200 ;
      RECT 0.6250 12.2000 99.6550 12.2800 ;
      RECT 0.0000 11.8600 99.6550 12.2000 ;
      RECT 0.0000 10.9200 100.2800 11.8600 ;
      RECT 0.6250 10.5800 100.2800 10.9200 ;
      RECT 0.6250 10.5000 99.6550 10.5800 ;
      RECT 0.0000 10.1600 99.6550 10.5000 ;
      RECT 0.0000 9.2200 100.2800 10.1600 ;
      RECT 0.6250 8.8000 100.2800 9.2200 ;
      RECT 0.0000 8.5400 100.2800 8.8000 ;
      RECT 0.0000 8.1200 99.6550 8.5400 ;
      RECT 0.0000 7.5200 100.2800 8.1200 ;
      RECT 0.6250 7.1000 100.2800 7.5200 ;
      RECT 0.0000 6.8400 100.2800 7.1000 ;
      RECT 0.0000 6.4200 99.6550 6.8400 ;
      RECT 0.0000 5.8200 100.2800 6.4200 ;
      RECT 0.6250 5.4000 100.2800 5.8200 ;
      RECT 0.0000 4.8000 100.2800 5.4000 ;
      RECT 0.0000 4.3800 99.6550 4.8000 ;
      RECT 0.0000 4.1200 100.2800 4.3800 ;
      RECT 0.6250 3.7000 100.2800 4.1200 ;
      RECT 0.0000 3.1000 100.2800 3.7000 ;
      RECT 0.0000 2.6800 99.6550 3.1000 ;
      RECT 0.0000 2.4200 100.2800 2.6800 ;
      RECT 0.6250 2.0000 100.2800 2.4200 ;
      RECT 0.0000 1.4000 100.2800 2.0000 ;
      RECT 0.0000 0.9800 99.6550 1.4000 ;
      RECT 0.0000 0.8600 100.2800 0.9800 ;
      RECT 98.0800 0.0000 100.2800 0.8600 ;
      RECT 97.1600 0.0000 97.4200 0.8600 ;
      RECT 96.2400 0.0000 96.5000 0.8600 ;
      RECT 95.3200 0.0000 95.5800 0.8600 ;
      RECT 94.4000 0.0000 94.6600 0.8600 ;
      RECT 93.4800 0.0000 93.7400 0.8600 ;
      RECT 92.5600 0.0000 92.8200 0.8600 ;
      RECT 91.6400 0.0000 91.9000 0.8600 ;
      RECT 90.7200 0.0000 90.9800 0.8600 ;
      RECT 89.8000 0.0000 90.0600 0.8600 ;
      RECT 88.8800 0.0000 89.1400 0.8600 ;
      RECT 87.9600 0.0000 88.2200 0.8600 ;
      RECT 87.0400 0.0000 87.3000 0.8600 ;
      RECT 86.1200 0.0000 86.3800 0.8600 ;
      RECT 85.2000 0.0000 85.4600 0.8600 ;
      RECT 84.2800 0.0000 84.5400 0.8600 ;
      RECT 82.9000 0.0000 83.6200 0.8600 ;
      RECT 0.0000 0.0000 82.2400 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 100.2800 30.2600 ;
      RECT 98.0200 25.7000 100.2800 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 100.2800 25.7000 ;
      RECT 95.0200 22.7000 100.2800 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 100.2800 22.7000 ;
      RECT 95.0200 20.2000 100.2800 21.2800 ;
      RECT 7.8600 20.2000 92.4200 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 100.2800 20.2000 ;
      RECT 98.0200 17.4800 100.2800 18.5600 ;
      RECT 4.8600 17.4800 95.4200 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 100.2800 17.4800 ;
      RECT 95.0200 14.7600 100.2800 15.8400 ;
      RECT 7.8600 14.7600 92.4200 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 100.2800 14.7600 ;
      RECT 98.0200 12.0400 100.2800 13.1200 ;
      RECT 4.8600 12.0400 95.4200 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 100.2800 12.0400 ;
      RECT 95.0200 9.3200 100.2800 10.4000 ;
      RECT 7.8600 9.3200 92.4200 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 100.2800 9.3200 ;
      RECT 98.0200 6.6000 100.2800 7.6800 ;
      RECT 4.8600 6.6000 95.4200 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 100.2800 6.6000 ;
      RECT 95.0200 3.7700 100.2800 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 100.2800 3.7700 ;
      RECT 98.0200 0.7700 100.2800 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 100.2800 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 100.2800 30.2600 ;
      RECT 4.8600 25.3000 95.4200 28.3000 ;
      RECT 95.0200 3.7700 95.4200 25.3000 ;
      RECT 7.8600 3.7700 92.4200 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 98.0200 0.7700 100.2800 28.3000 ;
      RECT 4.8600 0.7700 95.4200 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 100.2800 0.7700 ;
  END
END S_term_RAM_IO

END LIBRARY
