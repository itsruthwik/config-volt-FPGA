##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 01:31:30 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_single2
  CLASS BLOCK ;
  SIZE 240.1200 BY 30.2600 ;
  FOREIGN S_term_single2 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 29.5400 14.2200 30.2600 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8428 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.28 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.1856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.264 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 29.5400 12.8400 30.2600 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.322 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 29.5400 11.4600 30.2600 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.0884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.3645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 29.5400 10.5400 30.2600 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 29.5400 25.2600 30.2600 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.8656 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.63 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 29.5400 23.8800 30.2600 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.0208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 100.027 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.796 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 29.5400 22.5000 30.2600 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 29.5400 21.1200 30.2600 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.4648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.616 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 29.5400 19.7400 30.2600 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21295 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.427 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.12 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.5225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.086 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 29.5400 18.3600 30.2600 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.415 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.7398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 29.5400 16.9800 30.2600 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.576 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.644 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 29.5400 15.6000 30.2600 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.144 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 29.5400 35.8400 30.2600 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.002 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 29.5400 34.4600 30.2600 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.223 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 29.5400 33.5400 30.2600 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.3978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.208 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 29.5400 32.1600 30.2600 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.51 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 29.5400 30.7800 30.2600 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.611 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.6552 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 83.1985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.476 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 29.5400 29.4000 30.2600 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.725 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.032 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 29.5400 28.0200 30.2600 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.5944 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 72.8945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.262 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 29.5400 26.6400 30.2600 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1656 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.592 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 29.5400 57.4600 30.2600 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.6584 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 78.2145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 29.5400 56.5400 30.2600 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 29.5400 55.1600 30.2600 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 29.5400 53.7800 30.2600 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.997 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.472 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 29.5400 52.4000 30.2600 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4656 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.092 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 29.5400 51.0200 30.2600 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8272 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.1248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.136 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 29.5400 49.6400 30.2600 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.162 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 29.5400 48.2600 30.2600 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.939 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 29.5400 46.8800 30.2600 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.968 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 29.5400 45.5000 30.2600 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9627 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.5048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.496 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 29.5400 44.1200 30.2600 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.216 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 29.5400 42.7400 30.2600 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.596 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 29.5400 41.3600 30.2600 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.5272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.77 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 29.5400 39.9800 30.2600 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.8492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.084 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 29.5400 38.6000 30.2600 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.0678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.832 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 29.5400 37.2200 30.2600 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 29.5400 79.5400 30.2600 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 29.5400 78.1600 30.2600 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.7216 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 63.4935 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.416 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 29.5400 76.7800 30.2600 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 29.5400 75.4000 30.2600 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 29.5400 74.0200 30.2600 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.877 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 29.5400 72.6400 30.2600 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.64 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 29.5400 71.2600 30.2600 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.7004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3135 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 29.5400 69.8800 30.2600 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.6788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.424 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 29.5400 68.5000 30.2600 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 29.5400 67.1200 30.2600 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.726 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 29.5400 65.7400 30.2600 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.7636 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 58.7405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 29.5400 64.3600 30.2600 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.2744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.466 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 29.5400 62.9800 30.2600 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6822 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.293 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 29.5400 61.6000 30.2600 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.941 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 29.5400 60.2200 30.2600 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.63495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.747 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.5668 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 67.7565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.342 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 29.5400 58.8400 30.2600 ;
    END
  END NN4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.1176 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.4735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.512 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.1657 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.3805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 29.5400 84.6000 30.2600 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7921 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.217 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 29.5400 83.2200 30.2600 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8076 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.684 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 44.7204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 217.67 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 29.5400 81.8400 30.2600 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4108 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 30.4563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 146.349 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 29.5400 80.4600 30.2600 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7134 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.449 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.1255 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.6038 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 29.5400 106.2200 30.2600 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.407 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.043 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.9758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.431 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 29.5400 104.8400 30.2600 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1469 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.3805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 29.5400 103.4600 30.2600 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8374 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.951 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4814 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.217 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 29.5400 102.5400 30.2600 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.367 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.0252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 29.5400 101.1600 30.2600 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6082 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 31.2921 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 170.786 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 29.5400 99.7800 30.2600 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.988 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.4085 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 116.789 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 29.5400 98.4000 30.2600 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.03955 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.223 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.172 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.767 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.1604 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 29.5400 97.0200 30.2600 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.4452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.1485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.224 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.3896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.9245 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 29.5400 95.6400 30.2600 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1258 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.393 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.7192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.991 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 29.5400 94.2600 30.2600 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.568 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5374 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.451 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.3682 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.651 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 29.5400 92.8800 30.2600 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.486 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8701 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.8774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 29.5400 91.5000 30.2600 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.3128 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.4865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.608 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.80975 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.0252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 29.5400 90.1200 30.2600 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9792 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.849 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.082 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.174 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 30.0085 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 144.852 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 29.5400 88.7400 30.2600 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.7044 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4075 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.486 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2437 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.7704 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 29.5400 87.3600 30.2600 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.952 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.2563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.418 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 29.5400 85.9800 30.2600 ;
    END
  END S2END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.9695 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.3994 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 29.5400 149.4600 30.2600 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.009 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.3129 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 141.374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 29.5400 148.5400 30.2600 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 22.3412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.667 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 29.5400 147.1600 30.2600 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3695 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.3994 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 29.5400 145.7800 30.2600 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.86132 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.8585 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 29.5400 144.4000 30.2600 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.016 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.607 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 29.5400 143.0200 30.2600 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 56.2393 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 299.698 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 29.5400 141.6400 30.2600 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.618 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 29.5400 140.2600 30.2600 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.074 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.84497 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.2296 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 29.5400 138.8800 30.2600 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.046 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.055 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.802 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 29.5400 137.5000 30.2600 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.3154 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.8396 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 29.5400 136.1200 30.2600 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1284 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.5275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.5 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 29.5400 134.7400 30.2600 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.605 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.2356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 42.467 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 225.918 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 29.5400 133.3600 30.2600 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.42415 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.499 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.856 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.474 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.3645 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.3742 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 29.5400 131.9800 30.2600 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.468 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.6478 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 29.5400 130.6000 30.2600 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 104.339 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 551.267 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 29.5400 129.2200 30.2600 ;
    END
  END SS4END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.77945 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.917 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.33 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.1242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.8553 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 29.5400 127.8400 30.2600 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.834 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.5632 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.05 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 29.5400 126.4600 30.2600 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.95035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6475 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.5028 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.3333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 29.5400 125.5400 30.2600 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.17175 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.555 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3278 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.403 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.3204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.9969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 29.5400 124.1600 30.2600 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.87395 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.087 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6056 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.62 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.6349 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.9591 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 29.5400 122.7800 30.2600 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21635 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.431 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.452 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.7619 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.2044 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 29.5400 121.4000 30.2600 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.12115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.319 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.486 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.6487 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.7956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 29.5400 120.0200 30.2600 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.69 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2022 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.9874 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 29.5400 118.6400 30.2600 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.571 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.972 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.6698 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 29.5400 117.2600 30.2600 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.615 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.584 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.5406 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.5126 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 29.5400 115.8800 30.2600 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.69275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.815 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.5472 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.916 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.3428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 29.5400 114.5000 30.2600 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.322 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.0336 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.953 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 29.5400 113.1200 30.2600 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.628 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.4865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 113.079 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 29.5400 111.7400 30.2600 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 30.3827 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 164.579 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 29.5400 110.3600 30.2600 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.9168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 79.3211 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 414.83 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 29.5400 108.9800 30.2600 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.53975 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.635 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.6252 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.0485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.094 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.1947 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.9497 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 29.5400 107.6000 30.2600 ;
    END
  END S4END[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.411 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.66 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 21.5496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 107.671 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.202 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.29906 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.4717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.84 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.2948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 63.2657 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 323.252 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 61.306 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 79.1884 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 387.843 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.7228 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 78.5365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.29 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.1824 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.853 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.18 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.5752 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 72.7615 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.3428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3448 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8833 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0832 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 36.784 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.981 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.66 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 63.1855 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.966 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.07893 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.9465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4056 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.142 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5827 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 191.528 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.0502 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.1735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.93 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3632 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.0503 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.8728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.379 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.3484 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 103.214 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 550.179 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.089 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.9722 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.7835 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.862 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.3028 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.582 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.296 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.4025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.13975 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.3654 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 81.8129 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 435.201 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.8184 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.0145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.69 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.3506 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.9874 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.3068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0992 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.26 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.7607 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.9739 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 69.755 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.704 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.59088 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.5063 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8692 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.2685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.15 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 40.7739 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.972 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.178 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 59.4437 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 286.286 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.303 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9292 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.9748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.1448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 86.8934 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 448.755 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.683 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.08019 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.2736 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.75 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 29.4632 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.292 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.17138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.1541 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 43.0921 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 215.006 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7921 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.0912 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.141 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.8522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9273 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5406 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 32.1538 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 172.956 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.298 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.146 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.51289 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.1195 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.2028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.4316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 51.8582 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 275.921 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.8525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.1352 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8195 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.53616 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.8113 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.712 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6462 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.0786 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.791 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.653 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.542 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 51.2053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.481 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1896 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.787 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.0248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.936 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 28.6600 240.1200 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.483 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 26.6200 240.1200 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.3118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 188.8 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 24.9200 240.1200 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.168 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 22.8800 240.1200 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9955 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 21.1800 240.1200 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 19.1400 240.1200 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.727 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 17.4400 240.1200 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.25 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.906 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 15.7400 240.1200 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.352 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 13.7000 240.1200 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.187 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.4728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.992 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 12.0000 240.1200 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 10.3000 240.1200 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.9938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.104 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 8.2600 240.1200 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.85 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.157 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 6.5600 240.1200 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.5838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.584 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 4.5200 240.1200 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.712 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5452 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 2.8200 240.1200 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7988 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.65 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 1.1200 240.1200 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.0892 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.3685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 27.6250 240.1200 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.018 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.0125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 25.9250 240.1200 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.992 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.52 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 11.3768 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.847 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 24.2250 240.1200 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.824 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 22.5250 240.1200 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.066 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.2525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.856 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 20.8250 240.1200 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.2964 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.4045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.572 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 19.1250 240.1200 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.089 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.836 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 17.4250 240.1200 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.5752 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 72.7615 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.238 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 15.7250 240.1200 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.0592 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.2185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 14.0250 240.1200 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.9436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.6405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 12.3250 240.1200 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.5236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.5405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.576 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 10.6250 240.1200 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 17.8812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.369 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 8.9250 240.1200 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.4652 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.2485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.705 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 7.2250 240.1200 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8704 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.024 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.7708 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.7765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.024 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 5.5250 240.1200 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.24905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.293 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.1908 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 75.8765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.748 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.622 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 3.8250 240.1200 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.116 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.5025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 2.1250 240.1200 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6035 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.8899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 179.4400 0.0000 179.8200 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.227 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.4689 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.802 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 173.9200 0.0000 174.3000 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 35.8412 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 173.336 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 168.8600 0.0000 169.2400 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.917 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5921 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.2579 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 163.3400 0.0000 163.7200 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.9947 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.104 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 158.2800 0.0000 158.6600 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.845 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.6824 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 153.2200 0.0000 153.6000 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.953 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1443 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.3113 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 147.2400 0.0000 147.6200 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.251 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.911 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.1909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.085 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 142.1800 0.0000 142.5600 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.4525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.075 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 137.5800 0.0000 137.9600 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9754 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.651 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.6186 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.9654 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 132.0600 0.0000 132.4400 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.779 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.8311 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.028 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 127.0000 0.0000 127.3800 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.4626 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.77 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 121.4800 0.0000 121.8600 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.861 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5217 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.9057 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 116.4200 0.0000 116.8000 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.217 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.0047 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.349 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 111.3600 0.0000 111.7400 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.929 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.4651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 102.94 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 105.8400 0.0000 106.2200 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.491 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5846 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.0535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 100.7800 0.0000 101.1600 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.047 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7544 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.9717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 95.2600 0.0000 95.6400 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.1481 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.6226 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.2000 0.0000 90.5800 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.047 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.8437 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.0283 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 85.1400 0.0000 85.5200 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.8676 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.2107 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 80.0800 0.0000 80.4600 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.073 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.8000 29.5400 210.1800 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.333 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 206.5800 29.5400 206.9600 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.561 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 203.8200 29.5400 204.2000 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.3438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.304 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 201.0600 29.5400 201.4400 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.887 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 198.3000 29.5400 198.6800 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 195.0800 29.5400 195.4600 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.3200 29.5400 192.7000 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.085 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 189.5600 29.5400 189.9400 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5854 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 186.8000 29.5400 187.1800 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.071 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 184.0400 29.5400 184.4200 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.8200 29.5400 181.2000 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.286 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 178.0600 29.5400 178.4400 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.652 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 175.3000 29.5400 175.6800 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 172.5400 29.5400 172.9200 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.83 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 169.7800 29.5400 170.1600 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9306 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.427 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.5600 29.5400 166.9400 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.241 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 163.8000 29.5400 164.1800 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.069 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.0400 29.5400 161.4200 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 158.2800 29.5400 158.6600 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.44 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.5200 29.5400 155.9000 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 234.5600 6.0700 ;
        RECT 5.5600 23.0000 234.5600 25.0000 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 232.5600 15.0600 234.5600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 232.5600 9.6200 234.5600 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 232.5600 20.5000 234.5600 20.9800 ;
      LAYER met4 ;
        RECT 232.5600 4.0700 234.5600 25.0000 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 237.5600 3.0700 ;
        RECT 2.5600 26.0000 237.5600 28.0000 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 235.5600 6.9000 237.5600 7.3800 ;
        RECT 235.5600 12.3400 237.5600 12.8200 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 235.5600 17.7800 237.5600 18.2600 ;
      LAYER met4 ;
        RECT 235.5600 1.0700 237.5600 28.0000 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.6300 29.3700 240.1200 30.2600 ;
      RECT 148.7100 29.3700 148.9100 30.2600 ;
      RECT 147.3300 29.3700 147.9900 30.2600 ;
      RECT 145.9500 29.3700 146.6100 30.2600 ;
      RECT 144.5700 29.3700 145.2300 30.2600 ;
      RECT 143.1900 29.3700 143.8500 30.2600 ;
      RECT 141.8100 29.3700 142.4700 30.2600 ;
      RECT 140.4300 29.3700 141.0900 30.2600 ;
      RECT 139.0500 29.3700 139.7100 30.2600 ;
      RECT 137.6700 29.3700 138.3300 30.2600 ;
      RECT 136.2900 29.3700 136.9500 30.2600 ;
      RECT 134.9100 29.3700 135.5700 30.2600 ;
      RECT 133.5300 29.3700 134.1900 30.2600 ;
      RECT 132.1500 29.3700 132.8100 30.2600 ;
      RECT 130.7700 29.3700 131.4300 30.2600 ;
      RECT 129.3900 29.3700 130.0500 30.2600 ;
      RECT 128.0100 29.3700 128.6700 30.2600 ;
      RECT 126.6300 29.3700 127.2900 30.2600 ;
      RECT 125.7100 29.3700 125.9100 30.2600 ;
      RECT 124.3300 29.3700 124.9900 30.2600 ;
      RECT 122.9500 29.3700 123.6100 30.2600 ;
      RECT 121.5700 29.3700 122.2300 30.2600 ;
      RECT 120.1900 29.3700 120.8500 30.2600 ;
      RECT 118.8100 29.3700 119.4700 30.2600 ;
      RECT 117.4300 29.3700 118.0900 30.2600 ;
      RECT 116.0500 29.3700 116.7100 30.2600 ;
      RECT 114.6700 29.3700 115.3300 30.2600 ;
      RECT 113.2900 29.3700 113.9500 30.2600 ;
      RECT 111.9100 29.3700 112.5700 30.2600 ;
      RECT 110.5300 29.3700 111.1900 30.2600 ;
      RECT 109.1500 29.3700 109.8100 30.2600 ;
      RECT 107.7700 29.3700 108.4300 30.2600 ;
      RECT 106.3900 29.3700 107.0500 30.2600 ;
      RECT 105.0100 29.3700 105.6700 30.2600 ;
      RECT 103.6300 29.3700 104.2900 30.2600 ;
      RECT 102.7100 29.3700 102.9100 30.2600 ;
      RECT 101.3300 29.3700 101.9900 30.2600 ;
      RECT 99.9500 29.3700 100.6100 30.2600 ;
      RECT 98.5700 29.3700 99.2300 30.2600 ;
      RECT 97.1900 29.3700 97.8500 30.2600 ;
      RECT 95.8100 29.3700 96.4700 30.2600 ;
      RECT 94.4300 29.3700 95.0900 30.2600 ;
      RECT 93.0500 29.3700 93.7100 30.2600 ;
      RECT 91.6700 29.3700 92.3300 30.2600 ;
      RECT 90.2900 29.3700 90.9500 30.2600 ;
      RECT 88.9100 29.3700 89.5700 30.2600 ;
      RECT 87.5300 29.3700 88.1900 30.2600 ;
      RECT 86.1500 29.3700 86.8100 30.2600 ;
      RECT 84.7700 29.3700 85.4300 30.2600 ;
      RECT 83.3900 29.3700 84.0500 30.2600 ;
      RECT 82.0100 29.3700 82.6700 30.2600 ;
      RECT 80.6300 29.3700 81.2900 30.2600 ;
      RECT 79.7100 29.3700 79.9100 30.2600 ;
      RECT 78.3300 29.3700 78.9900 30.2600 ;
      RECT 76.9500 29.3700 77.6100 30.2600 ;
      RECT 75.5700 29.3700 76.2300 30.2600 ;
      RECT 74.1900 29.3700 74.8500 30.2600 ;
      RECT 72.8100 29.3700 73.4700 30.2600 ;
      RECT 71.4300 29.3700 72.0900 30.2600 ;
      RECT 70.0500 29.3700 70.7100 30.2600 ;
      RECT 68.6700 29.3700 69.3300 30.2600 ;
      RECT 67.2900 29.3700 67.9500 30.2600 ;
      RECT 65.9100 29.3700 66.5700 30.2600 ;
      RECT 64.5300 29.3700 65.1900 30.2600 ;
      RECT 63.1500 29.3700 63.8100 30.2600 ;
      RECT 61.7700 29.3700 62.4300 30.2600 ;
      RECT 60.3900 29.3700 61.0500 30.2600 ;
      RECT 59.0100 29.3700 59.6700 30.2600 ;
      RECT 57.6300 29.3700 58.2900 30.2600 ;
      RECT 56.7100 29.3700 56.9100 30.2600 ;
      RECT 55.3300 29.3700 55.9900 30.2600 ;
      RECT 53.9500 29.3700 54.6100 30.2600 ;
      RECT 52.5700 29.3700 53.2300 30.2600 ;
      RECT 51.1900 29.3700 51.8500 30.2600 ;
      RECT 49.8100 29.3700 50.4700 30.2600 ;
      RECT 48.4300 29.3700 49.0900 30.2600 ;
      RECT 47.0500 29.3700 47.7100 30.2600 ;
      RECT 45.6700 29.3700 46.3300 30.2600 ;
      RECT 44.2900 29.3700 44.9500 30.2600 ;
      RECT 42.9100 29.3700 43.5700 30.2600 ;
      RECT 41.5300 29.3700 42.1900 30.2600 ;
      RECT 40.1500 29.3700 40.8100 30.2600 ;
      RECT 38.7700 29.3700 39.4300 30.2600 ;
      RECT 37.3900 29.3700 38.0500 30.2600 ;
      RECT 36.0100 29.3700 36.6700 30.2600 ;
      RECT 34.6300 29.3700 35.2900 30.2600 ;
      RECT 33.7100 29.3700 33.9100 30.2600 ;
      RECT 32.3300 29.3700 32.9900 30.2600 ;
      RECT 30.9500 29.3700 31.6100 30.2600 ;
      RECT 29.5700 29.3700 30.2300 30.2600 ;
      RECT 28.1900 29.3700 28.8500 30.2600 ;
      RECT 26.8100 29.3700 27.4700 30.2600 ;
      RECT 25.4300 29.3700 26.0900 30.2600 ;
      RECT 24.0500 29.3700 24.7100 30.2600 ;
      RECT 22.6700 29.3700 23.3300 30.2600 ;
      RECT 21.2900 29.3700 21.9500 30.2600 ;
      RECT 19.9100 29.3700 20.5700 30.2600 ;
      RECT 18.5300 29.3700 19.1900 30.2600 ;
      RECT 17.1500 29.3700 17.8100 30.2600 ;
      RECT 15.7700 29.3700 16.4300 30.2600 ;
      RECT 14.3900 29.3700 15.0500 30.2600 ;
      RECT 13.0100 29.3700 13.6700 30.2600 ;
      RECT 11.6300 29.3700 12.2900 30.2600 ;
      RECT 10.7100 29.3700 10.9100 30.2600 ;
      RECT 0.0000 29.3700 9.9900 30.2600 ;
      RECT 0.0000 28.9850 240.1200 29.3700 ;
      RECT 0.5000 28.4750 240.1200 28.9850 ;
      RECT 0.0000 27.9650 240.1200 28.4750 ;
      RECT 0.0000 27.4550 239.6200 27.9650 ;
      RECT 0.0000 26.9450 240.1200 27.4550 ;
      RECT 0.5000 26.4350 240.1200 26.9450 ;
      RECT 0.0000 26.2650 240.1200 26.4350 ;
      RECT 0.0000 25.7550 239.6200 26.2650 ;
      RECT 0.0000 25.2450 240.1200 25.7550 ;
      RECT 0.5000 24.7350 240.1200 25.2450 ;
      RECT 0.0000 24.5650 240.1200 24.7350 ;
      RECT 0.0000 24.0550 239.6200 24.5650 ;
      RECT 0.0000 23.2050 240.1200 24.0550 ;
      RECT 0.5000 22.8650 240.1200 23.2050 ;
      RECT 0.5000 22.6950 239.6200 22.8650 ;
      RECT 0.0000 22.3550 239.6200 22.6950 ;
      RECT 0.0000 21.5050 240.1200 22.3550 ;
      RECT 0.5000 21.1650 240.1200 21.5050 ;
      RECT 0.5000 20.9950 239.6200 21.1650 ;
      RECT 0.0000 20.6550 239.6200 20.9950 ;
      RECT 0.0000 19.4650 240.1200 20.6550 ;
      RECT 0.5000 18.9550 239.6200 19.4650 ;
      RECT 0.0000 17.7650 240.1200 18.9550 ;
      RECT 0.5000 17.2550 239.6200 17.7650 ;
      RECT 0.0000 16.0650 240.1200 17.2550 ;
      RECT 0.5000 15.5550 239.6200 16.0650 ;
      RECT 0.0000 14.3650 240.1200 15.5550 ;
      RECT 0.0000 14.0250 239.6200 14.3650 ;
      RECT 0.5000 13.8550 239.6200 14.0250 ;
      RECT 0.5000 13.5150 240.1200 13.8550 ;
      RECT 0.0000 12.6650 240.1200 13.5150 ;
      RECT 0.0000 12.3250 239.6200 12.6650 ;
      RECT 0.5000 12.1550 239.6200 12.3250 ;
      RECT 0.5000 11.8150 240.1200 12.1550 ;
      RECT 0.0000 10.9650 240.1200 11.8150 ;
      RECT 0.0000 10.6250 239.6200 10.9650 ;
      RECT 0.5000 10.4550 239.6200 10.6250 ;
      RECT 0.5000 10.1150 240.1200 10.4550 ;
      RECT 0.0000 9.2650 240.1200 10.1150 ;
      RECT 0.0000 8.7550 239.6200 9.2650 ;
      RECT 0.0000 8.5850 240.1200 8.7550 ;
      RECT 0.5000 8.0750 240.1200 8.5850 ;
      RECT 0.0000 7.5650 240.1200 8.0750 ;
      RECT 0.0000 7.0550 239.6200 7.5650 ;
      RECT 0.0000 6.8850 240.1200 7.0550 ;
      RECT 0.5000 6.3750 240.1200 6.8850 ;
      RECT 0.0000 5.8650 240.1200 6.3750 ;
      RECT 0.0000 5.3550 239.6200 5.8650 ;
      RECT 0.0000 4.8450 240.1200 5.3550 ;
      RECT 0.5000 4.3350 240.1200 4.8450 ;
      RECT 0.0000 4.1650 240.1200 4.3350 ;
      RECT 0.0000 3.6550 239.6200 4.1650 ;
      RECT 0.0000 3.1450 240.1200 3.6550 ;
      RECT 0.5000 2.6350 240.1200 3.1450 ;
      RECT 0.0000 2.4650 240.1200 2.6350 ;
      RECT 0.0000 1.9550 239.6200 2.4650 ;
      RECT 0.0000 1.4450 240.1200 1.9550 ;
      RECT 0.5000 0.9350 240.1200 1.4450 ;
      RECT 0.0000 0.0000 240.1200 0.9350 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 240.1200 30.2600 ;
    LAYER met2 ;
      RECT 210.3200 29.4000 240.1200 30.2600 ;
      RECT 207.1000 29.4000 209.6600 30.2600 ;
      RECT 204.3400 29.4000 206.4400 30.2600 ;
      RECT 201.5800 29.4000 203.6800 30.2600 ;
      RECT 198.8200 29.4000 200.9200 30.2600 ;
      RECT 195.6000 29.4000 198.1600 30.2600 ;
      RECT 192.8400 29.4000 194.9400 30.2600 ;
      RECT 190.0800 29.4000 192.1800 30.2600 ;
      RECT 187.3200 29.4000 189.4200 30.2600 ;
      RECT 184.5600 29.4000 186.6600 30.2600 ;
      RECT 181.3400 29.4000 183.9000 30.2600 ;
      RECT 178.5800 29.4000 180.6800 30.2600 ;
      RECT 175.8200 29.4000 177.9200 30.2600 ;
      RECT 173.0600 29.4000 175.1600 30.2600 ;
      RECT 170.3000 29.4000 172.4000 30.2600 ;
      RECT 167.0800 29.4000 169.6400 30.2600 ;
      RECT 164.3200 29.4000 166.4200 30.2600 ;
      RECT 161.5600 29.4000 163.6600 30.2600 ;
      RECT 158.8000 29.4000 160.9000 30.2600 ;
      RECT 156.0400 29.4000 158.1400 30.2600 ;
      RECT 0.0000 29.4000 155.3800 30.2600 ;
      RECT 0.0000 28.9400 240.1200 29.4000 ;
      RECT 0.0000 28.5200 239.4950 28.9400 ;
      RECT 0.0000 27.9200 240.1200 28.5200 ;
      RECT 0.6250 27.5000 240.1200 27.9200 ;
      RECT 0.0000 26.9000 240.1200 27.5000 ;
      RECT 0.0000 26.4800 239.4950 26.9000 ;
      RECT 0.0000 26.2200 240.1200 26.4800 ;
      RECT 0.6250 25.8000 240.1200 26.2200 ;
      RECT 0.0000 25.2000 240.1200 25.8000 ;
      RECT 0.0000 24.7800 239.4950 25.2000 ;
      RECT 0.0000 24.5200 240.1200 24.7800 ;
      RECT 0.6250 24.1000 240.1200 24.5200 ;
      RECT 0.0000 23.1600 240.1200 24.1000 ;
      RECT 0.0000 22.8200 239.4950 23.1600 ;
      RECT 0.6250 22.7400 239.4950 22.8200 ;
      RECT 0.6250 22.4000 240.1200 22.7400 ;
      RECT 0.0000 21.4600 240.1200 22.4000 ;
      RECT 0.0000 21.1200 239.4950 21.4600 ;
      RECT 0.6250 21.0400 239.4950 21.1200 ;
      RECT 0.6250 20.7000 240.1200 21.0400 ;
      RECT 0.0000 19.4200 240.1200 20.7000 ;
      RECT 0.6250 19.0000 239.4950 19.4200 ;
      RECT 0.0000 17.7200 240.1200 19.0000 ;
      RECT 0.6250 17.3000 239.4950 17.7200 ;
      RECT 0.0000 16.0200 240.1200 17.3000 ;
      RECT 0.6250 15.6000 239.4950 16.0200 ;
      RECT 0.0000 14.3200 240.1200 15.6000 ;
      RECT 0.6250 13.9800 240.1200 14.3200 ;
      RECT 0.6250 13.9000 239.4950 13.9800 ;
      RECT 0.0000 13.5600 239.4950 13.9000 ;
      RECT 0.0000 12.6200 240.1200 13.5600 ;
      RECT 0.6250 12.2800 240.1200 12.6200 ;
      RECT 0.6250 12.2000 239.4950 12.2800 ;
      RECT 0.0000 11.8600 239.4950 12.2000 ;
      RECT 0.0000 10.9200 240.1200 11.8600 ;
      RECT 0.6250 10.5800 240.1200 10.9200 ;
      RECT 0.6250 10.5000 239.4950 10.5800 ;
      RECT 0.0000 10.1600 239.4950 10.5000 ;
      RECT 0.0000 9.2200 240.1200 10.1600 ;
      RECT 0.6250 8.8000 240.1200 9.2200 ;
      RECT 0.0000 8.5400 240.1200 8.8000 ;
      RECT 0.0000 8.1200 239.4950 8.5400 ;
      RECT 0.0000 7.5200 240.1200 8.1200 ;
      RECT 0.6250 7.1000 240.1200 7.5200 ;
      RECT 0.0000 6.8400 240.1200 7.1000 ;
      RECT 0.0000 6.4200 239.4950 6.8400 ;
      RECT 0.0000 5.8200 240.1200 6.4200 ;
      RECT 0.6250 5.4000 240.1200 5.8200 ;
      RECT 0.0000 4.8000 240.1200 5.4000 ;
      RECT 0.0000 4.3800 239.4950 4.8000 ;
      RECT 0.0000 4.1200 240.1200 4.3800 ;
      RECT 0.6250 3.7000 240.1200 4.1200 ;
      RECT 0.0000 3.1000 240.1200 3.7000 ;
      RECT 0.0000 2.6800 239.4950 3.1000 ;
      RECT 0.0000 2.4200 240.1200 2.6800 ;
      RECT 0.6250 2.0000 240.1200 2.4200 ;
      RECT 0.0000 1.4000 240.1200 2.0000 ;
      RECT 0.0000 0.9800 239.4950 1.4000 ;
      RECT 0.0000 0.8600 240.1200 0.9800 ;
      RECT 179.9600 0.0000 240.1200 0.8600 ;
      RECT 174.4400 0.0000 179.3000 0.8600 ;
      RECT 169.3800 0.0000 173.7800 0.8600 ;
      RECT 163.8600 0.0000 168.7200 0.8600 ;
      RECT 158.8000 0.0000 163.2000 0.8600 ;
      RECT 153.7400 0.0000 158.1400 0.8600 ;
      RECT 147.7600 0.0000 153.0800 0.8600 ;
      RECT 142.7000 0.0000 147.1000 0.8600 ;
      RECT 138.1000 0.0000 142.0400 0.8600 ;
      RECT 132.5800 0.0000 137.4400 0.8600 ;
      RECT 127.5200 0.0000 131.9200 0.8600 ;
      RECT 122.0000 0.0000 126.8600 0.8600 ;
      RECT 116.9400 0.0000 121.3400 0.8600 ;
      RECT 111.8800 0.0000 116.2800 0.8600 ;
      RECT 106.3600 0.0000 111.2200 0.8600 ;
      RECT 101.3000 0.0000 105.7000 0.8600 ;
      RECT 95.7800 0.0000 100.6400 0.8600 ;
      RECT 90.7200 0.0000 95.1200 0.8600 ;
      RECT 85.6600 0.0000 90.0600 0.8600 ;
      RECT 80.6000 0.0000 85.0000 0.8600 ;
      RECT 0.0000 0.0000 79.9400 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 240.1200 30.2600 ;
      RECT 237.8600 25.7000 240.1200 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 240.1200 25.7000 ;
      RECT 234.8600 22.7000 240.1200 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 240.1200 22.7000 ;
      RECT 234.8600 20.2000 240.1200 21.2800 ;
      RECT 7.8600 20.2000 232.2600 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 240.1200 20.2000 ;
      RECT 237.8600 17.4800 240.1200 18.5600 ;
      RECT 4.8600 17.4800 235.2600 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 240.1200 17.4800 ;
      RECT 234.8600 14.7600 240.1200 15.8400 ;
      RECT 7.8600 14.7600 232.2600 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 240.1200 14.7600 ;
      RECT 237.8600 12.0400 240.1200 13.1200 ;
      RECT 4.8600 12.0400 235.2600 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 240.1200 12.0400 ;
      RECT 234.8600 9.3200 240.1200 10.4000 ;
      RECT 7.8600 9.3200 232.2600 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 240.1200 9.3200 ;
      RECT 237.8600 6.6000 240.1200 7.6800 ;
      RECT 4.8600 6.6000 235.2600 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 240.1200 6.6000 ;
      RECT 234.8600 3.7700 240.1200 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 240.1200 3.7700 ;
      RECT 237.8600 0.7700 240.1200 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 240.1200 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 240.1200 30.2600 ;
      RECT 4.8600 25.3000 235.2600 28.3000 ;
      RECT 234.8600 3.7700 235.2600 25.3000 ;
      RECT 7.8600 3.7700 232.2600 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 237.8600 0.7700 240.1200 28.3000 ;
      RECT 4.8600 0.7700 235.2600 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 240.1200 0.7700 ;
  END
END S_term_single2

END LIBRARY
