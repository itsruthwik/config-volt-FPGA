##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 01:11:25 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO N_term_single2
  CLASS BLOCK ;
  SIZE 240.1200 BY 30.2600 ;
  FOREIGN N_term_single2 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.79 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 87.2116 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 465.88 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 0.0000 14.2200 0.7200 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.442 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 21.3248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 112.274 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 0.0000 12.8400 0.7200 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.743 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 39.6148 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 192.884 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 0.0000 11.4600 0.7200 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.1278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 25.2733 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.899 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 0.0000 10.5400 0.7200 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 60.3154 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 295.261 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 0.0000 25.2600 0.7200 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.385 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 29.0909 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.129 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 0.0000 23.8800 0.7200 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.03955 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.223 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.6992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 58.4185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.20975 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.0252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 0.0000 22.5000 0.7200 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.184 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 41.3846 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 201.733 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 0.0000 21.1200 0.7200 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.382 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.4814 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.8365 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 0.0000 19.7400 0.7200 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6229 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 149.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.0382 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 84.3311 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 455.025 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 0.0000 18.3600 0.7200 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.1708 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.7765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.4575 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.4245 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 0.0000 16.9800 0.7200 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.524 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.7318 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.6635 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 0.0000 15.6000 0.7200 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.2705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.106 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 38.9619 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 188.877 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 0.0000 35.8400 0.7200 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.001 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 88.0594 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 463.887 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 0.0000 34.4600 0.7200 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.491 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 32.7066 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 155.374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 0.0000 33.5400 0.7200 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.0116 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.9805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.382 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.08396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.1667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 0.0000 32.1600 0.7200 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8608 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.068 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 34.5871 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 167.745 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 0.0000 30.7800 0.7200 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.28815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.339 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 18.2267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 96.6132 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 0.0000 29.4000 0.7200 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.7532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.53 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 43.8223 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 214.346 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 0.0000 28.0200 0.7200 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 45.9544 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 222.299 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 0.0000 26.6400 0.7200 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.31 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 70.7173 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 376.89 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 0.0000 57.4600 0.7200 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.9418 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 138.714 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 0.0000 56.5400 0.7200 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.28815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.339 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9712 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.25 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.132 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6336 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.695 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 0.0000 55.1600 0.7200 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1217 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.1352 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 0.0000 53.7800 0.7200 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.228 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.3783 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.4182 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 0.0000 52.4000 0.7200 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4864 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.55 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.094 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.1887 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 0.0000 51.0200 0.7200 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.802 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6009 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.0723 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 0.0000 49.6400 0.7200 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 24.3305 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 130.792 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 0.0000 48.2600 0.7200 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.5405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.9848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 56.8255 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 299.044 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 0.0000 46.8800 0.7200 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.1101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 0.0000 45.5000 0.7200 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.09 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 45.8928 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 224.274 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 0.0000 44.1200 0.7200 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.2194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.861 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 49.2336 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 235.173 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 0.0000 42.7400 0.7200 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.521 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 44.4135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 210.582 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 0.0000 41.3600 0.7200 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.4772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 43.4525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 211.33 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 0.0000 39.9800 0.7200 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 18.267 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.012 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.5682 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.3931 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 0.0000 38.6000 0.7200 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.7432 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 68.6385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.249 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 31.6186 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 149.877 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 0.0000 37.2200 0.7200 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.8924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 59.3845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.69277 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.0157 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 0.0000 79.5400 0.7200 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.354 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.6925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.30535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.5031 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 0.0000 78.1600 0.7200 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.567 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.5818 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 0.0000 76.7800 0.7200 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 64.3752 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.409 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 0.0000 75.4000 0.7200 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 48.5513 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 257.654 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 0.0000 74.0200 0.7200 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.6108 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.818 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 36.6374 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 178.421 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 0.0000 72.6400 0.7200 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.2044 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 0.0000 71.2600 0.7200 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.0986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 70.8053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 377.695 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 0.0000 69.8800 0.7200 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.642 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.5091 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.3553 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 0.0000 68.5000 0.7200 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.5357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.2194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 62.2329 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 331.654 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 0.0000 67.1200 0.7200 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 24.9261 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 135.151 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 0.0000 65.7400 0.7200 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8424 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.964 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0965 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.0346 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 0.0000 64.3600 0.7200 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.2135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.204 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 0.0000 62.9800 0.7200 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.51935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.611 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.8548 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 74.1965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.286 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.7708 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.4057 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 0.0000 61.6000 0.7200 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9352 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5615 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1796 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.4245 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 0.0000 60.2200 0.7200 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.90535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.0786 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 0.0000 58.8400 0.7200 ;
    END
  END NN4END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.17555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6114 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.672 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 0.0000 84.6000 0.7200 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2608 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 0.0000 83.2200 0.7200 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.548 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 0.0000 81.8400 0.7200 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 0.0000 80.4600 0.7200 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 0.0000 106.2200 0.7200 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.62 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 0.0000 104.8400 0.7200 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6354 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 0.0000 103.4600 0.7200 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 0.0000 102.5400 0.7200 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 0.0000 101.1600 0.7200 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 0.0000 99.7800 0.7200 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5792 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7815 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 0.0000 98.4000 0.7200 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 0.0000 97.0200 0.7200 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.382 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 0.0000 95.6400 0.7200 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.402 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 0.0000 94.2600 0.7200 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 0.0000 92.8800 0.7200 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 0.0000 91.5000 0.7200 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 0.0000 90.1200 0.7200 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.46155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.543 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.183 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 0.0000 88.7400 0.7200 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2688 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 0.0000 87.3600 0.7200 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.9908 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.8765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.762 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 0.0000 85.9800 0.7200 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48835 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.751 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1158 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.225 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 0.0000 127.8400 0.7200 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.2548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.496 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 0.0000 126.4600 0.7200 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.676 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.3025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 0.0000 125.5400 0.7200 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 0.0000 124.1600 0.7200 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 0.0000 122.7800 0.7200 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4606 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.949 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 0.0000 121.4000 0.7200 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.05995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 0.0000 120.0200 0.7200 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.25075 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.295 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.2556 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.2005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 0.0000 118.6400 0.7200 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.581 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 0.0000 117.2600 0.7200 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.203 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 0.0000 115.8800 0.7200 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 0.0000 114.5000 0.7200 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 0.0000 113.1200 0.7200 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.999 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.638 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 0.0000 111.7400 0.7200 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.77095 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.907 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 0.0000 110.3600 0.7200 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 0.0000 108.9800 0.7200 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75395 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.887 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 0.0000 107.6000 0.7200 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5984 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 0.0000 149.4600 0.7200 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 0.0000 148.5400 0.7200 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.17555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 0.0000 147.1600 0.7200 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.106 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 0.0000 145.7800 0.7200 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4824 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4041 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.664 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 0.0000 144.4000 0.7200 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.559 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 0.0000 143.0200 0.7200 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 0.0000 141.6400 0.7200 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 0.0000 140.2600 0.7200 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 0.0000 138.8800 0.7200 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.12655 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8054 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 0.0000 137.5000 0.7200 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 0.0000 136.1200 0.7200 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7216 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.561 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.581 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 0.0000 134.7400 0.7200 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 0.0000 133.3600 0.7200 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.69275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.815 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.68 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 0.0000 131.9800 0.7200 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.03955 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.223 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.481 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 0.0000 130.6000 0.7200 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.172 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.624 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 0.0000 129.2200 0.7200 ;
    END
  END SS4BEG[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.1956 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.8635 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 43.8959 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 223.047 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.2292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.1716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 46.0821 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 240.494 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.91165 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.249 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.025 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.088 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 77.2462 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 379.755 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.34 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 36.8984 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 194.739 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6392 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.752 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.5464 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.6545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.618 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.0844 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.186 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 33.3267 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 161.868 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3736 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.616 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.5504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.6745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.63742 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.5283 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9078 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 62.9934 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 310.519 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.53805 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.633 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.9168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 69.5065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.966 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 2.71289 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.54088 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.88 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 81.4884 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.818 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9202 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.612 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.1625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.422 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.7821 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.915 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.7164 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 53.5045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 56.419 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 299.925 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.821 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 23.1148 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 122.937 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8296 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.976 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0992 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.26 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.2689 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.9434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.9004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.856 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.2261 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.2673 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.3068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.543 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 25.6858 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.047 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 79.4796 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 415.484 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.298 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7267 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.5063 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 78.3525 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.031 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.724 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2714 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.9119 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.1928 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.745 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.11 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 67.8664 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 334.204 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.254 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.5242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.692 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.063 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 40.5022 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 211.371 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.2564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 58.3827 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 313.748 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.2275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 68.3097 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 335.679 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.8798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 107.349 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 550.44 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 54.3557 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.097 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.493 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 27.9535 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.925 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6528 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.038 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.45503 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.5723 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 104.227 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 540.487 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5909 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.202 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 22.6318 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 125.022 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.433 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 28.6600 240.1200 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.248 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.7048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.896 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 26.6200 240.1200 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.9748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.336 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 24.9200 240.1200 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.494 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 22.8800 240.1200 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 21.1800 240.1200 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.541 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 19.1400 240.1200 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 17.4400 240.1200 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.147 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 15.7400 240.1200 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.915 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 13.7000 240.1200 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 12.0000 240.1200 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.4758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.008 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 10.3000 240.1200 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 8.2600 240.1200 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.9168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.36 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 6.5600 240.1200 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 4.5200 240.1200 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.079 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 2.8200 240.1200 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 1.1200 240.1200 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 22.8324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 114.048 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 27.6250 240.1200 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.358 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.166 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 25.9250 240.1200 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.089 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.8468 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.1195 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 24.2250 240.1200 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.1536 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 85.6905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 22.5250 240.1200 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.911 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4775 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 20.8250 240.1200 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.0228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.592 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 19.1250 240.1200 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6282 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.092 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.1536 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.6905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 17.4250 240.1200 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.6112 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 72.9785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 15.7250 240.1200 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.086 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.3525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.096 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 14.0250 240.1200 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.8352 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.0985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.647 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 12.3250 240.1200 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.3844 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.8445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.454 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 10.6250 240.1200 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7952 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.9536 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 64.6905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.337 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 8.9250 240.1200 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 16.1606 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.766 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 7.2250 240.1200 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6562 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.772 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2328 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.4548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 194.896 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 5.5250 240.1200 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.0212 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.0285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 3.8250 240.1200 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.1164 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.5045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.046 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 2.1250 240.1200 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.3148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 102.224 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 528.786 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.8000 0.0000 210.1800 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 34.7915 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 183.969 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 206.5800 0.0000 206.9600 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.013 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.3316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 75.5248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.233 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 203.8200 0.0000 204.2000 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.5706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 76.8204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.516 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 201.0600 0.0000 201.4400 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0514 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 23.3701 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 129.453 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 198.3000 0.0000 198.6800 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.232 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 49.7928 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.333 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 195.0800 0.0000 195.4600 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.8915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.7547 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.3200 0.0000 192.7000 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.797 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 19.5097 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 105.994 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 189.5600 0.0000 189.9400 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.475 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 29.7101 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 160.95 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 186.8000 0.0000 187.1800 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.533 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.0248 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.513 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 184.0400 0.0000 184.4200 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.769 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 40.3594 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 196.67 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 180.8200 0.0000 181.2000 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.627 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 40.4399 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 192.657 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 178.0600 0.0000 178.4400 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.991 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3796 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.2862 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 175.3000 0.0000 175.6800 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.497 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 31.8085 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 153.173 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 172.5400 0.0000 172.9200 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.993 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 59.828 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.44 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 169.7800 0.0000 170.1600 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.169 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.9582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.921 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 166.5600 0.0000 166.9400 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.545 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 38.5443 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 184.569 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 163.8000 0.0000 164.1800 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.427 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.294 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.0849 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 161.0400 0.0000 161.4200 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.1532 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 88.4079 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 479.358 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 158.2800 0.0000 158.6600 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.8128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 70.3072 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 367.871 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 155.5200 0.0000 155.9000 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.9436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.64 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.8000 29.5400 210.1800 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.0553 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 206.5800 29.5400 206.9600 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.013 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 203.8200 29.5400 204.2000 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.035 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 201.0600 29.5400 201.4400 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4302 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.033 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 198.3000 29.5400 198.6800 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.333 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 195.0800 29.5400 195.4600 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.951 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.3200 29.5400 192.7000 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.717 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 189.5600 29.5400 189.9400 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.8000 29.5400 187.1800 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 184.0400 29.5400 184.4200 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.559 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.8200 29.5400 181.2000 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.5256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 178.0600 29.5400 178.4400 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.429 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 175.3000 29.5400 175.6800 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.963 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 172.5400 29.5400 172.9200 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.763 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 169.7800 29.5400 170.1600 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.397 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.523 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.5600 29.5400 166.9400 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.107 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.8000 29.5400 164.1800 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.069 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.0400 29.5400 161.4200 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.342 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.8200 29.5400 158.2000 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.134 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.5200 29.5400 155.9000 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 234.5600 6.0700 ;
        RECT 5.5600 23.0000 234.5600 25.0000 ;
        RECT 232.5600 15.0600 234.5600 15.5400 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 232.5600 9.6200 234.5600 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 232.5600 20.5000 234.5600 20.9800 ;
      LAYER met4 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
        RECT 232.5600 4.0700 234.5600 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 237.5600 3.0700 ;
        RECT 2.5600 26.0000 237.5600 28.0000 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 235.5600 12.3400 237.5600 12.8200 ;
        RECT 235.5600 6.9000 237.5600 7.3800 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 235.5600 17.7800 237.5600 18.2600 ;
      LAYER met4 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
        RECT 235.5600 1.0700 237.5600 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.0000 28.9850 240.1200 30.2600 ;
      RECT 0.5000 28.4750 240.1200 28.9850 ;
      RECT 0.0000 27.9650 240.1200 28.4750 ;
      RECT 0.0000 27.4550 239.6200 27.9650 ;
      RECT 0.0000 26.9450 240.1200 27.4550 ;
      RECT 0.5000 26.4350 240.1200 26.9450 ;
      RECT 0.0000 26.2650 240.1200 26.4350 ;
      RECT 0.0000 25.7550 239.6200 26.2650 ;
      RECT 0.0000 25.2450 240.1200 25.7550 ;
      RECT 0.5000 24.7350 240.1200 25.2450 ;
      RECT 0.0000 24.5650 240.1200 24.7350 ;
      RECT 0.0000 24.0550 239.6200 24.5650 ;
      RECT 0.0000 23.2050 240.1200 24.0550 ;
      RECT 0.5000 22.8650 240.1200 23.2050 ;
      RECT 0.5000 22.6950 239.6200 22.8650 ;
      RECT 0.0000 22.3550 239.6200 22.6950 ;
      RECT 0.0000 21.5050 240.1200 22.3550 ;
      RECT 0.5000 21.1650 240.1200 21.5050 ;
      RECT 0.5000 20.9950 239.6200 21.1650 ;
      RECT 0.0000 20.6550 239.6200 20.9950 ;
      RECT 0.0000 19.4650 240.1200 20.6550 ;
      RECT 0.5000 18.9550 239.6200 19.4650 ;
      RECT 0.0000 17.7650 240.1200 18.9550 ;
      RECT 0.5000 17.2550 239.6200 17.7650 ;
      RECT 0.0000 16.0650 240.1200 17.2550 ;
      RECT 0.5000 15.5550 239.6200 16.0650 ;
      RECT 0.0000 14.3650 240.1200 15.5550 ;
      RECT 0.0000 14.0250 239.6200 14.3650 ;
      RECT 0.5000 13.8550 239.6200 14.0250 ;
      RECT 0.5000 13.5150 240.1200 13.8550 ;
      RECT 0.0000 12.6650 240.1200 13.5150 ;
      RECT 0.0000 12.3250 239.6200 12.6650 ;
      RECT 0.5000 12.1550 239.6200 12.3250 ;
      RECT 0.5000 11.8150 240.1200 12.1550 ;
      RECT 0.0000 10.9650 240.1200 11.8150 ;
      RECT 0.0000 10.6250 239.6200 10.9650 ;
      RECT 0.5000 10.4550 239.6200 10.6250 ;
      RECT 0.5000 10.1150 240.1200 10.4550 ;
      RECT 0.0000 9.2650 240.1200 10.1150 ;
      RECT 0.0000 8.7550 239.6200 9.2650 ;
      RECT 0.0000 8.5850 240.1200 8.7550 ;
      RECT 0.5000 8.0750 240.1200 8.5850 ;
      RECT 0.0000 7.5650 240.1200 8.0750 ;
      RECT 0.0000 7.0550 239.6200 7.5650 ;
      RECT 0.0000 6.8850 240.1200 7.0550 ;
      RECT 0.5000 6.3750 240.1200 6.8850 ;
      RECT 0.0000 5.8650 240.1200 6.3750 ;
      RECT 0.0000 5.3550 239.6200 5.8650 ;
      RECT 0.0000 4.8450 240.1200 5.3550 ;
      RECT 0.5000 4.3350 240.1200 4.8450 ;
      RECT 0.0000 4.1650 240.1200 4.3350 ;
      RECT 0.0000 3.6550 239.6200 4.1650 ;
      RECT 0.0000 3.1450 240.1200 3.6550 ;
      RECT 0.5000 2.6350 240.1200 3.1450 ;
      RECT 0.0000 2.4650 240.1200 2.6350 ;
      RECT 0.0000 1.9550 239.6200 2.4650 ;
      RECT 0.0000 1.4450 240.1200 1.9550 ;
      RECT 0.5000 0.9350 240.1200 1.4450 ;
      RECT 0.0000 0.8900 240.1200 0.9350 ;
      RECT 149.6300 0.0000 240.1200 0.8900 ;
      RECT 148.7100 0.0000 148.9100 0.8900 ;
      RECT 147.3300 0.0000 147.9900 0.8900 ;
      RECT 145.9500 0.0000 146.6100 0.8900 ;
      RECT 144.5700 0.0000 145.2300 0.8900 ;
      RECT 143.1900 0.0000 143.8500 0.8900 ;
      RECT 141.8100 0.0000 142.4700 0.8900 ;
      RECT 140.4300 0.0000 141.0900 0.8900 ;
      RECT 139.0500 0.0000 139.7100 0.8900 ;
      RECT 137.6700 0.0000 138.3300 0.8900 ;
      RECT 136.2900 0.0000 136.9500 0.8900 ;
      RECT 134.9100 0.0000 135.5700 0.8900 ;
      RECT 133.5300 0.0000 134.1900 0.8900 ;
      RECT 132.1500 0.0000 132.8100 0.8900 ;
      RECT 130.7700 0.0000 131.4300 0.8900 ;
      RECT 129.3900 0.0000 130.0500 0.8900 ;
      RECT 128.0100 0.0000 128.6700 0.8900 ;
      RECT 126.6300 0.0000 127.2900 0.8900 ;
      RECT 125.7100 0.0000 125.9100 0.8900 ;
      RECT 124.3300 0.0000 124.9900 0.8900 ;
      RECT 122.9500 0.0000 123.6100 0.8900 ;
      RECT 121.5700 0.0000 122.2300 0.8900 ;
      RECT 120.1900 0.0000 120.8500 0.8900 ;
      RECT 118.8100 0.0000 119.4700 0.8900 ;
      RECT 117.4300 0.0000 118.0900 0.8900 ;
      RECT 116.0500 0.0000 116.7100 0.8900 ;
      RECT 114.6700 0.0000 115.3300 0.8900 ;
      RECT 113.2900 0.0000 113.9500 0.8900 ;
      RECT 111.9100 0.0000 112.5700 0.8900 ;
      RECT 110.5300 0.0000 111.1900 0.8900 ;
      RECT 109.1500 0.0000 109.8100 0.8900 ;
      RECT 107.7700 0.0000 108.4300 0.8900 ;
      RECT 106.3900 0.0000 107.0500 0.8900 ;
      RECT 105.0100 0.0000 105.6700 0.8900 ;
      RECT 103.6300 0.0000 104.2900 0.8900 ;
      RECT 102.7100 0.0000 102.9100 0.8900 ;
      RECT 101.3300 0.0000 101.9900 0.8900 ;
      RECT 99.9500 0.0000 100.6100 0.8900 ;
      RECT 98.5700 0.0000 99.2300 0.8900 ;
      RECT 97.1900 0.0000 97.8500 0.8900 ;
      RECT 95.8100 0.0000 96.4700 0.8900 ;
      RECT 94.4300 0.0000 95.0900 0.8900 ;
      RECT 93.0500 0.0000 93.7100 0.8900 ;
      RECT 91.6700 0.0000 92.3300 0.8900 ;
      RECT 90.2900 0.0000 90.9500 0.8900 ;
      RECT 88.9100 0.0000 89.5700 0.8900 ;
      RECT 87.5300 0.0000 88.1900 0.8900 ;
      RECT 86.1500 0.0000 86.8100 0.8900 ;
      RECT 84.7700 0.0000 85.4300 0.8900 ;
      RECT 83.3900 0.0000 84.0500 0.8900 ;
      RECT 82.0100 0.0000 82.6700 0.8900 ;
      RECT 80.6300 0.0000 81.2900 0.8900 ;
      RECT 79.7100 0.0000 79.9100 0.8900 ;
      RECT 78.3300 0.0000 78.9900 0.8900 ;
      RECT 76.9500 0.0000 77.6100 0.8900 ;
      RECT 75.5700 0.0000 76.2300 0.8900 ;
      RECT 74.1900 0.0000 74.8500 0.8900 ;
      RECT 72.8100 0.0000 73.4700 0.8900 ;
      RECT 71.4300 0.0000 72.0900 0.8900 ;
      RECT 70.0500 0.0000 70.7100 0.8900 ;
      RECT 68.6700 0.0000 69.3300 0.8900 ;
      RECT 67.2900 0.0000 67.9500 0.8900 ;
      RECT 65.9100 0.0000 66.5700 0.8900 ;
      RECT 64.5300 0.0000 65.1900 0.8900 ;
      RECT 63.1500 0.0000 63.8100 0.8900 ;
      RECT 61.7700 0.0000 62.4300 0.8900 ;
      RECT 60.3900 0.0000 61.0500 0.8900 ;
      RECT 59.0100 0.0000 59.6700 0.8900 ;
      RECT 57.6300 0.0000 58.2900 0.8900 ;
      RECT 56.7100 0.0000 56.9100 0.8900 ;
      RECT 55.3300 0.0000 55.9900 0.8900 ;
      RECT 53.9500 0.0000 54.6100 0.8900 ;
      RECT 52.5700 0.0000 53.2300 0.8900 ;
      RECT 51.1900 0.0000 51.8500 0.8900 ;
      RECT 49.8100 0.0000 50.4700 0.8900 ;
      RECT 48.4300 0.0000 49.0900 0.8900 ;
      RECT 47.0500 0.0000 47.7100 0.8900 ;
      RECT 45.6700 0.0000 46.3300 0.8900 ;
      RECT 44.2900 0.0000 44.9500 0.8900 ;
      RECT 42.9100 0.0000 43.5700 0.8900 ;
      RECT 41.5300 0.0000 42.1900 0.8900 ;
      RECT 40.1500 0.0000 40.8100 0.8900 ;
      RECT 38.7700 0.0000 39.4300 0.8900 ;
      RECT 37.3900 0.0000 38.0500 0.8900 ;
      RECT 36.0100 0.0000 36.6700 0.8900 ;
      RECT 34.6300 0.0000 35.2900 0.8900 ;
      RECT 33.7100 0.0000 33.9100 0.8900 ;
      RECT 32.3300 0.0000 32.9900 0.8900 ;
      RECT 30.9500 0.0000 31.6100 0.8900 ;
      RECT 29.5700 0.0000 30.2300 0.8900 ;
      RECT 28.1900 0.0000 28.8500 0.8900 ;
      RECT 26.8100 0.0000 27.4700 0.8900 ;
      RECT 25.4300 0.0000 26.0900 0.8900 ;
      RECT 24.0500 0.0000 24.7100 0.8900 ;
      RECT 22.6700 0.0000 23.3300 0.8900 ;
      RECT 21.2900 0.0000 21.9500 0.8900 ;
      RECT 19.9100 0.0000 20.5700 0.8900 ;
      RECT 18.5300 0.0000 19.1900 0.8900 ;
      RECT 17.1500 0.0000 17.8100 0.8900 ;
      RECT 15.7700 0.0000 16.4300 0.8900 ;
      RECT 14.3900 0.0000 15.0500 0.8900 ;
      RECT 13.0100 0.0000 13.6700 0.8900 ;
      RECT 11.6300 0.0000 12.2900 0.8900 ;
      RECT 10.7100 0.0000 10.9100 0.8900 ;
      RECT 0.0000 0.0000 9.9900 0.8900 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 240.1200 30.2600 ;
    LAYER met2 ;
      RECT 210.3200 29.4000 240.1200 30.2600 ;
      RECT 207.1000 29.4000 209.6600 30.2600 ;
      RECT 204.3400 29.4000 206.4400 30.2600 ;
      RECT 201.5800 29.4000 203.6800 30.2600 ;
      RECT 198.8200 29.4000 200.9200 30.2600 ;
      RECT 195.6000 29.4000 198.1600 30.2600 ;
      RECT 192.8400 29.4000 194.9400 30.2600 ;
      RECT 190.0800 29.4000 192.1800 30.2600 ;
      RECT 187.3200 29.4000 189.4200 30.2600 ;
      RECT 184.5600 29.4000 186.6600 30.2600 ;
      RECT 181.3400 29.4000 183.9000 30.2600 ;
      RECT 178.5800 29.4000 180.6800 30.2600 ;
      RECT 175.8200 29.4000 177.9200 30.2600 ;
      RECT 173.0600 29.4000 175.1600 30.2600 ;
      RECT 170.3000 29.4000 172.4000 30.2600 ;
      RECT 167.0800 29.4000 169.6400 30.2600 ;
      RECT 164.3200 29.4000 166.4200 30.2600 ;
      RECT 161.5600 29.4000 163.6600 30.2600 ;
      RECT 158.3400 29.4000 160.9000 30.2600 ;
      RECT 156.0400 29.4000 157.6800 30.2600 ;
      RECT 0.0000 29.4000 155.3800 30.2600 ;
      RECT 0.0000 28.9400 240.1200 29.4000 ;
      RECT 0.0000 28.5200 239.4950 28.9400 ;
      RECT 0.0000 27.9200 240.1200 28.5200 ;
      RECT 0.6250 27.5000 240.1200 27.9200 ;
      RECT 0.0000 26.9000 240.1200 27.5000 ;
      RECT 0.0000 26.4800 239.4950 26.9000 ;
      RECT 0.0000 26.2200 240.1200 26.4800 ;
      RECT 0.6250 25.8000 240.1200 26.2200 ;
      RECT 0.0000 25.2000 240.1200 25.8000 ;
      RECT 0.0000 24.7800 239.4950 25.2000 ;
      RECT 0.0000 24.5200 240.1200 24.7800 ;
      RECT 0.6250 24.1000 240.1200 24.5200 ;
      RECT 0.0000 23.1600 240.1200 24.1000 ;
      RECT 0.0000 22.8200 239.4950 23.1600 ;
      RECT 0.6250 22.7400 239.4950 22.8200 ;
      RECT 0.6250 22.4000 240.1200 22.7400 ;
      RECT 0.0000 21.4600 240.1200 22.4000 ;
      RECT 0.0000 21.1200 239.4950 21.4600 ;
      RECT 0.6250 21.0400 239.4950 21.1200 ;
      RECT 0.6250 20.7000 240.1200 21.0400 ;
      RECT 0.0000 19.4200 240.1200 20.7000 ;
      RECT 0.6250 19.0000 239.4950 19.4200 ;
      RECT 0.0000 17.7200 240.1200 19.0000 ;
      RECT 0.6250 17.3000 239.4950 17.7200 ;
      RECT 0.0000 16.0200 240.1200 17.3000 ;
      RECT 0.6250 15.6000 239.4950 16.0200 ;
      RECT 0.0000 14.3200 240.1200 15.6000 ;
      RECT 0.6250 13.9800 240.1200 14.3200 ;
      RECT 0.6250 13.9000 239.4950 13.9800 ;
      RECT 0.0000 13.5600 239.4950 13.9000 ;
      RECT 0.0000 12.6200 240.1200 13.5600 ;
      RECT 0.6250 12.2800 240.1200 12.6200 ;
      RECT 0.6250 12.2000 239.4950 12.2800 ;
      RECT 0.0000 11.8600 239.4950 12.2000 ;
      RECT 0.0000 10.9200 240.1200 11.8600 ;
      RECT 0.6250 10.5800 240.1200 10.9200 ;
      RECT 0.6250 10.5000 239.4950 10.5800 ;
      RECT 0.0000 10.1600 239.4950 10.5000 ;
      RECT 0.0000 9.2200 240.1200 10.1600 ;
      RECT 0.6250 8.8000 240.1200 9.2200 ;
      RECT 0.0000 8.5400 240.1200 8.8000 ;
      RECT 0.0000 8.1200 239.4950 8.5400 ;
      RECT 0.0000 7.5200 240.1200 8.1200 ;
      RECT 0.6250 7.1000 240.1200 7.5200 ;
      RECT 0.0000 6.8400 240.1200 7.1000 ;
      RECT 0.0000 6.4200 239.4950 6.8400 ;
      RECT 0.0000 5.8200 240.1200 6.4200 ;
      RECT 0.6250 5.4000 240.1200 5.8200 ;
      RECT 0.0000 4.8000 240.1200 5.4000 ;
      RECT 0.0000 4.3800 239.4950 4.8000 ;
      RECT 0.0000 4.1200 240.1200 4.3800 ;
      RECT 0.6250 3.7000 240.1200 4.1200 ;
      RECT 0.0000 3.1000 240.1200 3.7000 ;
      RECT 0.0000 2.6800 239.4950 3.1000 ;
      RECT 0.0000 2.4200 240.1200 2.6800 ;
      RECT 0.6250 2.0000 240.1200 2.4200 ;
      RECT 0.0000 1.4000 240.1200 2.0000 ;
      RECT 0.0000 0.9800 239.4950 1.4000 ;
      RECT 0.0000 0.8600 240.1200 0.9800 ;
      RECT 210.3200 0.0000 240.1200 0.8600 ;
      RECT 207.1000 0.0000 209.6600 0.8600 ;
      RECT 204.3400 0.0000 206.4400 0.8600 ;
      RECT 201.5800 0.0000 203.6800 0.8600 ;
      RECT 198.8200 0.0000 200.9200 0.8600 ;
      RECT 195.6000 0.0000 198.1600 0.8600 ;
      RECT 192.8400 0.0000 194.9400 0.8600 ;
      RECT 190.0800 0.0000 192.1800 0.8600 ;
      RECT 187.3200 0.0000 189.4200 0.8600 ;
      RECT 184.5600 0.0000 186.6600 0.8600 ;
      RECT 181.3400 0.0000 183.9000 0.8600 ;
      RECT 178.5800 0.0000 180.6800 0.8600 ;
      RECT 175.8200 0.0000 177.9200 0.8600 ;
      RECT 173.0600 0.0000 175.1600 0.8600 ;
      RECT 170.3000 0.0000 172.4000 0.8600 ;
      RECT 167.0800 0.0000 169.6400 0.8600 ;
      RECT 164.3200 0.0000 166.4200 0.8600 ;
      RECT 161.5600 0.0000 163.6600 0.8600 ;
      RECT 158.8000 0.0000 160.9000 0.8600 ;
      RECT 156.0400 0.0000 158.1400 0.8600 ;
      RECT 0.0000 0.0000 155.3800 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 240.1200 30.2600 ;
      RECT 237.8600 25.7000 240.1200 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 240.1200 25.7000 ;
      RECT 234.8600 22.7000 240.1200 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 240.1200 22.7000 ;
      RECT 234.8600 20.2000 240.1200 21.2800 ;
      RECT 7.8600 20.2000 232.2600 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 240.1200 20.2000 ;
      RECT 237.8600 17.4800 240.1200 18.5600 ;
      RECT 4.8600 17.4800 235.2600 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 240.1200 17.4800 ;
      RECT 234.8600 14.7600 240.1200 15.8400 ;
      RECT 7.8600 14.7600 232.2600 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 240.1200 14.7600 ;
      RECT 237.8600 12.0400 240.1200 13.1200 ;
      RECT 4.8600 12.0400 235.2600 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 240.1200 12.0400 ;
      RECT 234.8600 9.3200 240.1200 10.4000 ;
      RECT 7.8600 9.3200 232.2600 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 240.1200 9.3200 ;
      RECT 237.8600 6.6000 240.1200 7.6800 ;
      RECT 4.8600 6.6000 235.2600 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 240.1200 6.6000 ;
      RECT 234.8600 3.7700 240.1200 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 240.1200 3.7700 ;
      RECT 237.8600 0.7700 240.1200 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 240.1200 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 240.1200 30.2600 ;
      RECT 4.8600 25.3000 235.2600 28.3000 ;
      RECT 234.8600 3.7700 235.2600 25.3000 ;
      RECT 7.8600 3.7700 232.2600 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 237.8600 0.7700 240.1200 28.3000 ;
      RECT 4.8600 0.7700 235.2600 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 240.1200 0.7700 ;
  END
END N_term_single2

END LIBRARY
