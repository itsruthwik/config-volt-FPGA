##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 02:01:49 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RAM_IO
  CLASS BLOCK ;
  SIZE 100.2800 BY 219.6400 ;
  FOREIGN RAM_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.358 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7545 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.5332 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.392 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 7.8600 218.9200 8.2400 219.6400 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.62 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.5164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 6.9400 218.9200 7.3200 219.6400 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.6868 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.455 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.0008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 6.0200 218.9200 6.4000 219.6400 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.517 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.8198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.176 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 5.1000 218.9200 5.4800 219.6400 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.6754 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.141 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 218.9200 16.9800 219.6400 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.0796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.032 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 218.9200 15.6000 219.6400 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21295 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.427 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.6556 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.2878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.672 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 14.3000 218.9200 14.6800 219.6400 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.5396 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.3800 218.9200 13.7600 219.6400 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.3586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.52 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 12.0000 218.9200 12.3800 219.6400 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.2817 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.0848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.256 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 218.9200 11.4600 219.6400 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77395 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.087 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.414 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 218.9200 10.5400 219.6400 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.04255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.3208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 9.2400 218.9200 9.6200 219.6400 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.432 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 218.9200 25.2600 219.6400 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.8376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.408 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.9600 218.9200 24.3400 219.6400 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.5956 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.904 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 22.5800 218.9200 22.9600 219.6400 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.758 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 21.6600 218.9200 22.0400 219.6400 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.853 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 218.9200 21.1200 219.6400 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.9078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 293.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 218.9200 19.7400 219.6400 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.368 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 18.4400 218.9200 18.8200 219.6400 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.318 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 17.5200 218.9200 17.9000 219.6400 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 41.4400 218.9200 41.8200 219.6400 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.6436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 40.5200 218.9200 40.9000 219.6400 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.471 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.4228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.392 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 218.9200 39.9800 219.6400 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.066 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.6800 218.9200 39.0600 219.6400 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.07 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.7248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 37.3000 218.9200 37.6800 219.6400 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.0688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.226 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.3800 218.9200 36.7600 219.6400 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 218.9200 35.8400 219.6400 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.1845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 218.9200 34.4600 219.6400 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.156 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 218.9200 33.5400 219.6400 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 32.2400 218.9200 32.6200 219.6400 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7545 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.4828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.3200 218.9200 31.7000 219.6400 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.9400 218.9200 30.3200 219.6400 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.46155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.543 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.4225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.844 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 218.9200 29.4000 219.6400 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.0728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.192 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 28.1000 218.9200 28.4800 219.6400 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.7200 218.9200 27.1000 219.6400 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.38 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 25.8000 218.9200 26.1800 219.6400 ;
    END
  END N4BEG[0]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.05995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1357 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4595 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1232 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 7.8600 0.0000 8.2400 0.7200 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.17815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.739 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1232 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.5088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.184 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 6.9400 0.0000 7.3200 0.7200 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1232 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 6.0200 0.0000 6.4000 0.7200 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.2264 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.031 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.9008 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.359 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.1232 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8894 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.877 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 5.1000 0.0000 5.4800 0.7200 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.6284 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 52.3204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 268.653 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 0.0000 16.9800 0.7200 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.1735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.009 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.89589 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.0303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 0.0000 15.6000 0.7200 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.63795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.97 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.624 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.91475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.0337 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 14.3000 0.0000 14.6800 0.7200 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.6028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 85.6912 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 454.42 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 13.3800 0.0000 13.7600 0.7200 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 41.2199 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.409 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 12.0000 0.0000 12.3800 0.7200 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.736 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.70788 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.0902 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 0.0000 11.4600 0.7200 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.4633 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.0798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.4257 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 95.3724 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 0.0000 10.5400 0.7200 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2998 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.317 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 0.956768 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 3.48013 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 9.2400 0.0000 9.6200 0.7200 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.23335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.8707 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.216 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 0.0000 25.2600 0.7200 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.531 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.5775 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.618 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 23.9600 0.0000 24.3400 0.7200 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5128 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.328 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.5800 0.0000 22.9600 0.7200 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.3728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 21.6600 0.0000 22.0400 0.7200 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.1908 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.5176 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.514 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 0.0000 21.1200 0.7200 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.498 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 0.0000 19.7400 0.7200 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2328 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.7896 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.83 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 18.4400 0.0000 18.8200 0.7200 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.5398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.016 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 17.5200 0.0000 17.9000 0.7200 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.6478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.33643 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 37.0384 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 41.4400 0.0000 41.8200 0.7200 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.702 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.97077 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.3912 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 40.5200 0.0000 40.9000 0.7200 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0098 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9715 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0377 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.3308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 61.1037 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.003 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 0.0000 39.9800 0.7200 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.676 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.3025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.1456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.9366 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 227.317 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 38.6800 0.0000 39.0600 0.7200 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.6508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.9937 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.599 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 37.3000 0.0000 37.6800 0.7200 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.3365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.5115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.9096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 56.2769 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.444 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 36.3800 0.0000 36.7600 0.7200 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.94418 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.6303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 0.0000 35.8400 0.7200 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4041 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.1706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.7267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 371.41 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 0.0000 34.4600 0.7200 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.40675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4056 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.954 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 14.3106 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 70.3219 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 0.0000 33.5400 0.7200 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3611 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.5918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 296.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 81.1692 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.391 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 32.2400 0.0000 32.6200 0.7200 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.40675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.9938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.0023 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 31.3200 0.0000 31.7000 0.7200 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.6944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.3428 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 425.098 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 29.9400 0.0000 30.3200 0.7200 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.182 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.8123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3477 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.9314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 0.0000 29.4000 0.7200 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9504 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.116 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 28.1000 0.0000 28.4800 0.7200 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9504 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.7308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.612 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.7200 0.0000 27.1000 0.7200 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7013 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.4028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.952 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 25.8000 0.0000 26.1800 0.7200 ;
    END
  END N4END[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.413 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3104 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.744 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 84.6400 0.7200 85.0200 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6362 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.073 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0779 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3104 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0567 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.768 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 82.9400 0.7200 83.3200 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7586 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.206 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.3104 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0977 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.32 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 81.5800 0.7200 81.9600 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.9549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.4855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.3104 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.008 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 80.2200 0.7200 80.6000 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3446 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.615 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.76 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 96.2000 0.7200 96.5800 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.199 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.887 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.168 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 94.8400 0.7200 95.2200 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3446 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.615 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.4939 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 93.4800 0.7200 93.8600 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6254 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.429 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 91.7800 0.7200 92.1600 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8678 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.194 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.9728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.992 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 90.4200 0.7200 90.8000 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.199 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.887 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4913 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.0844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 89.0600 0.7200 89.4400 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5378 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.581 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.562 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 87.3600 0.7200 87.7400 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8238 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.974 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.1686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.017 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 86.0000 0.7200 86.3800 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9074 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.429 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.8695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 108.1000 0.7200 108.4800 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7006 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.231 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.784 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 106.4000 0.7200 106.7800 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8602 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.193 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.882 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.3594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.328 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 105.0400 0.7200 105.4200 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.3616 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.536 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 103.6800 0.7200 104.0600 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.886 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 101.9800 0.7200 102.3600 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1106 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.0578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.112 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 100.6200 0.7200 101.0000 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.837 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.077 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.684 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 99.2600 0.7200 99.6400 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5018 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.364 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.8877 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 97.5600 0.7200 97.9400 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6102 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.906 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.7316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.176 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 131.5600 0.7200 131.9400 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.6305 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.632 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 129.8600 0.7200 130.2400 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7023 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4035 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.484 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 127.8200 0.7200 128.2000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8906 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.1255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.272 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 127.1400 0.7200 127.5200 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5714 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.4698 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.976 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 125.4400 0.7200 125.8200 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.6738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.064 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 124.0800 0.7200 124.4600 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1908 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.9416 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4955 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 122.7200 0.7200 123.1000 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7414 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.599 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9516 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.178 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 121.3600 0.7200 121.7400 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0666 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 119.6600 0.7200 120.0400 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2906 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 118.3000 0.7200 118.6800 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0158 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.971 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.96 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 116.9400 0.7200 117.3200 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9038 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.411 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.141 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 115.2400 0.7200 115.6200 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.7802 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.68 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 113.8800 0.7200 114.2600 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4062 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.923 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.3525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 112.5200 0.7200 112.9000 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3744 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.6343 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.922 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.144 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 110.8200 0.7200 111.2000 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0194 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.989 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.928 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 109.4600 0.7200 109.8400 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.282 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 149.2400 0.7200 149.6200 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3426 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.568 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.929 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.64 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 147.2000 0.7200 147.5800 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.664 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 146.1800 0.7200 146.5600 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4013 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 144.8200 0.7200 145.2000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.633 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.057 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.0363 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.3318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.24 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 142.7800 0.7200 143.1600 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9582 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.683 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.55 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6422 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.64 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 141.7600 0.7200 142.1400 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.848 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 139.7200 0.7200 140.1000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4478 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.094 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.824 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 138.3600 0.7200 138.7400 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0186 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8435 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.3068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.44 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 137.3400 0.7200 137.7200 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7955 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.512 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 135.9800 0.7200 136.3600 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6022 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.903 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.756 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.3226 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.033 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 134.2800 0.7200 134.6600 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4442 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.2492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 132.9200 0.7200 133.3000 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.3846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.992 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 45.5800 0.0000 45.9600 0.7200 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.9942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.735 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 44.6600 0.0000 45.0400 0.7200 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.5038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.824 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 0.0000 44.1200 0.7200 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0836 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3467 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.056 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.8200 0.0000 43.2000 0.7200 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 0.0000 62.9800 0.7200 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.472 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.3448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.976 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.6800 0.0000 62.0600 0.7200 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.3098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.456 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 60.3000 0.0000 60.6800 0.7200 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.0808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.3800 0.0000 59.7600 0.7200 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.1536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 193.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 0.0000 58.8400 0.7200 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.7228 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.378 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 57.5400 0.0000 57.9200 0.7200 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.6088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.808 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 0.0000 56.5400 0.7200 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.7258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.008 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 55.2400 0.0000 55.6200 0.7200 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.9108 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.48 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 54.3200 0.0000 54.7000 0.7200 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.466 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.9400 0.0000 53.3200 0.7200 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.34895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.53 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 0.0000 52.4000 0.7200 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.2758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 332.608 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 51.1000 0.0000 51.4800 0.7200 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.7508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 313.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 50.1800 0.0000 50.5600 0.7200 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.056 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 48.8000 0.0000 49.1800 0.7200 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.23335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.776 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 0.0000 48.2600 0.7200 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.3826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 46.9600 0.0000 47.3400 0.7200 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.5248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.936 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 0.0000 79.5400 0.7200 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 78.2400 0.0000 78.6200 0.7200 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.827 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.061 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 77.3200 0.0000 77.7000 0.7200 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.63795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.6508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 302.608 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 0.0000 76.7800 0.7200 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.8504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1375 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 0.0000 75.4000 0.7200 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.4614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 291.872 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 74.1000 0.0000 74.4800 0.7200 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.4588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 73.1800 0.0000 73.5600 0.7200 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.9456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.6135 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.7628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.4986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 0.0000 72.6400 0.7200 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.856 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 0.0000 71.2600 0.7200 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.9600 0.0000 70.3400 0.7200 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.63795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.739 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.0148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.216 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 69.0400 0.0000 69.4200 0.7200 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 315.888 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 67.6600 0.0000 68.0400 0.7200 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.222 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.0325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 0.0000 67.1200 0.7200 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.3576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.336 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.8200 0.0000 66.2000 0.7200 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.3576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.594 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 64.9000 0.0000 65.2800 0.7200 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.9948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 325.776 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 63.5200 0.0000 63.9000 0.7200 ;
    END
  END S4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9169 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.399 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 1.1268 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.502 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.5800 218.9200 45.9600 219.6400 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.2658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.888 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 44.6600 218.9200 45.0400 219.6400 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.432 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 218.9200 44.1200 219.6400 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1988 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.1285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1268 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.928 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 42.8200 218.9200 43.2000 219.6400 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.40675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.976 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.35205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.0613 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 218.9200 62.9800 219.6400 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.6418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 86.6063 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 458.568 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 61.6800 218.9200 62.0600 219.6400 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.4768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 61.056 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.886 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 60.3000 218.9200 60.6800 219.6400 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6132 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9515 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3186 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.249 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.51744 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.8882 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 59.3800 218.9200 59.7600 219.6400 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4315 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.67192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.6801 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.264 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.5491 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 117.659 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 218.9200 58.8400 219.6400 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.7356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 61.8823 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.288 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 57.5400 218.9200 57.9200 219.6400 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.473 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.6128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 31.1323 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.352 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 218.9200 56.5400 219.6400 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.2252 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.542 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.50626 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.9912 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 55.2400 218.9200 55.6200 219.6400 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.104 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 54.3200 218.9200 54.7000 219.6400 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.7858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 287.328 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.9400 218.9200 53.3200 219.6400 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.7338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.384 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 218.9200 52.4000 219.6400 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.07 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 51.1000 218.9200 51.4800 219.6400 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 50.1800 218.9200 50.5600 219.6400 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 16.6623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.9045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.077 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 48.8000 218.9200 49.1800 219.6400 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.38975 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.635 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.1796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 218.9200 48.2600 219.6400 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.7272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.924 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 46.9600 218.9200 47.3400 219.6400 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.05995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.8932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.77 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.41859 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.7892 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 218.9200 79.5400 219.6400 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.2352 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 46.0985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.89347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.0727 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 78.2400 218.9200 78.6200 219.6400 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.63771 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 6.79394 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.3200 218.9200 77.7000 219.6400 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.63795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.2896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.23151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.763 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 218.9200 76.7800 219.6400 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.3916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 42.071 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.87 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 218.9200 75.4000 219.6400 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.11775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.0506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 294.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.5908 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 428.897 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 74.1000 218.9200 74.4800 219.6400 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.59715 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.879 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0964 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.618 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.32512 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.231 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 73.1800 218.9200 73.5600 219.6400 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.23335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.38061 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.5084 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 218.9200 72.6400 219.6400 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.9688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.7191 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 417.282 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 218.9200 71.2600 219.6400 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8075 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6229 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.1884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 12.7581 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 67.1111 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 69.9600 218.9200 70.3400 219.6400 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.132 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.31475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.0202 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 69.0400 218.9200 69.4200 219.6400 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.35865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 5.39865 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 67.6600 218.9200 68.0400 219.6400 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5724 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.0505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.9848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.3318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.24 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 218.9200 67.1200 219.6400 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.1388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 278.544 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 65.8200 218.9200 66.2000 219.6400 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.56 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 64.9000 218.9200 65.2800 219.6400 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3752 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5724 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.8999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.4315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.954 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.928 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 63.5200 218.9200 63.9000 219.6400 ;
    END
  END S4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9818 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.801 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.737 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.224 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 13.9200 0.7200 14.3000 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.731 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.547 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 12.5600 0.7200 12.9400 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9378 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.581 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 11.2000 0.7200 11.5800 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7482 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.633 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.4314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.712 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 9.8400 0.7200 10.2200 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.38 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.5704 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.12 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 25.8200 0.7200 26.2000 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7123 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.4535 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.42 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 24.4600 0.7200 24.8400 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.481 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 22.7600 0.7200 23.1400 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.296 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 21.4000 0.7200 21.7800 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.481 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.38 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.6164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.032 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 20.0400 0.7200 20.4200 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 18.3400 0.7200 18.7200 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4986 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.348 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 16.9800 0.7200 17.3600 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3278 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.531 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.9278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.752 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 15.6200 0.7200 16.0000 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3754 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.769 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5301 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 37.7200 0.7200 38.1000 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3196 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.453 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.598 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 36.0200 0.7200 36.4000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.481 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.1388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.544 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 34.6600 0.7200 35.0400 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8938 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.3548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.696 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 33.3000 0.7200 33.6800 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.607 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.696 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 31.6000 0.7200 31.9800 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2802 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.293 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.592 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 30.2400 0.7200 30.6200 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5718 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.751 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.5048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.496 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 28.8800 0.7200 29.2600 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6646 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.178 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.0633 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.1455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 27.1800 0.7200 27.5600 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.673 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.6998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.536 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 61.1800 0.7200 61.5600 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.504 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 58.8000 0.7200 59.1800 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.275 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 58.1200 0.7200 58.5000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.945 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.3508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.008 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 56.7600 0.7200 57.1400 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.047 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 55.0600 0.7200 55.4400 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3414 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.599 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.632 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 53.7000 0.7200 54.0800 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.024 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 52.3400 0.7200 52.7200 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5718 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.751 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.991 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.8584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.656 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 50.6400 0.7200 51.0200 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.481 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 132.174 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 49.2800 0.7200 49.6600 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5766 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.738 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 47.9200 0.7200 48.3000 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.409 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.937 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 46.2200 0.7200 46.6000 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0702 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.243 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.2886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.48 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 44.8600 0.7200 45.2400 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.549 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.9726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.128 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 43.5000 0.7200 43.8800 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3611 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.368 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 41.8000 0.7200 42.1800 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5006 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.77 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 40.4400 0.7200 40.8200 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3414 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.599 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.5734 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.136 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 39.0800 0.7200 39.4600 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.695 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.33 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.622 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.824 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 78.5200 0.7200 78.9000 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6774 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.279 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.557 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 77.1600 0.7200 77.5400 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0534 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4913 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.7134 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.216 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 75.8000 0.7200 76.1800 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5042 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.413 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.3728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.792 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 74.1000 0.7200 74.4800 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0914 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.312 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.646 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 72.7400 0.7200 73.1200 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2158 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.971 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.696 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 71.3800 0.7200 71.7600 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.871 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.7171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.7918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.36 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 69.6800 0.7200 70.0600 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.0736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 69.0000 0.7200 69.3800 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.181 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.4318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.44 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 67.3000 0.7200 67.6800 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.2766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.416 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 65.6000 0.7200 65.9800 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6838 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.311 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 64.2400 0.7200 64.6200 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19805 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.7858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.328 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 62.5400 0.7200 62.9200 ;
    END
  END W6BEG[0]
  PIN RAM2FAB_D0_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5844 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.777 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.08 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 50.5401 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.952 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 45.2000 100.2800 45.5800 ;
    END
  END RAM2FAB_D0_I0
  PIN RAM2FAB_D0_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3387 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.481 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 44.9091 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 212.452 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 50.3028 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 238.952 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 48.2600 100.2800 48.6400 ;
    END
  END RAM2FAB_D0_I1
  PIN RAM2FAB_D0_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.0528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 91.594 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 473.097 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 52.3400 100.2800 52.7200 ;
    END
  END RAM2FAB_D0_I2
  PIN RAM2FAB_D0_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.4963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.3105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.1317 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 81.4647 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 414.028 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 54.3800 100.2800 54.7600 ;
    END
  END RAM2FAB_D0_I3
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.7206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 62.886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 337.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 14.2045 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 75.4134 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 80.5400 0.0000 80.9200 0.7200 ;
    END
  END UserCLK
  PIN RAM2FAB_D1_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.091 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 14.1313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.9834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 74.023 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 382.518 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 32.9600 100.2800 33.3400 ;
    END
  END RAM2FAB_D1_I0
  PIN RAM2FAB_D1_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6638 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.211 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.224 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 23.9056 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.077 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.318651 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 36.3600 100.2800 36.7400 ;
    END
  END RAM2FAB_D1_I1
  PIN RAM2FAB_D1_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9582 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.683 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.004 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 30.8214 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 142.188 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.318651 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 40.7800 100.2800 41.1600 ;
    END
  END RAM2FAB_D1_I2
  PIN RAM2FAB_D1_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.3646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.7308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 67.046 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.246 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 42.4800 100.2800 42.8600 ;
    END
  END RAM2FAB_D1_I3
  PIN RAM2FAB_D2_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.843 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.107 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.339 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 55.4845 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 288.935 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 21.4000 100.2800 21.7800 ;
    END
  END RAM2FAB_D2_I0
  PIN RAM2FAB_D2_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.819 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 54.2798 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.45 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 24.4600 100.2800 24.8400 ;
    END
  END RAM2FAB_D2_I1
  PIN RAM2FAB_D2_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2158 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.971 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 45.1567 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.694 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 27.5200 100.2800 27.9000 ;
    END
  END RAM2FAB_D2_I2
  PIN RAM2FAB_D2_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.463 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.4077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 43.7825 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.343 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 30.5800 100.2800 30.9600 ;
    END
  END RAM2FAB_D2_I3
  PIN RAM2FAB_D3_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4482 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 65.5163 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.141 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 9.8400 100.2800 10.2200 ;
    END
  END RAM2FAB_D3_I0
  PIN RAM2FAB_D3_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4416 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.026 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 21.4889 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 97.3968 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.163 LAYER met2  ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 34.504 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 161.536 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 12.5600 100.2800 12.9400 ;
    END
  END RAM2FAB_D3_I1
  PIN RAM2FAB_D3_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2498 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.942 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 36.4385 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.911 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 15.6200 100.2800 16.0000 ;
    END
  END RAM2FAB_D3_I2
  PIN RAM2FAB_D3_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.481 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.4741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.7275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.505 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.8906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 80.3167 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.028 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.636111 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 19.0200 100.2800 19.4000 ;
    END
  END RAM2FAB_D3_I3
  PIN FAB2RAM_D0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2498 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 140.0600 100.2800 140.4400 ;
    END
  END FAB2RAM_D0_O0
  PIN FAB2RAM_D0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7838 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.774 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.3938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.904 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 143.4600 100.2800 143.8400 ;
    END
  END FAB2RAM_D0_O1
  PIN FAB2RAM_D0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.661 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.16 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 144.1400 100.2800 144.5200 ;
    END
  END FAB2RAM_D0_O2
  PIN FAB2RAM_D0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6014 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9025 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 149.5800 100.2800 149.9600 ;
    END
  END FAB2RAM_D0_O3
  PIN FAB2RAM_D1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5196 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.453 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 128.8400 100.2800 129.2200 ;
    END
  END FAB2RAM_D1_O0
  PIN FAB2RAM_D1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.436 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.2987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.2045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.28 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 131.5600 100.2800 131.9400 ;
    END
  END FAB2RAM_D1_O1
  PIN FAB2RAM_D1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8818 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.264 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.117 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 134.6200 100.2800 135.0000 ;
    END
  END FAB2RAM_D1_O2
  PIN FAB2RAM_D1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3278 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.531 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.4478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.192 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 137.6800 100.2800 138.0600 ;
    END
  END FAB2RAM_D1_O3
  PIN FAB2RAM_D2_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.688 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 116.6000 100.2800 116.9800 ;
    END
  END FAB2RAM_D2_O0
  PIN FAB2RAM_D2_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2802 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.293 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5269 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.9818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 119.6600 100.2800 120.0400 ;
    END
  END FAB2RAM_D2_O1
  PIN FAB2RAM_D2_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1462 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.586 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.7888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.344 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 122.7200 100.2800 123.1000 ;
    END
  END FAB2RAM_D2_O2
  PIN FAB2RAM_D2_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8262 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.023 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.7978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.392 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 125.4400 100.2800 125.8200 ;
    END
  END FAB2RAM_D2_O3
  PIN FAB2RAM_D3_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.6262 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0265 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 105.0400 100.2800 105.4200 ;
    END
  END FAB2RAM_D3_O0
  PIN FAB2RAM_D3_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2792 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.278 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 107.7600 100.2800 108.1400 ;
    END
  END FAB2RAM_D3_O1
  PIN FAB2RAM_D3_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.311 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.447 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.496 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 110.8200 100.2800 111.2000 ;
    END
  END FAB2RAM_D3_O2
  PIN FAB2RAM_D3_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1854 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.188 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 113.8800 100.2800 114.2600 ;
    END
  END FAB2RAM_D3_O3
  PIN FAB2RAM_A0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8695 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.8918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.56 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 92.8000 100.2800 93.1800 ;
    END
  END FAB2RAM_A0_O0
  PIN FAB2RAM_A0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.475 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.23 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 95.8600 100.2800 96.2400 ;
    END
  END FAB2RAM_A0_O1
  PIN FAB2RAM_A0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.849 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.063 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 98.9200 100.2800 99.3000 ;
    END
  END FAB2RAM_A0_O2
  PIN FAB2RAM_A0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2498 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.784 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 101.9800 100.2800 102.3600 ;
    END
  END FAB2RAM_A0_O3
  PIN FAB2RAM_A1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2158 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.971 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.5578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.112 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 80.9000 100.2800 81.2800 ;
    END
  END FAB2RAM_A1_O0
  PIN FAB2RAM_A1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2802 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.293 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.722 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 84.3000 100.2800 84.6800 ;
    END
  END FAB2RAM_A1_O1
  PIN FAB2RAM_A1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.2658 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2615 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 87.3600 100.2800 87.7400 ;
    END
  END FAB2RAM_A1_O2
  PIN FAB2RAM_A1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1482 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.633 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.656 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 90.0800 100.2800 90.4600 ;
    END
  END FAB2RAM_A1_O3
  PIN FAB2RAM_C_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.409 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.937 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.551 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.9458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.848 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 69.0000 100.2800 69.3800 ;
    END
  END FAB2RAM_C_O0
  PIN FAB2RAM_C_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2498 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.127 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.2506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.944 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 70.7000 100.2800 71.0800 ;
    END
  END FAB2RAM_C_O1
  PIN FAB2RAM_C_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.9868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.4 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 75.1200 100.2800 75.5000 ;
    END
  END FAB2RAM_C_O2
  PIN FAB2RAM_C_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4714 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.212 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.8068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.44 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 78.1800 100.2800 78.5600 ;
    END
  END FAB2RAM_C_O3
  PIN Config_accessC_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5686 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.816 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 57.1000 100.2800 57.4800 ;
    END
  END Config_accessC_bit0
  PIN Config_accessC_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2602 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1965 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 60.1600 100.2800 60.5400 ;
    END
  END Config_accessC_bit1
  PIN Config_accessC_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.087 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.327 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.624 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 62.8800 100.2800 63.2600 ;
    END
  END Config_accessC_bit2
  PIN Config_accessC_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.3596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6935 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.5600 66.6200 100.2800 67.0000 ;
    END
  END Config_accessC_bit3
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.5125 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 45.0138 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 236.232 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 209.3100 0.7200 209.6900 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.1005 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 44.612 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.528 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.6587 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 207.4800 0.7200 207.8600 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.7156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.7442 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 51.4638 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 262.909 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.666038 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 205.6500 0.7200 206.0300 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.7326 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 181.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 63.3108 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.669 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 203.8200 0.7200 204.2000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.6986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 31.8394 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 158.39 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.496889 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 201.9900 0.7200 202.3700 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.3984 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 243.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 48.231 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.368 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 200.1600 0.7200 200.5400 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8516 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 35.75 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.014 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.898293 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 198.3300 0.7200 198.7100 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1811 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 31.0406 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 150.297 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643096 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 196.5000 0.7200 196.8800 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2429 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 38.0249 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 188.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.684338 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.0596 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.112 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 44.91 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 225.454 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 195.2800 0.7200 195.6600 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1482 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 26.6258 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.404 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.646721 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 193.4500 0.7200 193.8300 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.2106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 44.1779 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 222.791 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.666038 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 191.6200 0.7200 192.0000 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.3154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.1716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 28.9509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.148 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.666038 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 189.7900 0.7200 190.1700 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 73.4572 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 364 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.064 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.36 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 80.773 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.026 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 187.9600 0.7200 188.3400 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5169 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 38.4727 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.962 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.758281 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.901 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.824 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 41.0026 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 206.463 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 186.1300 0.7200 186.5100 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1012 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 21.8999 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 105.753 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 184.3000 0.7200 184.6800 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4433 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 22.7959 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 111.106 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 182.4700 0.7200 182.8500 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 26.1869 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 126.492 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 181.2500 0.7200 181.6300 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 27.2451 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 133.125 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.684338 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.5116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.336 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 52.2212 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 270.393 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.99413 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 179.4200 0.7200 179.8000 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.9277 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 188.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met3  ;
    ANTENNAMAXAREACAR 51.1314 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 256.596 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.897574 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4674 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.904 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 52.618 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.129 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.897574 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 177.5900 0.7200 177.9700 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.6944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 45.5028 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 231.761 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 175.7600 0.7200 176.1400 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.1386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 62.3718 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.496 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 173.9300 0.7200 174.3100 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.1763 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 64.3569 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.872 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 172.1000 0.7200 172.4800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 24.7998 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.669182 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 170.2700 0.7200 170.6500 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 46.0129 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 231.322 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.653459 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.6685 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.688 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 54.874 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.777 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 168.4400 0.7200 168.8200 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.4928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 38.6597 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 192.354 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.506709 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 167.2200 0.7200 167.6000 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13455 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 23.4159 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.542829 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6764 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.352 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 52.6317 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 264.389 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 165.3900 0.7200 165.7700 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 35.9607 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.309 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.843564 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 163.5600 0.7200 163.9400 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 60.9975 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 310.572 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.3694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 205.568 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 77.4474 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 398.704 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 161.7300 0.7200 162.1100 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.3873 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 33.1644 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.564 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 159.9000 0.7200 160.2800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 27.3143 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.128 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.499078 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 158.0700 0.7200 158.4500 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 24.9422 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 121.028 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.529452 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.4846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.712 LAYER met4  ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 42.1168 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.354 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 156.2400 0.7200 156.6200 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met4  ;
    ANTENNAMAXAREACAR 21.4844 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.344 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.607715 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 155.0200 0.7200 155.4000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.1224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 209.3100 100.2800 209.6900 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 207.4800 100.2800 207.8600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2066 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.3056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.904 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 205.6500 100.2800 206.0300 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.944 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 203.8200 100.2800 204.2000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.6168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 201.9900 100.2800 202.3700 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.8598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 293.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 200.1600 100.2800 200.5400 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.0516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.216 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 198.3300 100.2800 198.7100 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.5916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.2748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.936 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 196.5000 100.2800 196.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.552 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 195.2800 100.2800 195.6600 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 193.4500 100.2800 193.8300 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.68 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 191.6200 100.2800 192.0000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 189.7900 100.2800 190.1700 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 187.9600 100.2800 188.3400 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 186.1300 100.2800 186.5100 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.2424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.704 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 184.3000 100.2800 184.6800 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2132 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.352 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 182.4700 100.2800 182.8500 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.4544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 181.2500 100.2800 181.6300 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 179.4200 100.2800 179.8000 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.869 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.32 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 177.5900 100.2800 177.9700 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1542 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.704 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 175.7600 100.2800 176.1400 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.7708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.248 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 173.9300 100.2800 174.3100 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.432 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 172.1000 100.2800 172.4800 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1396 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.5116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.336 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 170.2700 100.2800 170.6500 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.2236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.304 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 168.4400 100.2800 168.8200 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 167.2200 100.2800 167.6000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 165.3900 100.2800 165.7700 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.2166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.096 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 163.5600 100.2800 163.9400 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.7934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.976 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 161.7300 100.2800 162.1100 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 159.9000 100.2800 160.2800 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.0154 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.16 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 157.4600 100.2800 157.8400 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.7506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.664 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 156.2400 100.2800 156.6200 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0346 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.5600 155.0200 100.2800 155.4000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.501 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 19.8316 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.2135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 97.2200 0.0000 97.3600 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.9255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.9648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 85.578 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 452.053 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 0.0000 96.9000 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.443 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.01279 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.6148 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 95.8400 0.0000 95.9800 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.85306 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8162 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 0.0000 95.0600 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.8025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.6588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.0276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 45.7877 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 242.401 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 94.4600 0.0000 94.6000 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.703 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.86242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.0761 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 0.0000 92.7600 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9786 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.667 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.05919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.7623 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.1600 0.0000 92.3000 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7306 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.545 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.58828 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.5603 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.2400 0.0000 91.3800 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.72444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.0822 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.3200 0.0000 90.4600 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.0292 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met4  ;
    ANTENNAMAXAREACAR 37.2137 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.541 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 0.0000 89.5400 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.4246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 43.3395 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.157 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.01366 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 88.9400 0.0000 89.0800 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.2176 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 124.124 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met2  ;
    ANTENNAMAXAREACAR 24.5944 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 113.987 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.528599 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.9496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.672 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 25.1526 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 117.681 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.593756 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 88.0200 0.0000 88.1600 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.3358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 20.4495 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 99.7891 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.505724 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 87.1000 0.0000 87.2400 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.9415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.431 LAYER met2  ;
    ANTENNAMAXAREACAR 19.2939 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.3498 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.492732 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 1.431 LAYER met3  ;
    ANTENNAMAXAREACAR 19.5252 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.9095 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.520685 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.416 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 25.4572 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.886 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 0.0000 86.7800 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.8205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.7195 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.544 LAYER met2  ;
    ANTENNAMAXAREACAR 18.5068 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.3583 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.763522 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAGATEAREA 2.544 LAYER met3  ;
    ANTENNAMAXAREACAR 18.6098 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 87.091 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.6957 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.176 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 27.2569 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.297 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 85.2600 0.0000 85.4000 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met2  ;
    ANTENNAMAXAREACAR 19.4896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.5791 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.506709 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.888 LAYER met3  ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 20.7517 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.7993 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.2646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.352 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 28.5445 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 134.121 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.825288 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 84.8000 0.0000 84.9400 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.0378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.5466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 27.2734 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 129.569 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732304 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 84.3400 0.0000 84.4800 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.405 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 43.8057 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 212.456 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.9902 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.816 LAYER met3  ;
    ANTENNAGATEAREA 4.8075 LAYER met3  ;
    ANTENNAMAXAREACAR 47.5478 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.803 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.598886 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.6057 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.696 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 48.2301 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 236.53 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 83.4200 0.0000 83.5600 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.429 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 25.2132 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 115.517 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.2968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.52 LAYER met3  ;
    ANTENNAGATEAREA 4.0125 LAYER met3  ;
    ANTENNAMAXAREACAR 26.7825 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 124.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.639951 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.1274 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.424 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 28.1312 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 136.332 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.645597 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.5000 0.0000 82.6400 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.7227 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.68847 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 14.6573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 65.4481 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.730398 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.9139 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.888 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 38.8208 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 194.234 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.0400 0.0000 82.1800 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.6436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 97.6800 218.9200 97.8200 219.6400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.455 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 218.9200 96.9000 219.6400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 32.941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 164.479 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.8400 218.9200 95.9800 219.6400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.3076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 218.9200 95.0600 219.6400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.141 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.0000 218.9200 94.1400 219.6400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0637 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.0395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.2634 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 93.5400 218.9200 93.6800 219.6400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.5897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.6695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.897 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.0308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 218.9200 92.7600 219.6400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0786 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.285 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.7000 218.9200 91.8400 219.6400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7209 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.3556 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 90.7800 218.9200 90.9200 219.6400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.7388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 89.8600 218.9200 90.0000 219.6400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0342 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.063 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 218.9200 89.5400 219.6400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.985 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.4800 218.9200 88.6200 219.6400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.7998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 87.1000 218.9200 87.2400 219.6400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.1808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 218.9200 86.7800 219.6400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.785 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 85.7200 218.9200 85.8600 219.6400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 85.2600 218.9200 85.4000 219.6400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.3400 218.9200 84.4800 219.6400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.852 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.4200 218.9200 83.5600 219.6400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.1288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.824 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 82.5000 218.9200 82.6400 219.6400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.819 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.0400 218.9200 82.1800 219.6400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 94.7200 6.9300 ;
        RECT 5.5600 212.0300 94.7200 213.5300 ;
        RECT 5.5600 12.3400 7.0600 12.8200 ;
        RECT 5.5600 17.7800 7.0600 18.2600 ;
        RECT 5.5600 23.2200 7.0600 23.7000 ;
        RECT 5.5600 28.6600 7.0600 29.1400 ;
        RECT 5.5600 34.1000 7.0600 34.5800 ;
        RECT 5.5600 39.5400 7.0600 40.0200 ;
        RECT 5.5600 44.9800 7.0600 45.4600 ;
        RECT 5.5600 50.4200 7.0600 50.9000 ;
        RECT 5.5600 55.8600 7.0600 56.3400 ;
        RECT 5.5600 61.3000 7.0600 61.7800 ;
        RECT 5.5600 66.7400 7.0600 67.2200 ;
        RECT 5.5600 72.1800 7.0600 72.6600 ;
        RECT 5.5600 77.6200 7.0600 78.1000 ;
        RECT 5.5600 83.0600 7.0600 83.5400 ;
        RECT 5.5600 88.5000 7.0600 88.9800 ;
        RECT 5.5600 93.9400 7.0600 94.4200 ;
        RECT 5.5600 99.3800 7.0600 99.8600 ;
        RECT 5.5600 104.8200 7.0600 105.3000 ;
        RECT 93.2200 12.3400 94.7200 12.8200 ;
        RECT 93.2200 17.7800 94.7200 18.2600 ;
        RECT 93.2200 23.2200 94.7200 23.7000 ;
        RECT 93.2200 28.6600 94.7200 29.1400 ;
        RECT 93.2200 34.1000 94.7200 34.5800 ;
        RECT 93.2200 39.5400 94.7200 40.0200 ;
        RECT 93.2200 44.9800 94.7200 45.4600 ;
        RECT 93.2200 50.4200 94.7200 50.9000 ;
        RECT 93.2200 55.8600 94.7200 56.3400 ;
        RECT 93.2200 61.3000 94.7200 61.7800 ;
        RECT 93.2200 66.7400 94.7200 67.2200 ;
        RECT 93.2200 72.1800 94.7200 72.6600 ;
        RECT 93.2200 77.6200 94.7200 78.1000 ;
        RECT 93.2200 83.0600 94.7200 83.5400 ;
        RECT 93.2200 88.5000 94.7200 88.9800 ;
        RECT 93.2200 93.9400 94.7200 94.4200 ;
        RECT 93.2200 99.3800 94.7200 99.8600 ;
        RECT 93.2200 104.8200 94.7200 105.3000 ;
        RECT 5.5600 164.6600 7.0600 165.1400 ;
        RECT 5.5600 110.2600 7.0600 110.7400 ;
        RECT 5.5600 115.7000 7.0600 116.1800 ;
        RECT 5.5600 121.1400 7.0600 121.6200 ;
        RECT 5.5600 126.5800 7.0600 127.0600 ;
        RECT 5.5600 132.0200 7.0600 132.5000 ;
        RECT 5.5600 137.4600 7.0600 137.9400 ;
        RECT 5.5600 142.9000 7.0600 143.3800 ;
        RECT 5.5600 148.3400 7.0600 148.8200 ;
        RECT 5.5600 153.7800 7.0600 154.2600 ;
        RECT 5.5600 159.2200 7.0600 159.7000 ;
        RECT 5.5600 191.8600 7.0600 192.3400 ;
        RECT 5.5600 170.1000 7.0600 170.5800 ;
        RECT 5.5600 175.5400 7.0600 176.0200 ;
        RECT 5.5600 180.9800 7.0600 181.4600 ;
        RECT 5.5600 186.4200 7.0600 186.9000 ;
        RECT 5.5600 197.3000 7.0600 197.7800 ;
        RECT 5.5600 202.7400 7.0600 203.2200 ;
        RECT 5.5600 208.1800 7.0600 208.6600 ;
        RECT 93.2200 164.6600 94.7200 165.1400 ;
        RECT 93.2200 110.2600 94.7200 110.7400 ;
        RECT 93.2200 115.7000 94.7200 116.1800 ;
        RECT 93.2200 121.1400 94.7200 121.6200 ;
        RECT 93.2200 126.5800 94.7200 127.0600 ;
        RECT 93.2200 132.0200 94.7200 132.5000 ;
        RECT 93.2200 137.4600 94.7200 137.9400 ;
        RECT 93.2200 142.9000 94.7200 143.3800 ;
        RECT 93.2200 148.3400 94.7200 148.8200 ;
        RECT 93.2200 153.7800 94.7200 154.2600 ;
        RECT 93.2200 159.2200 94.7200 159.7000 ;
        RECT 93.2200 191.8600 94.7200 192.3400 ;
        RECT 93.2200 170.1000 94.7200 170.5800 ;
        RECT 93.2200 175.5400 94.7200 176.0200 ;
        RECT 93.2200 180.9800 94.7200 181.4600 ;
        RECT 93.2200 186.4200 94.7200 186.9000 ;
        RECT 93.2200 197.3000 94.7200 197.7800 ;
        RECT 93.2200 202.7400 94.7200 203.2200 ;
        RECT 93.2200 208.1800 94.7200 208.6600 ;
      LAYER met4 ;
        RECT 93.2200 5.4300 94.7200 213.5300 ;
        RECT 5.5600 5.4300 7.0600 213.5300 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 3.0600 2.9300 97.2200 4.4300 ;
        RECT 3.0600 214.5300 97.2200 216.0300 ;
        RECT 3.0600 9.6200 4.5600 10.1000 ;
        RECT 3.0600 15.0600 4.5600 15.5400 ;
        RECT 3.0600 20.5000 4.5600 20.9800 ;
        RECT 3.0600 25.9400 4.5600 26.4200 ;
        RECT 3.0600 31.3800 4.5600 31.8600 ;
        RECT 3.0600 36.8200 4.5600 37.3000 ;
        RECT 3.0600 42.2600 4.5600 42.7400 ;
        RECT 3.0600 47.7000 4.5600 48.1800 ;
        RECT 3.0600 53.1400 4.5600 53.6200 ;
        RECT 3.0600 58.5800 4.5600 59.0600 ;
        RECT 3.0600 64.0200 4.5600 64.5000 ;
        RECT 3.0600 69.4600 4.5600 69.9400 ;
        RECT 3.0600 74.9000 4.5600 75.3800 ;
        RECT 3.0600 80.3400 4.5600 80.8200 ;
        RECT 3.0600 85.7800 4.5600 86.2600 ;
        RECT 3.0600 91.2200 4.5600 91.7000 ;
        RECT 3.0600 96.6600 4.5600 97.1400 ;
        RECT 3.0600 102.1000 4.5600 102.5800 ;
        RECT 3.0600 107.5400 4.5600 108.0200 ;
        RECT 95.7200 9.6200 97.2200 10.1000 ;
        RECT 95.7200 15.0600 97.2200 15.5400 ;
        RECT 95.7200 20.5000 97.2200 20.9800 ;
        RECT 95.7200 25.9400 97.2200 26.4200 ;
        RECT 95.7200 31.3800 97.2200 31.8600 ;
        RECT 95.7200 36.8200 97.2200 37.3000 ;
        RECT 95.7200 42.2600 97.2200 42.7400 ;
        RECT 95.7200 47.7000 97.2200 48.1800 ;
        RECT 95.7200 53.1400 97.2200 53.6200 ;
        RECT 95.7200 58.5800 97.2200 59.0600 ;
        RECT 95.7200 64.0200 97.2200 64.5000 ;
        RECT 95.7200 69.4600 97.2200 69.9400 ;
        RECT 95.7200 74.9000 97.2200 75.3800 ;
        RECT 95.7200 80.3400 97.2200 80.8200 ;
        RECT 95.7200 85.7800 97.2200 86.2600 ;
        RECT 95.7200 91.2200 97.2200 91.7000 ;
        RECT 95.7200 96.6600 97.2200 97.1400 ;
        RECT 95.7200 102.1000 97.2200 102.5800 ;
        RECT 95.7200 107.5400 97.2200 108.0200 ;
        RECT 3.0600 112.9800 4.5600 113.4600 ;
        RECT 3.0600 118.4200 4.5600 118.9000 ;
        RECT 3.0600 123.8600 4.5600 124.3400 ;
        RECT 3.0600 129.3000 4.5600 129.7800 ;
        RECT 3.0600 134.7400 4.5600 135.2200 ;
        RECT 3.0600 140.1800 4.5600 140.6600 ;
        RECT 3.0600 145.6200 4.5600 146.1000 ;
        RECT 3.0600 151.0600 4.5600 151.5400 ;
        RECT 3.0600 156.5000 4.5600 156.9800 ;
        RECT 3.0600 161.9400 4.5600 162.4200 ;
        RECT 3.0600 178.2600 4.5600 178.7400 ;
        RECT 3.0600 167.3800 4.5600 167.8600 ;
        RECT 3.0600 172.8200 4.5600 173.3000 ;
        RECT 3.0600 183.7000 4.5600 184.1800 ;
        RECT 3.0600 189.1400 4.5600 189.6200 ;
        RECT 3.0600 205.4600 4.5600 205.9400 ;
        RECT 3.0600 194.5800 4.5600 195.0600 ;
        RECT 3.0600 200.0200 4.5600 200.5000 ;
        RECT 95.7200 112.9800 97.2200 113.4600 ;
        RECT 95.7200 118.4200 97.2200 118.9000 ;
        RECT 95.7200 123.8600 97.2200 124.3400 ;
        RECT 95.7200 129.3000 97.2200 129.7800 ;
        RECT 95.7200 134.7400 97.2200 135.2200 ;
        RECT 95.7200 140.1800 97.2200 140.6600 ;
        RECT 95.7200 145.6200 97.2200 146.1000 ;
        RECT 95.7200 151.0600 97.2200 151.5400 ;
        RECT 95.7200 156.5000 97.2200 156.9800 ;
        RECT 95.7200 161.9400 97.2200 162.4200 ;
        RECT 95.7200 178.2600 97.2200 178.7400 ;
        RECT 95.7200 167.3800 97.2200 167.8600 ;
        RECT 95.7200 172.8200 97.2200 173.3000 ;
        RECT 95.7200 183.7000 97.2200 184.1800 ;
        RECT 95.7200 189.1400 97.2200 189.6200 ;
        RECT 95.7200 205.4600 97.2200 205.9400 ;
        RECT 95.7200 194.5800 97.2200 195.0600 ;
        RECT 95.7200 200.0200 97.2200 200.5000 ;
      LAYER met4 ;
        RECT 95.7200 2.9300 97.2200 216.0300 ;
        RECT 3.0600 2.9300 4.5600 216.0300 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 79.7100 218.7500 100.2800 219.6400 ;
      RECT 78.7900 218.7500 78.9900 219.6400 ;
      RECT 77.8700 218.7500 78.0700 219.6400 ;
      RECT 76.9500 218.7500 77.1500 219.6400 ;
      RECT 75.5700 218.7500 76.2300 219.6400 ;
      RECT 74.6500 218.7500 74.8500 219.6400 ;
      RECT 73.7300 218.7500 73.9300 219.6400 ;
      RECT 72.8100 218.7500 73.0100 219.6400 ;
      RECT 71.4300 218.7500 72.0900 219.6400 ;
      RECT 70.5100 218.7500 70.7100 219.6400 ;
      RECT 69.5900 218.7500 69.7900 219.6400 ;
      RECT 68.2100 218.7500 68.8700 219.6400 ;
      RECT 67.2900 218.7500 67.4900 219.6400 ;
      RECT 66.3700 218.7500 66.5700 219.6400 ;
      RECT 65.4500 218.7500 65.6500 219.6400 ;
      RECT 64.0700 218.7500 64.7300 219.6400 ;
      RECT 63.1500 218.7500 63.3500 219.6400 ;
      RECT 62.2300 218.7500 62.4300 219.6400 ;
      RECT 60.8500 218.7500 61.5100 219.6400 ;
      RECT 59.9300 218.7500 60.1300 219.6400 ;
      RECT 59.0100 218.7500 59.2100 219.6400 ;
      RECT 58.0900 218.7500 58.2900 219.6400 ;
      RECT 56.7100 218.7500 57.3700 219.6400 ;
      RECT 55.7900 218.7500 55.9900 219.6400 ;
      RECT 54.8700 218.7500 55.0700 219.6400 ;
      RECT 53.4900 218.7500 54.1500 219.6400 ;
      RECT 52.5700 218.7500 52.7700 219.6400 ;
      RECT 51.6500 218.7500 51.8500 219.6400 ;
      RECT 50.7300 218.7500 50.9300 219.6400 ;
      RECT 49.3500 218.7500 50.0100 219.6400 ;
      RECT 48.4300 218.7500 48.6300 219.6400 ;
      RECT 47.5100 218.7500 47.7100 219.6400 ;
      RECT 46.1300 218.7500 46.7900 219.6400 ;
      RECT 45.2100 218.7500 45.4100 219.6400 ;
      RECT 44.2900 218.7500 44.4900 219.6400 ;
      RECT 43.3700 218.7500 43.5700 219.6400 ;
      RECT 41.9900 218.7500 42.6500 219.6400 ;
      RECT 41.0700 218.7500 41.2700 219.6400 ;
      RECT 40.1500 218.7500 40.3500 219.6400 ;
      RECT 39.2300 218.7500 39.4300 219.6400 ;
      RECT 37.8500 218.7500 38.5100 219.6400 ;
      RECT 36.9300 218.7500 37.1300 219.6400 ;
      RECT 36.0100 218.7500 36.2100 219.6400 ;
      RECT 34.6300 218.7500 35.2900 219.6400 ;
      RECT 33.7100 218.7500 33.9100 219.6400 ;
      RECT 32.7900 218.7500 32.9900 219.6400 ;
      RECT 31.8700 218.7500 32.0700 219.6400 ;
      RECT 30.4900 218.7500 31.1500 219.6400 ;
      RECT 29.5700 218.7500 29.7700 219.6400 ;
      RECT 28.6500 218.7500 28.8500 219.6400 ;
      RECT 27.2700 218.7500 27.9300 219.6400 ;
      RECT 26.3500 218.7500 26.5500 219.6400 ;
      RECT 25.4300 218.7500 25.6300 219.6400 ;
      RECT 24.5100 218.7500 24.7100 219.6400 ;
      RECT 23.1300 218.7500 23.7900 219.6400 ;
      RECT 22.2100 218.7500 22.4100 219.6400 ;
      RECT 21.2900 218.7500 21.4900 219.6400 ;
      RECT 19.9100 218.7500 20.5700 219.6400 ;
      RECT 18.9900 218.7500 19.1900 219.6400 ;
      RECT 18.0700 218.7500 18.2700 219.6400 ;
      RECT 17.1500 218.7500 17.3500 219.6400 ;
      RECT 15.7700 218.7500 16.4300 219.6400 ;
      RECT 14.8500 218.7500 15.0500 219.6400 ;
      RECT 13.9300 218.7500 14.1300 219.6400 ;
      RECT 12.5500 218.7500 13.2100 219.6400 ;
      RECT 11.6300 218.7500 11.8300 219.6400 ;
      RECT 10.7100 218.7500 10.9100 219.6400 ;
      RECT 9.7900 218.7500 9.9900 219.6400 ;
      RECT 8.4100 218.7500 9.0700 219.6400 ;
      RECT 7.4900 218.7500 7.6900 219.6400 ;
      RECT 6.5700 218.7500 6.7700 219.6400 ;
      RECT 5.6500 218.7500 5.8500 219.6400 ;
      RECT 0.0000 218.7500 4.9300 219.6400 ;
      RECT 0.0000 0.8900 100.2800 218.7500 ;
      RECT 79.7100 0.0000 100.2800 0.8900 ;
      RECT 78.7900 0.0000 78.9900 0.8900 ;
      RECT 77.8700 0.0000 78.0700 0.8900 ;
      RECT 76.9500 0.0000 77.1500 0.8900 ;
      RECT 75.5700 0.0000 76.2300 0.8900 ;
      RECT 74.6500 0.0000 74.8500 0.8900 ;
      RECT 73.7300 0.0000 73.9300 0.8900 ;
      RECT 72.8100 0.0000 73.0100 0.8900 ;
      RECT 71.4300 0.0000 72.0900 0.8900 ;
      RECT 70.5100 0.0000 70.7100 0.8900 ;
      RECT 69.5900 0.0000 69.7900 0.8900 ;
      RECT 68.2100 0.0000 68.8700 0.8900 ;
      RECT 67.2900 0.0000 67.4900 0.8900 ;
      RECT 66.3700 0.0000 66.5700 0.8900 ;
      RECT 65.4500 0.0000 65.6500 0.8900 ;
      RECT 64.0700 0.0000 64.7300 0.8900 ;
      RECT 63.1500 0.0000 63.3500 0.8900 ;
      RECT 62.2300 0.0000 62.4300 0.8900 ;
      RECT 60.8500 0.0000 61.5100 0.8900 ;
      RECT 59.9300 0.0000 60.1300 0.8900 ;
      RECT 59.0100 0.0000 59.2100 0.8900 ;
      RECT 58.0900 0.0000 58.2900 0.8900 ;
      RECT 56.7100 0.0000 57.3700 0.8900 ;
      RECT 55.7900 0.0000 55.9900 0.8900 ;
      RECT 54.8700 0.0000 55.0700 0.8900 ;
      RECT 53.4900 0.0000 54.1500 0.8900 ;
      RECT 52.5700 0.0000 52.7700 0.8900 ;
      RECT 51.6500 0.0000 51.8500 0.8900 ;
      RECT 50.7300 0.0000 50.9300 0.8900 ;
      RECT 49.3500 0.0000 50.0100 0.8900 ;
      RECT 48.4300 0.0000 48.6300 0.8900 ;
      RECT 47.5100 0.0000 47.7100 0.8900 ;
      RECT 46.1300 0.0000 46.7900 0.8900 ;
      RECT 45.2100 0.0000 45.4100 0.8900 ;
      RECT 44.2900 0.0000 44.4900 0.8900 ;
      RECT 43.3700 0.0000 43.5700 0.8900 ;
      RECT 41.9900 0.0000 42.6500 0.8900 ;
      RECT 41.0700 0.0000 41.2700 0.8900 ;
      RECT 40.1500 0.0000 40.3500 0.8900 ;
      RECT 39.2300 0.0000 39.4300 0.8900 ;
      RECT 37.8500 0.0000 38.5100 0.8900 ;
      RECT 36.9300 0.0000 37.1300 0.8900 ;
      RECT 36.0100 0.0000 36.2100 0.8900 ;
      RECT 34.6300 0.0000 35.2900 0.8900 ;
      RECT 33.7100 0.0000 33.9100 0.8900 ;
      RECT 32.7900 0.0000 32.9900 0.8900 ;
      RECT 31.8700 0.0000 32.0700 0.8900 ;
      RECT 30.4900 0.0000 31.1500 0.8900 ;
      RECT 29.5700 0.0000 29.7700 0.8900 ;
      RECT 28.6500 0.0000 28.8500 0.8900 ;
      RECT 27.2700 0.0000 27.9300 0.8900 ;
      RECT 26.3500 0.0000 26.5500 0.8900 ;
      RECT 25.4300 0.0000 25.6300 0.8900 ;
      RECT 24.5100 0.0000 24.7100 0.8900 ;
      RECT 23.1300 0.0000 23.7900 0.8900 ;
      RECT 22.2100 0.0000 22.4100 0.8900 ;
      RECT 21.2900 0.0000 21.4900 0.8900 ;
      RECT 19.9100 0.0000 20.5700 0.8900 ;
      RECT 18.9900 0.0000 19.1900 0.8900 ;
      RECT 18.0700 0.0000 18.2700 0.8900 ;
      RECT 17.1500 0.0000 17.3500 0.8900 ;
      RECT 15.7700 0.0000 16.4300 0.8900 ;
      RECT 14.8500 0.0000 15.0500 0.8900 ;
      RECT 13.9300 0.0000 14.1300 0.8900 ;
      RECT 12.5500 0.0000 13.2100 0.8900 ;
      RECT 11.6300 0.0000 11.8300 0.8900 ;
      RECT 10.7100 0.0000 10.9100 0.8900 ;
      RECT 9.7900 0.0000 9.9900 0.8900 ;
      RECT 8.4100 0.0000 9.0700 0.8900 ;
      RECT 7.4900 0.0000 7.6900 0.8900 ;
      RECT 6.5700 0.0000 6.7700 0.8900 ;
      RECT 5.6500 0.0000 5.8500 0.8900 ;
      RECT 0.0000 0.0000 4.9300 0.8900 ;
    LAYER met1 ;
      RECT 0.0000 150.1000 100.2800 219.6400 ;
      RECT 0.0000 149.7600 99.4200 150.1000 ;
      RECT 0.8600 149.4400 99.4200 149.7600 ;
      RECT 0.8600 149.1000 100.2800 149.4400 ;
      RECT 0.0000 147.7200 100.2800 149.1000 ;
      RECT 0.8600 147.0600 100.2800 147.7200 ;
      RECT 0.0000 146.7000 100.2800 147.0600 ;
      RECT 0.8600 146.0400 100.2800 146.7000 ;
      RECT 0.0000 145.3400 100.2800 146.0400 ;
      RECT 0.8600 144.6800 100.2800 145.3400 ;
      RECT 0.0000 144.6600 100.2800 144.6800 ;
      RECT 0.0000 144.0000 99.4200 144.6600 ;
      RECT 0.0000 143.9800 100.2800 144.0000 ;
      RECT 0.0000 143.3200 99.4200 143.9800 ;
      RECT 0.0000 143.3000 100.2800 143.3200 ;
      RECT 0.8600 142.6400 100.2800 143.3000 ;
      RECT 0.0000 142.2800 100.2800 142.6400 ;
      RECT 0.8600 141.6200 100.2800 142.2800 ;
      RECT 0.0000 140.5800 100.2800 141.6200 ;
      RECT 0.0000 140.2400 99.4200 140.5800 ;
      RECT 0.8600 139.9200 99.4200 140.2400 ;
      RECT 0.8600 139.5800 100.2800 139.9200 ;
      RECT 0.0000 138.8800 100.2800 139.5800 ;
      RECT 0.8600 138.2200 100.2800 138.8800 ;
      RECT 0.0000 138.2000 100.2800 138.2200 ;
      RECT 0.0000 137.8600 99.4200 138.2000 ;
      RECT 0.8600 137.5400 99.4200 137.8600 ;
      RECT 0.8600 137.2000 100.2800 137.5400 ;
      RECT 0.0000 136.5000 100.2800 137.2000 ;
      RECT 0.8600 135.8400 100.2800 136.5000 ;
      RECT 0.0000 135.1400 100.2800 135.8400 ;
      RECT 0.0000 134.8000 99.4200 135.1400 ;
      RECT 0.8600 134.4800 99.4200 134.8000 ;
      RECT 0.8600 134.1400 100.2800 134.4800 ;
      RECT 0.0000 133.4400 100.2800 134.1400 ;
      RECT 0.8600 132.7800 100.2800 133.4400 ;
      RECT 0.0000 132.0800 100.2800 132.7800 ;
      RECT 0.8600 131.4200 99.4200 132.0800 ;
      RECT 0.0000 130.3800 100.2800 131.4200 ;
      RECT 0.8600 129.7200 100.2800 130.3800 ;
      RECT 0.0000 129.3600 100.2800 129.7200 ;
      RECT 0.0000 128.7000 99.4200 129.3600 ;
      RECT 0.0000 128.3400 100.2800 128.7000 ;
      RECT 0.8600 127.6800 100.2800 128.3400 ;
      RECT 0.0000 127.6600 100.2800 127.6800 ;
      RECT 0.8600 127.0000 100.2800 127.6600 ;
      RECT 0.0000 125.9600 100.2800 127.0000 ;
      RECT 0.8600 125.3000 99.4200 125.9600 ;
      RECT 0.0000 124.6000 100.2800 125.3000 ;
      RECT 0.8600 123.9400 100.2800 124.6000 ;
      RECT 0.0000 123.2400 100.2800 123.9400 ;
      RECT 0.8600 122.5800 99.4200 123.2400 ;
      RECT 0.0000 121.8800 100.2800 122.5800 ;
      RECT 0.8600 121.2200 100.2800 121.8800 ;
      RECT 0.0000 120.1800 100.2800 121.2200 ;
      RECT 0.8600 119.5200 99.4200 120.1800 ;
      RECT 0.0000 118.8200 100.2800 119.5200 ;
      RECT 0.8600 118.1600 100.2800 118.8200 ;
      RECT 0.0000 117.4600 100.2800 118.1600 ;
      RECT 0.8600 117.1200 100.2800 117.4600 ;
      RECT 0.8600 116.8000 99.4200 117.1200 ;
      RECT 0.0000 116.4600 99.4200 116.8000 ;
      RECT 0.0000 115.7600 100.2800 116.4600 ;
      RECT 0.8600 115.1000 100.2800 115.7600 ;
      RECT 0.0000 114.4000 100.2800 115.1000 ;
      RECT 0.8600 113.7400 99.4200 114.4000 ;
      RECT 0.0000 113.0400 100.2800 113.7400 ;
      RECT 0.8600 112.3800 100.2800 113.0400 ;
      RECT 0.0000 111.3400 100.2800 112.3800 ;
      RECT 0.8600 110.6800 99.4200 111.3400 ;
      RECT 0.0000 109.9800 100.2800 110.6800 ;
      RECT 0.8600 109.3200 100.2800 109.9800 ;
      RECT 0.0000 108.6200 100.2800 109.3200 ;
      RECT 0.8600 108.2800 100.2800 108.6200 ;
      RECT 0.8600 107.9600 99.4200 108.2800 ;
      RECT 0.0000 107.6200 99.4200 107.9600 ;
      RECT 0.0000 106.9200 100.2800 107.6200 ;
      RECT 0.8600 106.2600 100.2800 106.9200 ;
      RECT 0.0000 105.5600 100.2800 106.2600 ;
      RECT 0.8600 104.9000 99.4200 105.5600 ;
      RECT 0.0000 104.2000 100.2800 104.9000 ;
      RECT 0.8600 103.5400 100.2800 104.2000 ;
      RECT 0.0000 102.5000 100.2800 103.5400 ;
      RECT 0.8600 101.8400 99.4200 102.5000 ;
      RECT 0.0000 101.1400 100.2800 101.8400 ;
      RECT 0.8600 100.4800 100.2800 101.1400 ;
      RECT 0.0000 99.7800 100.2800 100.4800 ;
      RECT 0.8600 99.4400 100.2800 99.7800 ;
      RECT 0.8600 99.1200 99.4200 99.4400 ;
      RECT 0.0000 98.7800 99.4200 99.1200 ;
      RECT 0.0000 98.0800 100.2800 98.7800 ;
      RECT 0.8600 97.4200 100.2800 98.0800 ;
      RECT 0.0000 96.7200 100.2800 97.4200 ;
      RECT 0.8600 96.3800 100.2800 96.7200 ;
      RECT 0.8600 96.0600 99.4200 96.3800 ;
      RECT 0.0000 95.7200 99.4200 96.0600 ;
      RECT 0.0000 95.3600 100.2800 95.7200 ;
      RECT 0.8600 94.7000 100.2800 95.3600 ;
      RECT 0.0000 94.0000 100.2800 94.7000 ;
      RECT 0.8600 93.3400 100.2800 94.0000 ;
      RECT 0.0000 93.3200 100.2800 93.3400 ;
      RECT 0.0000 92.6600 99.4200 93.3200 ;
      RECT 0.0000 92.3000 100.2800 92.6600 ;
      RECT 0.8600 91.6400 100.2800 92.3000 ;
      RECT 0.0000 90.9400 100.2800 91.6400 ;
      RECT 0.8600 90.6000 100.2800 90.9400 ;
      RECT 0.8600 90.2800 99.4200 90.6000 ;
      RECT 0.0000 89.9400 99.4200 90.2800 ;
      RECT 0.0000 89.5800 100.2800 89.9400 ;
      RECT 0.8600 88.9200 100.2800 89.5800 ;
      RECT 0.0000 87.8800 100.2800 88.9200 ;
      RECT 0.8600 87.2200 99.4200 87.8800 ;
      RECT 0.0000 86.5200 100.2800 87.2200 ;
      RECT 0.8600 85.8600 100.2800 86.5200 ;
      RECT 0.0000 85.1600 100.2800 85.8600 ;
      RECT 0.8600 84.8200 100.2800 85.1600 ;
      RECT 0.8600 84.5000 99.4200 84.8200 ;
      RECT 0.0000 84.1600 99.4200 84.5000 ;
      RECT 0.0000 83.4600 100.2800 84.1600 ;
      RECT 0.8600 82.8000 100.2800 83.4600 ;
      RECT 0.0000 82.1000 100.2800 82.8000 ;
      RECT 0.8600 81.4400 100.2800 82.1000 ;
      RECT 0.0000 81.4200 100.2800 81.4400 ;
      RECT 0.0000 80.7600 99.4200 81.4200 ;
      RECT 0.0000 80.7400 100.2800 80.7600 ;
      RECT 0.8600 80.0800 100.2800 80.7400 ;
      RECT 0.0000 79.0400 100.2800 80.0800 ;
      RECT 0.8600 78.7000 100.2800 79.0400 ;
      RECT 0.8600 78.3800 99.4200 78.7000 ;
      RECT 0.0000 78.0400 99.4200 78.3800 ;
      RECT 0.0000 77.6800 100.2800 78.0400 ;
      RECT 0.8600 77.0200 100.2800 77.6800 ;
      RECT 0.0000 76.3200 100.2800 77.0200 ;
      RECT 0.8600 75.6600 100.2800 76.3200 ;
      RECT 0.0000 75.6400 100.2800 75.6600 ;
      RECT 0.0000 74.9800 99.4200 75.6400 ;
      RECT 0.0000 74.6200 100.2800 74.9800 ;
      RECT 0.8600 73.9600 100.2800 74.6200 ;
      RECT 0.0000 73.2600 100.2800 73.9600 ;
      RECT 0.8600 72.6000 100.2800 73.2600 ;
      RECT 0.0000 71.9000 100.2800 72.6000 ;
      RECT 0.8600 71.2400 100.2800 71.9000 ;
      RECT 0.0000 71.2200 100.2800 71.2400 ;
      RECT 0.0000 70.5600 99.4200 71.2200 ;
      RECT 0.0000 70.2000 100.2800 70.5600 ;
      RECT 0.8600 69.5400 100.2800 70.2000 ;
      RECT 0.0000 69.5200 100.2800 69.5400 ;
      RECT 0.8600 68.8600 99.4200 69.5200 ;
      RECT 0.0000 67.8200 100.2800 68.8600 ;
      RECT 0.8600 67.1600 100.2800 67.8200 ;
      RECT 0.0000 67.1400 100.2800 67.1600 ;
      RECT 0.0000 66.4800 99.4200 67.1400 ;
      RECT 0.0000 66.1200 100.2800 66.4800 ;
      RECT 0.8600 65.4600 100.2800 66.1200 ;
      RECT 0.0000 64.7600 100.2800 65.4600 ;
      RECT 0.8600 64.1000 100.2800 64.7600 ;
      RECT 0.0000 63.4000 100.2800 64.1000 ;
      RECT 0.0000 63.0600 99.4200 63.4000 ;
      RECT 0.8600 62.7400 99.4200 63.0600 ;
      RECT 0.8600 62.4000 100.2800 62.7400 ;
      RECT 0.0000 61.7000 100.2800 62.4000 ;
      RECT 0.8600 61.0400 100.2800 61.7000 ;
      RECT 0.0000 60.6800 100.2800 61.0400 ;
      RECT 0.0000 60.0200 99.4200 60.6800 ;
      RECT 0.0000 59.3200 100.2800 60.0200 ;
      RECT 0.8600 58.6600 100.2800 59.3200 ;
      RECT 0.0000 58.6400 100.2800 58.6600 ;
      RECT 0.8600 57.9800 100.2800 58.6400 ;
      RECT 0.0000 57.6200 100.2800 57.9800 ;
      RECT 0.0000 57.2800 99.4200 57.6200 ;
      RECT 0.8600 56.9600 99.4200 57.2800 ;
      RECT 0.8600 56.6200 100.2800 56.9600 ;
      RECT 0.0000 55.5800 100.2800 56.6200 ;
      RECT 0.8600 54.9200 100.2800 55.5800 ;
      RECT 0.0000 54.9000 100.2800 54.9200 ;
      RECT 0.0000 54.2400 99.4200 54.9000 ;
      RECT 0.0000 54.2200 100.2800 54.2400 ;
      RECT 0.8600 53.5600 100.2800 54.2200 ;
      RECT 0.0000 52.8600 100.2800 53.5600 ;
      RECT 0.8600 52.2000 99.4200 52.8600 ;
      RECT 0.0000 51.1600 100.2800 52.2000 ;
      RECT 0.8600 50.5000 100.2800 51.1600 ;
      RECT 0.0000 49.8000 100.2800 50.5000 ;
      RECT 0.8600 49.1400 100.2800 49.8000 ;
      RECT 0.0000 48.7800 100.2800 49.1400 ;
      RECT 0.0000 48.4400 99.4200 48.7800 ;
      RECT 0.8600 48.1200 99.4200 48.4400 ;
      RECT 0.8600 47.7800 100.2800 48.1200 ;
      RECT 0.0000 46.7400 100.2800 47.7800 ;
      RECT 0.8600 46.0800 100.2800 46.7400 ;
      RECT 0.0000 45.7200 100.2800 46.0800 ;
      RECT 0.0000 45.3800 99.4200 45.7200 ;
      RECT 0.8600 45.0600 99.4200 45.3800 ;
      RECT 0.8600 44.7200 100.2800 45.0600 ;
      RECT 0.0000 44.0200 100.2800 44.7200 ;
      RECT 0.8600 43.3600 100.2800 44.0200 ;
      RECT 0.0000 43.0000 100.2800 43.3600 ;
      RECT 0.0000 42.3400 99.4200 43.0000 ;
      RECT 0.0000 42.3200 100.2800 42.3400 ;
      RECT 0.8600 41.6600 100.2800 42.3200 ;
      RECT 0.0000 41.3000 100.2800 41.6600 ;
      RECT 0.0000 40.9600 99.4200 41.3000 ;
      RECT 0.8600 40.6400 99.4200 40.9600 ;
      RECT 0.8600 40.3000 100.2800 40.6400 ;
      RECT 0.0000 39.6000 100.2800 40.3000 ;
      RECT 0.8600 38.9400 100.2800 39.6000 ;
      RECT 0.0000 38.2400 100.2800 38.9400 ;
      RECT 0.8600 37.5800 100.2800 38.2400 ;
      RECT 0.0000 36.8800 100.2800 37.5800 ;
      RECT 0.0000 36.5400 99.4200 36.8800 ;
      RECT 0.8600 36.2200 99.4200 36.5400 ;
      RECT 0.8600 35.8800 100.2800 36.2200 ;
      RECT 0.0000 35.1800 100.2800 35.8800 ;
      RECT 0.8600 34.5200 100.2800 35.1800 ;
      RECT 0.0000 33.8200 100.2800 34.5200 ;
      RECT 0.8600 33.4800 100.2800 33.8200 ;
      RECT 0.8600 33.1600 99.4200 33.4800 ;
      RECT 0.0000 32.8200 99.4200 33.1600 ;
      RECT 0.0000 32.1200 100.2800 32.8200 ;
      RECT 0.8600 31.4600 100.2800 32.1200 ;
      RECT 0.0000 31.1000 100.2800 31.4600 ;
      RECT 0.0000 30.7600 99.4200 31.1000 ;
      RECT 0.8600 30.4400 99.4200 30.7600 ;
      RECT 0.8600 30.1000 100.2800 30.4400 ;
      RECT 0.0000 29.4000 100.2800 30.1000 ;
      RECT 0.8600 28.7400 100.2800 29.4000 ;
      RECT 0.0000 28.0400 100.2800 28.7400 ;
      RECT 0.0000 27.7000 99.4200 28.0400 ;
      RECT 0.8600 27.3800 99.4200 27.7000 ;
      RECT 0.8600 27.0400 100.2800 27.3800 ;
      RECT 0.0000 26.3400 100.2800 27.0400 ;
      RECT 0.8600 25.6800 100.2800 26.3400 ;
      RECT 0.0000 24.9800 100.2800 25.6800 ;
      RECT 0.8600 24.3200 99.4200 24.9800 ;
      RECT 0.0000 23.2800 100.2800 24.3200 ;
      RECT 0.8600 22.6200 100.2800 23.2800 ;
      RECT 0.0000 21.9200 100.2800 22.6200 ;
      RECT 0.8600 21.2600 99.4200 21.9200 ;
      RECT 0.0000 20.5600 100.2800 21.2600 ;
      RECT 0.8600 19.9000 100.2800 20.5600 ;
      RECT 0.0000 19.5400 100.2800 19.9000 ;
      RECT 0.0000 18.8800 99.4200 19.5400 ;
      RECT 0.0000 18.8600 100.2800 18.8800 ;
      RECT 0.8600 18.2000 100.2800 18.8600 ;
      RECT 0.0000 17.5000 100.2800 18.2000 ;
      RECT 0.8600 16.8400 100.2800 17.5000 ;
      RECT 0.0000 16.1400 100.2800 16.8400 ;
      RECT 0.8600 15.4800 99.4200 16.1400 ;
      RECT 0.0000 14.4400 100.2800 15.4800 ;
      RECT 0.8600 13.7800 100.2800 14.4400 ;
      RECT 0.0000 13.0800 100.2800 13.7800 ;
      RECT 0.8600 12.4200 99.4200 13.0800 ;
      RECT 0.0000 11.7200 100.2800 12.4200 ;
      RECT 0.8600 11.0600 100.2800 11.7200 ;
      RECT 0.0000 10.3600 100.2800 11.0600 ;
      RECT 0.8600 9.7000 99.4200 10.3600 ;
      RECT 0.0000 0.0000 100.2800 9.7000 ;
    LAYER met2 ;
      RECT 97.9600 218.7800 100.2800 219.6400 ;
      RECT 97.0400 218.7800 97.5400 219.6400 ;
      RECT 96.1200 218.7800 96.6200 219.6400 ;
      RECT 95.2000 218.7800 95.7000 219.6400 ;
      RECT 94.2800 218.7800 94.7800 219.6400 ;
      RECT 93.8200 218.7800 93.8600 219.6400 ;
      RECT 92.9000 218.7800 93.4000 219.6400 ;
      RECT 91.9800 218.7800 92.4800 219.6400 ;
      RECT 91.0600 218.7800 91.5600 219.6400 ;
      RECT 90.1400 218.7800 90.6400 219.6400 ;
      RECT 89.6800 218.7800 89.7200 219.6400 ;
      RECT 88.7600 218.7800 89.2600 219.6400 ;
      RECT 87.3800 218.7800 88.3400 219.6400 ;
      RECT 86.9200 218.7800 86.9600 219.6400 ;
      RECT 86.0000 218.7800 86.5000 219.6400 ;
      RECT 85.5400 218.7800 85.5800 219.6400 ;
      RECT 84.6200 218.7800 85.1200 219.6400 ;
      RECT 83.7000 218.7800 84.2000 219.6400 ;
      RECT 82.7800 218.7800 83.2800 219.6400 ;
      RECT 82.3200 218.7800 82.3600 219.6400 ;
      RECT 0.0000 218.7800 81.9000 219.6400 ;
      RECT 0.0000 0.8600 100.2800 218.7800 ;
      RECT 97.5000 0.0000 100.2800 0.8600 ;
      RECT 97.0400 0.0000 97.0800 0.8600 ;
      RECT 96.1200 0.0000 96.6200 0.8600 ;
      RECT 95.2000 0.0000 95.7000 0.8600 ;
      RECT 94.7400 0.0000 94.7800 0.8600 ;
      RECT 92.9000 0.0000 94.3200 0.8600 ;
      RECT 92.4400 0.0000 92.4800 0.8600 ;
      RECT 91.5200 0.0000 92.0200 0.8600 ;
      RECT 90.6000 0.0000 91.1000 0.8600 ;
      RECT 89.6800 0.0000 90.1800 0.8600 ;
      RECT 89.2200 0.0000 89.2600 0.8600 ;
      RECT 88.3000 0.0000 88.8000 0.8600 ;
      RECT 87.3800 0.0000 87.8800 0.8600 ;
      RECT 86.9200 0.0000 86.9600 0.8600 ;
      RECT 85.5400 0.0000 86.5000 0.8600 ;
      RECT 85.0800 0.0000 85.1200 0.8600 ;
      RECT 84.6200 0.0000 84.6600 0.8600 ;
      RECT 83.7000 0.0000 84.2000 0.8600 ;
      RECT 82.7800 0.0000 83.2800 0.8600 ;
      RECT 82.3200 0.0000 82.3600 0.8600 ;
      RECT 0.0000 0.0000 81.9000 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 216.3300 100.2800 219.6400 ;
      RECT 97.5200 214.2300 100.2800 216.3300 ;
      RECT 0.0000 214.2300 2.7600 216.3300 ;
      RECT 0.0000 213.8300 100.2800 214.2300 ;
      RECT 95.0200 211.7300 100.2800 213.8300 ;
      RECT 0.0000 211.7300 5.2600 213.8300 ;
      RECT 0.0000 209.9900 100.2800 211.7300 ;
      RECT 1.0200 209.0100 99.2600 209.9900 ;
      RECT 0.0000 208.9600 100.2800 209.0100 ;
      RECT 95.0200 208.1600 100.2800 208.9600 ;
      RECT 0.0000 208.1600 5.2600 208.9600 ;
      RECT 95.0200 207.8800 99.2600 208.1600 ;
      RECT 7.3600 207.8800 92.9200 208.9600 ;
      RECT 1.0200 207.8800 5.2600 208.1600 ;
      RECT 1.0200 207.1800 99.2600 207.8800 ;
      RECT 0.0000 206.3300 100.2800 207.1800 ;
      RECT 1.0200 206.2400 99.2600 206.3300 ;
      RECT 97.5200 205.3500 99.2600 206.2400 ;
      RECT 1.0200 205.3500 2.7600 206.2400 ;
      RECT 97.5200 205.1600 100.2800 205.3500 ;
      RECT 4.8600 205.1600 95.4200 206.2400 ;
      RECT 0.0000 205.1600 2.7600 205.3500 ;
      RECT 0.0000 204.5000 100.2800 205.1600 ;
      RECT 1.0200 203.5200 99.2600 204.5000 ;
      RECT 95.0200 202.6700 100.2800 203.5200 ;
      RECT 0.0000 202.6700 5.2600 203.5200 ;
      RECT 95.0200 202.4400 99.2600 202.6700 ;
      RECT 7.3600 202.4400 92.9200 203.5200 ;
      RECT 1.0200 202.4400 5.2600 202.6700 ;
      RECT 1.0200 201.6900 99.2600 202.4400 ;
      RECT 0.0000 200.8400 100.2800 201.6900 ;
      RECT 1.0200 200.8000 99.2600 200.8400 ;
      RECT 97.5200 199.8600 99.2600 200.8000 ;
      RECT 1.0200 199.8600 2.7600 200.8000 ;
      RECT 97.5200 199.7200 100.2800 199.8600 ;
      RECT 4.8600 199.7200 95.4200 200.8000 ;
      RECT 0.0000 199.7200 2.7600 199.8600 ;
      RECT 0.0000 199.0100 100.2800 199.7200 ;
      RECT 1.0200 198.0800 99.2600 199.0100 ;
      RECT 95.0200 198.0300 99.2600 198.0800 ;
      RECT 1.0200 198.0300 5.2600 198.0800 ;
      RECT 95.0200 197.1800 100.2800 198.0300 ;
      RECT 0.0000 197.1800 5.2600 198.0300 ;
      RECT 95.0200 197.0000 99.2600 197.1800 ;
      RECT 7.3600 197.0000 92.9200 198.0800 ;
      RECT 1.0200 197.0000 5.2600 197.1800 ;
      RECT 1.0200 196.2000 99.2600 197.0000 ;
      RECT 0.0000 195.9600 100.2800 196.2000 ;
      RECT 1.0200 195.3600 99.2600 195.9600 ;
      RECT 97.5200 194.9800 99.2600 195.3600 ;
      RECT 1.0200 194.9800 2.7600 195.3600 ;
      RECT 97.5200 194.2800 100.2800 194.9800 ;
      RECT 4.8600 194.2800 95.4200 195.3600 ;
      RECT 0.0000 194.2800 2.7600 194.9800 ;
      RECT 0.0000 194.1300 100.2800 194.2800 ;
      RECT 1.0200 193.1500 99.2600 194.1300 ;
      RECT 0.0000 192.6400 100.2800 193.1500 ;
      RECT 95.0200 192.3000 100.2800 192.6400 ;
      RECT 0.0000 192.3000 5.2600 192.6400 ;
      RECT 95.0200 191.5600 99.2600 192.3000 ;
      RECT 7.3600 191.5600 92.9200 192.6400 ;
      RECT 1.0200 191.5600 5.2600 192.3000 ;
      RECT 1.0200 191.3200 99.2600 191.5600 ;
      RECT 0.0000 190.4700 100.2800 191.3200 ;
      RECT 1.0200 189.9200 99.2600 190.4700 ;
      RECT 97.5200 189.4900 99.2600 189.9200 ;
      RECT 1.0200 189.4900 2.7600 189.9200 ;
      RECT 97.5200 188.8400 100.2800 189.4900 ;
      RECT 4.8600 188.8400 95.4200 189.9200 ;
      RECT 0.0000 188.8400 2.7600 189.4900 ;
      RECT 0.0000 188.6400 100.2800 188.8400 ;
      RECT 1.0200 187.6600 99.2600 188.6400 ;
      RECT 0.0000 187.2000 100.2800 187.6600 ;
      RECT 95.0200 186.8100 100.2800 187.2000 ;
      RECT 0.0000 186.8100 5.2600 187.2000 ;
      RECT 95.0200 186.1200 99.2600 186.8100 ;
      RECT 7.3600 186.1200 92.9200 187.2000 ;
      RECT 1.0200 186.1200 5.2600 186.8100 ;
      RECT 1.0200 185.8300 99.2600 186.1200 ;
      RECT 0.0000 184.9800 100.2800 185.8300 ;
      RECT 1.0200 184.4800 99.2600 184.9800 ;
      RECT 97.5200 184.0000 99.2600 184.4800 ;
      RECT 1.0200 184.0000 2.7600 184.4800 ;
      RECT 97.5200 183.4000 100.2800 184.0000 ;
      RECT 4.8600 183.4000 95.4200 184.4800 ;
      RECT 0.0000 183.4000 2.7600 184.0000 ;
      RECT 0.0000 183.1500 100.2800 183.4000 ;
      RECT 1.0200 182.1700 99.2600 183.1500 ;
      RECT 0.0000 181.9300 100.2800 182.1700 ;
      RECT 1.0200 181.7600 99.2600 181.9300 ;
      RECT 95.0200 180.9500 99.2600 181.7600 ;
      RECT 1.0200 180.9500 5.2600 181.7600 ;
      RECT 95.0200 180.6800 100.2800 180.9500 ;
      RECT 7.3600 180.6800 92.9200 181.7600 ;
      RECT 0.0000 180.6800 5.2600 180.9500 ;
      RECT 0.0000 180.1000 100.2800 180.6800 ;
      RECT 1.0200 179.1200 99.2600 180.1000 ;
      RECT 0.0000 179.0400 100.2800 179.1200 ;
      RECT 97.5200 178.2700 100.2800 179.0400 ;
      RECT 0.0000 178.2700 2.7600 179.0400 ;
      RECT 97.5200 177.9600 99.2600 178.2700 ;
      RECT 4.8600 177.9600 95.4200 179.0400 ;
      RECT 1.0200 177.9600 2.7600 178.2700 ;
      RECT 1.0200 177.2900 99.2600 177.9600 ;
      RECT 0.0000 176.4400 100.2800 177.2900 ;
      RECT 1.0200 176.3200 99.2600 176.4400 ;
      RECT 95.0200 175.4600 99.2600 176.3200 ;
      RECT 1.0200 175.4600 5.2600 176.3200 ;
      RECT 95.0200 175.2400 100.2800 175.4600 ;
      RECT 7.3600 175.2400 92.9200 176.3200 ;
      RECT 0.0000 175.2400 5.2600 175.4600 ;
      RECT 0.0000 174.6100 100.2800 175.2400 ;
      RECT 1.0200 173.6300 99.2600 174.6100 ;
      RECT 0.0000 173.6000 100.2800 173.6300 ;
      RECT 97.5200 172.7800 100.2800 173.6000 ;
      RECT 0.0000 172.7800 2.7600 173.6000 ;
      RECT 97.5200 172.5200 99.2600 172.7800 ;
      RECT 4.8600 172.5200 95.4200 173.6000 ;
      RECT 1.0200 172.5200 2.7600 172.7800 ;
      RECT 1.0200 171.8000 99.2600 172.5200 ;
      RECT 0.0000 170.9500 100.2800 171.8000 ;
      RECT 1.0200 170.8800 99.2600 170.9500 ;
      RECT 95.0200 169.9700 99.2600 170.8800 ;
      RECT 1.0200 169.9700 5.2600 170.8800 ;
      RECT 95.0200 169.8000 100.2800 169.9700 ;
      RECT 7.3600 169.8000 92.9200 170.8800 ;
      RECT 0.0000 169.8000 5.2600 169.9700 ;
      RECT 0.0000 169.1200 100.2800 169.8000 ;
      RECT 1.0200 168.1600 99.2600 169.1200 ;
      RECT 97.5200 168.1400 99.2600 168.1600 ;
      RECT 1.0200 168.1400 2.7600 168.1600 ;
      RECT 97.5200 167.9000 100.2800 168.1400 ;
      RECT 0.0000 167.9000 2.7600 168.1400 ;
      RECT 97.5200 167.0800 99.2600 167.9000 ;
      RECT 4.8600 167.0800 95.4200 168.1600 ;
      RECT 1.0200 167.0800 2.7600 167.9000 ;
      RECT 1.0200 166.9200 99.2600 167.0800 ;
      RECT 0.0000 166.0700 100.2800 166.9200 ;
      RECT 1.0200 165.4400 99.2600 166.0700 ;
      RECT 95.0200 165.0900 99.2600 165.4400 ;
      RECT 1.0200 165.0900 5.2600 165.4400 ;
      RECT 95.0200 164.3600 100.2800 165.0900 ;
      RECT 7.3600 164.3600 92.9200 165.4400 ;
      RECT 0.0000 164.3600 5.2600 165.0900 ;
      RECT 0.0000 164.2400 100.2800 164.3600 ;
      RECT 1.0200 163.2600 99.2600 164.2400 ;
      RECT 0.0000 162.7200 100.2800 163.2600 ;
      RECT 97.5200 162.4100 100.2800 162.7200 ;
      RECT 0.0000 162.4100 2.7600 162.7200 ;
      RECT 97.5200 161.6400 99.2600 162.4100 ;
      RECT 4.8600 161.6400 95.4200 162.7200 ;
      RECT 1.0200 161.6400 2.7600 162.4100 ;
      RECT 1.0200 161.4300 99.2600 161.6400 ;
      RECT 0.0000 160.5800 100.2800 161.4300 ;
      RECT 1.0200 160.0000 99.2600 160.5800 ;
      RECT 95.0200 159.6000 99.2600 160.0000 ;
      RECT 1.0200 159.6000 5.2600 160.0000 ;
      RECT 95.0200 158.9200 100.2800 159.6000 ;
      RECT 7.3600 158.9200 92.9200 160.0000 ;
      RECT 0.0000 158.9200 5.2600 159.6000 ;
      RECT 0.0000 158.7500 100.2800 158.9200 ;
      RECT 1.0200 158.1400 100.2800 158.7500 ;
      RECT 1.0200 157.7700 99.2600 158.1400 ;
      RECT 0.0000 157.2800 99.2600 157.7700 ;
      RECT 97.5200 157.1600 99.2600 157.2800 ;
      RECT 97.5200 156.9200 100.2800 157.1600 ;
      RECT 0.0000 156.9200 2.7600 157.2800 ;
      RECT 97.5200 156.2000 99.2600 156.9200 ;
      RECT 4.8600 156.2000 95.4200 157.2800 ;
      RECT 1.0200 156.2000 2.7600 156.9200 ;
      RECT 1.0200 155.9400 99.2600 156.2000 ;
      RECT 0.0000 155.7000 100.2800 155.9400 ;
      RECT 1.0200 154.7200 99.2600 155.7000 ;
      RECT 0.0000 154.5600 100.2800 154.7200 ;
      RECT 95.0200 153.4800 100.2800 154.5600 ;
      RECT 7.3600 153.4800 92.9200 154.5600 ;
      RECT 0.0000 153.4800 5.2600 154.5600 ;
      RECT 0.0000 151.8400 100.2800 153.4800 ;
      RECT 97.5200 150.7600 100.2800 151.8400 ;
      RECT 4.8600 150.7600 95.4200 151.8400 ;
      RECT 0.0000 150.7600 2.7600 151.8400 ;
      RECT 0.0000 149.1200 100.2800 150.7600 ;
      RECT 95.0200 148.0400 100.2800 149.1200 ;
      RECT 7.3600 148.0400 92.9200 149.1200 ;
      RECT 0.0000 148.0400 5.2600 149.1200 ;
      RECT 0.0000 146.4000 100.2800 148.0400 ;
      RECT 97.5200 145.3200 100.2800 146.4000 ;
      RECT 4.8600 145.3200 95.4200 146.4000 ;
      RECT 0.0000 145.3200 2.7600 146.4000 ;
      RECT 0.0000 143.6800 100.2800 145.3200 ;
      RECT 95.0200 142.6000 100.2800 143.6800 ;
      RECT 7.3600 142.6000 92.9200 143.6800 ;
      RECT 0.0000 142.6000 5.2600 143.6800 ;
      RECT 0.0000 140.9600 100.2800 142.6000 ;
      RECT 97.5200 139.8800 100.2800 140.9600 ;
      RECT 4.8600 139.8800 95.4200 140.9600 ;
      RECT 0.0000 139.8800 2.7600 140.9600 ;
      RECT 0.0000 138.2400 100.2800 139.8800 ;
      RECT 95.0200 137.1600 100.2800 138.2400 ;
      RECT 7.3600 137.1600 92.9200 138.2400 ;
      RECT 0.0000 137.1600 5.2600 138.2400 ;
      RECT 0.0000 135.5200 100.2800 137.1600 ;
      RECT 97.5200 134.4400 100.2800 135.5200 ;
      RECT 4.8600 134.4400 95.4200 135.5200 ;
      RECT 0.0000 134.4400 2.7600 135.5200 ;
      RECT 0.0000 132.8000 100.2800 134.4400 ;
      RECT 95.0200 131.7200 100.2800 132.8000 ;
      RECT 7.3600 131.7200 92.9200 132.8000 ;
      RECT 0.0000 131.7200 5.2600 132.8000 ;
      RECT 0.0000 130.0800 100.2800 131.7200 ;
      RECT 97.5200 129.0000 100.2800 130.0800 ;
      RECT 4.8600 129.0000 95.4200 130.0800 ;
      RECT 0.0000 129.0000 2.7600 130.0800 ;
      RECT 0.0000 127.3600 100.2800 129.0000 ;
      RECT 95.0200 126.2800 100.2800 127.3600 ;
      RECT 7.3600 126.2800 92.9200 127.3600 ;
      RECT 0.0000 126.2800 5.2600 127.3600 ;
      RECT 0.0000 124.6400 100.2800 126.2800 ;
      RECT 97.5200 123.5600 100.2800 124.6400 ;
      RECT 4.8600 123.5600 95.4200 124.6400 ;
      RECT 0.0000 123.5600 2.7600 124.6400 ;
      RECT 0.0000 121.9200 100.2800 123.5600 ;
      RECT 95.0200 120.8400 100.2800 121.9200 ;
      RECT 7.3600 120.8400 92.9200 121.9200 ;
      RECT 0.0000 120.8400 5.2600 121.9200 ;
      RECT 0.0000 119.2000 100.2800 120.8400 ;
      RECT 97.5200 118.1200 100.2800 119.2000 ;
      RECT 4.8600 118.1200 95.4200 119.2000 ;
      RECT 0.0000 118.1200 2.7600 119.2000 ;
      RECT 0.0000 116.4800 100.2800 118.1200 ;
      RECT 95.0200 115.4000 100.2800 116.4800 ;
      RECT 7.3600 115.4000 92.9200 116.4800 ;
      RECT 0.0000 115.4000 5.2600 116.4800 ;
      RECT 0.0000 113.7600 100.2800 115.4000 ;
      RECT 97.5200 112.6800 100.2800 113.7600 ;
      RECT 4.8600 112.6800 95.4200 113.7600 ;
      RECT 0.0000 112.6800 2.7600 113.7600 ;
      RECT 0.0000 111.0400 100.2800 112.6800 ;
      RECT 95.0200 109.9600 100.2800 111.0400 ;
      RECT 7.3600 109.9600 92.9200 111.0400 ;
      RECT 0.0000 109.9600 5.2600 111.0400 ;
      RECT 0.0000 108.3200 100.2800 109.9600 ;
      RECT 97.5200 107.2400 100.2800 108.3200 ;
      RECT 4.8600 107.2400 95.4200 108.3200 ;
      RECT 0.0000 107.2400 2.7600 108.3200 ;
      RECT 0.0000 105.6000 100.2800 107.2400 ;
      RECT 95.0200 104.5200 100.2800 105.6000 ;
      RECT 7.3600 104.5200 92.9200 105.6000 ;
      RECT 0.0000 104.5200 5.2600 105.6000 ;
      RECT 0.0000 102.8800 100.2800 104.5200 ;
      RECT 97.5200 101.8000 100.2800 102.8800 ;
      RECT 4.8600 101.8000 95.4200 102.8800 ;
      RECT 0.0000 101.8000 2.7600 102.8800 ;
      RECT 0.0000 100.1600 100.2800 101.8000 ;
      RECT 95.0200 99.0800 100.2800 100.1600 ;
      RECT 7.3600 99.0800 92.9200 100.1600 ;
      RECT 0.0000 99.0800 5.2600 100.1600 ;
      RECT 0.0000 97.4400 100.2800 99.0800 ;
      RECT 97.5200 96.3600 100.2800 97.4400 ;
      RECT 4.8600 96.3600 95.4200 97.4400 ;
      RECT 0.0000 96.3600 2.7600 97.4400 ;
      RECT 0.0000 94.7200 100.2800 96.3600 ;
      RECT 95.0200 93.6400 100.2800 94.7200 ;
      RECT 7.3600 93.6400 92.9200 94.7200 ;
      RECT 0.0000 93.6400 5.2600 94.7200 ;
      RECT 0.0000 92.0000 100.2800 93.6400 ;
      RECT 97.5200 90.9200 100.2800 92.0000 ;
      RECT 4.8600 90.9200 95.4200 92.0000 ;
      RECT 0.0000 90.9200 2.7600 92.0000 ;
      RECT 0.0000 89.2800 100.2800 90.9200 ;
      RECT 95.0200 88.2000 100.2800 89.2800 ;
      RECT 7.3600 88.2000 92.9200 89.2800 ;
      RECT 0.0000 88.2000 5.2600 89.2800 ;
      RECT 0.0000 86.5600 100.2800 88.2000 ;
      RECT 97.5200 85.4800 100.2800 86.5600 ;
      RECT 4.8600 85.4800 95.4200 86.5600 ;
      RECT 0.0000 85.4800 2.7600 86.5600 ;
      RECT 0.0000 83.8400 100.2800 85.4800 ;
      RECT 95.0200 82.7600 100.2800 83.8400 ;
      RECT 7.3600 82.7600 92.9200 83.8400 ;
      RECT 0.0000 82.7600 5.2600 83.8400 ;
      RECT 0.0000 81.1200 100.2800 82.7600 ;
      RECT 97.5200 80.0400 100.2800 81.1200 ;
      RECT 4.8600 80.0400 95.4200 81.1200 ;
      RECT 0.0000 80.0400 2.7600 81.1200 ;
      RECT 0.0000 78.4000 100.2800 80.0400 ;
      RECT 95.0200 77.3200 100.2800 78.4000 ;
      RECT 7.3600 77.3200 92.9200 78.4000 ;
      RECT 0.0000 77.3200 5.2600 78.4000 ;
      RECT 0.0000 75.6800 100.2800 77.3200 ;
      RECT 97.5200 74.6000 100.2800 75.6800 ;
      RECT 4.8600 74.6000 95.4200 75.6800 ;
      RECT 0.0000 74.6000 2.7600 75.6800 ;
      RECT 0.0000 72.9600 100.2800 74.6000 ;
      RECT 95.0200 71.8800 100.2800 72.9600 ;
      RECT 7.3600 71.8800 92.9200 72.9600 ;
      RECT 0.0000 71.8800 5.2600 72.9600 ;
      RECT 0.0000 70.2400 100.2800 71.8800 ;
      RECT 97.5200 69.1600 100.2800 70.2400 ;
      RECT 4.8600 69.1600 95.4200 70.2400 ;
      RECT 0.0000 69.1600 2.7600 70.2400 ;
      RECT 0.0000 67.5200 100.2800 69.1600 ;
      RECT 95.0200 66.4400 100.2800 67.5200 ;
      RECT 7.3600 66.4400 92.9200 67.5200 ;
      RECT 0.0000 66.4400 5.2600 67.5200 ;
      RECT 0.0000 64.8000 100.2800 66.4400 ;
      RECT 97.5200 63.7200 100.2800 64.8000 ;
      RECT 4.8600 63.7200 95.4200 64.8000 ;
      RECT 0.0000 63.7200 2.7600 64.8000 ;
      RECT 0.0000 62.0800 100.2800 63.7200 ;
      RECT 95.0200 61.0000 100.2800 62.0800 ;
      RECT 7.3600 61.0000 92.9200 62.0800 ;
      RECT 0.0000 61.0000 5.2600 62.0800 ;
      RECT 0.0000 59.3600 100.2800 61.0000 ;
      RECT 97.5200 58.2800 100.2800 59.3600 ;
      RECT 4.8600 58.2800 95.4200 59.3600 ;
      RECT 0.0000 58.2800 2.7600 59.3600 ;
      RECT 0.0000 56.6400 100.2800 58.2800 ;
      RECT 95.0200 55.5600 100.2800 56.6400 ;
      RECT 7.3600 55.5600 92.9200 56.6400 ;
      RECT 0.0000 55.5600 5.2600 56.6400 ;
      RECT 0.0000 53.9200 100.2800 55.5600 ;
      RECT 97.5200 52.8400 100.2800 53.9200 ;
      RECT 4.8600 52.8400 95.4200 53.9200 ;
      RECT 0.0000 52.8400 2.7600 53.9200 ;
      RECT 0.0000 51.2000 100.2800 52.8400 ;
      RECT 95.0200 50.1200 100.2800 51.2000 ;
      RECT 7.3600 50.1200 92.9200 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 100.2800 50.1200 ;
      RECT 97.5200 47.4000 100.2800 48.4800 ;
      RECT 4.8600 47.4000 95.4200 48.4800 ;
      RECT 0.0000 47.4000 2.7600 48.4800 ;
      RECT 0.0000 45.7600 100.2800 47.4000 ;
      RECT 95.0200 44.6800 100.2800 45.7600 ;
      RECT 7.3600 44.6800 92.9200 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 100.2800 44.6800 ;
      RECT 97.5200 41.9600 100.2800 43.0400 ;
      RECT 4.8600 41.9600 95.4200 43.0400 ;
      RECT 0.0000 41.9600 2.7600 43.0400 ;
      RECT 0.0000 40.3200 100.2800 41.9600 ;
      RECT 95.0200 39.2400 100.2800 40.3200 ;
      RECT 7.3600 39.2400 92.9200 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 100.2800 39.2400 ;
      RECT 97.5200 36.5200 100.2800 37.6000 ;
      RECT 4.8600 36.5200 95.4200 37.6000 ;
      RECT 0.0000 36.5200 2.7600 37.6000 ;
      RECT 0.0000 34.8800 100.2800 36.5200 ;
      RECT 95.0200 33.8000 100.2800 34.8800 ;
      RECT 7.3600 33.8000 92.9200 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 100.2800 33.8000 ;
      RECT 97.5200 31.0800 100.2800 32.1600 ;
      RECT 4.8600 31.0800 95.4200 32.1600 ;
      RECT 0.0000 31.0800 2.7600 32.1600 ;
      RECT 0.0000 29.4400 100.2800 31.0800 ;
      RECT 95.0200 28.3600 100.2800 29.4400 ;
      RECT 7.3600 28.3600 92.9200 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 100.2800 28.3600 ;
      RECT 97.5200 25.6400 100.2800 26.7200 ;
      RECT 4.8600 25.6400 95.4200 26.7200 ;
      RECT 0.0000 25.6400 2.7600 26.7200 ;
      RECT 0.0000 24.0000 100.2800 25.6400 ;
      RECT 95.0200 22.9200 100.2800 24.0000 ;
      RECT 7.3600 22.9200 92.9200 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 100.2800 22.9200 ;
      RECT 97.5200 20.2000 100.2800 21.2800 ;
      RECT 4.8600 20.2000 95.4200 21.2800 ;
      RECT 0.0000 20.2000 2.7600 21.2800 ;
      RECT 0.0000 18.5600 100.2800 20.2000 ;
      RECT 95.0200 17.4800 100.2800 18.5600 ;
      RECT 7.3600 17.4800 92.9200 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 100.2800 17.4800 ;
      RECT 97.5200 14.7600 100.2800 15.8400 ;
      RECT 4.8600 14.7600 95.4200 15.8400 ;
      RECT 0.0000 14.7600 2.7600 15.8400 ;
      RECT 0.0000 13.1200 100.2800 14.7600 ;
      RECT 95.0200 12.0400 100.2800 13.1200 ;
      RECT 7.3600 12.0400 92.9200 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 100.2800 12.0400 ;
      RECT 97.5200 9.3200 100.2800 10.4000 ;
      RECT 4.8600 9.3200 95.4200 10.4000 ;
      RECT 0.0000 9.3200 2.7600 10.4000 ;
      RECT 0.0000 7.2300 100.2800 9.3200 ;
      RECT 95.0200 5.1300 100.2800 7.2300 ;
      RECT 0.0000 5.1300 5.2600 7.2300 ;
      RECT 0.0000 4.7300 100.2800 5.1300 ;
      RECT 97.5200 2.6300 100.2800 4.7300 ;
      RECT 0.0000 2.6300 2.7600 4.7300 ;
      RECT 0.0000 1.0200 100.2800 2.6300 ;
      RECT 81.2200 0.0000 100.2800 1.0200 ;
      RECT 0.0000 0.0000 80.2400 1.0200 ;
    LAYER met4 ;
      RECT 0.0000 216.3300 100.2800 219.6400 ;
      RECT 4.8600 213.8300 95.4200 216.3300 ;
      RECT 95.0200 5.1300 95.4200 213.8300 ;
      RECT 7.3600 5.1300 92.9200 213.8300 ;
      RECT 4.8600 5.1300 5.2600 213.8300 ;
      RECT 97.5200 2.6300 100.2800 216.3300 ;
      RECT 4.8600 2.6300 95.4200 5.1300 ;
      RECT 0.0000 2.6300 2.7600 216.3300 ;
      RECT 0.0000 0.0000 100.2800 2.6300 ;
  END
END RAM_IO

END LIBRARY
