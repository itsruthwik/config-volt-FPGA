##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 00:32:58 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RegFile
  CLASS BLOCK ;
  SIZE 240.1200 BY 219.6400 ;
  FOREIGN RegFile 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.4456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.1505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.392 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 218.9200 14.2200 219.6400 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.712 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 218.9200 12.8400 219.6400 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.104 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 218.9200 11.4600 219.6400 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.8624 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.2345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.928 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 218.9200 10.5400 219.6400 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.358 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 218.9200 25.2600 219.6400 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.856 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 218.9200 23.8800 219.6400 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.46155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.543 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.0692 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.2685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.0548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.096 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 218.9200 22.5000 219.6400 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.1684 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.7275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 218.9200 21.1200 219.6400 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.4128 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.71 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 218.9200 19.7400 219.6400 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.1508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.6765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2209 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.4318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.44 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 218.9200 18.3600 219.6400 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.866 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 218.9200 16.9800 219.6400 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.8856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.31 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 218.9200 15.6000 219.6400 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.512 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 218.9200 35.8400 219.6400 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.5798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 218.9200 34.4600 219.6400 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.118 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 218.9200 33.5400 219.6400 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 218.9200 32.1600 219.6400 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.1 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 218.9200 30.7800 219.6400 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.844 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 218.9200 29.4000 219.6400 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 218.9200 28.0200 219.6400 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.226 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 218.9200 26.6400 219.6400 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 218.9200 57.4600 219.6400 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.2177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.7518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 218.9200 56.5400 219.6400 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.407 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.8288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.0665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.528 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 218.9200 55.1600 219.6400 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.8178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 218.9200 53.7800 219.6400 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 218.9200 52.4000 219.6400 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.9538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 218.9200 51.0200 219.6400 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.6668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.36 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 218.9200 49.6400 219.6400 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 218.9200 48.2600 219.6400 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.2718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 218.9200 46.8800 219.6400 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.8404 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.56 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 218.9200 45.5000 219.6400 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.724 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 218.9200 44.1200 219.6400 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.444 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 218.9200 42.7400 219.6400 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 218.9200 41.3600 219.6400 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.508 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 218.9200 39.9800 219.6400 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.198 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 218.9200 38.6000 219.6400 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 218.9200 37.2200 219.6400 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.2876 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 61.3235 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.8948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.238 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 218.9200 79.5400 219.6400 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0728 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.246 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 218.9200 78.1600 219.6400 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.952 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 218.9200 76.7800 219.6400 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.1516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.416 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 218.9200 75.4000 219.6400 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.65495 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.947 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.7486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 218.9200 74.0200 219.6400 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.6058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.368 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 218.9200 72.6400 219.6400 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.7038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 218.9200 71.2600 219.6400 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 218.9200 69.8800 219.6400 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.7298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.696 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 218.9200 68.5000 219.6400 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 218.9200 67.1200 219.6400 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.2268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.68 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 218.9200 65.7400 219.6400 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.0518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 278.08 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 218.9200 64.3600 219.6400 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.93 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.532 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 218.9200 62.9800 219.6400 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 218.9200 61.6000 219.6400 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.6598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 218.9200 60.2200 219.6400 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 218.9200 58.8400 219.6400 ;
    END
  END NN4BEG[0]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.1633 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 303.296 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 0.0000 14.2200 0.7200 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3412 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.1155 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 0.0000 12.8400 0.7200 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 21.4684 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 107.265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.2265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.3688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.104 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 0.0000 11.4600 0.7200 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9076 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.7775 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.416 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 0.0000 10.5400 0.7200 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.46155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.543 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5624 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.0473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.8295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 23.3677 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 115.145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.2034 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 146.898 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.8398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.616 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 37.0684 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 189.478 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 0.0000 25.2600 0.7200 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.69275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.815 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.1616 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.6225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.16 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.663 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.3846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 50.5847 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.11 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 0.0000 23.8800 0.7200 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.413 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.0624 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 337.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 96.9965 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 517.447 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.284714 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 0.0000 22.5000 0.7200 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.4446 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 355.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 100.021 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 532.023 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315017 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 0.0000 21.1200 0.7200 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.4661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.6405 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.5486 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.113 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 0.0000 19.7400 0.7200 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 80.1456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 428.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 142.948 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 761.694 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 0.0000 18.3600 0.7200 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.0296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 48.6207 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 259.545 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 0.0000 16.9800 0.7200 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.702 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.328 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.186 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4811 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 0.0000 15.6000 0.7200 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.3096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 322.592 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 0.0000 35.8400 0.7200 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 25.4748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 127.152 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.756 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.4789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.6635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 0.0000 34.4600 0.7200 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.13475 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.335 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 21.166 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 105.753 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.3468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 0.0000 33.5400 0.7200 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.4418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.16 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 0.0000 32.1600 0.7200 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.40375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.475 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.778 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.756 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.8633 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.4475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5048 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.8466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.456 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 0.0000 30.7800 0.7200 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5048 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.0434 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.976 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 0.0000 29.4000 0.7200 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.201 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5048 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.4106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.464 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 0.0000 28.0200 0.7200 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.6975 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 0.0000 26.6400 0.7200 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.3088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.69 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.603 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 0.0000 57.4600 0.7200 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.33 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.532 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.2264 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.7374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 0.0000 56.5400 0.7200 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.5058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 34.8481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.156 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 0.0000 55.1600 0.7200 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.4568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 296.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.7314 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.501 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 0.0000 53.7800 0.7200 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3272 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.518 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.78896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.5502 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 0.0000 52.4000 0.7200 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.87051 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.9643 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 0.0000 51.0200 0.7200 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.3828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.6215 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 416.877 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 0.0000 49.6400 0.7200 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.3708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 33.8846 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.962 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 0.0000 48.2600 0.7200 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6273 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.6878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.6139 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.376 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 0.0000 46.8800 0.7200 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.2238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 289.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.708 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.292 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 0.0000 45.5000 0.7200 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.6028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7091 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.74 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 0.0000 44.1200 0.7200 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.1738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 73.303 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 389.195 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 0.0000 42.7400 0.7200 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.8522 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 0.0000 41.3600 0.7200 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.2033 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 311.824 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 0.0000 39.9800 0.7200 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.553 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.4983 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 0.0000 38.6000 0.7200 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 67.7583 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 362.784 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 0.0000 37.2200 0.7200 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.9068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 29.6272 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 156.929 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 0.0000 79.5400 0.7200 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.4588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.176 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 15.8411 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.9017 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 0.0000 78.1600 0.7200 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.2468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.116 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.862 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.0061 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 0.0000 76.7800 0.7200 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.5768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.357 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.954 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 0.0000 75.4000 0.7200 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.0896 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.33 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.6815 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 0.0000 74.0200 0.7200 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.2238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 73.9143 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 392.356 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 0.0000 72.6400 0.7200 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.9068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 28.7568 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.787 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 0.0000 71.2600 0.7200 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.65865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.9051 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 0.0000 69.8800 0.7200 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.4048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7382 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 396.419 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 0.0000 68.5000 0.7200 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.2588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.5394 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 395.034 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 0.0000 67.1200 0.7200 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.866 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.84175 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.8141 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 0.0000 65.7400 0.7200 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.1628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 294.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.0298 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 414.92 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 0.0000 64.3600 0.7200 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.5581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.661 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.9732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 0.0000 62.9800 0.7200 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.4788 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.3165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.12 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 0.0000 61.6000 0.7200 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.6453 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 0.0000 60.2200 0.7200 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.63835 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.751 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.4905 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 0.0000 58.8400 0.7200 ;
    END
  END NN4END[0]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.9988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 84.6400 240.1200 85.0200 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6627 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.5498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 83.2800 240.1200 83.6600 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.2068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.24 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 81.5800 240.1200 81.9600 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.93 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.2046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 80.2200 240.1200 80.6000 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.9858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.728 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 96.5400 240.1200 96.9200 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.955 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 94.8400 240.1200 95.2200 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 93.4800 240.1200 93.8600 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 92.1200 240.1200 92.5000 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 90.4200 240.1200 90.8000 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.449 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 89.0600 240.1200 89.4400 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 194.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 87.7000 240.1200 88.0800 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 86.0000 240.1200 86.3800 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.258 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 108.1000 240.1200 108.4800 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.988 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 106.7400 240.1200 107.1200 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 105.3800 240.1200 105.7600 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 103.6800 240.1200 104.0600 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6333 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 102.3200 240.1200 102.7000 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 100.9600 240.1200 101.3400 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9556 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 99.2600 240.1200 99.6400 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.955 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 97.9000 240.1200 98.2800 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 131.9000 240.1200 132.2800 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 130.2000 240.1200 130.5800 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.0558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.768 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 128.8400 240.1200 129.2200 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.946 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 127.4800 240.1200 127.8600 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.925 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 125.7800 240.1200 126.1600 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 124.4200 240.1200 124.8000 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 123.0600 240.1200 123.4400 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.7258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 121.3600 240.1200 121.7400 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8542 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.104 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 120.0000 240.1200 120.3800 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.15 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 118.6400 240.1200 119.0200 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.705 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 116.9400 240.1200 117.3200 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.171 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 115.5800 240.1200 115.9600 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 114.2200 240.1200 114.6000 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.929 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 112.5200 240.1200 112.9000 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.9664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.584 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 111.1600 240.1200 111.5400 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 109.8000 240.1200 110.1800 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.552 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 149.5800 240.1200 149.9600 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.641 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.88 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 147.8800 240.1200 148.2600 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 146.5200 240.1200 146.9000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.9898 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 145.1600 240.1200 145.5400 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 143.4600 240.1200 143.8400 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.806 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 142.1000 240.1200 142.4800 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 140.7400 240.1200 141.1200 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 139.0400 240.1200 139.4200 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 137.6800 240.1200 138.0600 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.52 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 136.3200 240.1200 136.7000 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.845 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.084 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.8 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 134.6200 240.1200 135.0000 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.565 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 243.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 133.2600 240.1200 133.6400 ;
    END
  END E6BEG[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.6896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0844 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.6257 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.6400 0.7200 85.0200 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0844 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.8672 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.2800 0.7200 83.6600 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.7345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.5800 0.7200 81.9600 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.49 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.2200 0.7200 80.6000 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.8644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 45.5031 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.556 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.5400 0.7200 96.9200 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.577 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.123 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 68.669 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.607 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.8400 0.7200 95.2200 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 10.7896 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 59.6424 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.4800 0.7200 93.8600 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.627 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1254 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 8.44236 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.2855 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.1200 0.7200 92.5000 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.3645 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.5561 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.531 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.4200 0.7200 90.8000 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.0074 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 27.7316 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 147.471 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.0600 0.7200 89.4400 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 20.5698 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.115 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.7000 0.7200 88.0800 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.567 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.29926 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.4929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.0000 0.7200 86.3800 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.0484 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.1000 0.7200 108.4800 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8492 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.7400 0.7200 107.1200 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.3208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.3800 0.7200 105.7600 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 199.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.6800 0.7200 104.0600 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.555 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.71 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9684 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.576 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.3200 0.7200 102.7000 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.0866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 100.9600 0.7200 101.3400 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.323 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.2600 0.7200 99.6400 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6733 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.9000 0.7200 98.2800 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.152 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.7662 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 16.3131 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 91.431 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 131.9000 0.7200 132.2800 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.339 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6523 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 251.345 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.2000 0.7200 130.5800 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.393 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 53.4991 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 285.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.8400 0.7200 129.2200 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.73327 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.2916 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.4800 0.7200 127.8600 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.26364 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.6458 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.7800 0.7200 126.1600 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.591 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.25401 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.8889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.4200 0.7200 124.8000 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.27583 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.83906 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.0600 0.7200 123.4400 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 281.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 6.40552 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 34.4256 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.3600 0.7200 121.7400 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.115 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.6758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 34.1919 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 181.77 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.0000 0.7200 120.3800 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.318 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.53152 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.2828 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.6400 0.7200 119.0200 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.305 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.36404 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.4391 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 116.9400 0.7200 117.3200 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 48.0878 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 238.958 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.5800 0.7200 115.9600 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.2528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.152 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.2200 0.7200 114.6000 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.232 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.5200 0.7200 112.9000 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.1600 0.7200 111.5400 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6463 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.8000 0.7200 110.1800 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.45609 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.9057 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.5800 0.7200 149.9600 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.687 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.43946 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.8162 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 147.8800 0.7200 148.2600 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 66.841 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 356.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 4.89542 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 24.862 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.5200 0.7200 146.9000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.4648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 39.8294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 204.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.1600 0.7200 145.5400 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.735 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.3786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 26.5092 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 141.344 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.4600 0.7200 143.8400 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.122 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 7.40081 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 39.7259 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.1000 0.7200 142.4800 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.852 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.3578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.4303 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 389.688 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.7400 0.7200 141.1200 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.591 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.391 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 47.7273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.43 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.0400 0.7200 139.4200 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.43158 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.7832 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.6800 0.7200 138.0600 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.1928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 14.9259 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.464 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.3200 0.7200 136.7000 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.473 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.4552 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.5216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 298.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.6200 0.7200 135.0000 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.4552 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.2600 0.7200 133.6400 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.9985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.2784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.156 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 0.0000 84.6000 0.7200 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.632 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 0.0000 83.2200 0.7200 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.711 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4775 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.5344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.554 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 0.0000 81.8400 0.7200 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.9738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.664 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 0.0000 80.4600 0.7200 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8124 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.2724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.126 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 0.0000 106.2200 0.7200 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.5998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 0.0000 104.8400 0.7200 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.1164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 0.0000 103.4600 0.7200 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.726 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 0.0000 102.5400 0.7200 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.2628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.952 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 0.0000 101.1600 0.7200 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8424 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 0.0000 99.7800 0.7200 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.4838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.384 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 0.0000 98.4000 0.7200 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.6876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.202 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 0.0000 97.0200 0.7200 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 0.0000 95.6400 0.7200 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 0.0000 94.2600 0.7200 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2073 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.6718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.72 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 0.0000 92.8800 0.7200 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.6468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.116 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 0.0000 91.5000 0.7200 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.1438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.904 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 0.0000 90.1200 0.7200 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.8218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.52 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 0.0000 88.7400 0.7200 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.5032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.398 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 0.0000 87.3600 0.7200 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.1988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 0.0000 85.9800 0.7200 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.3948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 116.62 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 0.0000 127.8400 0.7200 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.222 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 0.0000 126.4600 0.7200 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.4658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 0.0000 125.5400 0.7200 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.3138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.144 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 0.0000 124.1600 0.7200 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 0.0000 122.7800 0.7200 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 0.0000 121.4000 0.7200 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.81 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 0.0000 120.0200 0.7200 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.8798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.496 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 0.0000 118.6400 0.7200 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.798 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 0.0000 117.2600 0.7200 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.9616 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.736 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 0.0000 115.8800 0.7200 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.9128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.672 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 0.0000 114.5000 0.7200 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 0.0000 113.1200 0.7200 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 0.0000 111.7400 0.7200 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.4898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 248.416 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 0.0000 110.3600 0.7200 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3193 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.2218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 0.0000 108.9800 0.7200 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.0148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 251.216 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 0.0000 107.6000 0.7200 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.4942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.353 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 0.0000 149.4600 0.7200 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.0206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.384 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 0.0000 148.5400 0.7200 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.1698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 0.0000 147.1600 0.7200 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.3558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.368 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 0.0000 145.7800 0.7200 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.322 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 0.0000 144.4000 0.7200 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6836 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.01 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 0.0000 143.0200 0.7200 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.1738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 0.0000 141.6400 0.7200 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 0.0000 140.2600 0.7200 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 0.0000 138.8800 0.7200 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.798 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 0.0000 137.5000 0.7200 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 0.0000 136.1200 0.7200 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.9298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.096 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 0.0000 134.7400 0.7200 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 0.0000 133.3600 0.7200 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.9318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.44 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 0.0000 131.9800 0.7200 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 0.0000 130.6000 0.7200 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.8358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.928 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 0.0000 129.2200 0.7200 ;
    END
  END SS4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.0858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.4073 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 218.9200 84.6000 219.6400 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 218.9200 83.2200 219.6400 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.7394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.688 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 218.9200 81.8400 219.6400 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.7231 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 185.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.5322 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.72 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 218.9200 80.4600 219.6400 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.5465 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 345.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 93.8193 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 498.645 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 218.9200 106.2200 219.6400 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.46 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1903 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 101.526 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 539.805 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 218.9200 104.8400 219.6400 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.4688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 44.8411 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 235.626 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 218.9200 103.4600 219.6400 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.8955 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 57.1797 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 304.292 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 218.9200 102.5400 219.6400 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75055 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.883 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7488 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.1044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.844 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 21.9108 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.405 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 218.9200 101.1600 219.6400 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.3236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 49.8097 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.251 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 218.9200 99.7800 219.6400 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.1134 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 52.4457 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.549 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 218.9200 98.4000 219.6400 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.8868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 73.0726 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 389.949 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 218.9200 97.0200 219.6400 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9042 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 218.9200 95.6400 219.6400 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.3684 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 66.7275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8665 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.769 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.416 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 218.9200 94.2600 219.6400 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.9512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 64.6415 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.784 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 218.9200 92.8800 219.6400 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4112 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.9785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.272 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 218.9200 91.5000 219.6400 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.891 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5192 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.3432 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 211.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 218.9200 90.1200 219.6400 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.9215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.3085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via2  ;
    ANTENNADIFFAREA 0.7488 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.5048 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.1196 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 218.9200 88.7400 219.6400 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1964 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8675 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.1444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 218.9200 87.3600 219.6400 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.134 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.1013 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 113.887 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 1.3212 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.6638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5084 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 218.9200 85.9800 219.6400 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.8948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.864 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 398.073 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 218.9200 127.8400 219.6400 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 21.4109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 105.704 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.1864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.13138 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.2673 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 218.9200 126.4600 219.6400 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.1643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.0605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.4758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 29.7208 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.127 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 218.9200 125.5400 219.6400 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.779 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.5596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.4034 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 218.9200 124.1600 219.6400 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.5761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.8835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.0316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.99327 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.7704 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 218.9200 122.7800 219.6400 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.106 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.412 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.66451 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.9279 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 218.9200 121.4000 219.6400 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.1056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.41 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.28458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.1192 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 218.9200 120.0200 219.6400 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.3855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.6618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 276 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.0812 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 218.9200 118.6400 219.6400 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.7228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.5121 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.188 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 218.9200 117.2600 219.6400 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.36 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.682 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.8963 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 218.9200 115.8800 219.6400 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6324 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.044 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.64727 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.9327 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 218.9200 114.5000 219.6400 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2324 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.044 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.96754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.4431 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 218.9200 113.1200 219.6400 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.07 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.6468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 218.9200 111.7400 219.6400 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.86615 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.019 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0578 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.146 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 1.1376 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.1496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.598 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 218.9200 110.3600 219.6400 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.894 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 93.45 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 1.1376 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.6916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.296 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 218.9200 108.9800 219.6400 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.7596 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.2196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 218.9200 107.6000 219.6400 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.7338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.1486 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.171 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 218.9200 149.4600 219.6400 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.8112 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.6825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.166 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.75354 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.2141 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 218.9200 148.5400 219.6400 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.493 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.11071 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.1589 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 218.9200 147.1600 219.6400 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.2908 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.3409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.5335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.1888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 34.4068 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 170.078 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 218.9200 145.7800 219.6400 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.9344 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 64.5575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.912 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.20943 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.3347 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 218.9200 144.4000 219.6400 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.6028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.3601 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 400.809 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 218.9200 143.0200 219.6400 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.5944 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.437 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.0118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.8916 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 121.356 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 218.9200 141.6400 219.6400 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.948 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.65387 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.8747 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 218.9200 140.2600 219.6400 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.5049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.3678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.436 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 375.276 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 218.9200 138.8800 219.6400 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.76 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.16054 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.4081 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 218.9200 137.5000 219.6400 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.3184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 52.3172 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 277.864 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 218.9200 136.1200 219.6400 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.71275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.015 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.438 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.8136 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.6734 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 218.9200 134.7400 219.6400 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.57715 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.679 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.3691 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.512 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 218.9200 133.3600 219.6400 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.82 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 218.9200 131.9800 219.6400 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.9475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.9965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.352 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 218.9200 130.6000 219.6400 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.271 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.7359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.6925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.84 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 218.9200 129.2200 219.6400 ;
    END
  END SS4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.4954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 13.9200 0.7200 14.3000 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.0258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.5600 0.7200 12.9400 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 11.2000 0.7200 11.5800 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.2122 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.8400 0.7200 10.2200 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.8200 0.7200 26.2000 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.4600 0.7200 24.8400 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.7600 0.7200 23.1400 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.4000 0.7200 21.7800 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.0400 0.7200 20.4200 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.925 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.3400 0.7200 18.7200 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.9800 0.7200 17.3600 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.829 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.6200 0.7200 16.0000 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.2896 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.152 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.7200 0.7200 38.1000 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 194.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.0200 0.7200 36.4000 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.7038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.224 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.6600 0.7200 35.0400 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2625 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 47.1228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 251.792 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.3000 0.7200 33.6800 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.6000 0.7200 31.9800 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.2400 0.7200 30.6200 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 28.8800 0.7200 29.2600 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.1800 0.7200 27.5600 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.8334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.1800 0.7200 61.5600 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.5052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.576 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.8200 0.7200 60.2000 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.1200 0.7200 58.5000 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4292 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.7600 0.7200 57.1400 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.4000 0.7200 55.7800 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.7000 0.7200 54.0800 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.3400 0.7200 52.7200 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.293 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 204.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7484 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 50.9800 0.7200 51.3600 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1226 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.387 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.2800 0.7200 49.6600 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.745 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 47.9200 0.7200 48.3000 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.389 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.5600 0.7200 46.9400 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6922 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.353 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.8600 0.7200 45.2400 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.5000 0.7200 43.8800 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0782 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.165 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.1400 0.7200 42.5200 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.759 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.4400 0.7200 40.8200 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.7832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.68 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.0800 0.7200 39.4600 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.5414 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.8600 0.7200 79.2400 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.585 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.384 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.5000 0.7200 77.8800 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 58.8498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 314.336 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.8000 0.7200 76.1800 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 50.362 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 269.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.4400 0.7200 74.8200 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.1874 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 199.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.0800 0.7200 73.4600 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.677 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.3800 0.7200 71.7600 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6446 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.115 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.0200 0.7200 70.4000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.6600 0.7200 69.0400 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 212.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 66.9600 0.7200 67.3400 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.6000 0.7200 65.9800 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.2400 0.7200 64.6200 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9638 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.711 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.5400 0.7200 62.9200 ;
    END
  END W6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.07 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.4955 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 13.9200 240.1200 14.3000 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.07 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2545 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 12.5600 240.1200 12.9400 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.691 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.0936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.44 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 11.2000 240.1200 11.5800 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.1405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.1418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 9.8400 240.1200 10.2200 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.1626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 33.1763 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.966 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 25.8200 240.1200 26.2000 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.4938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 41.4525 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 216.073 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 24.4600 240.1200 24.8400 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.9811 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 34.5508 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.452 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 22.7600 240.1200 23.1400 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.167 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.1985 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.7211 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.221 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 21.4000 240.1200 21.7800 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 261.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.6003 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 79.0823 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 422.141 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 20.0400 240.1200 20.4200 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.541 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.1527 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 211.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.3743 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.993 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 18.3400 240.1200 18.7200 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7632 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.6366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 102.053 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 28.7545 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 141.015 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 16.9800 240.1200 17.3600 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 69.6236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 371.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.1696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.0172 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 128.375 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 15.6200 240.1200 16.0000 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.665 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.8856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 37.7200 240.1200 38.1000 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 36.0200 240.1200 36.4000 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.1256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 34.6600 240.1200 35.0400 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.516 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.044 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 33.3000 240.1200 33.6800 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.4334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 31.6000 240.1200 31.9800 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.616 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3284 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.4597 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 30.2400 240.1200 30.6200 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.5118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 28.8800 240.1200 29.2600 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.2086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 27.1800 240.1200 27.5600 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.2798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 16.0879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 84.2222 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 61.1800 240.1200 61.5600 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.0936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 9.00525 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 48.2983 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 59.8200 240.1200 60.2000 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.5978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.1744 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 288.102 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 58.1200 240.1200 58.5000 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.62721 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.9003 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 56.7600 240.1200 57.1400 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.683 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.09684 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.103 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 55.4000 240.1200 55.7800 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.171 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.87609 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.8404 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 53.7000 240.1200 54.0800 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.837 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.49832 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.9515 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 52.3400 240.1200 52.7200 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.747 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 64.9515 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 341.378 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 50.9800 240.1200 51.3600 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.949 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.83852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8114 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 49.2800 240.1200 49.6600 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.36579 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.398 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 47.9200 240.1200 48.3000 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.886 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.3714 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.729 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.882 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 46.5600 240.1200 46.9400 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.139 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.20054 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.6215 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 44.8600 240.1200 45.2400 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 43.5000 240.1200 43.8800 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.54 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 42.1400 240.1200 42.5200 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.352 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 40.4400 240.1200 40.8200 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 39.0800 240.1200 39.4600 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.1248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.1976 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 95.5987 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 78.8600 240.1200 79.2400 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.8598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.5782 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.9226 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 77.5000 240.1200 77.8800 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.107 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.5029 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.1333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 75.8000 240.1200 76.1800 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.56539 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.4869 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 74.4400 240.1200 74.8200 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 70.51 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 376.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 1.99057 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 10.3347 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 73.0800 240.1200 73.4600 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.567 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.269 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.8489 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219.688 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 71.3800 240.1200 71.7600 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.07098 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.9737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 70.0200 240.1200 70.4000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.422 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.87057 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.9717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 68.6600 240.1200 69.0400 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.503 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.4032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.0015 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.337 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 66.9600 240.1200 67.3400 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.6504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.3727 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 215.626 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 65.6000 240.1200 65.9800 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.2556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.0592 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.6859 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 64.2400 240.1200 64.6200 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0592 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.3571 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 62.5400 240.1200 62.9200 ;
    END
  END W6END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9764 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 6.78902 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 35.324 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 89.5100 0.0000 89.8900 0.7200 ;
    END
  END UserCLK
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.4943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 120.754 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met2  ;
    ANTENNAMAXAREACAR 46.3471 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 226.259 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.319 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.968 LAYER met3  ;
    ANTENNAGATEAREA 1.272 LAYER met3  ;
    ANTENNAMAXAREACAR 49.7425 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.102 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.9397 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.496 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 62.6805 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 329.593 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 209.4200 0.7200 209.8000 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.22 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met2  ;
    ANTENNAMAXAREACAR 13.1994 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.2301 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.412011 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4559 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.368 LAYER met3  ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 13.7051 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 66.966 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.500752 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 66.639 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 357.28 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 61.4242 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.624 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 207.7200 0.7200 208.1000 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 82.7097 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 444.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 82.5453 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 427.162 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 206.0200 0.7200 206.4000 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.179 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 77.4972 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 417.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5599 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.135 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 204.3200 0.7200 204.7000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.6296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.031 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 90.7621 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 472.972 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 202.6200 0.7200 203.0000 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met3  ;
    ANTENNAMAXAREACAR 36.2455 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 179.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.494963 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.2818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.64 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 47.3294 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 239.574 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 200.9200 0.7200 201.3000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.4903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 110.345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.749 LAYER met2  ;
    ANTENNAMAXAREACAR 29.4187 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 141.763 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.48765 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.72 LAYER met3  ;
    ANTENNAGATEAREA 2.067 LAYER met3  ;
    ANTENNAMAXAREACAR 36.2349 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.666 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.594194 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 37.4016 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.055 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.594194 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 198.8800 0.7200 199.2600 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.3164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met3  ;
    ANTENNAMAXAREACAR 73.368 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 371.395 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.752291 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.3741 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.392 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 86.3148 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.942 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 197.1800 0.7200 197.5600 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.7494 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 87.7828 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 452.283 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 195.4800 0.7200 195.8600 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.26 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 82.0392 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 421.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 193.7800 0.7200 194.1600 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.655 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.1495 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 127.392 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 664.848 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 192.0800 0.7200 192.4600 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.271 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 60.8505 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 78.6617 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.728 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 190.0400 0.7200 190.4200 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.1968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 194.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 49.9026 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 246.547 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 188.3400 0.7200 188.7200 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.1248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.6437 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 70.9411 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 370.6 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 186.6400 0.7200 187.0200 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.37 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.2562 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 49.2935 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 253.184 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 184.9400 0.7200 185.3200 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9259 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.4195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.1112 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.0331 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 53.8554 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.699 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 183.2400 0.7200 183.6200 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3185 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.9695 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 22.9247 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.518 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.3579 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.704 LAYER met3  ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 39.7271 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 199.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.625157 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.8418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.96 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 43.2301 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.562 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.987781 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 181.2000 0.7200 181.5800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4725 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.8365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 23.9285 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.414 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 26.2136 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.58 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.2666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.048 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 46.3228 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.394 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 179.5000 0.7200 179.8800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 34.3289 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 164.28 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.4531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.472 LAYER met3  ;
    ANTENNAGATEAREA 1.113 LAYER met3  ;
    ANTENNAMAXAREACAR 67.0641 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 335.602 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.862354 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.0508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.408 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 72.0653 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.443 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.88144 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 177.8000 0.7200 178.1800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.319 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.3853 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 76.9267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 392.55 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 176.1000 0.7200 176.4800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.8697 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 73.6283 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 391.613 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.58113 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 174.4000 0.7200 174.7800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.522 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.5387 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 79.9866 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 402.577 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 172.3600 0.7200 172.7400 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 81.3195 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 428.45 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.793 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.248 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 99.3985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 525.708 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07574 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 170.6600 0.7200 171.0400 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9385 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 58.8887 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 288.563 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.0168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.36 LAYER met3  ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 121.887 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 630.45 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.8037 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.104 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 141.394 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 735.488 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 168.9600 0.7200 169.3400 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.808 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met2  ;
    ANTENNAMAXAREACAR 26.1752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.636164 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 44.8519 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 240.608 LAYER met3  ;
    ANTENNAGATEAREA 2.1735 LAYER met3  ;
    ANTENNAMAXAREACAR 46.811 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.635 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.734756 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.8186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.64 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5286 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 315.539 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 167.2600 0.7200 167.6400 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.378 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.322 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 31.7182 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 152.679 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.3053 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 227.968 LAYER met3  ;
    ANTENNAGATEAREA 1.431 LAYER met3  ;
    ANTENNAMAXAREACAR 61.2817 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.986 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.02383 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.888 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 73.1301 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 376.014 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 165.5600 0.7200 165.9400 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 24.2619 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 116.997 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.7288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.824 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8418 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.5345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.12 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 44.7125 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.836 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 163.5200 0.7200 163.9000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.73 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.263 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 26.4667 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.991 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.2166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.896 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 47.2475 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 240.035 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.8322 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.32 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 65.7795 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 344.46 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.72264 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 161.8200 0.7200 162.2000 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6254 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.816 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met2  ;
    ANTENNAMAXAREACAR 39.5394 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 192.025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.642228 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.1784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.536 LAYER met3  ;
    ANTENNAGATEAREA 1.908 LAYER met3  ;
    ANTENNAMAXAREACAR 53.2597 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 265.681 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.847379 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.933 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.328 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 63.202 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 319.544 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.847379 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 160.1200 0.7200 160.5000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.4926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 44.0891 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 221.33 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.0221 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.328 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 56.1988 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.583 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 158.4200 0.7200 158.8000 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.9868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 60.7524 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 309.425 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.653459 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.4593 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 115.856 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 68.8487 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 353.136 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 156.7200 0.7200 157.1000 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.103 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 87.6024 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.799 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 155.0200 0.7200 155.4000 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 209.4200 240.1200 209.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 207.7200 240.1200 208.1000 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.771 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 206.0200 240.1200 206.4000 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 204.3200 240.1200 204.7000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 202.6200 240.1200 203.0000 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 200.9200 240.1200 201.3000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.8808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.168 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 198.8800 240.1200 199.2600 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 197.1800 240.1200 197.5600 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.52 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 195.4800 240.1200 195.8600 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 193.7800 240.1200 194.1600 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.264 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 192.0800 240.1200 192.4600 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 190.0400 240.1200 190.4200 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 188.3400 240.1200 188.7200 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 186.6400 240.1200 187.0200 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.734 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 184.9400 240.1200 185.3200 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 183.2400 240.1200 183.6200 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 181.2000 240.1200 181.5800 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 179.5000 240.1200 179.8800 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 177.8000 240.1200 178.1800 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4844 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.196 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 176.1000 240.1200 176.4800 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 174.4000 240.1200 174.7800 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 172.3600 240.1200 172.7400 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 170.6600 240.1200 171.0400 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.52 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 168.9600 240.1200 169.3400 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.272 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 167.2600 240.1200 167.6400 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.8728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.792 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 165.5600 240.1200 165.9400 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 163.5200 240.1200 163.9000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 161.8200 240.1200 162.2000 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 160.1200 240.1200 160.5000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 158.4200 240.1200 158.8000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 156.7200 240.1200 157.1000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.491 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.4000 155.0200 240.1200 155.4000 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4446 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.86013 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.9259 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.8000 0.0000 210.1800 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.20391 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.4795 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 206.5800 0.0000 206.9600 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.58 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.92404 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.2256 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 203.8200 0.0000 204.2000 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.3848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 90.9273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 483.822 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 201.0600 0.0000 201.4400 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.989 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.12808 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.3502 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 197.8400 0.0000 198.2200 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.445 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.6606 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 84.4435 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 447.428 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 195.0800 0.0000 195.4600 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.653 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.03758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.8976 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.3200 0.0000 192.7000 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 59.0943 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.9665 LAYER met4  ;
    ANTENNAMAXAREACAR 48.029 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 240.453 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.718099 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 189.5600 0.0000 189.9400 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.6234 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 37.8708 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 183.775 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.720549 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 186.3400 0.0000 186.7200 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.7725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 30.1724 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 144.384 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.621898 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 183.5800 0.0000 183.9600 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.1144 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 47.1611 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 235.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 180.8200 0.0000 181.2000 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.9187 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 33.5587 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 170.077 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.763907 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 178.0600 0.0000 178.4400 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.7186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 79.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 29.5442 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.931 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.710084 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 174.8400 0.0000 175.2200 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.909 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 25.4541 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.0654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 252.88 LAYER met3  ;
    ANTENNAGATEAREA 3.816 LAYER met3  ;
    ANTENNAMAXAREACAR 37.7878 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 185.023 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.690147 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.1386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.68 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 43.491 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 215.618 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.690147 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 172.0800 0.0000 172.4600 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3243 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.2897 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 38.1505 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 193.195 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 169.3200 0.0000 169.7000 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.0915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met2  ;
    ANTENNAMAXAREACAR 25.4381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.261 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.677987 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAGATEAREA 1.272 LAYER met3  ;
    ANTENNAMAXAREACAR 25.5879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 122.412 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.709434 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 61.4955 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 331.264 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 136.255 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 705.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.59686 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 166.5600 0.0000 166.9400 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.8639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.622 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.908 LAYER met2  ;
    ANTENNAMAXAREACAR 28.5672 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 136.962 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.506709 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.553 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.352 LAYER met3  ;
    ANTENNAGATEAREA 4.9665 LAYER met3  ;
    ANTENNAMAXAREACAR 63.493 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 312.557 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.635308 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 64.5197 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.122 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.635308 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 163.3400 0.0000 163.7200 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.3519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 174.996 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.908 LAYER met2  ;
    ANTENNAMAXAREACAR 33.9062 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 163.623 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.485744 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.6463 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.704 LAYER met3  ;
    ANTENNAGATEAREA 3.5355 LAYER met3  ;
    ANTENNAMAXAREACAR 39.4631 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 193.521 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.59747 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.7674 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.504 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 43.5822 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 215.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 160.5800 0.0000 160.9600 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 20.5088 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.1069 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.9784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.68 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 31.4811 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 151.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.7402 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.496 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 37.9497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.217 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.898113 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.8200 0.0000 158.2000 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.9465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met2  ;
    ANTENNAMAXAREACAR 21.0314 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.4406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.496226 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 1.272 LAYER met3  ;
    ANTENNAMAXAREACAR 21.5086 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 102.353 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.824 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 39.69 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 198.483 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590338 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 155.0600 0.0000 155.4400 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.2195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.643 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.5638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.3400 218.9200 209.7200 219.6400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.541 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.8318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.24 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 206.1200 218.9200 206.5000 219.6400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.141 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 203.3600 218.9200 203.7400 219.6400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.927 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 200.1400 218.9200 200.5200 219.6400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.3718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 197.8400 218.9200 198.2200 219.6400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.091 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 195.0800 218.9200 195.4600 219.6400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.9928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 304.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 192.3200 218.9200 192.7000 219.6400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9878 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.831 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.6400 218.9200 189.0200 219.6400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3018 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.401 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.3400 218.9200 186.7200 219.6400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.429 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.5800 218.9200 183.9600 219.6400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3638 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.711 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.8200 218.9200 181.2000 219.6400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.221 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 178.0600 218.9200 178.4400 219.6400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.757 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 175.3000 218.9200 175.6800 219.6400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.617 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 172.0800 218.9200 172.4600 219.6400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.209 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 169.3200 218.9200 169.7000 219.6400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.5600 218.9200 166.9400 219.6400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.559 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.8000 218.9200 164.1800 219.6400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.759 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 160.5800 218.9200 160.9600 219.6400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.604 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 158.2800 218.9200 158.6600 219.6400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.271 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.5200 218.9200 155.9000 219.6400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 234.5600 8.4300 ;
        RECT 5.5600 210.5300 234.5600 213.5300 ;
        RECT 5.5600 12.3400 8.5600 12.8200 ;
        RECT 5.5600 17.7800 8.5600 18.2600 ;
        RECT 55.1200 17.7800 56.1200 18.2600 ;
        RECT 55.1200 12.3400 56.1200 12.8200 ;
        RECT 5.5600 23.2200 8.5600 23.7000 ;
        RECT 5.5600 34.1000 8.5600 34.5800 ;
        RECT 5.5600 28.6600 8.5600 29.1400 ;
        RECT 5.5600 39.5400 8.5600 40.0200 ;
        RECT 5.5600 44.9800 8.5600 45.4600 ;
        RECT 55.1200 34.1000 56.1200 34.5800 ;
        RECT 55.1200 28.6600 56.1200 29.1400 ;
        RECT 55.1200 23.2200 56.1200 23.7000 ;
        RECT 55.1200 44.9800 56.1200 45.4600 ;
        RECT 55.1200 39.5400 56.1200 40.0200 ;
        RECT 100.1200 17.7800 101.1200 18.2600 ;
        RECT 100.1200 12.3400 101.1200 12.8200 ;
        RECT 100.1200 34.1000 101.1200 34.5800 ;
        RECT 100.1200 28.6600 101.1200 29.1400 ;
        RECT 100.1200 23.2200 101.1200 23.7000 ;
        RECT 100.1200 44.9800 101.1200 45.4600 ;
        RECT 100.1200 39.5400 101.1200 40.0200 ;
        RECT 5.5600 55.8600 8.5600 56.3400 ;
        RECT 5.5600 50.4200 8.5600 50.9000 ;
        RECT 5.5600 61.3000 8.5600 61.7800 ;
        RECT 5.5600 72.1800 8.5600 72.6600 ;
        RECT 5.5600 66.7400 8.5600 67.2200 ;
        RECT 5.5600 77.6200 8.5600 78.1000 ;
        RECT 55.1200 61.3000 56.1200 61.7800 ;
        RECT 55.1200 55.8600 56.1200 56.3400 ;
        RECT 55.1200 50.4200 56.1200 50.9000 ;
        RECT 55.1200 77.6200 56.1200 78.1000 ;
        RECT 55.1200 72.1800 56.1200 72.6600 ;
        RECT 55.1200 66.7400 56.1200 67.2200 ;
        RECT 5.5600 83.0600 8.5600 83.5400 ;
        RECT 5.5600 93.9400 8.5600 94.4200 ;
        RECT 5.5600 88.5000 8.5600 88.9800 ;
        RECT 5.5600 99.3800 8.5600 99.8600 ;
        RECT 5.5600 104.8200 8.5600 105.3000 ;
        RECT 55.1200 93.9400 56.1200 94.4200 ;
        RECT 55.1200 88.5000 56.1200 88.9800 ;
        RECT 55.1200 83.0600 56.1200 83.5400 ;
        RECT 55.1200 104.8200 56.1200 105.3000 ;
        RECT 55.1200 99.3800 56.1200 99.8600 ;
        RECT 100.1200 61.3000 101.1200 61.7800 ;
        RECT 100.1200 55.8600 101.1200 56.3400 ;
        RECT 100.1200 50.4200 101.1200 50.9000 ;
        RECT 100.1200 77.6200 101.1200 78.1000 ;
        RECT 100.1200 72.1800 101.1200 72.6600 ;
        RECT 100.1200 66.7400 101.1200 67.2200 ;
        RECT 100.1200 93.9400 101.1200 94.4200 ;
        RECT 100.1200 88.5000 101.1200 88.9800 ;
        RECT 100.1200 83.0600 101.1200 83.5400 ;
        RECT 100.1200 104.8200 101.1200 105.3000 ;
        RECT 100.1200 99.3800 101.1200 99.8600 ;
        RECT 145.1200 17.7800 146.1200 18.2600 ;
        RECT 145.1200 12.3400 146.1200 12.8200 ;
        RECT 145.1200 34.1000 146.1200 34.5800 ;
        RECT 145.1200 28.6600 146.1200 29.1400 ;
        RECT 145.1200 23.2200 146.1200 23.7000 ;
        RECT 145.1200 44.9800 146.1200 45.4600 ;
        RECT 145.1200 39.5400 146.1200 40.0200 ;
        RECT 190.1200 17.7800 191.1200 18.2600 ;
        RECT 190.1200 12.3400 191.1200 12.8200 ;
        RECT 231.5600 17.7800 234.5600 18.2600 ;
        RECT 231.5600 12.3400 234.5600 12.8200 ;
        RECT 190.1200 34.1000 191.1200 34.5800 ;
        RECT 190.1200 28.6600 191.1200 29.1400 ;
        RECT 190.1200 23.2200 191.1200 23.7000 ;
        RECT 190.1200 44.9800 191.1200 45.4600 ;
        RECT 190.1200 39.5400 191.1200 40.0200 ;
        RECT 231.5600 23.2200 234.5600 23.7000 ;
        RECT 231.5600 28.6600 234.5600 29.1400 ;
        RECT 231.5600 34.1000 234.5600 34.5800 ;
        RECT 231.5600 44.9800 234.5600 45.4600 ;
        RECT 231.5600 39.5400 234.5600 40.0200 ;
        RECT 145.1200 61.3000 146.1200 61.7800 ;
        RECT 145.1200 55.8600 146.1200 56.3400 ;
        RECT 145.1200 50.4200 146.1200 50.9000 ;
        RECT 145.1200 77.6200 146.1200 78.1000 ;
        RECT 145.1200 72.1800 146.1200 72.6600 ;
        RECT 145.1200 66.7400 146.1200 67.2200 ;
        RECT 145.1200 93.9400 146.1200 94.4200 ;
        RECT 145.1200 88.5000 146.1200 88.9800 ;
        RECT 145.1200 83.0600 146.1200 83.5400 ;
        RECT 145.1200 104.8200 146.1200 105.3000 ;
        RECT 145.1200 99.3800 146.1200 99.8600 ;
        RECT 190.1200 61.3000 191.1200 61.7800 ;
        RECT 190.1200 55.8600 191.1200 56.3400 ;
        RECT 190.1200 50.4200 191.1200 50.9000 ;
        RECT 190.1200 77.6200 191.1200 78.1000 ;
        RECT 190.1200 72.1800 191.1200 72.6600 ;
        RECT 190.1200 66.7400 191.1200 67.2200 ;
        RECT 231.5600 55.8600 234.5600 56.3400 ;
        RECT 231.5600 50.4200 234.5600 50.9000 ;
        RECT 231.5600 61.3000 234.5600 61.7800 ;
        RECT 231.5600 77.6200 234.5600 78.1000 ;
        RECT 231.5600 72.1800 234.5600 72.6600 ;
        RECT 231.5600 66.7400 234.5600 67.2200 ;
        RECT 190.1200 93.9400 191.1200 94.4200 ;
        RECT 190.1200 88.5000 191.1200 88.9800 ;
        RECT 190.1200 83.0600 191.1200 83.5400 ;
        RECT 190.1200 104.8200 191.1200 105.3000 ;
        RECT 190.1200 99.3800 191.1200 99.8600 ;
        RECT 231.5600 83.0600 234.5600 83.5400 ;
        RECT 231.5600 88.5000 234.5600 88.9800 ;
        RECT 231.5600 93.9400 234.5600 94.4200 ;
        RECT 231.5600 104.8200 234.5600 105.3000 ;
        RECT 231.5600 99.3800 234.5600 99.8600 ;
        RECT 5.5600 115.7000 8.5600 116.1800 ;
        RECT 5.5600 110.2600 8.5600 110.7400 ;
        RECT 5.5600 121.1400 8.5600 121.6200 ;
        RECT 5.5600 132.0200 8.5600 132.5000 ;
        RECT 5.5600 126.5800 8.5600 127.0600 ;
        RECT 5.5600 137.4600 8.5600 137.9400 ;
        RECT 55.1200 121.1400 56.1200 121.6200 ;
        RECT 55.1200 115.7000 56.1200 116.1800 ;
        RECT 55.1200 110.2600 56.1200 110.7400 ;
        RECT 55.1200 137.4600 56.1200 137.9400 ;
        RECT 55.1200 132.0200 56.1200 132.5000 ;
        RECT 55.1200 126.5800 56.1200 127.0600 ;
        RECT 5.5600 142.9000 8.5600 143.3800 ;
        RECT 5.5600 153.7800 8.5600 154.2600 ;
        RECT 5.5600 148.3400 8.5600 148.8200 ;
        RECT 5.5600 159.2200 8.5600 159.7000 ;
        RECT 5.5600 164.6600 8.5600 165.1400 ;
        RECT 55.1200 153.7800 56.1200 154.2600 ;
        RECT 55.1200 148.3400 56.1200 148.8200 ;
        RECT 55.1200 142.9000 56.1200 143.3800 ;
        RECT 55.1200 164.6600 56.1200 165.1400 ;
        RECT 55.1200 159.2200 56.1200 159.7000 ;
        RECT 100.1200 121.1400 101.1200 121.6200 ;
        RECT 100.1200 115.7000 101.1200 116.1800 ;
        RECT 100.1200 110.2600 101.1200 110.7400 ;
        RECT 100.1200 137.4600 101.1200 137.9400 ;
        RECT 100.1200 132.0200 101.1200 132.5000 ;
        RECT 100.1200 126.5800 101.1200 127.0600 ;
        RECT 100.1200 153.7800 101.1200 154.2600 ;
        RECT 100.1200 148.3400 101.1200 148.8200 ;
        RECT 100.1200 142.9000 101.1200 143.3800 ;
        RECT 100.1200 164.6600 101.1200 165.1400 ;
        RECT 100.1200 159.2200 101.1200 159.7000 ;
        RECT 5.5600 175.5400 8.5600 176.0200 ;
        RECT 5.5600 170.1000 8.5600 170.5800 ;
        RECT 5.5600 180.9800 8.5600 181.4600 ;
        RECT 5.5600 191.8600 8.5600 192.3400 ;
        RECT 5.5600 186.4200 8.5600 186.9000 ;
        RECT 5.5600 197.3000 8.5600 197.7800 ;
        RECT 55.1200 180.9800 56.1200 181.4600 ;
        RECT 55.1200 175.5400 56.1200 176.0200 ;
        RECT 55.1200 170.1000 56.1200 170.5800 ;
        RECT 55.1200 197.3000 56.1200 197.7800 ;
        RECT 55.1200 191.8600 56.1200 192.3400 ;
        RECT 55.1200 186.4200 56.1200 186.9000 ;
        RECT 5.5600 202.7400 8.5600 203.2200 ;
        RECT 5.5600 208.1800 8.5600 208.6600 ;
        RECT 55.1200 208.1800 56.1200 208.6600 ;
        RECT 55.1200 202.7400 56.1200 203.2200 ;
        RECT 100.1200 180.9800 101.1200 181.4600 ;
        RECT 100.1200 175.5400 101.1200 176.0200 ;
        RECT 100.1200 170.1000 101.1200 170.5800 ;
        RECT 100.1200 197.3000 101.1200 197.7800 ;
        RECT 100.1200 191.8600 101.1200 192.3400 ;
        RECT 100.1200 186.4200 101.1200 186.9000 ;
        RECT 100.1200 208.1800 101.1200 208.6600 ;
        RECT 100.1200 202.7400 101.1200 203.2200 ;
        RECT 145.1200 121.1400 146.1200 121.6200 ;
        RECT 145.1200 115.7000 146.1200 116.1800 ;
        RECT 145.1200 110.2600 146.1200 110.7400 ;
        RECT 145.1200 137.4600 146.1200 137.9400 ;
        RECT 145.1200 132.0200 146.1200 132.5000 ;
        RECT 145.1200 126.5800 146.1200 127.0600 ;
        RECT 145.1200 153.7800 146.1200 154.2600 ;
        RECT 145.1200 148.3400 146.1200 148.8200 ;
        RECT 145.1200 142.9000 146.1200 143.3800 ;
        RECT 145.1200 164.6600 146.1200 165.1400 ;
        RECT 145.1200 159.2200 146.1200 159.7000 ;
        RECT 190.1200 121.1400 191.1200 121.6200 ;
        RECT 190.1200 115.7000 191.1200 116.1800 ;
        RECT 190.1200 110.2600 191.1200 110.7400 ;
        RECT 190.1200 137.4600 191.1200 137.9400 ;
        RECT 190.1200 132.0200 191.1200 132.5000 ;
        RECT 190.1200 126.5800 191.1200 127.0600 ;
        RECT 231.5600 115.7000 234.5600 116.1800 ;
        RECT 231.5600 110.2600 234.5600 110.7400 ;
        RECT 231.5600 121.1400 234.5600 121.6200 ;
        RECT 231.5600 137.4600 234.5600 137.9400 ;
        RECT 231.5600 132.0200 234.5600 132.5000 ;
        RECT 231.5600 126.5800 234.5600 127.0600 ;
        RECT 190.1200 153.7800 191.1200 154.2600 ;
        RECT 190.1200 148.3400 191.1200 148.8200 ;
        RECT 190.1200 142.9000 191.1200 143.3800 ;
        RECT 190.1200 164.6600 191.1200 165.1400 ;
        RECT 190.1200 159.2200 191.1200 159.7000 ;
        RECT 231.5600 142.9000 234.5600 143.3800 ;
        RECT 231.5600 148.3400 234.5600 148.8200 ;
        RECT 231.5600 153.7800 234.5600 154.2600 ;
        RECT 231.5600 164.6600 234.5600 165.1400 ;
        RECT 231.5600 159.2200 234.5600 159.7000 ;
        RECT 145.1200 180.9800 146.1200 181.4600 ;
        RECT 145.1200 175.5400 146.1200 176.0200 ;
        RECT 145.1200 170.1000 146.1200 170.5800 ;
        RECT 145.1200 197.3000 146.1200 197.7800 ;
        RECT 145.1200 191.8600 146.1200 192.3400 ;
        RECT 145.1200 186.4200 146.1200 186.9000 ;
        RECT 145.1200 208.1800 146.1200 208.6600 ;
        RECT 145.1200 202.7400 146.1200 203.2200 ;
        RECT 190.1200 180.9800 191.1200 181.4600 ;
        RECT 190.1200 175.5400 191.1200 176.0200 ;
        RECT 190.1200 170.1000 191.1200 170.5800 ;
        RECT 190.1200 197.3000 191.1200 197.7800 ;
        RECT 190.1200 191.8600 191.1200 192.3400 ;
        RECT 190.1200 186.4200 191.1200 186.9000 ;
        RECT 231.5600 175.5400 234.5600 176.0200 ;
        RECT 231.5600 170.1000 234.5600 170.5800 ;
        RECT 231.5600 180.9800 234.5600 181.4600 ;
        RECT 231.5600 197.3000 234.5600 197.7800 ;
        RECT 231.5600 191.8600 234.5600 192.3400 ;
        RECT 231.5600 186.4200 234.5600 186.9000 ;
        RECT 190.1200 208.1800 191.1200 208.6600 ;
        RECT 190.1200 202.7400 191.1200 203.2200 ;
        RECT 231.5600 208.1800 234.5600 208.6600 ;
        RECT 231.5600 202.7400 234.5600 203.2200 ;
      LAYER met4 ;
        RECT 5.5600 5.4300 8.5600 213.5300 ;
        RECT 231.5600 5.4300 234.5600 213.5300 ;
        RECT 55.1200 5.4300 56.1200 213.5300 ;
        RECT 100.1200 5.4300 101.1200 213.5300 ;
        RECT 145.1200 5.4300 146.1200 213.5300 ;
        RECT 190.1200 5.4300 191.1200 213.5300 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 1.5600 1.4300 238.5600 4.4300 ;
        RECT 1.5600 214.5300 238.5600 217.5300 ;
        RECT 12.3200 9.6200 13.3200 10.1000 ;
        RECT 1.5600 9.6200 4.5600 10.1000 ;
        RECT 12.3200 15.0600 13.3200 15.5400 ;
        RECT 1.5600 15.0600 4.5600 15.5400 ;
        RECT 57.3200 15.0600 58.3200 15.5400 ;
        RECT 57.3200 9.6200 58.3200 10.1000 ;
        RECT 1.5600 20.5000 4.5600 20.9800 ;
        RECT 1.5600 25.9400 4.5600 26.4200 ;
        RECT 12.3200 20.5000 13.3200 20.9800 ;
        RECT 12.3200 25.9400 13.3200 26.4200 ;
        RECT 12.3200 31.3800 13.3200 31.8600 ;
        RECT 1.5600 31.3800 4.5600 31.8600 ;
        RECT 12.3200 42.2600 13.3200 42.7400 ;
        RECT 1.5600 42.2600 4.5600 42.7400 ;
        RECT 12.3200 36.8200 13.3200 37.3000 ;
        RECT 1.5600 36.8200 4.5600 37.3000 ;
        RECT 12.3200 47.7000 13.3200 48.1800 ;
        RECT 1.5600 47.7000 4.5600 48.1800 ;
        RECT 57.3200 31.3800 58.3200 31.8600 ;
        RECT 57.3200 25.9400 58.3200 26.4200 ;
        RECT 57.3200 20.5000 58.3200 20.9800 ;
        RECT 57.3200 47.7000 58.3200 48.1800 ;
        RECT 57.3200 42.2600 58.3200 42.7400 ;
        RECT 57.3200 36.8200 58.3200 37.3000 ;
        RECT 102.3200 15.0600 103.3200 15.5400 ;
        RECT 102.3200 9.6200 103.3200 10.1000 ;
        RECT 102.3200 31.3800 103.3200 31.8600 ;
        RECT 102.3200 25.9400 103.3200 26.4200 ;
        RECT 102.3200 20.5000 103.3200 20.9800 ;
        RECT 102.3200 47.7000 103.3200 48.1800 ;
        RECT 102.3200 42.2600 103.3200 42.7400 ;
        RECT 102.3200 36.8200 103.3200 37.3000 ;
        RECT 12.3200 53.1400 13.3200 53.6200 ;
        RECT 1.5600 53.1400 4.5600 53.6200 ;
        RECT 1.5600 58.5800 4.5600 59.0600 ;
        RECT 1.5600 64.0200 4.5600 64.5000 ;
        RECT 12.3200 58.5800 13.3200 59.0600 ;
        RECT 12.3200 64.0200 13.3200 64.5000 ;
        RECT 12.3200 69.4600 13.3200 69.9400 ;
        RECT 1.5600 69.4600 4.5600 69.9400 ;
        RECT 12.3200 74.9000 13.3200 75.3800 ;
        RECT 1.5600 74.9000 4.5600 75.3800 ;
        RECT 57.3200 64.0200 58.3200 64.5000 ;
        RECT 57.3200 58.5800 58.3200 59.0600 ;
        RECT 57.3200 53.1400 58.3200 53.6200 ;
        RECT 57.3200 74.9000 58.3200 75.3800 ;
        RECT 57.3200 69.4600 58.3200 69.9400 ;
        RECT 1.5600 80.3400 4.5600 80.8200 ;
        RECT 1.5600 85.7800 4.5600 86.2600 ;
        RECT 12.3200 80.3400 13.3200 80.8200 ;
        RECT 12.3200 85.7800 13.3200 86.2600 ;
        RECT 12.3200 91.2200 13.3200 91.7000 ;
        RECT 1.5600 91.2200 4.5600 91.7000 ;
        RECT 12.3200 102.1000 13.3200 102.5800 ;
        RECT 1.5600 102.1000 4.5600 102.5800 ;
        RECT 12.3200 96.6600 13.3200 97.1400 ;
        RECT 1.5600 96.6600 4.5600 97.1400 ;
        RECT 12.3200 107.5400 13.3200 108.0200 ;
        RECT 1.5600 107.5400 4.5600 108.0200 ;
        RECT 57.3200 91.2200 58.3200 91.7000 ;
        RECT 57.3200 85.7800 58.3200 86.2600 ;
        RECT 57.3200 80.3400 58.3200 80.8200 ;
        RECT 57.3200 107.5400 58.3200 108.0200 ;
        RECT 57.3200 102.1000 58.3200 102.5800 ;
        RECT 57.3200 96.6600 58.3200 97.1400 ;
        RECT 102.3200 64.0200 103.3200 64.5000 ;
        RECT 102.3200 58.5800 103.3200 59.0600 ;
        RECT 102.3200 53.1400 103.3200 53.6200 ;
        RECT 102.3200 74.9000 103.3200 75.3800 ;
        RECT 102.3200 69.4600 103.3200 69.9400 ;
        RECT 102.3200 91.2200 103.3200 91.7000 ;
        RECT 102.3200 85.7800 103.3200 86.2600 ;
        RECT 102.3200 80.3400 103.3200 80.8200 ;
        RECT 102.3200 107.5400 103.3200 108.0200 ;
        RECT 102.3200 102.1000 103.3200 102.5800 ;
        RECT 102.3200 96.6600 103.3200 97.1400 ;
        RECT 147.3200 15.0600 148.3200 15.5400 ;
        RECT 147.3200 9.6200 148.3200 10.1000 ;
        RECT 147.3200 31.3800 148.3200 31.8600 ;
        RECT 147.3200 25.9400 148.3200 26.4200 ;
        RECT 147.3200 20.5000 148.3200 20.9800 ;
        RECT 147.3200 47.7000 148.3200 48.1800 ;
        RECT 147.3200 42.2600 148.3200 42.7400 ;
        RECT 147.3200 36.8200 148.3200 37.3000 ;
        RECT 192.3200 15.0600 193.3200 15.5400 ;
        RECT 192.3200 9.6200 193.3200 10.1000 ;
        RECT 235.5600 15.0600 238.5600 15.5400 ;
        RECT 235.5600 9.6200 238.5600 10.1000 ;
        RECT 192.3200 31.3800 193.3200 31.8600 ;
        RECT 192.3200 25.9400 193.3200 26.4200 ;
        RECT 192.3200 20.5000 193.3200 20.9800 ;
        RECT 192.3200 47.7000 193.3200 48.1800 ;
        RECT 192.3200 42.2600 193.3200 42.7400 ;
        RECT 192.3200 36.8200 193.3200 37.3000 ;
        RECT 235.5600 25.9400 238.5600 26.4200 ;
        RECT 235.5600 20.5000 238.5600 20.9800 ;
        RECT 235.5600 31.3800 238.5600 31.8600 ;
        RECT 235.5600 47.7000 238.5600 48.1800 ;
        RECT 235.5600 42.2600 238.5600 42.7400 ;
        RECT 235.5600 36.8200 238.5600 37.3000 ;
        RECT 147.3200 64.0200 148.3200 64.5000 ;
        RECT 147.3200 58.5800 148.3200 59.0600 ;
        RECT 147.3200 53.1400 148.3200 53.6200 ;
        RECT 147.3200 74.9000 148.3200 75.3800 ;
        RECT 147.3200 69.4600 148.3200 69.9400 ;
        RECT 147.3200 91.2200 148.3200 91.7000 ;
        RECT 147.3200 85.7800 148.3200 86.2600 ;
        RECT 147.3200 80.3400 148.3200 80.8200 ;
        RECT 147.3200 107.5400 148.3200 108.0200 ;
        RECT 147.3200 102.1000 148.3200 102.5800 ;
        RECT 147.3200 96.6600 148.3200 97.1400 ;
        RECT 192.3200 64.0200 193.3200 64.5000 ;
        RECT 192.3200 58.5800 193.3200 59.0600 ;
        RECT 192.3200 53.1400 193.3200 53.6200 ;
        RECT 192.3200 74.9000 193.3200 75.3800 ;
        RECT 192.3200 69.4600 193.3200 69.9400 ;
        RECT 235.5600 53.1400 238.5600 53.6200 ;
        RECT 235.5600 64.0200 238.5600 64.5000 ;
        RECT 235.5600 58.5800 238.5600 59.0600 ;
        RECT 235.5600 74.9000 238.5600 75.3800 ;
        RECT 235.5600 69.4600 238.5600 69.9400 ;
        RECT 192.3200 91.2200 193.3200 91.7000 ;
        RECT 192.3200 85.7800 193.3200 86.2600 ;
        RECT 192.3200 80.3400 193.3200 80.8200 ;
        RECT 192.3200 107.5400 193.3200 108.0200 ;
        RECT 192.3200 102.1000 193.3200 102.5800 ;
        RECT 192.3200 96.6600 193.3200 97.1400 ;
        RECT 235.5600 85.7800 238.5600 86.2600 ;
        RECT 235.5600 80.3400 238.5600 80.8200 ;
        RECT 235.5600 91.2200 238.5600 91.7000 ;
        RECT 235.5600 107.5400 238.5600 108.0200 ;
        RECT 235.5600 102.1000 238.5600 102.5800 ;
        RECT 235.5600 96.6600 238.5600 97.1400 ;
        RECT 12.3200 112.9800 13.3200 113.4600 ;
        RECT 1.5600 112.9800 4.5600 113.4600 ;
        RECT 1.5600 118.4200 4.5600 118.9000 ;
        RECT 1.5600 123.8600 4.5600 124.3400 ;
        RECT 12.3200 118.4200 13.3200 118.9000 ;
        RECT 12.3200 123.8600 13.3200 124.3400 ;
        RECT 12.3200 129.3000 13.3200 129.7800 ;
        RECT 1.5600 129.3000 4.5600 129.7800 ;
        RECT 12.3200 134.7400 13.3200 135.2200 ;
        RECT 1.5600 134.7400 4.5600 135.2200 ;
        RECT 57.3200 123.8600 58.3200 124.3400 ;
        RECT 57.3200 118.4200 58.3200 118.9000 ;
        RECT 57.3200 112.9800 58.3200 113.4600 ;
        RECT 57.3200 134.7400 58.3200 135.2200 ;
        RECT 57.3200 129.3000 58.3200 129.7800 ;
        RECT 1.5600 140.1800 4.5600 140.6600 ;
        RECT 1.5600 145.6200 4.5600 146.1000 ;
        RECT 12.3200 140.1800 13.3200 140.6600 ;
        RECT 12.3200 145.6200 13.3200 146.1000 ;
        RECT 12.3200 151.0600 13.3200 151.5400 ;
        RECT 1.5600 151.0600 4.5600 151.5400 ;
        RECT 12.3200 161.9400 13.3200 162.4200 ;
        RECT 1.5600 161.9400 4.5600 162.4200 ;
        RECT 12.3200 156.5000 13.3200 156.9800 ;
        RECT 1.5600 156.5000 4.5600 156.9800 ;
        RECT 12.3200 167.3800 13.3200 167.8600 ;
        RECT 1.5600 167.3800 4.5600 167.8600 ;
        RECT 57.3200 151.0600 58.3200 151.5400 ;
        RECT 57.3200 145.6200 58.3200 146.1000 ;
        RECT 57.3200 140.1800 58.3200 140.6600 ;
        RECT 57.3200 167.3800 58.3200 167.8600 ;
        RECT 57.3200 161.9400 58.3200 162.4200 ;
        RECT 57.3200 156.5000 58.3200 156.9800 ;
        RECT 102.3200 123.8600 103.3200 124.3400 ;
        RECT 102.3200 118.4200 103.3200 118.9000 ;
        RECT 102.3200 112.9800 103.3200 113.4600 ;
        RECT 102.3200 134.7400 103.3200 135.2200 ;
        RECT 102.3200 129.3000 103.3200 129.7800 ;
        RECT 102.3200 151.0600 103.3200 151.5400 ;
        RECT 102.3200 145.6200 103.3200 146.1000 ;
        RECT 102.3200 140.1800 103.3200 140.6600 ;
        RECT 102.3200 167.3800 103.3200 167.8600 ;
        RECT 102.3200 161.9400 103.3200 162.4200 ;
        RECT 102.3200 156.5000 103.3200 156.9800 ;
        RECT 12.3200 172.8200 13.3200 173.3000 ;
        RECT 1.5600 172.8200 4.5600 173.3000 ;
        RECT 1.5600 178.2600 4.5600 178.7400 ;
        RECT 1.5600 183.7000 4.5600 184.1800 ;
        RECT 12.3200 178.2600 13.3200 178.7400 ;
        RECT 12.3200 183.7000 13.3200 184.1800 ;
        RECT 12.3200 189.1400 13.3200 189.6200 ;
        RECT 1.5600 189.1400 4.5600 189.6200 ;
        RECT 12.3200 194.5800 13.3200 195.0600 ;
        RECT 1.5600 194.5800 4.5600 195.0600 ;
        RECT 57.3200 183.7000 58.3200 184.1800 ;
        RECT 57.3200 178.2600 58.3200 178.7400 ;
        RECT 57.3200 172.8200 58.3200 173.3000 ;
        RECT 57.3200 194.5800 58.3200 195.0600 ;
        RECT 57.3200 189.1400 58.3200 189.6200 ;
        RECT 1.5600 200.0200 4.5600 200.5000 ;
        RECT 1.5600 205.4600 4.5600 205.9400 ;
        RECT 12.3200 200.0200 13.3200 200.5000 ;
        RECT 12.3200 205.4600 13.3200 205.9400 ;
        RECT 57.3200 205.4600 58.3200 205.9400 ;
        RECT 57.3200 200.0200 58.3200 200.5000 ;
        RECT 102.3200 183.7000 103.3200 184.1800 ;
        RECT 102.3200 178.2600 103.3200 178.7400 ;
        RECT 102.3200 172.8200 103.3200 173.3000 ;
        RECT 102.3200 194.5800 103.3200 195.0600 ;
        RECT 102.3200 189.1400 103.3200 189.6200 ;
        RECT 102.3200 205.4600 103.3200 205.9400 ;
        RECT 102.3200 200.0200 103.3200 200.5000 ;
        RECT 147.3200 123.8600 148.3200 124.3400 ;
        RECT 147.3200 118.4200 148.3200 118.9000 ;
        RECT 147.3200 112.9800 148.3200 113.4600 ;
        RECT 147.3200 134.7400 148.3200 135.2200 ;
        RECT 147.3200 129.3000 148.3200 129.7800 ;
        RECT 147.3200 151.0600 148.3200 151.5400 ;
        RECT 147.3200 145.6200 148.3200 146.1000 ;
        RECT 147.3200 140.1800 148.3200 140.6600 ;
        RECT 147.3200 167.3800 148.3200 167.8600 ;
        RECT 147.3200 161.9400 148.3200 162.4200 ;
        RECT 147.3200 156.5000 148.3200 156.9800 ;
        RECT 192.3200 123.8600 193.3200 124.3400 ;
        RECT 192.3200 118.4200 193.3200 118.9000 ;
        RECT 192.3200 112.9800 193.3200 113.4600 ;
        RECT 192.3200 134.7400 193.3200 135.2200 ;
        RECT 192.3200 129.3000 193.3200 129.7800 ;
        RECT 235.5600 112.9800 238.5600 113.4600 ;
        RECT 235.5600 123.8600 238.5600 124.3400 ;
        RECT 235.5600 118.4200 238.5600 118.9000 ;
        RECT 235.5600 134.7400 238.5600 135.2200 ;
        RECT 235.5600 129.3000 238.5600 129.7800 ;
        RECT 192.3200 151.0600 193.3200 151.5400 ;
        RECT 192.3200 145.6200 193.3200 146.1000 ;
        RECT 192.3200 140.1800 193.3200 140.6600 ;
        RECT 192.3200 167.3800 193.3200 167.8600 ;
        RECT 192.3200 161.9400 193.3200 162.4200 ;
        RECT 192.3200 156.5000 193.3200 156.9800 ;
        RECT 235.5600 145.6200 238.5600 146.1000 ;
        RECT 235.5600 140.1800 238.5600 140.6600 ;
        RECT 235.5600 151.0600 238.5600 151.5400 ;
        RECT 235.5600 167.3800 238.5600 167.8600 ;
        RECT 235.5600 161.9400 238.5600 162.4200 ;
        RECT 235.5600 156.5000 238.5600 156.9800 ;
        RECT 147.3200 183.7000 148.3200 184.1800 ;
        RECT 147.3200 178.2600 148.3200 178.7400 ;
        RECT 147.3200 172.8200 148.3200 173.3000 ;
        RECT 147.3200 194.5800 148.3200 195.0600 ;
        RECT 147.3200 189.1400 148.3200 189.6200 ;
        RECT 147.3200 205.4600 148.3200 205.9400 ;
        RECT 147.3200 200.0200 148.3200 200.5000 ;
        RECT 192.3200 183.7000 193.3200 184.1800 ;
        RECT 192.3200 178.2600 193.3200 178.7400 ;
        RECT 192.3200 172.8200 193.3200 173.3000 ;
        RECT 192.3200 194.5800 193.3200 195.0600 ;
        RECT 192.3200 189.1400 193.3200 189.6200 ;
        RECT 235.5600 172.8200 238.5600 173.3000 ;
        RECT 235.5600 183.7000 238.5600 184.1800 ;
        RECT 235.5600 178.2600 238.5600 178.7400 ;
        RECT 235.5600 194.5800 238.5600 195.0600 ;
        RECT 235.5600 189.1400 238.5600 189.6200 ;
        RECT 192.3200 205.4600 193.3200 205.9400 ;
        RECT 192.3200 200.0200 193.3200 200.5000 ;
        RECT 235.5600 205.4600 238.5600 205.9400 ;
        RECT 235.5600 200.0200 238.5600 200.5000 ;
      LAYER met4 ;
        RECT 1.5600 1.4300 4.5600 217.5300 ;
        RECT 235.5600 1.4300 238.5600 217.5300 ;
        RECT 12.3200 1.4300 13.3200 217.5300 ;
        RECT 57.3200 1.4300 58.3200 217.5300 ;
        RECT 102.3200 1.4300 103.3200 217.5300 ;
        RECT 147.3200 1.4300 148.3200 217.5300 ;
        RECT 192.3200 1.4300 193.3200 217.5300 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.6300 218.7500 240.1200 219.6400 ;
      RECT 148.7100 218.7500 148.9100 219.6400 ;
      RECT 147.3300 218.7500 147.9900 219.6400 ;
      RECT 145.9500 218.7500 146.6100 219.6400 ;
      RECT 144.5700 218.7500 145.2300 219.6400 ;
      RECT 143.1900 218.7500 143.8500 219.6400 ;
      RECT 141.8100 218.7500 142.4700 219.6400 ;
      RECT 140.4300 218.7500 141.0900 219.6400 ;
      RECT 139.0500 218.7500 139.7100 219.6400 ;
      RECT 137.6700 218.7500 138.3300 219.6400 ;
      RECT 136.2900 218.7500 136.9500 219.6400 ;
      RECT 134.9100 218.7500 135.5700 219.6400 ;
      RECT 133.5300 218.7500 134.1900 219.6400 ;
      RECT 132.1500 218.7500 132.8100 219.6400 ;
      RECT 130.7700 218.7500 131.4300 219.6400 ;
      RECT 129.3900 218.7500 130.0500 219.6400 ;
      RECT 128.0100 218.7500 128.6700 219.6400 ;
      RECT 126.6300 218.7500 127.2900 219.6400 ;
      RECT 125.7100 218.7500 125.9100 219.6400 ;
      RECT 124.3300 218.7500 124.9900 219.6400 ;
      RECT 122.9500 218.7500 123.6100 219.6400 ;
      RECT 121.5700 218.7500 122.2300 219.6400 ;
      RECT 120.1900 218.7500 120.8500 219.6400 ;
      RECT 118.8100 218.7500 119.4700 219.6400 ;
      RECT 117.4300 218.7500 118.0900 219.6400 ;
      RECT 116.0500 218.7500 116.7100 219.6400 ;
      RECT 114.6700 218.7500 115.3300 219.6400 ;
      RECT 113.2900 218.7500 113.9500 219.6400 ;
      RECT 111.9100 218.7500 112.5700 219.6400 ;
      RECT 110.5300 218.7500 111.1900 219.6400 ;
      RECT 109.1500 218.7500 109.8100 219.6400 ;
      RECT 107.7700 218.7500 108.4300 219.6400 ;
      RECT 106.3900 218.7500 107.0500 219.6400 ;
      RECT 105.0100 218.7500 105.6700 219.6400 ;
      RECT 103.6300 218.7500 104.2900 219.6400 ;
      RECT 102.7100 218.7500 102.9100 219.6400 ;
      RECT 101.3300 218.7500 101.9900 219.6400 ;
      RECT 99.9500 218.7500 100.6100 219.6400 ;
      RECT 98.5700 218.7500 99.2300 219.6400 ;
      RECT 97.1900 218.7500 97.8500 219.6400 ;
      RECT 95.8100 218.7500 96.4700 219.6400 ;
      RECT 94.4300 218.7500 95.0900 219.6400 ;
      RECT 93.0500 218.7500 93.7100 219.6400 ;
      RECT 91.6700 218.7500 92.3300 219.6400 ;
      RECT 90.2900 218.7500 90.9500 219.6400 ;
      RECT 88.9100 218.7500 89.5700 219.6400 ;
      RECT 87.5300 218.7500 88.1900 219.6400 ;
      RECT 86.1500 218.7500 86.8100 219.6400 ;
      RECT 84.7700 218.7500 85.4300 219.6400 ;
      RECT 83.3900 218.7500 84.0500 219.6400 ;
      RECT 82.0100 218.7500 82.6700 219.6400 ;
      RECT 80.6300 218.7500 81.2900 219.6400 ;
      RECT 79.7100 218.7500 79.9100 219.6400 ;
      RECT 78.3300 218.7500 78.9900 219.6400 ;
      RECT 76.9500 218.7500 77.6100 219.6400 ;
      RECT 75.5700 218.7500 76.2300 219.6400 ;
      RECT 74.1900 218.7500 74.8500 219.6400 ;
      RECT 72.8100 218.7500 73.4700 219.6400 ;
      RECT 71.4300 218.7500 72.0900 219.6400 ;
      RECT 70.0500 218.7500 70.7100 219.6400 ;
      RECT 68.6700 218.7500 69.3300 219.6400 ;
      RECT 67.2900 218.7500 67.9500 219.6400 ;
      RECT 65.9100 218.7500 66.5700 219.6400 ;
      RECT 64.5300 218.7500 65.1900 219.6400 ;
      RECT 63.1500 218.7500 63.8100 219.6400 ;
      RECT 61.7700 218.7500 62.4300 219.6400 ;
      RECT 60.3900 218.7500 61.0500 219.6400 ;
      RECT 59.0100 218.7500 59.6700 219.6400 ;
      RECT 57.6300 218.7500 58.2900 219.6400 ;
      RECT 56.7100 218.7500 56.9100 219.6400 ;
      RECT 55.3300 218.7500 55.9900 219.6400 ;
      RECT 53.9500 218.7500 54.6100 219.6400 ;
      RECT 52.5700 218.7500 53.2300 219.6400 ;
      RECT 51.1900 218.7500 51.8500 219.6400 ;
      RECT 49.8100 218.7500 50.4700 219.6400 ;
      RECT 48.4300 218.7500 49.0900 219.6400 ;
      RECT 47.0500 218.7500 47.7100 219.6400 ;
      RECT 45.6700 218.7500 46.3300 219.6400 ;
      RECT 44.2900 218.7500 44.9500 219.6400 ;
      RECT 42.9100 218.7500 43.5700 219.6400 ;
      RECT 41.5300 218.7500 42.1900 219.6400 ;
      RECT 40.1500 218.7500 40.8100 219.6400 ;
      RECT 38.7700 218.7500 39.4300 219.6400 ;
      RECT 37.3900 218.7500 38.0500 219.6400 ;
      RECT 36.0100 218.7500 36.6700 219.6400 ;
      RECT 34.6300 218.7500 35.2900 219.6400 ;
      RECT 33.7100 218.7500 33.9100 219.6400 ;
      RECT 32.3300 218.7500 32.9900 219.6400 ;
      RECT 30.9500 218.7500 31.6100 219.6400 ;
      RECT 29.5700 218.7500 30.2300 219.6400 ;
      RECT 28.1900 218.7500 28.8500 219.6400 ;
      RECT 26.8100 218.7500 27.4700 219.6400 ;
      RECT 25.4300 218.7500 26.0900 219.6400 ;
      RECT 24.0500 218.7500 24.7100 219.6400 ;
      RECT 22.6700 218.7500 23.3300 219.6400 ;
      RECT 21.2900 218.7500 21.9500 219.6400 ;
      RECT 19.9100 218.7500 20.5700 219.6400 ;
      RECT 18.5300 218.7500 19.1900 219.6400 ;
      RECT 17.1500 218.7500 17.8100 219.6400 ;
      RECT 15.7700 218.7500 16.4300 219.6400 ;
      RECT 14.3900 218.7500 15.0500 219.6400 ;
      RECT 13.0100 218.7500 13.6700 219.6400 ;
      RECT 11.6300 218.7500 12.2900 219.6400 ;
      RECT 10.7100 218.7500 10.9100 219.6400 ;
      RECT 0.0000 218.7500 9.9900 219.6400 ;
      RECT 0.0000 0.8900 240.1200 218.7500 ;
      RECT 149.6300 0.0000 240.1200 0.8900 ;
      RECT 148.7100 0.0000 148.9100 0.8900 ;
      RECT 147.3300 0.0000 147.9900 0.8900 ;
      RECT 145.9500 0.0000 146.6100 0.8900 ;
      RECT 144.5700 0.0000 145.2300 0.8900 ;
      RECT 143.1900 0.0000 143.8500 0.8900 ;
      RECT 141.8100 0.0000 142.4700 0.8900 ;
      RECT 140.4300 0.0000 141.0900 0.8900 ;
      RECT 139.0500 0.0000 139.7100 0.8900 ;
      RECT 137.6700 0.0000 138.3300 0.8900 ;
      RECT 136.2900 0.0000 136.9500 0.8900 ;
      RECT 134.9100 0.0000 135.5700 0.8900 ;
      RECT 133.5300 0.0000 134.1900 0.8900 ;
      RECT 132.1500 0.0000 132.8100 0.8900 ;
      RECT 130.7700 0.0000 131.4300 0.8900 ;
      RECT 129.3900 0.0000 130.0500 0.8900 ;
      RECT 128.0100 0.0000 128.6700 0.8900 ;
      RECT 126.6300 0.0000 127.2900 0.8900 ;
      RECT 125.7100 0.0000 125.9100 0.8900 ;
      RECT 124.3300 0.0000 124.9900 0.8900 ;
      RECT 122.9500 0.0000 123.6100 0.8900 ;
      RECT 121.5700 0.0000 122.2300 0.8900 ;
      RECT 120.1900 0.0000 120.8500 0.8900 ;
      RECT 118.8100 0.0000 119.4700 0.8900 ;
      RECT 117.4300 0.0000 118.0900 0.8900 ;
      RECT 116.0500 0.0000 116.7100 0.8900 ;
      RECT 114.6700 0.0000 115.3300 0.8900 ;
      RECT 113.2900 0.0000 113.9500 0.8900 ;
      RECT 111.9100 0.0000 112.5700 0.8900 ;
      RECT 110.5300 0.0000 111.1900 0.8900 ;
      RECT 109.1500 0.0000 109.8100 0.8900 ;
      RECT 107.7700 0.0000 108.4300 0.8900 ;
      RECT 106.3900 0.0000 107.0500 0.8900 ;
      RECT 105.0100 0.0000 105.6700 0.8900 ;
      RECT 103.6300 0.0000 104.2900 0.8900 ;
      RECT 102.7100 0.0000 102.9100 0.8900 ;
      RECT 101.3300 0.0000 101.9900 0.8900 ;
      RECT 99.9500 0.0000 100.6100 0.8900 ;
      RECT 98.5700 0.0000 99.2300 0.8900 ;
      RECT 97.1900 0.0000 97.8500 0.8900 ;
      RECT 95.8100 0.0000 96.4700 0.8900 ;
      RECT 94.4300 0.0000 95.0900 0.8900 ;
      RECT 93.0500 0.0000 93.7100 0.8900 ;
      RECT 91.6700 0.0000 92.3300 0.8900 ;
      RECT 90.2900 0.0000 90.9500 0.8900 ;
      RECT 88.9100 0.0000 89.5700 0.8900 ;
      RECT 87.5300 0.0000 88.1900 0.8900 ;
      RECT 86.1500 0.0000 86.8100 0.8900 ;
      RECT 84.7700 0.0000 85.4300 0.8900 ;
      RECT 83.3900 0.0000 84.0500 0.8900 ;
      RECT 82.0100 0.0000 82.6700 0.8900 ;
      RECT 80.6300 0.0000 81.2900 0.8900 ;
      RECT 79.7100 0.0000 79.9100 0.8900 ;
      RECT 78.3300 0.0000 78.9900 0.8900 ;
      RECT 76.9500 0.0000 77.6100 0.8900 ;
      RECT 75.5700 0.0000 76.2300 0.8900 ;
      RECT 74.1900 0.0000 74.8500 0.8900 ;
      RECT 72.8100 0.0000 73.4700 0.8900 ;
      RECT 71.4300 0.0000 72.0900 0.8900 ;
      RECT 70.0500 0.0000 70.7100 0.8900 ;
      RECT 68.6700 0.0000 69.3300 0.8900 ;
      RECT 67.2900 0.0000 67.9500 0.8900 ;
      RECT 65.9100 0.0000 66.5700 0.8900 ;
      RECT 64.5300 0.0000 65.1900 0.8900 ;
      RECT 63.1500 0.0000 63.8100 0.8900 ;
      RECT 61.7700 0.0000 62.4300 0.8900 ;
      RECT 60.3900 0.0000 61.0500 0.8900 ;
      RECT 59.0100 0.0000 59.6700 0.8900 ;
      RECT 57.6300 0.0000 58.2900 0.8900 ;
      RECT 56.7100 0.0000 56.9100 0.8900 ;
      RECT 55.3300 0.0000 55.9900 0.8900 ;
      RECT 53.9500 0.0000 54.6100 0.8900 ;
      RECT 52.5700 0.0000 53.2300 0.8900 ;
      RECT 51.1900 0.0000 51.8500 0.8900 ;
      RECT 49.8100 0.0000 50.4700 0.8900 ;
      RECT 48.4300 0.0000 49.0900 0.8900 ;
      RECT 47.0500 0.0000 47.7100 0.8900 ;
      RECT 45.6700 0.0000 46.3300 0.8900 ;
      RECT 44.2900 0.0000 44.9500 0.8900 ;
      RECT 42.9100 0.0000 43.5700 0.8900 ;
      RECT 41.5300 0.0000 42.1900 0.8900 ;
      RECT 40.1500 0.0000 40.8100 0.8900 ;
      RECT 38.7700 0.0000 39.4300 0.8900 ;
      RECT 37.3900 0.0000 38.0500 0.8900 ;
      RECT 36.0100 0.0000 36.6700 0.8900 ;
      RECT 34.6300 0.0000 35.2900 0.8900 ;
      RECT 33.7100 0.0000 33.9100 0.8900 ;
      RECT 32.3300 0.0000 32.9900 0.8900 ;
      RECT 30.9500 0.0000 31.6100 0.8900 ;
      RECT 29.5700 0.0000 30.2300 0.8900 ;
      RECT 28.1900 0.0000 28.8500 0.8900 ;
      RECT 26.8100 0.0000 27.4700 0.8900 ;
      RECT 25.4300 0.0000 26.0900 0.8900 ;
      RECT 24.0500 0.0000 24.7100 0.8900 ;
      RECT 22.6700 0.0000 23.3300 0.8900 ;
      RECT 21.2900 0.0000 21.9500 0.8900 ;
      RECT 19.9100 0.0000 20.5700 0.8900 ;
      RECT 18.5300 0.0000 19.1900 0.8900 ;
      RECT 17.1500 0.0000 17.8100 0.8900 ;
      RECT 15.7700 0.0000 16.4300 0.8900 ;
      RECT 14.3900 0.0000 15.0500 0.8900 ;
      RECT 13.0100 0.0000 13.6700 0.8900 ;
      RECT 11.6300 0.0000 12.2900 0.8900 ;
      RECT 10.7100 0.0000 10.9100 0.8900 ;
      RECT 0.0000 0.0000 9.9900 0.8900 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 240.1200 219.6400 ;
    LAYER met2 ;
      RECT 209.8600 218.7800 240.1200 219.6400 ;
      RECT 206.6400 218.7800 209.2000 219.6400 ;
      RECT 203.8800 218.7800 205.9800 219.6400 ;
      RECT 200.6600 218.7800 203.2200 219.6400 ;
      RECT 198.3600 218.7800 200.0000 219.6400 ;
      RECT 195.6000 218.7800 197.7000 219.6400 ;
      RECT 192.8400 218.7800 194.9400 219.6400 ;
      RECT 189.1600 218.7800 192.1800 219.6400 ;
      RECT 186.8600 218.7800 188.5000 219.6400 ;
      RECT 184.1000 218.7800 186.2000 219.6400 ;
      RECT 181.3400 218.7800 183.4400 219.6400 ;
      RECT 178.5800 218.7800 180.6800 219.6400 ;
      RECT 175.8200 218.7800 177.9200 219.6400 ;
      RECT 172.6000 218.7800 175.1600 219.6400 ;
      RECT 169.8400 218.7800 171.9400 219.6400 ;
      RECT 167.0800 218.7800 169.1800 219.6400 ;
      RECT 164.3200 218.7800 166.4200 219.6400 ;
      RECT 161.1000 218.7800 163.6600 219.6400 ;
      RECT 158.8000 218.7800 160.4400 219.6400 ;
      RECT 156.0400 218.7800 158.1400 219.6400 ;
      RECT 0.0000 218.7800 155.3800 219.6400 ;
      RECT 0.0000 209.9400 240.1200 218.7800 ;
      RECT 0.8600 209.2800 239.2600 209.9400 ;
      RECT 0.0000 208.2400 240.1200 209.2800 ;
      RECT 0.8600 207.5800 239.2600 208.2400 ;
      RECT 0.0000 206.5400 240.1200 207.5800 ;
      RECT 0.8600 205.8800 239.2600 206.5400 ;
      RECT 0.0000 204.8400 240.1200 205.8800 ;
      RECT 0.8600 204.1800 239.2600 204.8400 ;
      RECT 0.0000 203.1400 240.1200 204.1800 ;
      RECT 0.8600 202.4800 239.2600 203.1400 ;
      RECT 0.0000 201.4400 240.1200 202.4800 ;
      RECT 0.8600 200.7800 239.2600 201.4400 ;
      RECT 0.0000 199.4000 240.1200 200.7800 ;
      RECT 0.8600 198.7400 239.2600 199.4000 ;
      RECT 0.0000 197.7000 240.1200 198.7400 ;
      RECT 0.8600 197.0400 239.2600 197.7000 ;
      RECT 0.0000 196.0000 240.1200 197.0400 ;
      RECT 0.8600 195.3400 239.2600 196.0000 ;
      RECT 0.0000 194.3000 240.1200 195.3400 ;
      RECT 0.8600 193.6400 239.2600 194.3000 ;
      RECT 0.0000 192.6000 240.1200 193.6400 ;
      RECT 0.8600 191.9400 239.2600 192.6000 ;
      RECT 0.0000 190.5600 240.1200 191.9400 ;
      RECT 0.8600 189.9000 239.2600 190.5600 ;
      RECT 0.0000 188.8600 240.1200 189.9000 ;
      RECT 0.8600 188.2000 239.2600 188.8600 ;
      RECT 0.0000 187.1600 240.1200 188.2000 ;
      RECT 0.8600 186.5000 239.2600 187.1600 ;
      RECT 0.0000 185.4600 240.1200 186.5000 ;
      RECT 0.8600 184.8000 239.2600 185.4600 ;
      RECT 0.0000 183.7600 240.1200 184.8000 ;
      RECT 0.8600 183.1000 239.2600 183.7600 ;
      RECT 0.0000 181.7200 240.1200 183.1000 ;
      RECT 0.8600 181.0600 239.2600 181.7200 ;
      RECT 0.0000 180.0200 240.1200 181.0600 ;
      RECT 0.8600 179.3600 239.2600 180.0200 ;
      RECT 0.0000 178.3200 240.1200 179.3600 ;
      RECT 0.8600 177.6600 239.2600 178.3200 ;
      RECT 0.0000 176.6200 240.1200 177.6600 ;
      RECT 0.8600 175.9600 239.2600 176.6200 ;
      RECT 0.0000 174.9200 240.1200 175.9600 ;
      RECT 0.8600 174.2600 239.2600 174.9200 ;
      RECT 0.0000 172.8800 240.1200 174.2600 ;
      RECT 0.8600 172.2200 239.2600 172.8800 ;
      RECT 0.0000 171.1800 240.1200 172.2200 ;
      RECT 0.8600 170.5200 239.2600 171.1800 ;
      RECT 0.0000 169.4800 240.1200 170.5200 ;
      RECT 0.8600 168.8200 239.2600 169.4800 ;
      RECT 0.0000 167.7800 240.1200 168.8200 ;
      RECT 0.8600 167.1200 239.2600 167.7800 ;
      RECT 0.0000 166.0800 240.1200 167.1200 ;
      RECT 0.8600 165.4200 239.2600 166.0800 ;
      RECT 0.0000 164.0400 240.1200 165.4200 ;
      RECT 0.8600 163.3800 239.2600 164.0400 ;
      RECT 0.0000 162.3400 240.1200 163.3800 ;
      RECT 0.8600 161.6800 239.2600 162.3400 ;
      RECT 0.0000 160.6400 240.1200 161.6800 ;
      RECT 0.8600 159.9800 239.2600 160.6400 ;
      RECT 0.0000 158.9400 240.1200 159.9800 ;
      RECT 0.8600 158.2800 239.2600 158.9400 ;
      RECT 0.0000 157.2400 240.1200 158.2800 ;
      RECT 0.8600 156.5800 239.2600 157.2400 ;
      RECT 0.0000 155.5400 240.1200 156.5800 ;
      RECT 0.8600 154.8800 239.2600 155.5400 ;
      RECT 0.0000 150.1000 240.1200 154.8800 ;
      RECT 0.8600 149.4400 239.2600 150.1000 ;
      RECT 0.0000 148.4000 240.1200 149.4400 ;
      RECT 0.8600 147.7400 239.2600 148.4000 ;
      RECT 0.0000 147.0400 240.1200 147.7400 ;
      RECT 0.8600 146.3800 239.2600 147.0400 ;
      RECT 0.0000 145.6800 240.1200 146.3800 ;
      RECT 0.8600 145.0200 239.2600 145.6800 ;
      RECT 0.0000 143.9800 240.1200 145.0200 ;
      RECT 0.8600 143.3200 239.2600 143.9800 ;
      RECT 0.0000 142.6200 240.1200 143.3200 ;
      RECT 0.8600 141.9600 239.2600 142.6200 ;
      RECT 0.0000 141.2600 240.1200 141.9600 ;
      RECT 0.8600 140.6000 239.2600 141.2600 ;
      RECT 0.0000 139.5600 240.1200 140.6000 ;
      RECT 0.8600 138.9000 239.2600 139.5600 ;
      RECT 0.0000 138.2000 240.1200 138.9000 ;
      RECT 0.8600 137.5400 239.2600 138.2000 ;
      RECT 0.0000 136.8400 240.1200 137.5400 ;
      RECT 0.8600 136.1800 239.2600 136.8400 ;
      RECT 0.0000 135.1400 240.1200 136.1800 ;
      RECT 0.8600 134.4800 239.2600 135.1400 ;
      RECT 0.0000 133.7800 240.1200 134.4800 ;
      RECT 0.8600 133.1200 239.2600 133.7800 ;
      RECT 0.0000 132.4200 240.1200 133.1200 ;
      RECT 0.8600 131.7600 239.2600 132.4200 ;
      RECT 0.0000 130.7200 240.1200 131.7600 ;
      RECT 0.8600 130.0600 239.2600 130.7200 ;
      RECT 0.0000 129.3600 240.1200 130.0600 ;
      RECT 0.8600 128.7000 239.2600 129.3600 ;
      RECT 0.0000 128.0000 240.1200 128.7000 ;
      RECT 0.8600 127.3400 239.2600 128.0000 ;
      RECT 0.0000 126.3000 240.1200 127.3400 ;
      RECT 0.8600 125.6400 239.2600 126.3000 ;
      RECT 0.0000 124.9400 240.1200 125.6400 ;
      RECT 0.8600 124.2800 239.2600 124.9400 ;
      RECT 0.0000 123.5800 240.1200 124.2800 ;
      RECT 0.8600 122.9200 239.2600 123.5800 ;
      RECT 0.0000 121.8800 240.1200 122.9200 ;
      RECT 0.8600 121.2200 239.2600 121.8800 ;
      RECT 0.0000 120.5200 240.1200 121.2200 ;
      RECT 0.8600 119.8600 239.2600 120.5200 ;
      RECT 0.0000 119.1600 240.1200 119.8600 ;
      RECT 0.8600 118.5000 239.2600 119.1600 ;
      RECT 0.0000 117.4600 240.1200 118.5000 ;
      RECT 0.8600 116.8000 239.2600 117.4600 ;
      RECT 0.0000 116.1000 240.1200 116.8000 ;
      RECT 0.8600 115.4400 239.2600 116.1000 ;
      RECT 0.0000 114.7400 240.1200 115.4400 ;
      RECT 0.8600 114.0800 239.2600 114.7400 ;
      RECT 0.0000 113.0400 240.1200 114.0800 ;
      RECT 0.8600 112.3800 239.2600 113.0400 ;
      RECT 0.0000 111.6800 240.1200 112.3800 ;
      RECT 0.8600 111.0200 239.2600 111.6800 ;
      RECT 0.0000 110.3200 240.1200 111.0200 ;
      RECT 0.8600 109.6600 239.2600 110.3200 ;
      RECT 0.0000 108.6200 240.1200 109.6600 ;
      RECT 0.8600 107.9600 239.2600 108.6200 ;
      RECT 0.0000 107.2600 240.1200 107.9600 ;
      RECT 0.8600 106.6000 239.2600 107.2600 ;
      RECT 0.0000 105.9000 240.1200 106.6000 ;
      RECT 0.8600 105.2400 239.2600 105.9000 ;
      RECT 0.0000 104.2000 240.1200 105.2400 ;
      RECT 0.8600 103.5400 239.2600 104.2000 ;
      RECT 0.0000 102.8400 240.1200 103.5400 ;
      RECT 0.8600 102.1800 239.2600 102.8400 ;
      RECT 0.0000 101.4800 240.1200 102.1800 ;
      RECT 0.8600 100.8200 239.2600 101.4800 ;
      RECT 0.0000 99.7800 240.1200 100.8200 ;
      RECT 0.8600 99.1200 239.2600 99.7800 ;
      RECT 0.0000 98.4200 240.1200 99.1200 ;
      RECT 0.8600 97.7600 239.2600 98.4200 ;
      RECT 0.0000 97.0600 240.1200 97.7600 ;
      RECT 0.8600 96.4000 239.2600 97.0600 ;
      RECT 0.0000 95.3600 240.1200 96.4000 ;
      RECT 0.8600 94.7000 239.2600 95.3600 ;
      RECT 0.0000 94.0000 240.1200 94.7000 ;
      RECT 0.8600 93.3400 239.2600 94.0000 ;
      RECT 0.0000 92.6400 240.1200 93.3400 ;
      RECT 0.8600 91.9800 239.2600 92.6400 ;
      RECT 0.0000 90.9400 240.1200 91.9800 ;
      RECT 0.8600 90.2800 239.2600 90.9400 ;
      RECT 0.0000 89.5800 240.1200 90.2800 ;
      RECT 0.8600 88.9200 239.2600 89.5800 ;
      RECT 0.0000 88.2200 240.1200 88.9200 ;
      RECT 0.8600 87.5600 239.2600 88.2200 ;
      RECT 0.0000 86.5200 240.1200 87.5600 ;
      RECT 0.8600 85.8600 239.2600 86.5200 ;
      RECT 0.0000 85.1600 240.1200 85.8600 ;
      RECT 0.8600 84.5000 239.2600 85.1600 ;
      RECT 0.0000 83.8000 240.1200 84.5000 ;
      RECT 0.8600 83.1400 239.2600 83.8000 ;
      RECT 0.0000 82.1000 240.1200 83.1400 ;
      RECT 0.8600 81.4400 239.2600 82.1000 ;
      RECT 0.0000 80.7400 240.1200 81.4400 ;
      RECT 0.8600 80.0800 239.2600 80.7400 ;
      RECT 0.0000 79.3800 240.1200 80.0800 ;
      RECT 0.8600 78.7200 239.2600 79.3800 ;
      RECT 0.0000 78.0200 240.1200 78.7200 ;
      RECT 0.8600 77.3600 239.2600 78.0200 ;
      RECT 0.0000 76.3200 240.1200 77.3600 ;
      RECT 0.8600 75.6600 239.2600 76.3200 ;
      RECT 0.0000 74.9600 240.1200 75.6600 ;
      RECT 0.8600 74.3000 239.2600 74.9600 ;
      RECT 0.0000 73.6000 240.1200 74.3000 ;
      RECT 0.8600 72.9400 239.2600 73.6000 ;
      RECT 0.0000 71.9000 240.1200 72.9400 ;
      RECT 0.8600 71.2400 239.2600 71.9000 ;
      RECT 0.0000 70.5400 240.1200 71.2400 ;
      RECT 0.8600 69.8800 239.2600 70.5400 ;
      RECT 0.0000 69.1800 240.1200 69.8800 ;
      RECT 0.8600 68.5200 239.2600 69.1800 ;
      RECT 0.0000 67.4800 240.1200 68.5200 ;
      RECT 0.8600 66.8200 239.2600 67.4800 ;
      RECT 0.0000 66.1200 240.1200 66.8200 ;
      RECT 0.8600 65.4600 239.2600 66.1200 ;
      RECT 0.0000 64.7600 240.1200 65.4600 ;
      RECT 0.8600 64.1000 239.2600 64.7600 ;
      RECT 0.0000 63.0600 240.1200 64.1000 ;
      RECT 0.8600 62.4000 239.2600 63.0600 ;
      RECT 0.0000 61.7000 240.1200 62.4000 ;
      RECT 0.8600 61.0400 239.2600 61.7000 ;
      RECT 0.0000 60.3400 240.1200 61.0400 ;
      RECT 0.8600 59.6800 239.2600 60.3400 ;
      RECT 0.0000 58.6400 240.1200 59.6800 ;
      RECT 0.8600 57.9800 239.2600 58.6400 ;
      RECT 0.0000 57.2800 240.1200 57.9800 ;
      RECT 0.8600 56.6200 239.2600 57.2800 ;
      RECT 0.0000 55.9200 240.1200 56.6200 ;
      RECT 0.8600 55.2600 239.2600 55.9200 ;
      RECT 0.0000 54.2200 240.1200 55.2600 ;
      RECT 0.8600 53.5600 239.2600 54.2200 ;
      RECT 0.0000 52.8600 240.1200 53.5600 ;
      RECT 0.8600 52.2000 239.2600 52.8600 ;
      RECT 0.0000 51.5000 240.1200 52.2000 ;
      RECT 0.8600 50.8400 239.2600 51.5000 ;
      RECT 0.0000 49.8000 240.1200 50.8400 ;
      RECT 0.8600 49.1400 239.2600 49.8000 ;
      RECT 0.0000 48.4400 240.1200 49.1400 ;
      RECT 0.8600 47.7800 239.2600 48.4400 ;
      RECT 0.0000 47.0800 240.1200 47.7800 ;
      RECT 0.8600 46.4200 239.2600 47.0800 ;
      RECT 0.0000 45.3800 240.1200 46.4200 ;
      RECT 0.8600 44.7200 239.2600 45.3800 ;
      RECT 0.0000 44.0200 240.1200 44.7200 ;
      RECT 0.8600 43.3600 239.2600 44.0200 ;
      RECT 0.0000 42.6600 240.1200 43.3600 ;
      RECT 0.8600 42.0000 239.2600 42.6600 ;
      RECT 0.0000 40.9600 240.1200 42.0000 ;
      RECT 0.8600 40.3000 239.2600 40.9600 ;
      RECT 0.0000 39.6000 240.1200 40.3000 ;
      RECT 0.8600 38.9400 239.2600 39.6000 ;
      RECT 0.0000 38.2400 240.1200 38.9400 ;
      RECT 0.8600 37.5800 239.2600 38.2400 ;
      RECT 0.0000 36.5400 240.1200 37.5800 ;
      RECT 0.8600 35.8800 239.2600 36.5400 ;
      RECT 0.0000 35.1800 240.1200 35.8800 ;
      RECT 0.8600 34.5200 239.2600 35.1800 ;
      RECT 0.0000 33.8200 240.1200 34.5200 ;
      RECT 0.8600 33.1600 239.2600 33.8200 ;
      RECT 0.0000 32.1200 240.1200 33.1600 ;
      RECT 0.8600 31.4600 239.2600 32.1200 ;
      RECT 0.0000 30.7600 240.1200 31.4600 ;
      RECT 0.8600 30.1000 239.2600 30.7600 ;
      RECT 0.0000 29.4000 240.1200 30.1000 ;
      RECT 0.8600 28.7400 239.2600 29.4000 ;
      RECT 0.0000 27.7000 240.1200 28.7400 ;
      RECT 0.8600 27.0400 239.2600 27.7000 ;
      RECT 0.0000 26.3400 240.1200 27.0400 ;
      RECT 0.8600 25.6800 239.2600 26.3400 ;
      RECT 0.0000 24.9800 240.1200 25.6800 ;
      RECT 0.8600 24.3200 239.2600 24.9800 ;
      RECT 0.0000 23.2800 240.1200 24.3200 ;
      RECT 0.8600 22.6200 239.2600 23.2800 ;
      RECT 0.0000 21.9200 240.1200 22.6200 ;
      RECT 0.8600 21.2600 239.2600 21.9200 ;
      RECT 0.0000 20.5600 240.1200 21.2600 ;
      RECT 0.8600 19.9000 239.2600 20.5600 ;
      RECT 0.0000 18.8600 240.1200 19.9000 ;
      RECT 0.8600 18.2000 239.2600 18.8600 ;
      RECT 0.0000 17.5000 240.1200 18.2000 ;
      RECT 0.8600 16.8400 239.2600 17.5000 ;
      RECT 0.0000 16.1400 240.1200 16.8400 ;
      RECT 0.8600 15.4800 239.2600 16.1400 ;
      RECT 0.0000 14.4400 240.1200 15.4800 ;
      RECT 0.8600 13.7800 239.2600 14.4400 ;
      RECT 0.0000 13.0800 240.1200 13.7800 ;
      RECT 0.8600 12.4200 239.2600 13.0800 ;
      RECT 0.0000 11.7200 240.1200 12.4200 ;
      RECT 0.8600 11.0600 239.2600 11.7200 ;
      RECT 0.0000 10.3600 240.1200 11.0600 ;
      RECT 0.8600 9.7000 239.2600 10.3600 ;
      RECT 0.0000 0.8600 240.1200 9.7000 ;
      RECT 210.3200 0.0000 240.1200 0.8600 ;
      RECT 207.1000 0.0000 209.6600 0.8600 ;
      RECT 204.3400 0.0000 206.4400 0.8600 ;
      RECT 201.5800 0.0000 203.6800 0.8600 ;
      RECT 198.3600 0.0000 200.9200 0.8600 ;
      RECT 195.6000 0.0000 197.7000 0.8600 ;
      RECT 192.8400 0.0000 194.9400 0.8600 ;
      RECT 190.0800 0.0000 192.1800 0.8600 ;
      RECT 186.8600 0.0000 189.4200 0.8600 ;
      RECT 184.1000 0.0000 186.2000 0.8600 ;
      RECT 181.3400 0.0000 183.4400 0.8600 ;
      RECT 178.5800 0.0000 180.6800 0.8600 ;
      RECT 175.3600 0.0000 177.9200 0.8600 ;
      RECT 172.6000 0.0000 174.7000 0.8600 ;
      RECT 169.8400 0.0000 171.9400 0.8600 ;
      RECT 167.0800 0.0000 169.1800 0.8600 ;
      RECT 163.8600 0.0000 166.4200 0.8600 ;
      RECT 161.1000 0.0000 163.2000 0.8600 ;
      RECT 158.3400 0.0000 160.4400 0.8600 ;
      RECT 155.5800 0.0000 157.6800 0.8600 ;
      RECT 0.0000 0.0000 154.9200 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 217.8300 240.1200 219.6400 ;
      RECT 238.8600 214.2300 240.1200 217.8300 ;
      RECT 0.0000 214.2300 1.2600 217.8300 ;
      RECT 0.0000 213.8300 240.1200 214.2300 ;
      RECT 234.8600 210.2300 240.1200 213.8300 ;
      RECT 0.0000 210.2300 5.2600 213.8300 ;
      RECT 0.0000 208.9600 240.1200 210.2300 ;
      RECT 234.8600 207.8800 240.1200 208.9600 ;
      RECT 191.4200 207.8800 231.2600 208.9600 ;
      RECT 146.4200 207.8800 189.8200 208.9600 ;
      RECT 101.4200 207.8800 144.8200 208.9600 ;
      RECT 56.4200 207.8800 99.8200 208.9600 ;
      RECT 8.8600 207.8800 54.8200 208.9600 ;
      RECT 0.0000 207.8800 5.2600 208.9600 ;
      RECT 0.0000 206.2400 240.1200 207.8800 ;
      RECT 238.8600 205.1600 240.1200 206.2400 ;
      RECT 193.6200 205.1600 235.2600 206.2400 ;
      RECT 148.6200 205.1600 192.0200 206.2400 ;
      RECT 103.6200 205.1600 147.0200 206.2400 ;
      RECT 58.6200 205.1600 102.0200 206.2400 ;
      RECT 13.6200 205.1600 57.0200 206.2400 ;
      RECT 4.8600 205.1600 12.0200 206.2400 ;
      RECT 0.0000 205.1600 1.2600 206.2400 ;
      RECT 0.0000 203.5200 240.1200 205.1600 ;
      RECT 234.8600 202.4400 240.1200 203.5200 ;
      RECT 191.4200 202.4400 231.2600 203.5200 ;
      RECT 146.4200 202.4400 189.8200 203.5200 ;
      RECT 101.4200 202.4400 144.8200 203.5200 ;
      RECT 56.4200 202.4400 99.8200 203.5200 ;
      RECT 8.8600 202.4400 54.8200 203.5200 ;
      RECT 0.0000 202.4400 5.2600 203.5200 ;
      RECT 0.0000 200.8000 240.1200 202.4400 ;
      RECT 238.8600 199.7200 240.1200 200.8000 ;
      RECT 193.6200 199.7200 235.2600 200.8000 ;
      RECT 148.6200 199.7200 192.0200 200.8000 ;
      RECT 103.6200 199.7200 147.0200 200.8000 ;
      RECT 58.6200 199.7200 102.0200 200.8000 ;
      RECT 13.6200 199.7200 57.0200 200.8000 ;
      RECT 4.8600 199.7200 12.0200 200.8000 ;
      RECT 0.0000 199.7200 1.2600 200.8000 ;
      RECT 0.0000 198.0800 240.1200 199.7200 ;
      RECT 234.8600 197.0000 240.1200 198.0800 ;
      RECT 191.4200 197.0000 231.2600 198.0800 ;
      RECT 146.4200 197.0000 189.8200 198.0800 ;
      RECT 101.4200 197.0000 144.8200 198.0800 ;
      RECT 56.4200 197.0000 99.8200 198.0800 ;
      RECT 8.8600 197.0000 54.8200 198.0800 ;
      RECT 0.0000 197.0000 5.2600 198.0800 ;
      RECT 0.0000 195.3600 240.1200 197.0000 ;
      RECT 238.8600 194.2800 240.1200 195.3600 ;
      RECT 193.6200 194.2800 235.2600 195.3600 ;
      RECT 148.6200 194.2800 192.0200 195.3600 ;
      RECT 103.6200 194.2800 147.0200 195.3600 ;
      RECT 58.6200 194.2800 102.0200 195.3600 ;
      RECT 13.6200 194.2800 57.0200 195.3600 ;
      RECT 4.8600 194.2800 12.0200 195.3600 ;
      RECT 0.0000 194.2800 1.2600 195.3600 ;
      RECT 0.0000 192.6400 240.1200 194.2800 ;
      RECT 234.8600 191.5600 240.1200 192.6400 ;
      RECT 191.4200 191.5600 231.2600 192.6400 ;
      RECT 146.4200 191.5600 189.8200 192.6400 ;
      RECT 101.4200 191.5600 144.8200 192.6400 ;
      RECT 56.4200 191.5600 99.8200 192.6400 ;
      RECT 8.8600 191.5600 54.8200 192.6400 ;
      RECT 0.0000 191.5600 5.2600 192.6400 ;
      RECT 0.0000 189.9200 240.1200 191.5600 ;
      RECT 238.8600 188.8400 240.1200 189.9200 ;
      RECT 193.6200 188.8400 235.2600 189.9200 ;
      RECT 148.6200 188.8400 192.0200 189.9200 ;
      RECT 103.6200 188.8400 147.0200 189.9200 ;
      RECT 58.6200 188.8400 102.0200 189.9200 ;
      RECT 13.6200 188.8400 57.0200 189.9200 ;
      RECT 4.8600 188.8400 12.0200 189.9200 ;
      RECT 0.0000 188.8400 1.2600 189.9200 ;
      RECT 0.0000 187.2000 240.1200 188.8400 ;
      RECT 234.8600 186.1200 240.1200 187.2000 ;
      RECT 191.4200 186.1200 231.2600 187.2000 ;
      RECT 146.4200 186.1200 189.8200 187.2000 ;
      RECT 101.4200 186.1200 144.8200 187.2000 ;
      RECT 56.4200 186.1200 99.8200 187.2000 ;
      RECT 8.8600 186.1200 54.8200 187.2000 ;
      RECT 0.0000 186.1200 5.2600 187.2000 ;
      RECT 0.0000 184.4800 240.1200 186.1200 ;
      RECT 238.8600 183.4000 240.1200 184.4800 ;
      RECT 193.6200 183.4000 235.2600 184.4800 ;
      RECT 148.6200 183.4000 192.0200 184.4800 ;
      RECT 103.6200 183.4000 147.0200 184.4800 ;
      RECT 58.6200 183.4000 102.0200 184.4800 ;
      RECT 13.6200 183.4000 57.0200 184.4800 ;
      RECT 4.8600 183.4000 12.0200 184.4800 ;
      RECT 0.0000 183.4000 1.2600 184.4800 ;
      RECT 0.0000 181.7600 240.1200 183.4000 ;
      RECT 234.8600 180.6800 240.1200 181.7600 ;
      RECT 191.4200 180.6800 231.2600 181.7600 ;
      RECT 146.4200 180.6800 189.8200 181.7600 ;
      RECT 101.4200 180.6800 144.8200 181.7600 ;
      RECT 56.4200 180.6800 99.8200 181.7600 ;
      RECT 8.8600 180.6800 54.8200 181.7600 ;
      RECT 0.0000 180.6800 5.2600 181.7600 ;
      RECT 0.0000 179.0400 240.1200 180.6800 ;
      RECT 238.8600 177.9600 240.1200 179.0400 ;
      RECT 193.6200 177.9600 235.2600 179.0400 ;
      RECT 148.6200 177.9600 192.0200 179.0400 ;
      RECT 103.6200 177.9600 147.0200 179.0400 ;
      RECT 58.6200 177.9600 102.0200 179.0400 ;
      RECT 13.6200 177.9600 57.0200 179.0400 ;
      RECT 4.8600 177.9600 12.0200 179.0400 ;
      RECT 0.0000 177.9600 1.2600 179.0400 ;
      RECT 0.0000 176.3200 240.1200 177.9600 ;
      RECT 234.8600 175.2400 240.1200 176.3200 ;
      RECT 191.4200 175.2400 231.2600 176.3200 ;
      RECT 146.4200 175.2400 189.8200 176.3200 ;
      RECT 101.4200 175.2400 144.8200 176.3200 ;
      RECT 56.4200 175.2400 99.8200 176.3200 ;
      RECT 8.8600 175.2400 54.8200 176.3200 ;
      RECT 0.0000 175.2400 5.2600 176.3200 ;
      RECT 0.0000 173.6000 240.1200 175.2400 ;
      RECT 238.8600 172.5200 240.1200 173.6000 ;
      RECT 193.6200 172.5200 235.2600 173.6000 ;
      RECT 148.6200 172.5200 192.0200 173.6000 ;
      RECT 103.6200 172.5200 147.0200 173.6000 ;
      RECT 58.6200 172.5200 102.0200 173.6000 ;
      RECT 13.6200 172.5200 57.0200 173.6000 ;
      RECT 4.8600 172.5200 12.0200 173.6000 ;
      RECT 0.0000 172.5200 1.2600 173.6000 ;
      RECT 0.0000 170.8800 240.1200 172.5200 ;
      RECT 234.8600 169.8000 240.1200 170.8800 ;
      RECT 191.4200 169.8000 231.2600 170.8800 ;
      RECT 146.4200 169.8000 189.8200 170.8800 ;
      RECT 101.4200 169.8000 144.8200 170.8800 ;
      RECT 56.4200 169.8000 99.8200 170.8800 ;
      RECT 8.8600 169.8000 54.8200 170.8800 ;
      RECT 0.0000 169.8000 5.2600 170.8800 ;
      RECT 0.0000 168.1600 240.1200 169.8000 ;
      RECT 238.8600 167.0800 240.1200 168.1600 ;
      RECT 193.6200 167.0800 235.2600 168.1600 ;
      RECT 148.6200 167.0800 192.0200 168.1600 ;
      RECT 103.6200 167.0800 147.0200 168.1600 ;
      RECT 58.6200 167.0800 102.0200 168.1600 ;
      RECT 13.6200 167.0800 57.0200 168.1600 ;
      RECT 4.8600 167.0800 12.0200 168.1600 ;
      RECT 0.0000 167.0800 1.2600 168.1600 ;
      RECT 0.0000 165.4400 240.1200 167.0800 ;
      RECT 234.8600 164.3600 240.1200 165.4400 ;
      RECT 191.4200 164.3600 231.2600 165.4400 ;
      RECT 146.4200 164.3600 189.8200 165.4400 ;
      RECT 101.4200 164.3600 144.8200 165.4400 ;
      RECT 56.4200 164.3600 99.8200 165.4400 ;
      RECT 8.8600 164.3600 54.8200 165.4400 ;
      RECT 0.0000 164.3600 5.2600 165.4400 ;
      RECT 0.0000 162.7200 240.1200 164.3600 ;
      RECT 238.8600 161.6400 240.1200 162.7200 ;
      RECT 193.6200 161.6400 235.2600 162.7200 ;
      RECT 148.6200 161.6400 192.0200 162.7200 ;
      RECT 103.6200 161.6400 147.0200 162.7200 ;
      RECT 58.6200 161.6400 102.0200 162.7200 ;
      RECT 13.6200 161.6400 57.0200 162.7200 ;
      RECT 4.8600 161.6400 12.0200 162.7200 ;
      RECT 0.0000 161.6400 1.2600 162.7200 ;
      RECT 0.0000 160.0000 240.1200 161.6400 ;
      RECT 234.8600 158.9200 240.1200 160.0000 ;
      RECT 191.4200 158.9200 231.2600 160.0000 ;
      RECT 146.4200 158.9200 189.8200 160.0000 ;
      RECT 101.4200 158.9200 144.8200 160.0000 ;
      RECT 56.4200 158.9200 99.8200 160.0000 ;
      RECT 8.8600 158.9200 54.8200 160.0000 ;
      RECT 0.0000 158.9200 5.2600 160.0000 ;
      RECT 0.0000 157.2800 240.1200 158.9200 ;
      RECT 238.8600 156.2000 240.1200 157.2800 ;
      RECT 193.6200 156.2000 235.2600 157.2800 ;
      RECT 148.6200 156.2000 192.0200 157.2800 ;
      RECT 103.6200 156.2000 147.0200 157.2800 ;
      RECT 58.6200 156.2000 102.0200 157.2800 ;
      RECT 13.6200 156.2000 57.0200 157.2800 ;
      RECT 4.8600 156.2000 12.0200 157.2800 ;
      RECT 0.0000 156.2000 1.2600 157.2800 ;
      RECT 0.0000 154.5600 240.1200 156.2000 ;
      RECT 234.8600 153.4800 240.1200 154.5600 ;
      RECT 191.4200 153.4800 231.2600 154.5600 ;
      RECT 146.4200 153.4800 189.8200 154.5600 ;
      RECT 101.4200 153.4800 144.8200 154.5600 ;
      RECT 56.4200 153.4800 99.8200 154.5600 ;
      RECT 8.8600 153.4800 54.8200 154.5600 ;
      RECT 0.0000 153.4800 5.2600 154.5600 ;
      RECT 0.0000 151.8400 240.1200 153.4800 ;
      RECT 238.8600 150.7600 240.1200 151.8400 ;
      RECT 193.6200 150.7600 235.2600 151.8400 ;
      RECT 148.6200 150.7600 192.0200 151.8400 ;
      RECT 103.6200 150.7600 147.0200 151.8400 ;
      RECT 58.6200 150.7600 102.0200 151.8400 ;
      RECT 13.6200 150.7600 57.0200 151.8400 ;
      RECT 4.8600 150.7600 12.0200 151.8400 ;
      RECT 0.0000 150.7600 1.2600 151.8400 ;
      RECT 0.0000 149.1200 240.1200 150.7600 ;
      RECT 234.8600 148.0400 240.1200 149.1200 ;
      RECT 191.4200 148.0400 231.2600 149.1200 ;
      RECT 146.4200 148.0400 189.8200 149.1200 ;
      RECT 101.4200 148.0400 144.8200 149.1200 ;
      RECT 56.4200 148.0400 99.8200 149.1200 ;
      RECT 8.8600 148.0400 54.8200 149.1200 ;
      RECT 0.0000 148.0400 5.2600 149.1200 ;
      RECT 0.0000 146.4000 240.1200 148.0400 ;
      RECT 238.8600 145.3200 240.1200 146.4000 ;
      RECT 193.6200 145.3200 235.2600 146.4000 ;
      RECT 148.6200 145.3200 192.0200 146.4000 ;
      RECT 103.6200 145.3200 147.0200 146.4000 ;
      RECT 58.6200 145.3200 102.0200 146.4000 ;
      RECT 13.6200 145.3200 57.0200 146.4000 ;
      RECT 4.8600 145.3200 12.0200 146.4000 ;
      RECT 0.0000 145.3200 1.2600 146.4000 ;
      RECT 0.0000 143.6800 240.1200 145.3200 ;
      RECT 234.8600 142.6000 240.1200 143.6800 ;
      RECT 191.4200 142.6000 231.2600 143.6800 ;
      RECT 146.4200 142.6000 189.8200 143.6800 ;
      RECT 101.4200 142.6000 144.8200 143.6800 ;
      RECT 56.4200 142.6000 99.8200 143.6800 ;
      RECT 8.8600 142.6000 54.8200 143.6800 ;
      RECT 0.0000 142.6000 5.2600 143.6800 ;
      RECT 0.0000 140.9600 240.1200 142.6000 ;
      RECT 238.8600 139.8800 240.1200 140.9600 ;
      RECT 193.6200 139.8800 235.2600 140.9600 ;
      RECT 148.6200 139.8800 192.0200 140.9600 ;
      RECT 103.6200 139.8800 147.0200 140.9600 ;
      RECT 58.6200 139.8800 102.0200 140.9600 ;
      RECT 13.6200 139.8800 57.0200 140.9600 ;
      RECT 4.8600 139.8800 12.0200 140.9600 ;
      RECT 0.0000 139.8800 1.2600 140.9600 ;
      RECT 0.0000 138.2400 240.1200 139.8800 ;
      RECT 234.8600 137.1600 240.1200 138.2400 ;
      RECT 191.4200 137.1600 231.2600 138.2400 ;
      RECT 146.4200 137.1600 189.8200 138.2400 ;
      RECT 101.4200 137.1600 144.8200 138.2400 ;
      RECT 56.4200 137.1600 99.8200 138.2400 ;
      RECT 8.8600 137.1600 54.8200 138.2400 ;
      RECT 0.0000 137.1600 5.2600 138.2400 ;
      RECT 0.0000 135.5200 240.1200 137.1600 ;
      RECT 238.8600 134.4400 240.1200 135.5200 ;
      RECT 193.6200 134.4400 235.2600 135.5200 ;
      RECT 148.6200 134.4400 192.0200 135.5200 ;
      RECT 103.6200 134.4400 147.0200 135.5200 ;
      RECT 58.6200 134.4400 102.0200 135.5200 ;
      RECT 13.6200 134.4400 57.0200 135.5200 ;
      RECT 4.8600 134.4400 12.0200 135.5200 ;
      RECT 0.0000 134.4400 1.2600 135.5200 ;
      RECT 0.0000 132.8000 240.1200 134.4400 ;
      RECT 234.8600 131.7200 240.1200 132.8000 ;
      RECT 191.4200 131.7200 231.2600 132.8000 ;
      RECT 146.4200 131.7200 189.8200 132.8000 ;
      RECT 101.4200 131.7200 144.8200 132.8000 ;
      RECT 56.4200 131.7200 99.8200 132.8000 ;
      RECT 8.8600 131.7200 54.8200 132.8000 ;
      RECT 0.0000 131.7200 5.2600 132.8000 ;
      RECT 0.0000 130.0800 240.1200 131.7200 ;
      RECT 238.8600 129.0000 240.1200 130.0800 ;
      RECT 193.6200 129.0000 235.2600 130.0800 ;
      RECT 148.6200 129.0000 192.0200 130.0800 ;
      RECT 103.6200 129.0000 147.0200 130.0800 ;
      RECT 58.6200 129.0000 102.0200 130.0800 ;
      RECT 13.6200 129.0000 57.0200 130.0800 ;
      RECT 4.8600 129.0000 12.0200 130.0800 ;
      RECT 0.0000 129.0000 1.2600 130.0800 ;
      RECT 0.0000 127.3600 240.1200 129.0000 ;
      RECT 234.8600 126.2800 240.1200 127.3600 ;
      RECT 191.4200 126.2800 231.2600 127.3600 ;
      RECT 146.4200 126.2800 189.8200 127.3600 ;
      RECT 101.4200 126.2800 144.8200 127.3600 ;
      RECT 56.4200 126.2800 99.8200 127.3600 ;
      RECT 8.8600 126.2800 54.8200 127.3600 ;
      RECT 0.0000 126.2800 5.2600 127.3600 ;
      RECT 0.0000 124.6400 240.1200 126.2800 ;
      RECT 238.8600 123.5600 240.1200 124.6400 ;
      RECT 193.6200 123.5600 235.2600 124.6400 ;
      RECT 148.6200 123.5600 192.0200 124.6400 ;
      RECT 103.6200 123.5600 147.0200 124.6400 ;
      RECT 58.6200 123.5600 102.0200 124.6400 ;
      RECT 13.6200 123.5600 57.0200 124.6400 ;
      RECT 4.8600 123.5600 12.0200 124.6400 ;
      RECT 0.0000 123.5600 1.2600 124.6400 ;
      RECT 0.0000 121.9200 240.1200 123.5600 ;
      RECT 234.8600 120.8400 240.1200 121.9200 ;
      RECT 191.4200 120.8400 231.2600 121.9200 ;
      RECT 146.4200 120.8400 189.8200 121.9200 ;
      RECT 101.4200 120.8400 144.8200 121.9200 ;
      RECT 56.4200 120.8400 99.8200 121.9200 ;
      RECT 8.8600 120.8400 54.8200 121.9200 ;
      RECT 0.0000 120.8400 5.2600 121.9200 ;
      RECT 0.0000 119.2000 240.1200 120.8400 ;
      RECT 238.8600 118.1200 240.1200 119.2000 ;
      RECT 193.6200 118.1200 235.2600 119.2000 ;
      RECT 148.6200 118.1200 192.0200 119.2000 ;
      RECT 103.6200 118.1200 147.0200 119.2000 ;
      RECT 58.6200 118.1200 102.0200 119.2000 ;
      RECT 13.6200 118.1200 57.0200 119.2000 ;
      RECT 4.8600 118.1200 12.0200 119.2000 ;
      RECT 0.0000 118.1200 1.2600 119.2000 ;
      RECT 0.0000 116.4800 240.1200 118.1200 ;
      RECT 234.8600 115.4000 240.1200 116.4800 ;
      RECT 191.4200 115.4000 231.2600 116.4800 ;
      RECT 146.4200 115.4000 189.8200 116.4800 ;
      RECT 101.4200 115.4000 144.8200 116.4800 ;
      RECT 56.4200 115.4000 99.8200 116.4800 ;
      RECT 8.8600 115.4000 54.8200 116.4800 ;
      RECT 0.0000 115.4000 5.2600 116.4800 ;
      RECT 0.0000 113.7600 240.1200 115.4000 ;
      RECT 238.8600 112.6800 240.1200 113.7600 ;
      RECT 193.6200 112.6800 235.2600 113.7600 ;
      RECT 148.6200 112.6800 192.0200 113.7600 ;
      RECT 103.6200 112.6800 147.0200 113.7600 ;
      RECT 58.6200 112.6800 102.0200 113.7600 ;
      RECT 13.6200 112.6800 57.0200 113.7600 ;
      RECT 4.8600 112.6800 12.0200 113.7600 ;
      RECT 0.0000 112.6800 1.2600 113.7600 ;
      RECT 0.0000 111.0400 240.1200 112.6800 ;
      RECT 234.8600 109.9600 240.1200 111.0400 ;
      RECT 191.4200 109.9600 231.2600 111.0400 ;
      RECT 146.4200 109.9600 189.8200 111.0400 ;
      RECT 101.4200 109.9600 144.8200 111.0400 ;
      RECT 56.4200 109.9600 99.8200 111.0400 ;
      RECT 8.8600 109.9600 54.8200 111.0400 ;
      RECT 0.0000 109.9600 5.2600 111.0400 ;
      RECT 0.0000 108.3200 240.1200 109.9600 ;
      RECT 238.8600 107.2400 240.1200 108.3200 ;
      RECT 193.6200 107.2400 235.2600 108.3200 ;
      RECT 148.6200 107.2400 192.0200 108.3200 ;
      RECT 103.6200 107.2400 147.0200 108.3200 ;
      RECT 58.6200 107.2400 102.0200 108.3200 ;
      RECT 13.6200 107.2400 57.0200 108.3200 ;
      RECT 4.8600 107.2400 12.0200 108.3200 ;
      RECT 0.0000 107.2400 1.2600 108.3200 ;
      RECT 0.0000 105.6000 240.1200 107.2400 ;
      RECT 234.8600 104.5200 240.1200 105.6000 ;
      RECT 191.4200 104.5200 231.2600 105.6000 ;
      RECT 146.4200 104.5200 189.8200 105.6000 ;
      RECT 101.4200 104.5200 144.8200 105.6000 ;
      RECT 56.4200 104.5200 99.8200 105.6000 ;
      RECT 8.8600 104.5200 54.8200 105.6000 ;
      RECT 0.0000 104.5200 5.2600 105.6000 ;
      RECT 0.0000 102.8800 240.1200 104.5200 ;
      RECT 238.8600 101.8000 240.1200 102.8800 ;
      RECT 193.6200 101.8000 235.2600 102.8800 ;
      RECT 148.6200 101.8000 192.0200 102.8800 ;
      RECT 103.6200 101.8000 147.0200 102.8800 ;
      RECT 58.6200 101.8000 102.0200 102.8800 ;
      RECT 13.6200 101.8000 57.0200 102.8800 ;
      RECT 4.8600 101.8000 12.0200 102.8800 ;
      RECT 0.0000 101.8000 1.2600 102.8800 ;
      RECT 0.0000 100.1600 240.1200 101.8000 ;
      RECT 234.8600 99.0800 240.1200 100.1600 ;
      RECT 191.4200 99.0800 231.2600 100.1600 ;
      RECT 146.4200 99.0800 189.8200 100.1600 ;
      RECT 101.4200 99.0800 144.8200 100.1600 ;
      RECT 56.4200 99.0800 99.8200 100.1600 ;
      RECT 8.8600 99.0800 54.8200 100.1600 ;
      RECT 0.0000 99.0800 5.2600 100.1600 ;
      RECT 0.0000 97.4400 240.1200 99.0800 ;
      RECT 238.8600 96.3600 240.1200 97.4400 ;
      RECT 193.6200 96.3600 235.2600 97.4400 ;
      RECT 148.6200 96.3600 192.0200 97.4400 ;
      RECT 103.6200 96.3600 147.0200 97.4400 ;
      RECT 58.6200 96.3600 102.0200 97.4400 ;
      RECT 13.6200 96.3600 57.0200 97.4400 ;
      RECT 4.8600 96.3600 12.0200 97.4400 ;
      RECT 0.0000 96.3600 1.2600 97.4400 ;
      RECT 0.0000 94.7200 240.1200 96.3600 ;
      RECT 234.8600 93.6400 240.1200 94.7200 ;
      RECT 191.4200 93.6400 231.2600 94.7200 ;
      RECT 146.4200 93.6400 189.8200 94.7200 ;
      RECT 101.4200 93.6400 144.8200 94.7200 ;
      RECT 56.4200 93.6400 99.8200 94.7200 ;
      RECT 8.8600 93.6400 54.8200 94.7200 ;
      RECT 0.0000 93.6400 5.2600 94.7200 ;
      RECT 0.0000 92.0000 240.1200 93.6400 ;
      RECT 238.8600 90.9200 240.1200 92.0000 ;
      RECT 193.6200 90.9200 235.2600 92.0000 ;
      RECT 148.6200 90.9200 192.0200 92.0000 ;
      RECT 103.6200 90.9200 147.0200 92.0000 ;
      RECT 58.6200 90.9200 102.0200 92.0000 ;
      RECT 13.6200 90.9200 57.0200 92.0000 ;
      RECT 4.8600 90.9200 12.0200 92.0000 ;
      RECT 0.0000 90.9200 1.2600 92.0000 ;
      RECT 0.0000 89.2800 240.1200 90.9200 ;
      RECT 234.8600 88.2000 240.1200 89.2800 ;
      RECT 191.4200 88.2000 231.2600 89.2800 ;
      RECT 146.4200 88.2000 189.8200 89.2800 ;
      RECT 101.4200 88.2000 144.8200 89.2800 ;
      RECT 56.4200 88.2000 99.8200 89.2800 ;
      RECT 8.8600 88.2000 54.8200 89.2800 ;
      RECT 0.0000 88.2000 5.2600 89.2800 ;
      RECT 0.0000 86.5600 240.1200 88.2000 ;
      RECT 238.8600 85.4800 240.1200 86.5600 ;
      RECT 193.6200 85.4800 235.2600 86.5600 ;
      RECT 148.6200 85.4800 192.0200 86.5600 ;
      RECT 103.6200 85.4800 147.0200 86.5600 ;
      RECT 58.6200 85.4800 102.0200 86.5600 ;
      RECT 13.6200 85.4800 57.0200 86.5600 ;
      RECT 4.8600 85.4800 12.0200 86.5600 ;
      RECT 0.0000 85.4800 1.2600 86.5600 ;
      RECT 0.0000 83.8400 240.1200 85.4800 ;
      RECT 234.8600 82.7600 240.1200 83.8400 ;
      RECT 191.4200 82.7600 231.2600 83.8400 ;
      RECT 146.4200 82.7600 189.8200 83.8400 ;
      RECT 101.4200 82.7600 144.8200 83.8400 ;
      RECT 56.4200 82.7600 99.8200 83.8400 ;
      RECT 8.8600 82.7600 54.8200 83.8400 ;
      RECT 0.0000 82.7600 5.2600 83.8400 ;
      RECT 0.0000 81.1200 240.1200 82.7600 ;
      RECT 238.8600 80.0400 240.1200 81.1200 ;
      RECT 193.6200 80.0400 235.2600 81.1200 ;
      RECT 148.6200 80.0400 192.0200 81.1200 ;
      RECT 103.6200 80.0400 147.0200 81.1200 ;
      RECT 58.6200 80.0400 102.0200 81.1200 ;
      RECT 13.6200 80.0400 57.0200 81.1200 ;
      RECT 4.8600 80.0400 12.0200 81.1200 ;
      RECT 0.0000 80.0400 1.2600 81.1200 ;
      RECT 0.0000 78.4000 240.1200 80.0400 ;
      RECT 234.8600 77.3200 240.1200 78.4000 ;
      RECT 191.4200 77.3200 231.2600 78.4000 ;
      RECT 146.4200 77.3200 189.8200 78.4000 ;
      RECT 101.4200 77.3200 144.8200 78.4000 ;
      RECT 56.4200 77.3200 99.8200 78.4000 ;
      RECT 8.8600 77.3200 54.8200 78.4000 ;
      RECT 0.0000 77.3200 5.2600 78.4000 ;
      RECT 0.0000 75.6800 240.1200 77.3200 ;
      RECT 238.8600 74.6000 240.1200 75.6800 ;
      RECT 193.6200 74.6000 235.2600 75.6800 ;
      RECT 148.6200 74.6000 192.0200 75.6800 ;
      RECT 103.6200 74.6000 147.0200 75.6800 ;
      RECT 58.6200 74.6000 102.0200 75.6800 ;
      RECT 13.6200 74.6000 57.0200 75.6800 ;
      RECT 4.8600 74.6000 12.0200 75.6800 ;
      RECT 0.0000 74.6000 1.2600 75.6800 ;
      RECT 0.0000 72.9600 240.1200 74.6000 ;
      RECT 234.8600 71.8800 240.1200 72.9600 ;
      RECT 191.4200 71.8800 231.2600 72.9600 ;
      RECT 146.4200 71.8800 189.8200 72.9600 ;
      RECT 101.4200 71.8800 144.8200 72.9600 ;
      RECT 56.4200 71.8800 99.8200 72.9600 ;
      RECT 8.8600 71.8800 54.8200 72.9600 ;
      RECT 0.0000 71.8800 5.2600 72.9600 ;
      RECT 0.0000 70.2400 240.1200 71.8800 ;
      RECT 238.8600 69.1600 240.1200 70.2400 ;
      RECT 193.6200 69.1600 235.2600 70.2400 ;
      RECT 148.6200 69.1600 192.0200 70.2400 ;
      RECT 103.6200 69.1600 147.0200 70.2400 ;
      RECT 58.6200 69.1600 102.0200 70.2400 ;
      RECT 13.6200 69.1600 57.0200 70.2400 ;
      RECT 4.8600 69.1600 12.0200 70.2400 ;
      RECT 0.0000 69.1600 1.2600 70.2400 ;
      RECT 0.0000 67.5200 240.1200 69.1600 ;
      RECT 234.8600 66.4400 240.1200 67.5200 ;
      RECT 191.4200 66.4400 231.2600 67.5200 ;
      RECT 146.4200 66.4400 189.8200 67.5200 ;
      RECT 101.4200 66.4400 144.8200 67.5200 ;
      RECT 56.4200 66.4400 99.8200 67.5200 ;
      RECT 8.8600 66.4400 54.8200 67.5200 ;
      RECT 0.0000 66.4400 5.2600 67.5200 ;
      RECT 0.0000 64.8000 240.1200 66.4400 ;
      RECT 238.8600 63.7200 240.1200 64.8000 ;
      RECT 193.6200 63.7200 235.2600 64.8000 ;
      RECT 148.6200 63.7200 192.0200 64.8000 ;
      RECT 103.6200 63.7200 147.0200 64.8000 ;
      RECT 58.6200 63.7200 102.0200 64.8000 ;
      RECT 13.6200 63.7200 57.0200 64.8000 ;
      RECT 4.8600 63.7200 12.0200 64.8000 ;
      RECT 0.0000 63.7200 1.2600 64.8000 ;
      RECT 0.0000 62.0800 240.1200 63.7200 ;
      RECT 234.8600 61.0000 240.1200 62.0800 ;
      RECT 191.4200 61.0000 231.2600 62.0800 ;
      RECT 146.4200 61.0000 189.8200 62.0800 ;
      RECT 101.4200 61.0000 144.8200 62.0800 ;
      RECT 56.4200 61.0000 99.8200 62.0800 ;
      RECT 8.8600 61.0000 54.8200 62.0800 ;
      RECT 0.0000 61.0000 5.2600 62.0800 ;
      RECT 0.0000 59.3600 240.1200 61.0000 ;
      RECT 238.8600 58.2800 240.1200 59.3600 ;
      RECT 193.6200 58.2800 235.2600 59.3600 ;
      RECT 148.6200 58.2800 192.0200 59.3600 ;
      RECT 103.6200 58.2800 147.0200 59.3600 ;
      RECT 58.6200 58.2800 102.0200 59.3600 ;
      RECT 13.6200 58.2800 57.0200 59.3600 ;
      RECT 4.8600 58.2800 12.0200 59.3600 ;
      RECT 0.0000 58.2800 1.2600 59.3600 ;
      RECT 0.0000 56.6400 240.1200 58.2800 ;
      RECT 234.8600 55.5600 240.1200 56.6400 ;
      RECT 191.4200 55.5600 231.2600 56.6400 ;
      RECT 146.4200 55.5600 189.8200 56.6400 ;
      RECT 101.4200 55.5600 144.8200 56.6400 ;
      RECT 56.4200 55.5600 99.8200 56.6400 ;
      RECT 8.8600 55.5600 54.8200 56.6400 ;
      RECT 0.0000 55.5600 5.2600 56.6400 ;
      RECT 0.0000 53.9200 240.1200 55.5600 ;
      RECT 238.8600 52.8400 240.1200 53.9200 ;
      RECT 193.6200 52.8400 235.2600 53.9200 ;
      RECT 148.6200 52.8400 192.0200 53.9200 ;
      RECT 103.6200 52.8400 147.0200 53.9200 ;
      RECT 58.6200 52.8400 102.0200 53.9200 ;
      RECT 13.6200 52.8400 57.0200 53.9200 ;
      RECT 4.8600 52.8400 12.0200 53.9200 ;
      RECT 0.0000 52.8400 1.2600 53.9200 ;
      RECT 0.0000 51.2000 240.1200 52.8400 ;
      RECT 234.8600 50.1200 240.1200 51.2000 ;
      RECT 191.4200 50.1200 231.2600 51.2000 ;
      RECT 146.4200 50.1200 189.8200 51.2000 ;
      RECT 101.4200 50.1200 144.8200 51.2000 ;
      RECT 56.4200 50.1200 99.8200 51.2000 ;
      RECT 8.8600 50.1200 54.8200 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 240.1200 50.1200 ;
      RECT 238.8600 47.4000 240.1200 48.4800 ;
      RECT 193.6200 47.4000 235.2600 48.4800 ;
      RECT 148.6200 47.4000 192.0200 48.4800 ;
      RECT 103.6200 47.4000 147.0200 48.4800 ;
      RECT 58.6200 47.4000 102.0200 48.4800 ;
      RECT 13.6200 47.4000 57.0200 48.4800 ;
      RECT 4.8600 47.4000 12.0200 48.4800 ;
      RECT 0.0000 47.4000 1.2600 48.4800 ;
      RECT 0.0000 45.7600 240.1200 47.4000 ;
      RECT 234.8600 44.6800 240.1200 45.7600 ;
      RECT 191.4200 44.6800 231.2600 45.7600 ;
      RECT 146.4200 44.6800 189.8200 45.7600 ;
      RECT 101.4200 44.6800 144.8200 45.7600 ;
      RECT 56.4200 44.6800 99.8200 45.7600 ;
      RECT 8.8600 44.6800 54.8200 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 240.1200 44.6800 ;
      RECT 238.8600 41.9600 240.1200 43.0400 ;
      RECT 193.6200 41.9600 235.2600 43.0400 ;
      RECT 148.6200 41.9600 192.0200 43.0400 ;
      RECT 103.6200 41.9600 147.0200 43.0400 ;
      RECT 58.6200 41.9600 102.0200 43.0400 ;
      RECT 13.6200 41.9600 57.0200 43.0400 ;
      RECT 4.8600 41.9600 12.0200 43.0400 ;
      RECT 0.0000 41.9600 1.2600 43.0400 ;
      RECT 0.0000 40.3200 240.1200 41.9600 ;
      RECT 234.8600 39.2400 240.1200 40.3200 ;
      RECT 191.4200 39.2400 231.2600 40.3200 ;
      RECT 146.4200 39.2400 189.8200 40.3200 ;
      RECT 101.4200 39.2400 144.8200 40.3200 ;
      RECT 56.4200 39.2400 99.8200 40.3200 ;
      RECT 8.8600 39.2400 54.8200 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 240.1200 39.2400 ;
      RECT 238.8600 36.5200 240.1200 37.6000 ;
      RECT 193.6200 36.5200 235.2600 37.6000 ;
      RECT 148.6200 36.5200 192.0200 37.6000 ;
      RECT 103.6200 36.5200 147.0200 37.6000 ;
      RECT 58.6200 36.5200 102.0200 37.6000 ;
      RECT 13.6200 36.5200 57.0200 37.6000 ;
      RECT 4.8600 36.5200 12.0200 37.6000 ;
      RECT 0.0000 36.5200 1.2600 37.6000 ;
      RECT 0.0000 34.8800 240.1200 36.5200 ;
      RECT 234.8600 33.8000 240.1200 34.8800 ;
      RECT 191.4200 33.8000 231.2600 34.8800 ;
      RECT 146.4200 33.8000 189.8200 34.8800 ;
      RECT 101.4200 33.8000 144.8200 34.8800 ;
      RECT 56.4200 33.8000 99.8200 34.8800 ;
      RECT 8.8600 33.8000 54.8200 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 240.1200 33.8000 ;
      RECT 238.8600 31.0800 240.1200 32.1600 ;
      RECT 193.6200 31.0800 235.2600 32.1600 ;
      RECT 148.6200 31.0800 192.0200 32.1600 ;
      RECT 103.6200 31.0800 147.0200 32.1600 ;
      RECT 58.6200 31.0800 102.0200 32.1600 ;
      RECT 13.6200 31.0800 57.0200 32.1600 ;
      RECT 4.8600 31.0800 12.0200 32.1600 ;
      RECT 0.0000 31.0800 1.2600 32.1600 ;
      RECT 0.0000 29.4400 240.1200 31.0800 ;
      RECT 234.8600 28.3600 240.1200 29.4400 ;
      RECT 191.4200 28.3600 231.2600 29.4400 ;
      RECT 146.4200 28.3600 189.8200 29.4400 ;
      RECT 101.4200 28.3600 144.8200 29.4400 ;
      RECT 56.4200 28.3600 99.8200 29.4400 ;
      RECT 8.8600 28.3600 54.8200 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 240.1200 28.3600 ;
      RECT 238.8600 25.6400 240.1200 26.7200 ;
      RECT 193.6200 25.6400 235.2600 26.7200 ;
      RECT 148.6200 25.6400 192.0200 26.7200 ;
      RECT 103.6200 25.6400 147.0200 26.7200 ;
      RECT 58.6200 25.6400 102.0200 26.7200 ;
      RECT 13.6200 25.6400 57.0200 26.7200 ;
      RECT 4.8600 25.6400 12.0200 26.7200 ;
      RECT 0.0000 25.6400 1.2600 26.7200 ;
      RECT 0.0000 24.0000 240.1200 25.6400 ;
      RECT 234.8600 22.9200 240.1200 24.0000 ;
      RECT 191.4200 22.9200 231.2600 24.0000 ;
      RECT 146.4200 22.9200 189.8200 24.0000 ;
      RECT 101.4200 22.9200 144.8200 24.0000 ;
      RECT 56.4200 22.9200 99.8200 24.0000 ;
      RECT 8.8600 22.9200 54.8200 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 240.1200 22.9200 ;
      RECT 238.8600 20.2000 240.1200 21.2800 ;
      RECT 193.6200 20.2000 235.2600 21.2800 ;
      RECT 148.6200 20.2000 192.0200 21.2800 ;
      RECT 103.6200 20.2000 147.0200 21.2800 ;
      RECT 58.6200 20.2000 102.0200 21.2800 ;
      RECT 13.6200 20.2000 57.0200 21.2800 ;
      RECT 4.8600 20.2000 12.0200 21.2800 ;
      RECT 0.0000 20.2000 1.2600 21.2800 ;
      RECT 0.0000 18.5600 240.1200 20.2000 ;
      RECT 234.8600 17.4800 240.1200 18.5600 ;
      RECT 191.4200 17.4800 231.2600 18.5600 ;
      RECT 146.4200 17.4800 189.8200 18.5600 ;
      RECT 101.4200 17.4800 144.8200 18.5600 ;
      RECT 56.4200 17.4800 99.8200 18.5600 ;
      RECT 8.8600 17.4800 54.8200 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 240.1200 17.4800 ;
      RECT 238.8600 14.7600 240.1200 15.8400 ;
      RECT 193.6200 14.7600 235.2600 15.8400 ;
      RECT 148.6200 14.7600 192.0200 15.8400 ;
      RECT 103.6200 14.7600 147.0200 15.8400 ;
      RECT 58.6200 14.7600 102.0200 15.8400 ;
      RECT 13.6200 14.7600 57.0200 15.8400 ;
      RECT 4.8600 14.7600 12.0200 15.8400 ;
      RECT 0.0000 14.7600 1.2600 15.8400 ;
      RECT 0.0000 13.1200 240.1200 14.7600 ;
      RECT 234.8600 12.0400 240.1200 13.1200 ;
      RECT 191.4200 12.0400 231.2600 13.1200 ;
      RECT 146.4200 12.0400 189.8200 13.1200 ;
      RECT 101.4200 12.0400 144.8200 13.1200 ;
      RECT 56.4200 12.0400 99.8200 13.1200 ;
      RECT 8.8600 12.0400 54.8200 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 240.1200 12.0400 ;
      RECT 238.8600 9.3200 240.1200 10.4000 ;
      RECT 193.6200 9.3200 235.2600 10.4000 ;
      RECT 148.6200 9.3200 192.0200 10.4000 ;
      RECT 103.6200 9.3200 147.0200 10.4000 ;
      RECT 58.6200 9.3200 102.0200 10.4000 ;
      RECT 13.6200 9.3200 57.0200 10.4000 ;
      RECT 4.8600 9.3200 12.0200 10.4000 ;
      RECT 0.0000 9.3200 1.2600 10.4000 ;
      RECT 0.0000 8.7300 240.1200 9.3200 ;
      RECT 234.8600 5.1300 240.1200 8.7300 ;
      RECT 0.0000 5.1300 5.2600 8.7300 ;
      RECT 0.0000 4.7300 240.1200 5.1300 ;
      RECT 238.8600 1.1300 240.1200 4.7300 ;
      RECT 0.0000 1.1300 1.2600 4.7300 ;
      RECT 0.0000 0.0000 240.1200 1.1300 ;
    LAYER met4 ;
      RECT 0.0000 217.8300 240.1200 219.6400 ;
      RECT 193.6200 213.8300 235.2600 217.8300 ;
      RECT 148.6200 213.8300 192.0200 217.8300 ;
      RECT 103.6200 213.8300 147.0200 217.8300 ;
      RECT 58.6200 213.8300 102.0200 217.8300 ;
      RECT 13.6200 213.8300 57.0200 217.8300 ;
      RECT 4.8600 213.8300 12.0200 217.8300 ;
      RECT 234.8600 5.1300 235.2600 213.8300 ;
      RECT 193.6200 5.1300 231.2600 213.8300 ;
      RECT 191.4200 5.1300 192.0200 213.8300 ;
      RECT 148.6200 5.1300 189.8200 213.8300 ;
      RECT 146.4200 5.1300 147.0200 213.8300 ;
      RECT 103.6200 5.1300 144.8200 213.8300 ;
      RECT 101.4200 5.1300 102.0200 213.8300 ;
      RECT 58.6200 5.1300 99.8200 213.8300 ;
      RECT 56.4200 5.1300 57.0200 213.8300 ;
      RECT 13.6200 5.1300 54.8200 213.8300 ;
      RECT 8.8600 5.1300 12.0200 213.8300 ;
      RECT 4.8600 5.1300 5.2600 213.8300 ;
      RECT 238.8600 1.1300 240.1200 217.8300 ;
      RECT 193.6200 1.1300 235.2600 5.1300 ;
      RECT 148.6200 1.1300 192.0200 5.1300 ;
      RECT 103.6200 1.1300 147.0200 5.1300 ;
      RECT 58.6200 1.1300 102.0200 5.1300 ;
      RECT 13.6200 1.1300 57.0200 5.1300 ;
      RECT 4.8600 1.1300 12.0200 5.1300 ;
      RECT 0.0000 1.1300 1.2600 217.8300 ;
      RECT 0.0000 1.0200 240.1200 1.1300 ;
      RECT 90.1900 0.0000 240.1200 1.0200 ;
      RECT 0.0000 0.0000 89.2100 1.0200 ;
    LAYER met5 ;
      RECT 0.0000 0.0000 240.1200 219.6400 ;
  END
END RegFile

END LIBRARY
