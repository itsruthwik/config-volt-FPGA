##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 01:17:29 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO N_term_RAM_IO
  CLASS BLOCK ;
  SIZE 100.2800 BY 30.2600 ;
  FOREIGN N_term_RAM_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.34855 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.763 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 46.1437 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 243.868 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 7.8600 0.0000 8.2400 0.7200 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.66055 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.483 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.3884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 44.5381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 218.242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 6.9400 0.0000 7.3200 0.7200 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.31415 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.899 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.4739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.9214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 6.0200 0.0000 6.4000 0.7200 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.40675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.785 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 11.923 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 56.1635 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 5.1000 0.0000 5.4800 0.7200 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.2628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.897 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 38.2418 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 202.931 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 0.0000 16.9800 0.7200 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.902 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 39.6236 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 192.928 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 0.0000 15.6000 0.7200 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.714 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2009 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.9811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 14.3000 0.0000 14.6800 0.7200 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4836 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.572 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.0248 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.2956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 13.3800 0.0000 13.7600 0.7200 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.05995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5232 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 61.9462 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.72 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 12.0000 0.0000 12.3800 0.7200 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 21.055 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 114.447 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 0.0000 11.4600 0.7200 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.46455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7242 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 5.38082 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 23.4528 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 0.0000 10.5400 0.7200 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.79095 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.107 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.783 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 18.2097 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 87.5975 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 9.2400 0.0000 9.6200 0.7200 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.606 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.84 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 0.0000 25.2600 0.7200 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.40375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.475 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.8656 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.418 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.2739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.9214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 23.9600 0.0000 24.3400 0.7200 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.9128 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.328 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 45.7871 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 223.745 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 22.5800 0.0000 22.9600 0.7200 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6229 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 47.3777 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.082 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 21.6600 0.0000 22.0400 0.7200 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1852 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.7481 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 113.55 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 0.0000 21.1200 0.7200 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.50283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.4906 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 0.0000 19.7400 0.7200 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.20975 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.0252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 18.4400 0.0000 18.8200 0.7200 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.5404 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.6245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0072 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.0126 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 17.5200 0.0000 17.9000 0.7200 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.568 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.084 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5846 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.4748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 41.4400 0.0000 41.8200 0.7200 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75055 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.883 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.61226 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.0377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 40.5200 0.0000 40.9000 0.7200 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 48.8645 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.204 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 0.0000 39.9800 0.7200 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.37201 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.4119 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 38.6800 0.0000 39.0600 0.7200 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.494 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.4465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 37.3000 0.0000 37.6800 0.7200 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.10157 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.4843 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 36.3800 0.0000 36.7600 0.7200 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.07642 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.934 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 0.0000 35.8400 0.7200 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.39088 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.5063 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 0.0000 34.4600 0.7200 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.37 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.9267 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.186 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 0.0000 33.5400 0.7200 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.36195 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.3616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 32.2400 0.0000 32.6200 0.7200 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.31 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.5 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 31.3200 0.0000 31.7000 0.7200 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.014 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 46.4877 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 214.173 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 29.9400 0.0000 30.3200 0.7200 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.608 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5619 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.3365 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 0.0000 29.4000 0.7200 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.28019 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.9528 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 28.1000 0.0000 28.4800 0.7200 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.59 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 32.6852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 158.236 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 26.7200 0.0000 27.1000 0.7200 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 46.167 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 226.387 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 25.8000 0.0000 26.1800 0.7200 ;
    END
  END N4END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.5800 0.0000 45.9600 0.7200 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.17555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.238 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 44.6600 0.0000 45.0400 0.7200 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.142 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 0.0000 44.1200 0.7200 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 42.8200 0.0000 43.2000 0.7200 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.89 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 0.0000 62.9800 0.7200 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.5065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.6800 0.0000 62.0600 0.7200 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 60.3000 0.0000 60.6800 0.7200 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 59.3800 0.0000 59.7600 0.7200 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.17555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 0.0000 58.8400 0.7200 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.3398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.616 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 57.5400 0.0000 57.9200 0.7200 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 0.0000 56.5400 0.7200 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.778 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.228 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 55.2400 0.0000 55.6200 0.7200 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.074 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 54.3200 0.0000 54.7000 0.7200 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.80835 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.951 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4738 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.2915 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.9400 0.0000 53.3200 0.7200 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 0.0000 52.4000 0.7200 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.63 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 51.1000 0.0000 51.4800 0.7200 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.1800 0.0000 50.5600 0.7200 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 48.8000 0.0000 49.1800 0.7200 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 0.0000 48.2600 0.7200 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.68 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 46.9600 0.0000 47.3400 0.7200 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.17555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 0.0000 79.5400 0.7200 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 78.2400 0.0000 78.6200 0.7200 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.3200 0.0000 77.7000 0.7200 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.1928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.832 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 0.0000 76.7800 0.7200 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 0.0000 75.4000 0.7200 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.942 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 74.1000 0.0000 74.4800 0.7200 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.048 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.1800 0.0000 73.5600 0.7200 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 0.0000 72.6400 0.7200 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.084 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 0.0000 71.2600 0.7200 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.9600 0.0000 70.3400 0.7200 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.0400 0.0000 69.4200 0.7200 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 67.6600 0.0000 68.0400 0.7200 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 0.0000 67.1200 0.7200 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.8200 0.0000 66.2000 0.7200 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01915 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.199 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 64.9000 0.0000 65.2800 0.7200 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96135 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6229 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 63.5200 0.0000 63.9000 0.7200 ;
    END
  END S4BEG[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.34 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.512 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8362 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.7327 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.5704 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.7005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.0063 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.75 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.5041 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.4969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.618 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.9619 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.3616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.9959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 115.531 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4828 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.568 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.7272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.55 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.3695 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.0818 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.002 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.31038 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.1038 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.658 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.7934 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.0346 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2372 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.4452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.1485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.442 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.2421 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.207 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 33.0582 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.358 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.312 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.6261 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.9403 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3616 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 75.7425 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.962 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.68 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 39.1978 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.308 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.34 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.1348 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.5595 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.66384 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.8805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.72505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.853 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.934 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 46.2997 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.179 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.493 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9871 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.8176 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.31 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.4245 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.592 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.40975 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.3459 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.608 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9066 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.4057 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.2026 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 43.5274 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.421 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.5818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 59.0808 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.255 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 54.4934 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.818 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.242 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 65.9991 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.34 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.8688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 80.4821 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 421.277 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 11.2019 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 63.2233 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.594 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 33.9393 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.531 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 50.9752 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.138 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.022 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.5041 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.942 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.7645 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.9528 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.386 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.4324 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.233 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.37 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 22.5299 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 119.069 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.087 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 28.6600 100.2800 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.421 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 26.6200 100.2800 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.381 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.5198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.576 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 24.9200 100.2800 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 22.8800 100.2800 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.919 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 21.1800 100.2800 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 19.1400 100.2800 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.3285 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 17.4400 100.2800 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 15.7400 100.2800 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 13.7000 100.2800 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.9498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.536 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 12.0000 100.2800 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.2706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.384 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 10.3000 100.2800 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 8.2600 100.2800 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.4796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 6.5600 100.2800 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4345 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 4.5200 100.2800 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 2.8200 100.2800 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 1.1200 100.2800 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 27.6250 100.2800 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7825 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 25.9250 100.2800 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.653 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 58.1875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 24.2250 100.2800 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.617 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 57.9705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.486 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 22.5250 100.2800 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5984 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.704 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.5472 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.238 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 20.8250 100.2800 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.698 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 19.1250 100.2800 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.521 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2824 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.375 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 17.4250 100.2800 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.312 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 15.7250 100.2800 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.62 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.9956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 14.0250 100.2800 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8874 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.044 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.3468 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.697 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 12.3250 100.2800 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 10.6250 100.2800 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.907 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.8586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.52 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 8.9250 100.2800 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.4706 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2755 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.286 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 7.2250 100.2800 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7438 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.228 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.6356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.141 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 5.5250 100.2800 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2708 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.2395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.538 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 3.8250 100.2800 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5406 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.636 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.28 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 2.1250 100.2800 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.878 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.6362 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.311 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 97.5600 0.0000 97.9400 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.353 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.1858 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.4811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 96.6400 0.0000 97.0200 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.547 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 32.9016 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 159.381 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 95.7200 0.0000 96.1000 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.215 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1079 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.6698 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.8000 0.0000 95.1800 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.7448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 74.3689 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 392.547 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 93.8800 0.0000 94.2600 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.523 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.1909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.9600 0.0000 93.3400 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1158 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 33.5242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 162.176 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.0400 0.0000 92.4200 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.259 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 28.1921 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 136.575 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.1200 0.0000 91.5000 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.569 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.6978 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.1038 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.2000 0.0000 90.5800 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.451 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.5884 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.557 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 89.2800 0.0000 89.6600 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5682 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.7138 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 88.3600 0.0000 88.7400 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.127 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3915 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.701 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 87.4400 0.0000 87.8200 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9793 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 87.1802 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 463.242 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.5200 0.0000 86.9000 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.917 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5783 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.7642 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 85.6000 0.0000 85.9800 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0193 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.63 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 42.3575 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 228.327 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 84.6800 0.0000 85.0600 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.357 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 40.289 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 196.318 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 83.7600 0.0000 84.1400 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.1928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 69.0657 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 364.874 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 82.3800 0.0000 82.7600 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.237 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.5600 29.5400 97.9400 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.333 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.6400 29.5400 97.0200 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.96 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 95.7200 29.5400 96.1000 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.8000 29.5400 95.1800 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9142 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.345 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 93.8800 29.5400 94.2600 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.037 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 92.9600 29.5400 93.3400 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.0400 29.5400 92.4200 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.686 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.1200 29.5400 91.5000 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.747 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.2000 29.5400 90.5800 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.201 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.2800 29.5400 89.6600 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.3600 29.5400 88.7400 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1378 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.463 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 87.4400 29.5400 87.8200 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.691 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.5200 29.5400 86.9000 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6354 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.069 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 85.6000 29.5400 85.9800 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.011 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.6800 29.5400 85.0600 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.011 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.7600 29.5400 84.1400 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.465 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.3800 29.5400 82.7600 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 94.7200 6.0700 ;
        RECT 5.5600 23.0000 94.7200 25.0000 ;
        RECT 92.7200 15.0600 94.7200 15.5400 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 92.7200 9.6200 94.7200 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 92.7200 20.5000 94.7200 20.9800 ;
      LAYER met4 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
        RECT 92.7200 4.0700 94.7200 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 97.7200 3.0700 ;
        RECT 2.5600 26.0000 97.7200 28.0000 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 95.7200 12.3400 97.7200 12.8200 ;
        RECT 95.7200 6.9000 97.7200 7.3800 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 95.7200 17.7800 97.7200 18.2600 ;
      LAYER met4 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
        RECT 95.7200 1.0700 97.7200 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.0000 28.9850 100.2800 30.2600 ;
      RECT 0.5000 28.4750 100.2800 28.9850 ;
      RECT 0.0000 27.9650 100.2800 28.4750 ;
      RECT 0.0000 27.4550 99.7800 27.9650 ;
      RECT 0.0000 26.9450 100.2800 27.4550 ;
      RECT 0.5000 26.4350 100.2800 26.9450 ;
      RECT 0.0000 26.2650 100.2800 26.4350 ;
      RECT 0.0000 25.7550 99.7800 26.2650 ;
      RECT 0.0000 25.2450 100.2800 25.7550 ;
      RECT 0.5000 24.7350 100.2800 25.2450 ;
      RECT 0.0000 24.5650 100.2800 24.7350 ;
      RECT 0.0000 24.0550 99.7800 24.5650 ;
      RECT 0.0000 23.2050 100.2800 24.0550 ;
      RECT 0.5000 22.8650 100.2800 23.2050 ;
      RECT 0.5000 22.6950 99.7800 22.8650 ;
      RECT 0.0000 22.3550 99.7800 22.6950 ;
      RECT 0.0000 21.5050 100.2800 22.3550 ;
      RECT 0.5000 21.1650 100.2800 21.5050 ;
      RECT 0.5000 20.9950 99.7800 21.1650 ;
      RECT 0.0000 20.6550 99.7800 20.9950 ;
      RECT 0.0000 19.4650 100.2800 20.6550 ;
      RECT 0.5000 18.9550 99.7800 19.4650 ;
      RECT 0.0000 17.7650 100.2800 18.9550 ;
      RECT 0.5000 17.2550 99.7800 17.7650 ;
      RECT 0.0000 16.0650 100.2800 17.2550 ;
      RECT 0.5000 15.5550 99.7800 16.0650 ;
      RECT 0.0000 14.3650 100.2800 15.5550 ;
      RECT 0.0000 14.0250 99.7800 14.3650 ;
      RECT 0.5000 13.8550 99.7800 14.0250 ;
      RECT 0.5000 13.5150 100.2800 13.8550 ;
      RECT 0.0000 12.6650 100.2800 13.5150 ;
      RECT 0.0000 12.3250 99.7800 12.6650 ;
      RECT 0.5000 12.1550 99.7800 12.3250 ;
      RECT 0.5000 11.8150 100.2800 12.1550 ;
      RECT 0.0000 10.9650 100.2800 11.8150 ;
      RECT 0.0000 10.6250 99.7800 10.9650 ;
      RECT 0.5000 10.4550 99.7800 10.6250 ;
      RECT 0.5000 10.1150 100.2800 10.4550 ;
      RECT 0.0000 9.2650 100.2800 10.1150 ;
      RECT 0.0000 8.7550 99.7800 9.2650 ;
      RECT 0.0000 8.5850 100.2800 8.7550 ;
      RECT 0.5000 8.0750 100.2800 8.5850 ;
      RECT 0.0000 7.5650 100.2800 8.0750 ;
      RECT 0.0000 7.0550 99.7800 7.5650 ;
      RECT 0.0000 6.8850 100.2800 7.0550 ;
      RECT 0.5000 6.3750 100.2800 6.8850 ;
      RECT 0.0000 5.8650 100.2800 6.3750 ;
      RECT 0.0000 5.3550 99.7800 5.8650 ;
      RECT 0.0000 4.8450 100.2800 5.3550 ;
      RECT 0.5000 4.3350 100.2800 4.8450 ;
      RECT 0.0000 4.1650 100.2800 4.3350 ;
      RECT 0.0000 3.6550 99.7800 4.1650 ;
      RECT 0.0000 3.1450 100.2800 3.6550 ;
      RECT 0.5000 2.6350 100.2800 3.1450 ;
      RECT 0.0000 2.4650 100.2800 2.6350 ;
      RECT 0.0000 1.9550 99.7800 2.4650 ;
      RECT 0.0000 1.4450 100.2800 1.9550 ;
      RECT 0.5000 0.9350 100.2800 1.4450 ;
      RECT 0.0000 0.8900 100.2800 0.9350 ;
      RECT 79.7100 0.0000 100.2800 0.8900 ;
      RECT 78.7900 0.0000 78.9900 0.8900 ;
      RECT 77.8700 0.0000 78.0700 0.8900 ;
      RECT 76.9500 0.0000 77.1500 0.8900 ;
      RECT 75.5700 0.0000 76.2300 0.8900 ;
      RECT 74.6500 0.0000 74.8500 0.8900 ;
      RECT 73.7300 0.0000 73.9300 0.8900 ;
      RECT 72.8100 0.0000 73.0100 0.8900 ;
      RECT 71.4300 0.0000 72.0900 0.8900 ;
      RECT 70.5100 0.0000 70.7100 0.8900 ;
      RECT 69.5900 0.0000 69.7900 0.8900 ;
      RECT 68.2100 0.0000 68.8700 0.8900 ;
      RECT 67.2900 0.0000 67.4900 0.8900 ;
      RECT 66.3700 0.0000 66.5700 0.8900 ;
      RECT 65.4500 0.0000 65.6500 0.8900 ;
      RECT 64.0700 0.0000 64.7300 0.8900 ;
      RECT 63.1500 0.0000 63.3500 0.8900 ;
      RECT 62.2300 0.0000 62.4300 0.8900 ;
      RECT 60.8500 0.0000 61.5100 0.8900 ;
      RECT 59.9300 0.0000 60.1300 0.8900 ;
      RECT 59.0100 0.0000 59.2100 0.8900 ;
      RECT 58.0900 0.0000 58.2900 0.8900 ;
      RECT 56.7100 0.0000 57.3700 0.8900 ;
      RECT 55.7900 0.0000 55.9900 0.8900 ;
      RECT 54.8700 0.0000 55.0700 0.8900 ;
      RECT 53.4900 0.0000 54.1500 0.8900 ;
      RECT 52.5700 0.0000 52.7700 0.8900 ;
      RECT 51.6500 0.0000 51.8500 0.8900 ;
      RECT 50.7300 0.0000 50.9300 0.8900 ;
      RECT 49.3500 0.0000 50.0100 0.8900 ;
      RECT 48.4300 0.0000 48.6300 0.8900 ;
      RECT 47.5100 0.0000 47.7100 0.8900 ;
      RECT 46.1300 0.0000 46.7900 0.8900 ;
      RECT 45.2100 0.0000 45.4100 0.8900 ;
      RECT 44.2900 0.0000 44.4900 0.8900 ;
      RECT 43.3700 0.0000 43.5700 0.8900 ;
      RECT 41.9900 0.0000 42.6500 0.8900 ;
      RECT 41.0700 0.0000 41.2700 0.8900 ;
      RECT 40.1500 0.0000 40.3500 0.8900 ;
      RECT 39.2300 0.0000 39.4300 0.8900 ;
      RECT 37.8500 0.0000 38.5100 0.8900 ;
      RECT 36.9300 0.0000 37.1300 0.8900 ;
      RECT 36.0100 0.0000 36.2100 0.8900 ;
      RECT 34.6300 0.0000 35.2900 0.8900 ;
      RECT 33.7100 0.0000 33.9100 0.8900 ;
      RECT 32.7900 0.0000 32.9900 0.8900 ;
      RECT 31.8700 0.0000 32.0700 0.8900 ;
      RECT 30.4900 0.0000 31.1500 0.8900 ;
      RECT 29.5700 0.0000 29.7700 0.8900 ;
      RECT 28.6500 0.0000 28.8500 0.8900 ;
      RECT 27.2700 0.0000 27.9300 0.8900 ;
      RECT 26.3500 0.0000 26.5500 0.8900 ;
      RECT 25.4300 0.0000 25.6300 0.8900 ;
      RECT 24.5100 0.0000 24.7100 0.8900 ;
      RECT 23.1300 0.0000 23.7900 0.8900 ;
      RECT 22.2100 0.0000 22.4100 0.8900 ;
      RECT 21.2900 0.0000 21.4900 0.8900 ;
      RECT 19.9100 0.0000 20.5700 0.8900 ;
      RECT 18.9900 0.0000 19.1900 0.8900 ;
      RECT 18.0700 0.0000 18.2700 0.8900 ;
      RECT 17.1500 0.0000 17.3500 0.8900 ;
      RECT 15.7700 0.0000 16.4300 0.8900 ;
      RECT 14.8500 0.0000 15.0500 0.8900 ;
      RECT 13.9300 0.0000 14.1300 0.8900 ;
      RECT 12.5500 0.0000 13.2100 0.8900 ;
      RECT 11.6300 0.0000 11.8300 0.8900 ;
      RECT 10.7100 0.0000 10.9100 0.8900 ;
      RECT 9.7900 0.0000 9.9900 0.8900 ;
      RECT 8.4100 0.0000 9.0700 0.8900 ;
      RECT 7.4900 0.0000 7.6900 0.8900 ;
      RECT 6.5700 0.0000 6.7700 0.8900 ;
      RECT 5.6500 0.0000 5.8500 0.8900 ;
      RECT 0.0000 0.0000 4.9300 0.8900 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 100.2800 30.2600 ;
    LAYER met2 ;
      RECT 98.0800 29.4000 100.2800 30.2600 ;
      RECT 97.1600 29.4000 97.4200 30.2600 ;
      RECT 96.2400 29.4000 96.5000 30.2600 ;
      RECT 95.3200 29.4000 95.5800 30.2600 ;
      RECT 94.4000 29.4000 94.6600 30.2600 ;
      RECT 93.4800 29.4000 93.7400 30.2600 ;
      RECT 92.5600 29.4000 92.8200 30.2600 ;
      RECT 91.6400 29.4000 91.9000 30.2600 ;
      RECT 90.7200 29.4000 90.9800 30.2600 ;
      RECT 89.8000 29.4000 90.0600 30.2600 ;
      RECT 88.8800 29.4000 89.1400 30.2600 ;
      RECT 87.9600 29.4000 88.2200 30.2600 ;
      RECT 87.0400 29.4000 87.3000 30.2600 ;
      RECT 86.1200 29.4000 86.3800 30.2600 ;
      RECT 85.2000 29.4000 85.4600 30.2600 ;
      RECT 84.2800 29.4000 84.5400 30.2600 ;
      RECT 82.9000 29.4000 83.6200 30.2600 ;
      RECT 0.0000 29.4000 82.2400 30.2600 ;
      RECT 0.0000 28.9400 100.2800 29.4000 ;
      RECT 0.0000 28.5200 99.6550 28.9400 ;
      RECT 0.0000 27.9200 100.2800 28.5200 ;
      RECT 0.6250 27.5000 100.2800 27.9200 ;
      RECT 0.0000 26.9000 100.2800 27.5000 ;
      RECT 0.0000 26.4800 99.6550 26.9000 ;
      RECT 0.0000 26.2200 100.2800 26.4800 ;
      RECT 0.6250 25.8000 100.2800 26.2200 ;
      RECT 0.0000 25.2000 100.2800 25.8000 ;
      RECT 0.0000 24.7800 99.6550 25.2000 ;
      RECT 0.0000 24.5200 100.2800 24.7800 ;
      RECT 0.6250 24.1000 100.2800 24.5200 ;
      RECT 0.0000 23.1600 100.2800 24.1000 ;
      RECT 0.0000 22.8200 99.6550 23.1600 ;
      RECT 0.6250 22.7400 99.6550 22.8200 ;
      RECT 0.6250 22.4000 100.2800 22.7400 ;
      RECT 0.0000 21.4600 100.2800 22.4000 ;
      RECT 0.0000 21.1200 99.6550 21.4600 ;
      RECT 0.6250 21.0400 99.6550 21.1200 ;
      RECT 0.6250 20.7000 100.2800 21.0400 ;
      RECT 0.0000 19.4200 100.2800 20.7000 ;
      RECT 0.6250 19.0000 99.6550 19.4200 ;
      RECT 0.0000 17.7200 100.2800 19.0000 ;
      RECT 0.6250 17.3000 99.6550 17.7200 ;
      RECT 0.0000 16.0200 100.2800 17.3000 ;
      RECT 0.6250 15.6000 99.6550 16.0200 ;
      RECT 0.0000 14.3200 100.2800 15.6000 ;
      RECT 0.6250 13.9800 100.2800 14.3200 ;
      RECT 0.6250 13.9000 99.6550 13.9800 ;
      RECT 0.0000 13.5600 99.6550 13.9000 ;
      RECT 0.0000 12.6200 100.2800 13.5600 ;
      RECT 0.6250 12.2800 100.2800 12.6200 ;
      RECT 0.6250 12.2000 99.6550 12.2800 ;
      RECT 0.0000 11.8600 99.6550 12.2000 ;
      RECT 0.0000 10.9200 100.2800 11.8600 ;
      RECT 0.6250 10.5800 100.2800 10.9200 ;
      RECT 0.6250 10.5000 99.6550 10.5800 ;
      RECT 0.0000 10.1600 99.6550 10.5000 ;
      RECT 0.0000 9.2200 100.2800 10.1600 ;
      RECT 0.6250 8.8000 100.2800 9.2200 ;
      RECT 0.0000 8.5400 100.2800 8.8000 ;
      RECT 0.0000 8.1200 99.6550 8.5400 ;
      RECT 0.0000 7.5200 100.2800 8.1200 ;
      RECT 0.6250 7.1000 100.2800 7.5200 ;
      RECT 0.0000 6.8400 100.2800 7.1000 ;
      RECT 0.0000 6.4200 99.6550 6.8400 ;
      RECT 0.0000 5.8200 100.2800 6.4200 ;
      RECT 0.6250 5.4000 100.2800 5.8200 ;
      RECT 0.0000 4.8000 100.2800 5.4000 ;
      RECT 0.0000 4.3800 99.6550 4.8000 ;
      RECT 0.0000 4.1200 100.2800 4.3800 ;
      RECT 0.6250 3.7000 100.2800 4.1200 ;
      RECT 0.0000 3.1000 100.2800 3.7000 ;
      RECT 0.0000 2.6800 99.6550 3.1000 ;
      RECT 0.0000 2.4200 100.2800 2.6800 ;
      RECT 0.6250 2.0000 100.2800 2.4200 ;
      RECT 0.0000 1.4000 100.2800 2.0000 ;
      RECT 0.0000 0.9800 99.6550 1.4000 ;
      RECT 0.0000 0.8600 100.2800 0.9800 ;
      RECT 98.0800 0.0000 100.2800 0.8600 ;
      RECT 97.1600 0.0000 97.4200 0.8600 ;
      RECT 96.2400 0.0000 96.5000 0.8600 ;
      RECT 95.3200 0.0000 95.5800 0.8600 ;
      RECT 94.4000 0.0000 94.6600 0.8600 ;
      RECT 93.4800 0.0000 93.7400 0.8600 ;
      RECT 92.5600 0.0000 92.8200 0.8600 ;
      RECT 91.6400 0.0000 91.9000 0.8600 ;
      RECT 90.7200 0.0000 90.9800 0.8600 ;
      RECT 89.8000 0.0000 90.0600 0.8600 ;
      RECT 88.8800 0.0000 89.1400 0.8600 ;
      RECT 87.9600 0.0000 88.2200 0.8600 ;
      RECT 87.0400 0.0000 87.3000 0.8600 ;
      RECT 86.1200 0.0000 86.3800 0.8600 ;
      RECT 85.2000 0.0000 85.4600 0.8600 ;
      RECT 84.2800 0.0000 84.5400 0.8600 ;
      RECT 82.9000 0.0000 83.6200 0.8600 ;
      RECT 0.0000 0.0000 82.2400 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 100.2800 30.2600 ;
      RECT 98.0200 25.7000 100.2800 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 100.2800 25.7000 ;
      RECT 95.0200 22.7000 100.2800 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 100.2800 22.7000 ;
      RECT 95.0200 20.2000 100.2800 21.2800 ;
      RECT 7.8600 20.2000 92.4200 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 100.2800 20.2000 ;
      RECT 98.0200 17.4800 100.2800 18.5600 ;
      RECT 4.8600 17.4800 95.4200 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 100.2800 17.4800 ;
      RECT 95.0200 14.7600 100.2800 15.8400 ;
      RECT 7.8600 14.7600 92.4200 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 100.2800 14.7600 ;
      RECT 98.0200 12.0400 100.2800 13.1200 ;
      RECT 4.8600 12.0400 95.4200 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 100.2800 12.0400 ;
      RECT 95.0200 9.3200 100.2800 10.4000 ;
      RECT 7.8600 9.3200 92.4200 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 100.2800 9.3200 ;
      RECT 98.0200 6.6000 100.2800 7.6800 ;
      RECT 4.8600 6.6000 95.4200 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 100.2800 6.6000 ;
      RECT 95.0200 3.7700 100.2800 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 100.2800 3.7700 ;
      RECT 98.0200 0.7700 100.2800 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 100.2800 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 100.2800 30.2600 ;
      RECT 4.8600 25.3000 95.4200 28.3000 ;
      RECT 95.0200 3.7700 95.4200 25.3000 ;
      RECT 7.8600 3.7700 92.4200 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 98.0200 0.7700 100.2800 28.3000 ;
      RECT 4.8600 0.7700 95.4200 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 100.2800 0.7700 ;
  END
END N_term_RAM_IO

END LIBRARY
