##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Fri Jun 18 17:53:36 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DSP
  CLASS BLOCK ;
  SIZE 210.2200 BY 449.8200 ;
  FOREIGN DSP 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN top_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.902 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3955 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.5841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.7495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.36 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 449.1000 14.2200 449.8200 ;
    END
  END top_N1BEG[3]
  PIN top_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0372 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0715 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7656 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.592 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 449.1000 12.8400 449.8200 ;
    END
  END top_N1BEG[2]
  PIN top_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1075 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.3344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.436 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 449.1000 11.4600 449.8200 ;
    END
  END top_N1BEG[1]
  PIN top_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.00215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 35.4996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 177.38 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 449.1000 10.5400 449.8200 ;
    END
  END top_N1BEG[0]
  PIN top_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 75.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 403.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 449.1000 25.2600 449.8200 ;
    END
  END top_N2BEG[7]
  PIN top_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.0614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 503.072 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 449.1000 23.8800 449.8200 ;
    END
  END top_N2BEG[6]
  PIN top_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.1826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 455.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 449.1000 22.5000 449.8200 ;
    END
  END top_N2BEG[5]
  PIN top_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.334 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6501 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.2228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 486.992 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 449.1000 21.1200 449.8200 ;
    END
  END top_N2BEG[4]
  PIN top_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 32.9781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 164.602 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 449.1000 19.7400 449.8200 ;
    END
  END top_N2BEG[3]
  PIN top_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.372 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.786 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 449.1000 18.3600 449.8200 ;
    END
  END top_N2BEG[2]
  PIN top_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 34.1276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 170.52 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 449.1000 16.9800 449.8200 ;
    END
  END top_N2BEG[1]
  PIN top_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 33.8952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 169.358 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 449.1000 15.6000 449.8200 ;
    END
  END top_N2BEG[0]
  PIN top_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 29.534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 147.434 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 449.1000 35.8400 449.8200 ;
    END
  END top_N2BEGb[7]
  PIN top_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.8318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.24 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 449.1000 34.4600 449.8200 ;
    END
  END top_N2BEGb[6]
  PIN top_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 30.076 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 150.262 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 449.1000 33.5400 449.8200 ;
    END
  END top_N2BEGb[5]
  PIN top_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.4588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 333.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 449.1000 32.1600 449.8200 ;
    END
  END top_N2BEGb[4]
  PIN top_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.3508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.008 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 449.1000 30.7800 449.8200 ;
    END
  END top_N2BEGb[3]
  PIN top_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.1698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 449.1000 29.4000 449.8200 ;
    END
  END top_N2BEGb[2]
  PIN top_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.608 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.9625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 123.662 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 449.1000 28.0200 449.8200 ;
    END
  END top_N2BEGb[1]
  PIN top_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1912 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.8785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.1888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.826 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 449.1000 26.6400 449.8200 ;
    END
  END top_N2BEGb[0]
  PIN top_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.3019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.3385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.0448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 315.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 449.1000 57.4600 449.8200 ;
    END
  END top_N4BEG[15]
  PIN top_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 103.778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 553.952 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 449.1000 56.5400 449.8200 ;
    END
  END top_N4BEG[14]
  PIN top_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6742 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2935 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 105.965 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 565.616 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 449.1000 55.1600 449.8200 ;
    END
  END top_N4BEG[13]
  PIN top_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4909 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.0918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 480.96 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 449.1000 53.7800 449.8200 ;
    END
  END top_N4BEG[12]
  PIN top_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 449.1000 52.4000 449.8200 ;
    END
  END top_N4BEG[11]
  PIN top_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.74 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.582 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 449.1000 51.0200 449.8200 ;
    END
  END top_N4BEG[10]
  PIN top_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 449.1000 49.6400 449.8200 ;
    END
  END top_N4BEG[9]
  PIN top_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 449.1000 48.2600 449.8200 ;
    END
  END top_N4BEG[8]
  PIN top_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 116.38 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 621.632 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 449.1000 46.8800 449.8200 ;
    END
  END top_N4BEG[7]
  PIN top_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.952 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 449.1000 45.5000 449.8200 ;
    END
  END top_N4BEG[6]
  PIN top_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.8276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 426.688 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 449.1000 44.1200 449.8200 ;
    END
  END top_N4BEG[5]
  PIN top_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5553 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.5156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 473.024 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 449.1000 42.7400 449.8200 ;
    END
  END top_N4BEG[4]
  PIN top_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 449.1000 41.3600 449.8200 ;
    END
  END top_N4BEG[3]
  PIN top_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 449.1000 39.9800 449.8200 ;
    END
  END top_N4BEG[2]
  PIN top_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 449.1000 38.6000 449.8200 ;
    END
  END top_N4BEG[1]
  PIN top_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 120.152 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 641.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 449.1000 37.2200 449.8200 ;
    END
  END top_N4BEG[0]
  PIN top_NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4265 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 98.9238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 528.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 449.1000 79.5400 449.8200 ;
    END
  END top_NN4BEG[15]
  PIN top_NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 105.695 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 564.176 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 449.1000 78.1600 449.8200 ;
    END
  END top_NN4BEG[14]
  PIN top_NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.7102 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 416.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 449.1000 76.7800 449.8200 ;
    END
  END top_NN4BEG[13]
  PIN top_NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7994 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9195 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.4088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 311.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 449.1000 75.4000 449.8200 ;
    END
  END top_NN4BEG[12]
  PIN top_NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 449.1000 74.0200 449.8200 ;
    END
  END top_NN4BEG[11]
  PIN top_NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.692 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 449.1000 72.6400 449.8200 ;
    END
  END top_NN4BEG[10]
  PIN top_NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 449.1000 71.2600 449.8200 ;
    END
  END top_NN4BEG[9]
  PIN top_NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.798 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 449.1000 69.8800 449.8200 ;
    END
  END top_NN4BEG[8]
  PIN top_NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 95.7564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 512.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 449.1000 68.5000 449.8200 ;
    END
  END top_NN4BEG[7]
  PIN top_NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 120.242 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 641.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 449.1000 67.1200 449.8200 ;
    END
  END top_NN4BEG[6]
  PIN top_NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.25 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.132 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 449.1000 65.7400 449.8200 ;
    END
  END top_NN4BEG[5]
  PIN top_NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.25 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.132 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 449.1000 64.3600 449.8200 ;
    END
  END top_NN4BEG[4]
  PIN top_NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 449.1000 62.9800 449.8200 ;
    END
  END top_NN4BEG[3]
  PIN top_NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 449.1000 61.6000 449.8200 ;
    END
  END top_NN4BEG[2]
  PIN top_NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 449.1000 60.2200 449.8200 ;
    END
  END top_NN4BEG[1]
  PIN top_NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 449.1000 58.8400 449.8200 ;
    END
  END top_NN4BEG[0]
  PIN top_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.242 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.8298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 449.1000 84.6000 449.8200 ;
    END
  END top_S1END[3]
  PIN top_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.5781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.7195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.4273 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 366.352 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 449.1000 83.2200 449.8200 ;
    END
  END top_S1END[2]
  PIN top_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.7902 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 486.096 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 449.1000 81.8400 449.8200 ;
    END
  END top_S1END[1]
  PIN top_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.3544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 122.197 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 652.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 449.1000 80.4600 449.8200 ;
    END
  END top_S1END[0]
  PIN top_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1268 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.5565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8792 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 76.6647 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 411.216 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 449.1000 106.2200 449.8200 ;
    END
  END top_S2MID[7]
  PIN top_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.8474 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.264 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 449.1000 104.8400 449.8200 ;
    END
  END top_S2MID[6]
  PIN top_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6608 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.4195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.625 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.352 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 449.1000 103.4600 449.8200 ;
    END
  END top_S2MID[5]
  PIN top_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 73.7733 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 394.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 449.1000 102.5400 449.8200 ;
    END
  END top_S2MID[4]
  PIN top_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7596 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 22.8801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 113.565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7596 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8828 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 449.1000 101.1600 449.8200 ;
    END
  END top_S2MID[3]
  PIN top_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.7806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 342.976 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 449.1000 99.7800 449.8200 ;
    END
  END top_S2MID[2]
  PIN top_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7073 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.2475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1268 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.4594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 449.1000 98.4000 449.8200 ;
    END
  END top_S2MID[1]
  PIN top_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.5752 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.7985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 28.4987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 141.46 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.6992 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.9598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.256 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 449.1000 97.0200 449.8200 ;
    END
  END top_S2MID[0]
  PIN top_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.2994 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 96.2745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.271 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.76 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 449.1000 95.6400 449.8200 ;
    END
  END top_S2END[7]
  PIN top_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.4328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 312.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 449.1000 94.2600 449.8200 ;
    END
  END top_S2END[6]
  PIN top_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.102 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.1138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 459.744 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 449.1000 92.8800 449.8200 ;
    END
  END top_S2END[5]
  PIN top_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.2174 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.904 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 449.1000 91.5000 449.8200 ;
    END
  END top_S2END[4]
  PIN top_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 114.814 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 613.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 449.1000 90.1200 449.8200 ;
    END
  END top_S2END[3]
  PIN top_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.581 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 536.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 449.1000 88.7400 449.8200 ;
    END
  END top_S2END[2]
  PIN top_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84575 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.995 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.2434 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 449.1000 87.3600 449.8200 ;
    END
  END top_S2END[1]
  PIN top_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5852 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6977 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 108.136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 578.608 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 449.1000 85.9800 449.8200 ;
    END
  END top_S2END[0]
  PIN top_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.378 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 61.7015 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.9157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.1715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.5684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 15.9032 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 84.536 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 449.1000 127.8400 449.8200 ;
    END
  END top_S4END[15]
  PIN top_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.404 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.0738 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.9744 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 449.1000 126.4600 449.8200 ;
    END
  END top_S4END[14]
  PIN top_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.5612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.3192 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 32.3759 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.339 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 449.1000 125.5400 449.8200 ;
    END
  END top_S4END[13]
  PIN top_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.866 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.14788 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.3448 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 449.1000 124.1600 449.8200 ;
    END
  END top_S4END[12]
  PIN top_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.5812 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 39.692 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 200.603 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 449.1000 122.7800 449.8200 ;
    END
  END top_S4END[11]
  PIN top_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.5699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.3245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.197 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.8836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.4283 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 127.135 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 449.1000 121.4000 449.8200 ;
    END
  END top_S4END[10]
  PIN top_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.176 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.08067 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.0088 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 449.1000 120.0200 449.8200 ;
    END
  END top_S4END[9]
  PIN top_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90355 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.063 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.2628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 66.1255 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.4279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.6145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.3244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.84997 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.9158 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 449.1000 118.6400 449.8200 ;
    END
  END top_S4END[8]
  PIN top_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9504 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.35 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.954 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 449.1000 117.2600 449.8200 ;
    END
  END top_S4END[7]
  PIN top_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.4795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 106.46 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 449.1000 115.8800 449.8200 ;
    END
  END top_S4END[6]
  PIN top_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.5921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.6815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 449.1000 114.5000 449.8200 ;
    END
  END top_S4END[5]
  PIN top_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4799 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0196 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 449.1000 113.1200 449.8200 ;
    END
  END top_S4END[4]
  PIN top_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 95.8056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 511.904 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 449.1000 111.7400 449.8200 ;
    END
  END top_S4END[3]
  PIN top_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.2794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 461.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 449.1000 110.3600 449.8200 ;
    END
  END top_S4END[2]
  PIN top_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.9036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 469.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 449.1000 108.9800 449.8200 ;
    END
  END top_S4END[1]
  PIN top_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.6208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.448 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 449.1000 107.6000 449.8200 ;
    END
  END top_S4END[0]
  PIN top_SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.176 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7655 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.1304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 56.604 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 301.942 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 449.1000 149.4600 449.8200 ;
    END
  END top_SS4END[15]
  PIN top_SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.7221 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.2035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.2088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.7436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 88.9766 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 466.341 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 449.1000 148.5400 449.8200 ;
    END
  END top_SS4END[14]
  PIN top_SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.0298 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.0715 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 43.4389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 216.906 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.4418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.1631 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 373.483 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 449.1000 147.1600 449.8200 ;
    END
  END top_SS4END[13]
  PIN top_SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8768 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.136 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.94141 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.4034 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 449.1000 145.7800 449.8200 ;
    END
  END top_SS4END[12]
  PIN top_SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.662 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.3666 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.4384 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 449.1000 144.4000 449.8200 ;
    END
  END top_SS4END[11]
  PIN top_SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.0873 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.2655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 40.4131 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 204.512 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 449.1000 143.0200 449.8200 ;
    END
  END top_SS4END[10]
  PIN top_SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.3624 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.6975 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.53 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.7476 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 100.008 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 449.1000 141.6400 449.8200 ;
    END
  END top_SS4END[9]
  PIN top_SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.48 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 52.788 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 283.624 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 449.1000 140.2600 449.8200 ;
    END
  END top_SS4END[8]
  PIN top_SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.2126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 199.408 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 449.1000 138.8800 449.8200 ;
    END
  END top_SS4END[7]
  PIN top_SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.925 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.5475 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.7082 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.144 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.9247 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.064 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 449.1000 137.5000 449.8200 ;
    END
  END top_SS4END[6]
  PIN top_SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53935 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.811 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.0185 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.9215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.0968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 449.1000 136.1200 449.8200 ;
    END
  END top_SS4END[5]
  PIN top_SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.1292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 115.066 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 449.1000 134.7400 449.8200 ;
    END
  END top_SS4END[4]
  PIN top_SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 70.4643 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 377.216 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 449.1000 133.3600 449.8200 ;
    END
  END top_SS4END[3]
  PIN top_SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 73.1514 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 391.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 449.1000 131.9800 449.8200 ;
    END
  END top_SS4END[2]
  PIN top_SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.2586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 466.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 449.1000 130.6000 449.8200 ;
    END
  END top_SS4END[1]
  PIN top_SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.36595 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.607 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.887 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 547.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 449.1000 129.2200 449.8200 ;
    END
  END top_SS4END[0]
  PIN top_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.559 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.5418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 291.36 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 314.8200 210.2200 315.2000 ;
    END
  END top_E1BEG[3]
  PIN top_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.52 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.4176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 313.4600 210.2200 313.8400 ;
    END
  END top_E1BEG[2]
  PIN top_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 311.7600 210.2200 312.1400 ;
    END
  END top_E1BEG[1]
  PIN top_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 310.4000 210.2200 310.7800 ;
    END
  END top_E1BEG[0]
  PIN top_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.951 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.7208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 249.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 326.7200 210.2200 327.1000 ;
    END
  END top_E2BEG[7]
  PIN top_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4538 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.161 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 325.0200 210.2200 325.4000 ;
    END
  END top_E2BEG[6]
  PIN top_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 323.6600 210.2200 324.0400 ;
    END
  END top_E2BEG[5]
  PIN top_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.81 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 322.3000 210.2200 322.6800 ;
    END
  END top_E2BEG[4]
  PIN top_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.8108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 320.6000 210.2200 320.9800 ;
    END
  END top_E2BEG[3]
  PIN top_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.177 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 319.2400 210.2200 319.6200 ;
    END
  END top_E2BEG[2]
  PIN top_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.616 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 317.8800 210.2200 318.2600 ;
    END
  END top_E2BEG[1]
  PIN top_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.3645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 316.1800 210.2200 316.5600 ;
    END
  END top_E2BEG[0]
  PIN top_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.877 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 338.2800 210.2200 338.6600 ;
    END
  END top_E2BEGb[7]
  PIN top_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 336.9200 210.2200 337.3000 ;
    END
  END top_E2BEGb[6]
  PIN top_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.216 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 335.5600 210.2200 335.9400 ;
    END
  END top_E2BEGb[5]
  PIN top_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 333.8600 210.2200 334.2400 ;
    END
  END top_E2BEGb[4]
  PIN top_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 332.5000 210.2200 332.8800 ;
    END
  END top_E2BEGb[3]
  PIN top_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 331.1400 210.2200 331.5200 ;
    END
  END top_E2BEGb[2]
  PIN top_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 329.4400 210.2200 329.8200 ;
    END
  END top_E2BEGb[1]
  PIN top_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 328.0800 210.2200 328.4600 ;
    END
  END top_E2BEGb[0]
  PIN top_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.2782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 494.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 362.0800 210.2200 362.4600 ;
    END
  END top_EE4BEG[15]
  PIN top_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.9675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.5354 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 360.3800 210.2200 360.7600 ;
    END
  END top_EE4BEG[14]
  PIN top_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.69 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.1598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 422.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 359.0200 210.2200 359.4000 ;
    END
  END top_EE4BEG[13]
  PIN top_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.3789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 156.734 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.6838 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 357.6600 210.2200 358.0400 ;
    END
  END top_EE4BEG[12]
  PIN top_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 355.9600 210.2200 356.3400 ;
    END
  END top_EE4BEG[11]
  PIN top_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 354.6000 210.2200 354.9800 ;
    END
  END top_EE4BEG[10]
  PIN top_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.92 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 353.2400 210.2200 353.6200 ;
    END
  END top_EE4BEG[9]
  PIN top_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.044 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 351.5400 210.2200 351.9200 ;
    END
  END top_EE4BEG[8]
  PIN top_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 350.1800 210.2200 350.5600 ;
    END
  END top_EE4BEG[7]
  PIN top_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.9418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.16 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 348.8200 210.2200 349.2000 ;
    END
  END top_EE4BEG[6]
  PIN top_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.544 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 347.1200 210.2200 347.5000 ;
    END
  END top_EE4BEG[5]
  PIN top_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.627 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 345.7600 210.2200 346.1400 ;
    END
  END top_EE4BEG[4]
  PIN top_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 344.4000 210.2200 344.7800 ;
    END
  END top_EE4BEG[3]
  PIN top_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.025 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 342.7000 210.2200 343.0800 ;
    END
  END top_EE4BEG[2]
  PIN top_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.9536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.36 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 341.3400 210.2200 341.7200 ;
    END
  END top_EE4BEG[1]
  PIN top_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5018 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.401 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 339.9800 210.2200 340.3600 ;
    END
  END top_EE4BEG[0]
  PIN top_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2873 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 104.595 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 560.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 379.7600 210.2200 380.1400 ;
    END
  END top_E6BEG[11]
  PIN top_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 87.7368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 468.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 378.0600 210.2200 378.4400 ;
    END
  END top_E6BEG[10]
  PIN top_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.056 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 376.7000 210.2200 377.0800 ;
    END
  END top_E6BEG[9]
  PIN top_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.0758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 230.208 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 375.3400 210.2200 375.7200 ;
    END
  END top_E6BEG[8]
  PIN top_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.993 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 251.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 373.6400 210.2200 374.0200 ;
    END
  END top_E6BEG[7]
  PIN top_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.9688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.304 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 372.2800 210.2200 372.6600 ;
    END
  END top_E6BEG[6]
  PIN top_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.219 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 370.9200 210.2200 371.3000 ;
    END
  END top_E6BEG[5]
  PIN top_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.323 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 369.2200 210.2200 369.6000 ;
    END
  END top_E6BEG[4]
  PIN top_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.8358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.928 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 367.8600 210.2200 368.2400 ;
    END
  END top_E6BEG[3]
  PIN top_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 240.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 366.5000 210.2200 366.8800 ;
    END
  END top_E6BEG[2]
  PIN top_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.114 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 54.0678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 288.832 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 364.8000 210.2200 365.1800 ;
    END
  END top_E6BEG[1]
  PIN top_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 363.4400 210.2200 363.8200 ;
    END
  END top_E6BEG[0]
  PIN top_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.5155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.0691 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 314.8200 0.7200 315.2000 ;
    END
  END top_E1END[3]
  PIN top_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.9837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 174.64 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.1878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.3014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.352 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 313.4600 0.7200 313.8400 ;
    END
  END top_E1END[2]
  PIN top_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.3201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.3215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.3056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.904 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 311.7600 0.7200 312.1400 ;
    END
  END top_E1END[1]
  PIN top_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.2891 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 328.752 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 310.4000 0.7200 310.7800 ;
    END
  END top_E1END[0]
  PIN top_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.093 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 182.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.4647 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 97.8858 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 520.549 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 326.7200 0.7200 327.1000 ;
    END
  END top_E2MID[7]
  PIN top_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.2624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 284.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 73.2828 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 389.572 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.7236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 324.8 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 155.065 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 827.013 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 325.0200 0.7200 325.4000 ;
    END
  END top_E2MID[6]
  PIN top_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4333 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.723 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.7287 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 81.2617 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.671 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 323.6600 0.7200 324.0400 ;
    END
  END top_E2MID[5]
  PIN top_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.9514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 293.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 77.4945 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 410.007 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.9648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.616 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 135.36 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 719.254 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 322.3000 0.7200 322.6800 ;
    END
  END top_E2MID[4]
  PIN top_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.3994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 290.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 76.4416 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 405.786 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.1198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.776 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 131.822 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 701.78 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 320.6000 0.7200 320.9800 ;
    END
  END top_E2MID[3]
  PIN top_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 51.6814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 276.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 73.8918 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 390.525 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.7046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.032 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 128.713 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 684.171 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 319.2400 0.7200 319.6200 ;
    END
  END top_E2MID[2]
  PIN top_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 41.0704 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.648 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 317.8800 0.7200 318.2600 ;
    END
  END top_E2MID[1]
  PIN top_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.8217 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 276.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 70.7881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 376.457 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 316.1800 0.7200 316.5600 ;
    END
  END top_E2MID[0]
  PIN top_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.01 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.2743 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 413.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 338.2800 0.7200 338.6600 ;
    END
  END top_E2END[7]
  PIN top_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.5348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1448 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.7003 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.808 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 336.9200 0.7200 337.3000 ;
    END
  END top_E2END[6]
  PIN top_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.2855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.02 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1448 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.6664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 335.5600 0.7200 335.9400 ;
    END
  END top_E2END[5]
  PIN top_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 74.6817 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 398.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 333.8600 0.7200 334.2400 ;
    END
  END top_E2END[4]
  PIN top_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.7544 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 458.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 332.5000 0.7200 332.8800 ;
    END
  END top_E2END[3]
  PIN top_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 32.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 159.754 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0309 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.332 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 331.1400 0.7200 331.5200 ;
    END
  END top_E2END[2]
  PIN top_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.0579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.928 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1864 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.072 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 329.4400 0.7200 329.8200 ;
    END
  END top_E2END[1]
  PIN top_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.189 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.4068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.64 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 328.0800 0.7200 328.4600 ;
    END
  END top_E2END[0]
  PIN top_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.7388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 18.365 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 100.689 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 362.0800 0.7200 362.4600 ;
    END
  END top_EE4END[15]
  PIN top_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 286.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 5.18842 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 27.6067 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 360.3800 0.7200 360.7600 ;
    END
  END top_EE4END[14]
  PIN top_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.887 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 7.4932 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 38.3609 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 359.0200 0.7200 359.4000 ;
    END
  END top_EE4END[13]
  PIN top_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 303.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.57926 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 19.1589 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 357.6600 0.7200 358.0400 ;
    END
  END top_EE4END[12]
  PIN top_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.389 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.98869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.5623 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 355.9600 0.7200 356.3400 ;
    END
  END top_EE4END[11]
  PIN top_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 15.4549 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 81.7737 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 354.6000 0.7200 354.9800 ;
    END
  END top_EE4END[10]
  PIN top_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.1728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 30.3481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 161.951 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 353.2400 0.7200 353.6200 ;
    END
  END top_EE4END[9]
  PIN top_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 41.422 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 221.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 17.971 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 96.1313 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 351.5400 0.7200 351.9200 ;
    END
  END top_EE4END[8]
  PIN top_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6374 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 37.3079 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.44 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 350.1800 0.7200 350.5600 ;
    END
  END top_EE4END[7]
  PIN top_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.442 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4882 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 8.66222 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 47.2956 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 348.8200 0.7200 349.2000 ;
    END
  END top_EE4END[6]
  PIN top_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.685 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 7.52114 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 37.7805 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 347.1200 0.7200 347.5000 ;
    END
  END top_EE4END[5]
  PIN top_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2611 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.5192 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.092 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 345.7600 0.7200 346.1400 ;
    END
  END top_EE4END[4]
  PIN top_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.3871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 101.539 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 344.4000 0.7200 344.7800 ;
    END
  END top_EE4END[3]
  PIN top_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.923 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.5684 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 342.7000 0.7200 343.0800 ;
    END
  END top_EE4END[2]
  PIN top_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.674 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.4428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.832 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 341.3400 0.7200 341.7200 ;
    END
  END top_EE4END[1]
  PIN top_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7545 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.942 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.3347 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 487.584 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 339.9800 0.7200 340.3600 ;
    END
  END top_EE4END[0]
  PIN top_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.521 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 253.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 6.29616 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 33.5367 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 379.7600 0.7200 380.1400 ;
    END
  END top_E6END[11]
  PIN top_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.5348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.4341 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 53.3737 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 378.0600 0.7200 378.4400 ;
    END
  END top_E6END[10]
  PIN top_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6922 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.353 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.54128 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.3253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 376.7000 0.7200 377.0800 ;
    END
  END top_E6END[9]
  PIN top_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.729 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 2.92155 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 13.9205 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 375.3400 0.7200 375.7200 ;
    END
  END top_E6END[8]
  PIN top_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.442 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 35.3805 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.018 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 373.6400 0.7200 374.0200 ;
    END
  END top_E6END[7]
  PIN top_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.9758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 32.9089 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 173.331 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 372.2800 0.7200 372.6600 ;
    END
  END top_E6END[6]
  PIN top_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.6118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 56.312 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 296.368 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 370.9200 0.7200 371.3000 ;
    END
  END top_E6END[5]
  PIN top_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 8.87636 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 45.6593 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 369.2200 0.7200 369.6000 ;
    END
  END top_E6END[4]
  PIN top_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.39044 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.571 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 367.8600 0.7200 368.2400 ;
    END
  END top_E6END[3]
  PIN top_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 214.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.8877 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.69 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 366.5000 0.7200 366.8800 ;
    END
  END top_E6END[2]
  PIN top_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.2716 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.1108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 364.8000 0.7200 365.1800 ;
    END
  END top_E6END[1]
  PIN top_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.2752 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.9526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 363.4400 0.7200 363.8200 ;
    END
  END top_E6END[0]
  PIN top_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.104 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 244.1000 0.7200 244.4800 ;
    END
  END top_W1BEG[3]
  PIN top_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 242.7400 0.7200 243.1200 ;
    END
  END top_W1BEG[2]
  PIN top_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 241.3800 0.7200 241.7600 ;
    END
  END top_W1BEG[1]
  PIN top_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.6858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.128 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 240.0200 0.7200 240.4000 ;
    END
  END top_W1BEG[0]
  PIN top_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 256.0000 0.7200 256.3800 ;
    END
  END top_W2BEG[7]
  PIN top_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.9888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.744 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 254.6400 0.7200 255.0200 ;
    END
  END top_W2BEG[6]
  PIN top_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.7388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.744 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 252.9400 0.7200 253.3200 ;
    END
  END top_W2BEG[5]
  PIN top_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.687 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 251.5800 0.7200 251.9600 ;
    END
  END top_W2BEG[4]
  PIN top_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.044 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 250.2200 0.7200 250.6000 ;
    END
  END top_W2BEG[3]
  PIN top_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 248.5200 0.7200 248.9000 ;
    END
  END top_W2BEG[2]
  PIN top_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.184 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 247.1600 0.7200 247.5400 ;
    END
  END top_W2BEG[1]
  PIN top_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 245.8000 0.7200 246.1800 ;
    END
  END top_W2BEG[0]
  PIN top_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.3913 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 267.9000 0.7200 268.2800 ;
    END
  END top_W2BEGb[7]
  PIN top_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 266.2000 0.7200 266.5800 ;
    END
  END top_W2BEGb[6]
  PIN top_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.2908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.688 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 264.8400 0.7200 265.2200 ;
    END
  END top_W2BEGb[5]
  PIN top_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.8968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.92 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 263.4800 0.7200 263.8600 ;
    END
  END top_W2BEGb[4]
  PIN top_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.8658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 197.088 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 261.7800 0.7200 262.1600 ;
    END
  END top_W2BEGb[3]
  PIN top_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.8608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.728 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 260.4200 0.7200 260.8000 ;
    END
  END top_W2BEGb[2]
  PIN top_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 259.0600 0.7200 259.4400 ;
    END
  END top_W2BEGb[1]
  PIN top_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 257.3600 0.7200 257.7400 ;
    END
  END top_W2BEGb[0]
  PIN top_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.2695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.5098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 205.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 291.3600 0.7200 291.7400 ;
    END
  END top_WW4BEG[15]
  PIN top_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.9728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 330.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 290.0000 0.7200 290.3800 ;
    END
  END top_WW4BEG[14]
  PIN top_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.647 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.4198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 288.3000 0.7200 288.6800 ;
    END
  END top_WW4BEG[13]
  PIN top_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.69 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.6866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 313.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 286.9400 0.7200 287.3200 ;
    END
  END top_WW4BEG[12]
  PIN top_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 285.5800 0.7200 285.9600 ;
    END
  END top_WW4BEG[11]
  PIN top_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.965 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 283.8800 0.7200 284.2600 ;
    END
  END top_WW4BEG[10]
  PIN top_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 281.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 282.5200 0.7200 282.9000 ;
    END
  END top_WW4BEG[9]
  PIN top_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.3078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 281.1600 0.7200 281.5400 ;
    END
  END top_WW4BEG[8]
  PIN top_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 279.4600 0.7200 279.8400 ;
    END
  END top_WW4BEG[7]
  PIN top_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 278.1000 0.7200 278.4800 ;
    END
  END top_WW4BEG[6]
  PIN top_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 276.7400 0.7200 277.1200 ;
    END
  END top_WW4BEG[5]
  PIN top_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.0348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.656 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 275.0400 0.7200 275.4200 ;
    END
  END top_WW4BEG[4]
  PIN top_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.0068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 197.84 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 273.6800 0.7200 274.0600 ;
    END
  END top_WW4BEG[3]
  PIN top_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 272.3200 0.7200 272.7000 ;
    END
  END top_WW4BEG[2]
  PIN top_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 270.6200 0.7200 271.0000 ;
    END
  END top_WW4BEG[1]
  PIN top_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.997 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 269.2600 0.7200 269.6400 ;
    END
  END top_WW4BEG[0]
  PIN top_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.621 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 309.0400 0.7200 309.4200 ;
    END
  END top_W6BEG[11]
  PIN top_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.1615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.8292 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 307.6800 0.7200 308.0600 ;
    END
  END top_W6BEG[10]
  PIN top_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 305.9800 0.7200 306.3600 ;
    END
  END top_W6BEG[9]
  PIN top_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 46.7568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 249.84 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 304.6200 0.7200 305.0000 ;
    END
  END top_W6BEG[8]
  PIN top_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.1518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.28 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 303.2600 0.7200 303.6400 ;
    END
  END top_W6BEG[7]
  PIN top_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 301.5600 0.7200 301.9400 ;
    END
  END top_W6BEG[6]
  PIN top_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.8348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.256 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 300.2000 0.7200 300.5800 ;
    END
  END top_W6BEG[5]
  PIN top_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 48.1758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 257.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 298.8400 0.7200 299.2200 ;
    END
  END top_W6BEG[4]
  PIN top_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.305 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 297.1400 0.7200 297.5200 ;
    END
  END top_W6BEG[3]
  PIN top_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 295.7800 0.7200 296.1600 ;
    END
  END top_W6BEG[2]
  PIN top_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 210.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 294.4200 0.7200 294.8000 ;
    END
  END top_W6BEG[1]
  PIN top_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 46.3908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 247.888 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 292.7200 0.7200 293.1000 ;
    END
  END top_W6BEG[0]
  PIN top_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.0154 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 244.1000 210.2200 244.4800 ;
    END
  END top_W1END[3]
  PIN top_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.192 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 242.7400 210.2200 243.1200 ;
    END
  END top_W1END[2]
  PIN top_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.082 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.8321 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 241.3800 210.2200 241.7600 ;
    END
  END top_W1END[1]
  PIN top_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.7456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.9438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 240.0200 210.2200 240.4000 ;
    END
  END top_W1END[0]
  PIN top_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.4044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 60.029 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 318.787 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.5818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.24 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 99.8698 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 531.904 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 256.0000 210.2200 256.3800 ;
    END
  END top_W2MID[7]
  PIN top_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.3712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 98.2967 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 525.632 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 254.6400 210.2200 255.0200 ;
    END
  END top_W2MID[6]
  PIN top_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.7076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 53.6648 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 280.094 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 252.9400 210.2200 253.3200 ;
    END
  END top_W2MID[5]
  PIN top_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.739 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 38.9933 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.667 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.284714 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 251.5800 210.2200 251.9600 ;
    END
  END top_W2MID[4]
  PIN top_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.2245 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 41.1749 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 217.442 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 250.2200 210.2200 250.6000 ;
    END
  END top_W2MID[3]
  PIN top_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.2977 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.2904 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 288.326 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 248.5200 210.2200 248.9000 ;
    END
  END top_W2MID[2]
  PIN top_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.163 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.1144 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 57.8368 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 308.102 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 247.1600 210.2200 247.5400 ;
    END
  END top_W2MID[1]
  PIN top_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 58.4806 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 312.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 85.9185 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 455.63 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 88.5432 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 470.261 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 245.8000 210.2200 246.1800 ;
    END
  END top_W2MID[0]
  PIN top_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.357 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.6575 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 48.9573 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 263.693 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 267.9000 210.2200 268.2800 ;
    END
  END top_W2END[7]
  PIN top_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.421 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.7736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 330.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 266.2000 210.2200 266.5800 ;
    END
  END top_W2END[6]
  PIN top_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.407 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.9798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 264.8400 210.2200 265.2200 ;
    END
  END top_W2END[5]
  PIN top_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.8415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 58.9807 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 315.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.3176 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 67.5358 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361.903 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 263.4800 210.2200 263.8600 ;
    END
  END top_W2END[4]
  PIN top_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 278.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.3568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 366.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 100.685 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 538.597 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 261.7800 210.2200 262.1600 ;
    END
  END top_W2END[3]
  PIN top_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.5436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 260.4200 210.2200 260.8000 ;
    END
  END top_W2END[2]
  PIN top_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.5325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.4022 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.36 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 259.0600 210.2200 259.4400 ;
    END
  END top_W2END[1]
  PIN top_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.571 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.4253 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.261 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 257.3600 210.2200 257.7400 ;
    END
  END top_W2END[0]
  PIN top_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.373 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.785 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.296 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 291.3600 210.2200 291.7400 ;
    END
  END top_WW4END[15]
  PIN top_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.6718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 190.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 50.1593 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 265.942 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 290.0000 210.2200 290.3800 ;
    END
  END top_WW4END[14]
  PIN top_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.829 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.50976 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.1677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 288.3000 210.2200 288.6800 ;
    END
  END top_WW4END[13]
  PIN top_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.29481 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.0929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 286.9400 210.2200 287.3200 ;
    END
  END top_WW4END[12]
  PIN top_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.4638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 242.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 64.2638 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 340.897 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 285.5800 210.2200 285.9600 ;
    END
  END top_WW4END[11]
  PIN top_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 57.73 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 308.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.6369 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 19.5205 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 283.8800 210.2200 284.2600 ;
    END
  END top_WW4END[10]
  PIN top_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.2468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 204.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 20.0249 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 105.902 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 282.5200 210.2200 282.9000 ;
    END
  END top_WW4END[9]
  PIN top_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.4758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 44.421 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 234.941 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 281.1600 210.2200 281.5400 ;
    END
  END top_WW4END[8]
  PIN top_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.3068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.4463 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.78 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 279.4600 210.2200 279.8400 ;
    END
  END top_WW4END[7]
  PIN top_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 56.0527 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.555 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 278.1000 210.2200 278.4800 ;
    END
  END top_WW4END[6]
  PIN top_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.6168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.9603 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 125.98 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 276.7400 210.2200 277.1200 ;
    END
  END top_WW4END[5]
  PIN top_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.5388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.3762 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 96.6774 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 275.0400 210.2200 275.4200 ;
    END
  END top_WW4END[4]
  PIN top_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.9608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 273.6800 210.2200 274.0600 ;
    END
  END top_WW4END[3]
  PIN top_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.187 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.6068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 272.3200 210.2200 272.7000 ;
    END
  END top_WW4END[2]
  PIN top_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.675 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.0418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 349.712 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 270.6200 210.2200 271.0000 ;
    END
  END top_WW4END[1]
  PIN top_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.3513 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 269.2600 210.2200 269.6400 ;
    END
  END top_WW4END[0]
  PIN top_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.861 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.73643 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 20.1273 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 309.0400 210.2200 309.4200 ;
    END
  END top_W6END[11]
  PIN top_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.6768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.8222 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.9697 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 307.6800 210.2200 308.0600 ;
    END
  END top_W6END[10]
  PIN top_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.8648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 32.2232 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 169.201 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 305.9800 210.2200 306.3600 ;
    END
  END top_W6END[9]
  PIN top_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 57.3872 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.271 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 304.6200 210.2200 305.0000 ;
    END
  END top_W6END[8]
  PIN top_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.1048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 43.7248 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 229.352 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 303.2600 210.2200 303.6400 ;
    END
  END top_W6END[7]
  PIN top_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.5578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.6535 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 113.97 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 301.5600 210.2200 301.9400 ;
    END
  END top_W6END[6]
  PIN top_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.6868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 25.4261 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 134.329 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 300.2000 210.2200 300.5800 ;
    END
  END top_W6END[5]
  PIN top_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 61.591 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 328.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 2.67906 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 13.9091 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 298.8400 210.2200 299.2200 ;
    END
  END top_W6END[4]
  PIN top_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.17104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.4741 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 297.1400 210.2200 297.5200 ;
    END
  END top_W6END[3]
  PIN top_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.498 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.55582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.3845 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 295.7800 210.2200 296.1600 ;
    END
  END top_W6END[2]
  PIN top_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.2253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.7295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.3168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.9044 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3266 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 294.4200 210.2200 294.8000 ;
    END
  END top_W6END[1]
  PIN top_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7136 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.7447 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 321.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 292.7200 210.2200 293.1000 ;
    END
  END top_W6END[0]
  PIN bot_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 84.6400 210.2200 85.0200 ;
    END
  END bot_E1BEG[3]
  PIN bot_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.8924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 331.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 83.2800 210.2200 83.6600 ;
    END
  END bot_E1BEG[2]
  PIN bot_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.1798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 348.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 81.5800 210.2200 81.9600 ;
    END
  END bot_E1BEG[1]
  PIN bot_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.3285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.7316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 80.2200 210.2200 80.6000 ;
    END
  END bot_E1BEG[0]
  PIN bot_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.808 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 96.5400 210.2200 96.9200 ;
    END
  END bot_E2BEG[7]
  PIN bot_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 94.8400 210.2200 95.2200 ;
    END
  END bot_E2BEG[6]
  PIN bot_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.8265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.3338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.584 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 93.4800 210.2200 93.8600 ;
    END
  END bot_E2BEG[5]
  PIN bot_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.2388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 321.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 92.1200 210.2200 92.5000 ;
    END
  END bot_E2BEG[4]
  PIN bot_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.3026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.888 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 90.4200 210.2200 90.8000 ;
    END
  END bot_E2BEG[3]
  PIN bot_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.2075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.432 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 89.0600 210.2200 89.4400 ;
    END
  END bot_E2BEG[2]
  PIN bot_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.7224 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 357.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 87.7000 210.2200 88.0800 ;
    END
  END bot_E2BEG[1]
  PIN bot_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 86.0000 210.2200 86.3800 ;
    END
  END bot_E2BEG[0]
  PIN bot_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 108.1000 210.2200 108.4800 ;
    END
  END bot_E2BEGb[7]
  PIN bot_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 106.7400 210.2200 107.1200 ;
    END
  END bot_E2BEGb[6]
  PIN bot_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 105.3800 210.2200 105.7600 ;
    END
  END bot_E2BEGb[5]
  PIN bot_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.389 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 103.6800 210.2200 104.0600 ;
    END
  END bot_E2BEGb[4]
  PIN bot_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6333 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 102.3200 210.2200 102.7000 ;
    END
  END bot_E2BEGb[3]
  PIN bot_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.7108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.928 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 100.9600 210.2200 101.3400 ;
    END
  END bot_E2BEGb[2]
  PIN bot_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0602 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 99.2600 210.2200 99.6400 ;
    END
  END bot_E2BEGb[1]
  PIN bot_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.1358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.528 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 97.9000 210.2200 98.2800 ;
    END
  END bot_E2BEGb[0]
  PIN bot_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.5658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.488 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 131.9000 210.2200 132.2800 ;
    END
  END bot_EE4BEG[15]
  PIN bot_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.472 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.1394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 199.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 130.2000 210.2200 130.5800 ;
    END
  END bot_EE4BEG[14]
  PIN bot_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.067 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.0956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 422.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 128.8400 210.2200 129.2200 ;
    END
  END bot_EE4BEG[13]
  PIN bot_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.7155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.6074 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 127.4800 210.2200 127.8600 ;
    END
  END bot_EE4BEG[12]
  PIN bot_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.254 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 125.7800 210.2200 126.1600 ;
    END
  END bot_EE4BEG[11]
  PIN bot_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.4 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 124.4200 210.2200 124.8000 ;
    END
  END bot_EE4BEG[10]
  PIN bot_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.122 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 123.0600 210.2200 123.4400 ;
    END
  END bot_EE4BEG[9]
  PIN bot_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.7668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.56 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 121.3600 210.2200 121.7400 ;
    END
  END bot_EE4BEG[8]
  PIN bot_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.657 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 233.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 120.0000 210.2200 120.3800 ;
    END
  END bot_EE4BEG[7]
  PIN bot_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 190.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 118.6400 210.2200 119.0200 ;
    END
  END bot_EE4BEG[6]
  PIN bot_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.097 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 116.9400 210.2200 117.3200 ;
    END
  END bot_EE4BEG[5]
  PIN bot_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.171 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 115.5800 210.2200 115.9600 ;
    END
  END bot_EE4BEG[4]
  PIN bot_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.448 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 114.2200 210.2200 114.6000 ;
    END
  END bot_EE4BEG[3]
  PIN bot_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 112.5200 210.2200 112.9000 ;
    END
  END bot_EE4BEG[2]
  PIN bot_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.012 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 111.1600 210.2200 111.5400 ;
    END
  END bot_EE4BEG[1]
  PIN bot_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.2118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 209.6 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 109.8000 210.2200 110.1800 ;
    END
  END bot_EE4BEG[0]
  PIN bot_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.2136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 338.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 149.5800 210.2200 149.9600 ;
    END
  END bot_E6BEG[11]
  PIN bot_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.1314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 418.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 147.8800 210.2200 148.2600 ;
    END
  END bot_E6BEG[10]
  PIN bot_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 146.5200 210.2200 146.9000 ;
    END
  END bot_E6BEG[9]
  PIN bot_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 225.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 145.1600 210.2200 145.5400 ;
    END
  END bot_E6BEG[8]
  PIN bot_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 143.4600 210.2200 143.8400 ;
    END
  END bot_E6BEG[7]
  PIN bot_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 142.1000 210.2200 142.4800 ;
    END
  END bot_E6BEG[6]
  PIN bot_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 59.8608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 319.728 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 140.7400 210.2200 141.1200 ;
    END
  END bot_E6BEG[5]
  PIN bot_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 139.0400 210.2200 139.4200 ;
    END
  END bot_E6BEG[4]
  PIN bot_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 59.1258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 315.808 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 137.6800 210.2200 138.0600 ;
    END
  END bot_E6BEG[3]
  PIN bot_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.2028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.552 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 136.3200 210.2200 136.7000 ;
    END
  END bot_E6BEG[2]
  PIN bot_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.0808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 134.6200 210.2200 135.0000 ;
    END
  END bot_E6BEG[1]
  PIN bot_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.64 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 133.2600 210.2200 133.6400 ;
    END
  END bot_E6BEG[0]
  PIN bot_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.0495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.5908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.584 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.6400 0.7200 85.0200 ;
    END
  END bot_E1END[3]
  PIN bot_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.7306 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.2800 0.7200 83.6600 ;
    END
  END bot_E1END[2]
  PIN bot_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.4045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 131.743 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.413 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.5800 0.7200 81.9600 ;
    END
  END bot_E1END[1]
  PIN bot_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.577 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 67.0425 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 358.496 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.2200 0.7200 80.6000 ;
    END
  END bot_E1END[0]
  PIN bot_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7354 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 27.0484 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 143.948 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.5400 0.7200 96.9200 ;
    END
  END bot_E2MID[7]
  PIN bot_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.589 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.242 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 95.4503 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 509.042 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.8400 0.7200 95.2200 ;
    END
  END bot_E2MID[6]
  PIN bot_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 66.6774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 357.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 95.5922 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 507.984 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.4800 0.7200 93.8600 ;
    END
  END bot_E2MID[5]
  PIN bot_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 67.0023 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.749 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.1200 0.7200 92.5000 ;
    END
  END bot_E2MID[4]
  PIN bot_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7632 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.598 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.977 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.9933 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.35 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.4200 0.7200 90.8000 ;
    END
  END bot_E2MID[3]
  PIN bot_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8251 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.2712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.7852 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 405.013 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.0600 0.7200 89.4400 ;
    END
  END bot_E2MID[2]
  PIN bot_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.0988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.2486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 217.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 58.9564 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.69 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.7000 0.7200 88.0800 ;
    END
  END bot_E2MID[1]
  PIN bot_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.049 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7596 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.8366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.9071 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 434.338 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.0000 0.7200 86.3800 ;
    END
  END bot_E2MID[0]
  PIN bot_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.3711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 176.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.3607 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.408 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.1000 0.7200 108.4800 ;
    END
  END bot_E2END[7]
  PIN bot_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1448 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.1426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.368 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.7400 0.7200 107.1200 ;
    END
  END bot_E2END[6]
  PIN bot_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 162.578 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1448 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.0134 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.3800 0.7200 105.7600 ;
    END
  END bot_E2END[5]
  PIN bot_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.2525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.2038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 332.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.6800 0.7200 104.0600 ;
    END
  END bot_E2END[4]
  PIN bot_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.8746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.272 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.3200 0.7200 102.7000 ;
    END
  END bot_E2END[3]
  PIN bot_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.332 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.9216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 357.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 100.9600 0.7200 101.3400 ;
    END
  END bot_E2END[2]
  PIN bot_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.1702 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 333.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.2600 0.7200 99.6400 ;
    END
  END bot_E2END[1]
  PIN bot_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7632 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 31.0456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.196 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.9000 0.7200 98.2800 ;
    END
  END bot_E2END[0]
  PIN bot_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.5108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.2582 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.9306 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 131.9000 0.7200 132.2800 ;
    END
  END bot_EE4END[15]
  PIN bot_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.5668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 59.2071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.821 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.2000 0.7200 130.5800 ;
    END
  END bot_EE4END[14]
  PIN bot_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 13.143 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 70.0155 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.8400 0.7200 129.2200 ;
    END
  END bot_EE4END[13]
  PIN bot_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.0578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 262.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 67.8794 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 360.026 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.4800 0.7200 127.8600 ;
    END
  END bot_EE4END[12]
  PIN bot_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.13165 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.9859 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.7800 0.7200 126.1600 ;
    END
  END bot_EE4END[11]
  PIN bot_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.933 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.65758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.7542 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.4200 0.7200 124.8000 ;
    END
  END bot_EE4END[10]
  PIN bot_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.5578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 22.1811 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.45 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.0600 0.7200 123.4400 ;
    END
  END bot_EE4END[9]
  PIN bot_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 41.956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 224.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 18.5286 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 98.9185 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.3600 0.7200 121.7400 ;
    END
  END bot_EE4END[8]
  PIN bot_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 183.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 17.7491 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 94.3946 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.0000 0.7200 120.3800 ;
    END
  END bot_EE4END[7]
  PIN bot_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 53.0872 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.091 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.6400 0.7200 119.0200 ;
    END
  END bot_EE4END[6]
  PIN bot_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.361 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.05953 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.7576 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 116.9400 0.7200 117.3200 ;
    END
  END bot_EE4END[5]
  PIN bot_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.6378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 31.7696 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 167.729 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.5800 0.7200 115.9600 ;
    END
  END bot_EE4END[4]
  PIN bot_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.7155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.2200 0.7200 114.6000 ;
    END
  END bot_EE4END[3]
  PIN bot_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.6379 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.5200 0.7200 112.9000 ;
    END
  END bot_EE4END[2]
  PIN bot_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.6655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 133.038 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.3104 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.1600 0.7200 111.5400 ;
    END
  END bot_EE4END[1]
  PIN bot_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.9515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.75 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.8958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.8000 0.7200 110.1800 ;
    END
  END bot_EE4END[0]
  PIN bot_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.6504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 16.5709 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 88.6209 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.5800 0.7200 149.9600 ;
    END
  END bot_E6END[11]
  PIN bot_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.5231 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.2343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 147.8800 0.7200 148.2600 ;
    END
  END bot_E6END[10]
  PIN bot_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.627 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 9.98828 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 54.035 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.5200 0.7200 146.9000 ;
    END
  END bot_E6END[9]
  PIN bot_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.0668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 246.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 66.5071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 352.469 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.1600 0.7200 145.5400 ;
    END
  END bot_E6END[8]
  PIN bot_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.62391 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.7448 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.4600 0.7200 143.8400 ;
    END
  END bot_E6END[7]
  PIN bot_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.0328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 52.3734 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 277.048 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.1000 0.7200 142.4800 ;
    END
  END bot_E6END[6]
  PIN bot_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.96195 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.1374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.7400 0.7200 141.1200 ;
    END
  END bot_E6END[5]
  PIN bot_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7211 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 296.647 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.0400 0.7200 139.4200 ;
    END
  END bot_E6END[4]
  PIN bot_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.907 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 49.0377 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.754 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.6800 0.7200 138.0600 ;
    END
  END bot_E6END[3]
  PIN bot_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.662 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 16.1437 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 85.7785 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.3200 0.7200 136.7000 ;
    END
  END bot_E6END[2]
  PIN bot_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.7935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.8864 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.5279 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.2644 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.9694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.6200 0.7200 135.0000 ;
    END
  END bot_E6END[1]
  PIN bot_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.655 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 72.1644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 386.288 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.2600 0.7200 133.6400 ;
    END
  END bot_E6END[0]
  PIN bot_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 172.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 13.9200 0.7200 14.3000 ;
    END
  END bot_W1BEG[3]
  PIN bot_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.5600 0.7200 12.9400 ;
    END
  END bot_W1BEG[2]
  PIN bot_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.1318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.84 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 11.2000 0.7200 11.5800 ;
    END
  END bot_W1BEG[1]
  PIN bot_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.0102 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 481.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.8400 0.7200 10.2200 ;
    END
  END bot_W1BEG[0]
  PIN bot_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.245 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.8200 0.7200 26.2000 ;
    END
  END bot_W2BEG[7]
  PIN bot_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.1896 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 337.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.4600 0.7200 24.8400 ;
    END
  END bot_W2BEG[6]
  PIN bot_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 29.7792 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 148.778 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.7600 0.7200 23.1400 ;
    END
  END bot_W2BEG[5]
  PIN bot_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.925 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.4000 0.7200 21.7800 ;
    END
  END bot_W2BEG[4]
  PIN bot_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.2148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.616 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.0400 0.7200 20.4200 ;
    END
  END bot_W2BEG[3]
  PIN bot_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.9178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.3400 0.7200 18.7200 ;
    END
  END bot_W2BEG[2]
  PIN bot_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.219 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.9800 0.7200 17.3600 ;
    END
  END bot_W2BEG[1]
  PIN bot_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.687 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.6200 0.7200 16.0000 ;
    END
  END bot_W2BEG[0]
  PIN bot_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.8438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 186.304 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.7200 0.7200 38.1000 ;
    END
  END bot_W2BEGb[7]
  PIN bot_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.8648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.416 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.0200 0.7200 36.4000 ;
    END
  END bot_W2BEGb[6]
  PIN bot_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.5518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.08 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.6600 0.7200 35.0400 ;
    END
  END bot_W2BEGb[5]
  PIN bot_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.1418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.56 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.3000 0.7200 33.6800 ;
    END
  END bot_W2BEGb[4]
  PIN bot_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.6000 0.7200 31.9800 ;
    END
  END bot_W2BEGb[3]
  PIN bot_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.2400 0.7200 30.6200 ;
    END
  END bot_W2BEGb[2]
  PIN bot_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 28.8800 0.7200 29.2600 ;
    END
  END bot_W2BEGb[1]
  PIN bot_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.1800 0.7200 27.5600 ;
    END
  END bot_W2BEGb[0]
  PIN bot_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 162.768 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.1800 0.7200 61.5600 ;
    END
  END bot_WW4BEG[15]
  PIN bot_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.0267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.7365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.471 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.8200 0.7200 60.2000 ;
    END
  END bot_WW4BEG[14]
  PIN bot_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.2205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.615 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.1200 0.7200 58.5000 ;
    END
  END bot_WW4BEG[13]
  PIN bot_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.5228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.7600 0.7200 57.1400 ;
    END
  END bot_WW4BEG[12]
  PIN bot_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 44.4558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 237.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.4000 0.7200 55.7800 ;
    END
  END bot_WW4BEG[11]
  PIN bot_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.8588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.384 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.7000 0.7200 54.0800 ;
    END
  END bot_WW4BEG[10]
  PIN bot_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.825 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.3400 0.7200 52.7200 ;
    END
  END bot_WW4BEG[9]
  PIN bot_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 47.2638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 252.544 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 50.9800 0.7200 51.3600 ;
    END
  END bot_WW4BEG[8]
  PIN bot_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.4708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.648 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.2800 0.7200 49.6600 ;
    END
  END bot_WW4BEG[7]
  PIN bot_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.449 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.437 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 47.9200 0.7200 48.3000 ;
    END
  END bot_WW4BEG[6]
  PIN bot_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.65 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.901 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.5600 0.7200 46.9400 ;
    END
  END bot_WW4BEG[5]
  PIN bot_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.8600 0.7200 45.2400 ;
    END
  END bot_WW4BEG[4]
  PIN bot_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.185 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.5000 0.7200 43.8800 ;
    END
  END bot_WW4BEG[3]
  PIN bot_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.1400 0.7200 42.5200 ;
    END
  END bot_WW4BEG[2]
  PIN bot_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.4400 0.7200 40.8200 ;
    END
  END bot_WW4BEG[1]
  PIN bot_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.9778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 288.352 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.0800 0.7200 39.4600 ;
    END
  END bot_WW4BEG[0]
  PIN bot_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.7456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.584 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.8600 0.7200 79.2400 ;
    END
  END bot_W6BEG[11]
  PIN bot_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.7136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 506.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.5000 0.7200 77.8800 ;
    END
  END bot_W6BEG[10]
  PIN bot_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.28 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.8000 0.7200 76.1800 ;
    END
  END bot_W6BEG[9]
  PIN bot_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.8188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.504 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.4400 0.7200 74.8200 ;
    END
  END bot_W6BEG[8]
  PIN bot_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.4588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.584 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.0800 0.7200 73.4600 ;
    END
  END bot_W6BEG[7]
  PIN bot_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.9988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.3800 0.7200 71.7600 ;
    END
  END bot_W6BEG[6]
  PIN bot_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.42 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.0200 0.7200 70.4000 ;
    END
  END bot_W6BEG[5]
  PIN bot_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 42.1578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 225.312 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.6600 0.7200 69.0400 ;
    END
  END bot_W6BEG[4]
  PIN bot_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.9528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.552 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 66.9600 0.7200 67.3400 ;
    END
  END bot_W6BEG[3]
  PIN bot_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.057 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.7398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.416 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.6000 0.7200 65.9800 ;
    END
  END bot_W6BEG[2]
  PIN bot_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.6 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.2400 0.7200 64.6200 ;
    END
  END bot_W6BEG[1]
  PIN bot_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.8838 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.184 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.5400 0.7200 62.9200 ;
    END
  END bot_W6BEG[0]
  PIN bot_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7632 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.0685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.7064 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.7225 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.3246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 13.9200 210.2200 14.3000 ;
    END
  END bot_W1END[3]
  PIN bot_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.8258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 12.5600 210.2200 12.9400 ;
    END
  END bot_W1END[2]
  PIN bot_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8896 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.051 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.4178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.0086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.32 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 11.2000 210.2200 11.5800 ;
    END
  END bot_W1END[1]
  PIN bot_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.5928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 373.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 9.8400 210.2200 10.2200 ;
    END
  END bot_W1END[0]
  PIN bot_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.6607 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 302.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 90.5969 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 482.548 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 25.8200 210.2200 26.2000 ;
    END
  END bot_W2MID[7]
  PIN bot_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.56 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.546 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 344.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 88.6527 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 472.905 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 24.4600 210.2200 24.8400 ;
    END
  END bot_W2MID[6]
  PIN bot_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.2514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.6222 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 100.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.1094 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 471.328 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 138.288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 735.081 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 22.7600 210.2200 23.1400 ;
    END
  END bot_W2MID[5]
  PIN bot_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.261 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 535.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 198.664 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1059.26 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 21.4000 210.2200 21.7800 ;
    END
  END bot_W2MID[4]
  PIN bot_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 59.359 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 317.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.0755 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 310.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 81.5453 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 435.353 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 20.0400 210.2200 20.4200 ;
    END
  END bot_W2MID[3]
  PIN bot_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.087 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.629 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 537.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 153.973 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 820.603 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 18.3400 210.2200 18.7200 ;
    END
  END bot_W2MID[2]
  PIN bot_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4193 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.075 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.0605 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 310.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 91.255 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 486.163 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 16.9800 210.2200 17.3600 ;
    END
  END bot_W2MID[1]
  PIN bot_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.69495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.5455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.86316 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.0754 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.2836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.12 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 89.7064 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 475.173 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 15.6200 210.2200 16.0000 ;
    END
  END bot_W2MID[0]
  PIN bot_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.0264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 174.79 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.8003 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 304.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.855 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 19.0213 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.447 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 37.7200 210.2200 38.1000 ;
    END
  END bot_W2END[7]
  PIN bot_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.5925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.5078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.512 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 36.0200 210.2200 36.4000 ;
    END
  END bot_W2END[6]
  PIN bot_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 103.712 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 554.544 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 34.6600 210.2200 35.0400 ;
    END
  END bot_W2END[5]
  PIN bot_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6065 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.01737 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.171 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.04296 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.6027 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via3  ;
    ANTENNADIFFAREA 1.3176 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.342 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 588.96 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 156.651 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 832.815 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 33.3000 210.2200 33.6800 ;
    END
  END bot_W2END[4]
  PIN bot_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.9735 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 124.47 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 34.0427 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 168.534 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNADIFFAREA 0.9396 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.1916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.616 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 73.358 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 379.465 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.6937 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.556 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 31.6000 210.2200 31.9800 ;
    END
  END bot_W2END[3]
  PIN bot_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.4099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 231.878 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1268 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.6858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 196.128 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 30.2400 210.2200 30.6200 ;
    END
  END bot_W2END[2]
  PIN bot_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.2956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 477.184 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 28.8800 210.2200 29.2600 ;
    END
  END bot_W2END[1]
  PIN bot_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.83717 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.5744 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.51327 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.4754 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.9916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 368.896 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 99.4312 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 529.305 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 27.1800 210.2200 27.5600 ;
    END
  END bot_W2END[0]
  PIN bot_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.8248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 26.1044 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.692 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 61.1800 210.2200 61.5600 ;
    END
  END bot_WW4END[15]
  PIN bot_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.3168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 258.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 66.4527 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 353.122 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 59.8200 210.2200 60.2000 ;
    END
  END bot_WW4END[14]
  PIN bot_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.0108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 25.3609 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 134.149 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 58.1200 210.2200 58.5000 ;
    END
  END bot_WW4END[13]
  PIN bot_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.26532 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 9.77306 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 56.7600 210.2200 57.1400 ;
    END
  END bot_WW4END[12]
  PIN bot_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.973 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 7.18397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 39.7077 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 55.4000 210.2200 55.7800 ;
    END
  END bot_WW4END[11]
  PIN bot_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.689 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 3.40781 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 18.4721 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 53.7000 210.2200 54.0800 ;
    END
  END bot_WW4END[10]
  PIN bot_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9302 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.543 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.27852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.0114 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 52.3400 210.2200 52.7200 ;
    END
  END bot_WW4END[9]
  PIN bot_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.9348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 14.3096 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 78.3933 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 50.9800 210.2200 51.3600 ;
    END
  END bot_WW4END[8]
  PIN bot_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.8278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.552 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 42.27 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 223.908 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 49.2800 210.2200 49.6600 ;
    END
  END bot_WW4END[7]
  PIN bot_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 50.3508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 269.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 72.8784 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 384.873 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 47.9200 210.2200 48.3000 ;
    END
  END bot_WW4END[6]
  PIN bot_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 199.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9652 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 31.2265 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.737 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 46.5600 210.2200 46.9400 ;
    END
  END bot_WW4END[5]
  PIN bot_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.509 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.95313 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.3165 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 44.8600 210.2200 45.2400 ;
    END
  END bot_WW4END[4]
  PIN bot_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.9625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.2229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8542 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.104 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 43.5000 210.2200 43.8800 ;
    END
  END bot_WW4END[3]
  PIN bot_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.102 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 538.8 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 42.1400 210.2200 42.5200 ;
    END
  END bot_WW4END[2]
  PIN bot_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 84.8394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 453.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 40.4400 210.2200 40.8200 ;
    END
  END bot_WW4END[1]
  PIN bot_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.2614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 39.0800 210.2200 39.4600 ;
    END
  END bot_WW4END[0]
  PIN bot_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.7648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 191.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 55.351 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 291.942 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 78.8600 210.2200 79.2400 ;
    END
  END bot_W6END[11]
  PIN bot_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.1888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 41.3825 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 219.253 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 77.5000 210.2200 77.8800 ;
    END
  END bot_W6END[10]
  PIN bot_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.7758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 46.2878 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.861 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 75.8000 210.2200 76.1800 ;
    END
  END bot_W6END[9]
  PIN bot_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.8528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 47.3108 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 250.022 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 74.4400 210.2200 74.8200 ;
    END
  END bot_W6END[8]
  PIN bot_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 17.901 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 94.532 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 73.0800 210.2200 73.4600 ;
    END
  END bot_W6END[7]
  PIN bot_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.1338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 16.6137 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 86.2384 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 71.3800 210.2200 71.7600 ;
    END
  END bot_W6END[6]
  PIN bot_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.07582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 3.98451 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 70.0200 210.2200 70.4000 ;
    END
  END bot_W6END[5]
  PIN bot_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.3928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 34.7554 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 183.446 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 68.6600 210.2200 69.0400 ;
    END
  END bot_W6END[4]
  PIN bot_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.2638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 28.997 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.25 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 66.9600 210.2200 67.3400 ;
    END
  END bot_W6END[3]
  PIN bot_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.0268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 33.1519 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.265 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 65.6000 210.2200 65.9800 ;
    END
  END bot_W6END[2]
  PIN bot_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8601 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.0215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8972 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 64.2400 210.2200 64.6200 ;
    END
  END bot_W6END[1]
  PIN bot_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.2265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7064 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.9224 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 62.5400 210.2200 62.9200 ;
    END
  END bot_W6END[0]
  PIN bot_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.8548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 415.696 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.2200 0.0000 84.6000 0.7200 ;
    END
  END bot_S1BEG[3]
  PIN bot_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.3845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 95.3676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 509.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.8400 0.0000 83.2200 0.7200 ;
    END
  END bot_S1BEG[2]
  PIN bot_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 67.2525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2333 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.1218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.12 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.4600 0.0000 81.8400 0.7200 ;
    END
  END bot_S1BEG[1]
  PIN bot_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.9586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 416.72 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.0800 0.0000 80.4600 0.7200 ;
    END
  END bot_S1BEG[0]
  PIN bot_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.273 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.9538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 105.8400 0.0000 106.2200 0.7200 ;
    END
  END bot_S2BEG[7]
  PIN bot_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.7428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.432 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.4600 0.0000 104.8400 0.7200 ;
    END
  END bot_S2BEG[6]
  PIN bot_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.63795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.4525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.9735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 103.0800 0.0000 103.4600 0.7200 ;
    END
  END bot_S2BEG[5]
  PIN bot_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.539 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.127 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 104.272 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 557.056 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 102.1600 0.0000 102.5400 0.7200 ;
    END
  END bot_S2BEG[4]
  PIN bot_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.9558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 100.7800 0.0000 101.1600 0.7200 ;
    END
  END bot_S2BEG[3]
  PIN bot_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.2538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 353.824 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.4000 0.0000 99.7800 0.7200 ;
    END
  END bot_S2BEG[2]
  PIN bot_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.9556 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 480.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 98.0200 0.0000 98.4000 0.7200 ;
    END
  END bot_S2BEG[1]
  PIN bot_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 73.5978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 392.992 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 96.6400 0.0000 97.0200 0.7200 ;
    END
  END bot_S2BEG[0]
  PIN bot_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 95.2600 0.0000 95.6400 0.7200 ;
    END
  END bot_S2BEGb[7]
  PIN bot_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.2616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.19 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 93.8800 0.0000 94.2600 0.7200 ;
    END
  END bot_S2BEGb[6]
  PIN bot_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.9828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.5000 0.0000 92.8800 0.7200 ;
    END
  END bot_S2BEGb[5]
  PIN bot_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.602 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.156 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 91.1200 0.0000 91.5000 0.7200 ;
    END
  END bot_S2BEGb[4]
  PIN bot_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.9476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 139.384 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 89.7400 0.0000 90.1200 0.7200 ;
    END
  END bot_S2BEGb[3]
  PIN bot_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.5388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.344 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.3600 0.0000 88.7400 0.7200 ;
    END
  END bot_S2BEGb[2]
  PIN bot_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.5048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.17 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 86.9800 0.0000 87.3600 0.7200 ;
    END
  END bot_S2BEGb[1]
  PIN bot_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.5858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.928 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 85.6000 0.0000 85.9800 0.7200 ;
    END
  END bot_S2BEGb[0]
  PIN bot_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.1126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 492.208 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 127.4600 0.0000 127.8400 0.7200 ;
    END
  END bot_S4BEG[15]
  PIN bot_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 72.2046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 386.032 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 126.0800 0.0000 126.4600 0.7200 ;
    END
  END bot_S4BEG[14]
  PIN bot_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.9126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 421.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 125.1600 0.0000 125.5400 0.7200 ;
    END
  END bot_S4BEG[13]
  PIN bot_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 84.6258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 451.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 123.7800 0.0000 124.1600 0.7200 ;
    END
  END bot_S4BEG[12]
  PIN bot_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 122.4000 0.0000 122.7800 0.7200 ;
    END
  END bot_S4BEG[11]
  PIN bot_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 121.0200 0.0000 121.4000 0.7200 ;
    END
  END bot_S4BEG[10]
  PIN bot_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 119.6400 0.0000 120.0200 0.7200 ;
    END
  END bot_S4BEG[9]
  PIN bot_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.098 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 118.2600 0.0000 118.6400 0.7200 ;
    END
  END bot_S4BEG[8]
  PIN bot_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.798 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 116.8800 0.0000 117.2600 0.7200 ;
    END
  END bot_S4BEG[7]
  PIN bot_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 99.6312 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 533.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 115.5000 0.0000 115.8800 0.7200 ;
    END
  END bot_S4BEG[6]
  PIN bot_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 114.1200 0.0000 114.5000 0.7200 ;
    END
  END bot_S4BEG[5]
  PIN bot_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 125.101 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 668.144 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 112.7400 0.0000 113.1200 0.7200 ;
    END
  END bot_S4BEG[4]
  PIN bot_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.048 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.3600 0.0000 111.7400 0.7200 ;
    END
  END bot_S4BEG[3]
  PIN bot_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 109.9800 0.0000 110.3600 0.7200 ;
    END
  END bot_S4BEG[2]
  PIN bot_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 123.088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 657.408 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.6000 0.0000 108.9800 0.7200 ;
    END
  END bot_S4BEG[1]
  PIN bot_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 107.2200 0.0000 107.6000 0.7200 ;
    END
  END bot_S4BEG[0]
  PIN bot_SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 114.232 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 610.176 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 149.0800 0.0000 149.4600 0.7200 ;
    END
  END bot_SS4BEG[15]
  PIN bot_SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.55 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.1976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 487.328 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 148.1600 0.0000 148.5400 0.7200 ;
    END
  END bot_SS4BEG[14]
  PIN bot_SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.925 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 597.872 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 146.7800 0.0000 147.1600 0.7200 ;
    END
  END bot_SS4BEG[13]
  PIN bot_SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.68 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.505 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.0386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 470.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 145.4000 0.0000 145.7800 0.7200 ;
    END
  END bot_SS4BEG[12]
  PIN bot_SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 144.0200 0.0000 144.4000 0.7200 ;
    END
  END bot_SS4BEG[11]
  PIN bot_SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1988 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 142.6400 0.0000 143.0200 0.7200 ;
    END
  END bot_SS4BEG[10]
  PIN bot_SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 141.2600 0.0000 141.6400 0.7200 ;
    END
  END bot_SS4BEG[9]
  PIN bot_SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 139.8800 0.0000 140.2600 0.7200 ;
    END
  END bot_SS4BEG[8]
  PIN bot_SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 138.5000 0.0000 138.8800 0.7200 ;
    END
  END bot_SS4BEG[7]
  PIN bot_SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 137.1200 0.0000 137.5000 0.7200 ;
    END
  END bot_SS4BEG[6]
  PIN bot_SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 135.7400 0.0000 136.1200 0.7200 ;
    END
  END bot_SS4BEG[5]
  PIN bot_SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.002 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 115.522 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 617.056 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 134.3600 0.0000 134.7400 0.7200 ;
    END
  END bot_SS4BEG[4]
  PIN bot_SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.859 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3119 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 117.487 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 627.536 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 132.9800 0.0000 133.3600 0.7200 ;
    END
  END bot_SS4BEG[3]
  PIN bot_SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 131.6000 0.0000 131.9800 0.7200 ;
    END
  END bot_SS4BEG[2]
  PIN bot_SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 130.2200 0.0000 130.6000 0.7200 ;
    END
  END bot_SS4BEG[1]
  PIN bot_SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.67235 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 128.8400 0.0000 129.2200 0.7200 ;
    END
  END bot_SS4BEG[0]
  PIN bot_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 23.3253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 116.456 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.744 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.8400 0.0000 14.2200 0.7200 ;
    END
  END bot_N1END[3]
  PIN bot_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5635 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 38.2612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 189.812 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 12.4600 0.0000 12.8400 0.7200 ;
    END
  END bot_N1END[2]
  PIN bot_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 109.077 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 583.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 11.0800 0.0000 11.4600 0.7200 ;
    END
  END bot_N1END[1]
  PIN bot_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.8214 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.731 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9516 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.3092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.396 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.1600 0.0000 10.5400 0.7200 ;
    END
  END bot_N1END[0]
  PIN bot_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8864 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.0016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.616 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.8800 0.0000 25.2600 0.7200 ;
    END
  END bot_N2MID[7]
  PIN bot_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75055 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.883 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.3644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.7445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9504 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.6115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9504 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.4658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 248.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.5000 0.0000 23.8800 0.7200 ;
    END
  END bot_N2MID[6]
  PIN bot_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.946 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.6525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.4645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.6992 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7157 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.616 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 22.1200 0.0000 22.5000 0.7200 ;
    END
  END bot_N2MID[5]
  PIN bot_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3014 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 81.1806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 433.904 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.7400 0.0000 21.1200 0.7200 ;
    END
  END bot_N2MID[4]
  PIN bot_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.6839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.9045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.2423 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8792 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.7528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 367.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.3600 0.0000 19.7400 0.7200 ;
    END
  END bot_N2MID[3]
  PIN bot_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.7213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.2095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5682 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5048 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.1206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 17.9800 0.0000 18.3600 0.7200 ;
    END
  END bot_N2MID[2]
  PIN bot_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.471 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 20.0269 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.9635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1864 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.072 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.6000 0.0000 16.9800 0.7200 ;
    END
  END bot_N2MID[1]
  PIN bot_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.3248 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.2455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.907 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.8864 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.592 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 15.2200 0.0000 15.6000 0.7200 ;
    END
  END bot_N2MID[0]
  PIN bot_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20995 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.4116 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 46.9805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.0784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 220.496 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.4600 0.0000 35.8400 0.7200 ;
    END
  END bot_N2END[7]
  PIN bot_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.78795 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.927 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.4536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.36 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.0800 0.0000 34.4600 0.7200 ;
    END
  END bot_N2END[6]
  PIN bot_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07695 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.267 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.7111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 143.384 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.2546 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.1600 0.0000 33.5400 0.7200 ;
    END
  END bot_N2END[5]
  PIN bot_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.42375 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.675 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4166 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0055 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 122.021 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 652.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.7800 0.0000 32.1600 0.7200 ;
    END
  END bot_N2END[4]
  PIN bot_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.7308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 356.368 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.4000 0.0000 30.7800 0.7200 ;
    END
  END bot_N2END[3]
  PIN bot_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7663 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.6686 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 425.84 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 29.0200 0.0000 29.4000 0.7200 ;
    END
  END bot_N2END[2]
  PIN bot_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 96.7824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 517.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.6400 0.0000 28.0200 0.7200 ;
    END
  END bot_N2END[1]
  PIN bot_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3248 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 75.4278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 402.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.2600 0.0000 26.6400 0.7200 ;
    END
  END bot_N2END[0]
  PIN bot_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6128 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.946 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.4338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.7744 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 57.0800 0.0000 57.4600 0.7200 ;
    END
  END bot_N4END[15]
  PIN bot_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 15.9191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.3065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.5136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 12.2048 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 61.3461 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 56.1600 0.0000 56.5400 0.7200 ;
    END
  END bot_N4END[14]
  PIN bot_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.28 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.37791 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.4949 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 54.7800 0.0000 55.1600 0.7200 ;
    END
  END bot_N4END[13]
  PIN bot_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38335 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.338 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.27919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.0013 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 53.4000 0.0000 53.7800 0.7200 ;
    END
  END bot_N4END[12]
  PIN bot_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.06 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 34.3046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 170.933 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 48.3542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.741 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 52.0200 0.0000 52.4000 0.7200 ;
    END
  END bot_N4END[11]
  PIN bot_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.9848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 22.3521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 111.472 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.3612 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 11.3329 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 59.8923 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 50.6400 0.0000 51.0200 0.7200 ;
    END
  END bot_N4END[10]
  PIN bot_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.3568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.7803 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.038 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 49.2600 0.0000 49.6400 0.7200 ;
    END
  END bot_N4END[9]
  PIN bot_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.46155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.543 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.433 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.82949 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.8438 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 47.8800 0.0000 48.2600 0.7200 ;
    END
  END bot_N4END[8]
  PIN bot_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.2951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.6165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3209 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 46.5000 0.0000 46.8800 0.7200 ;
    END
  END bot_N4END[7]
  PIN bot_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.29 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.774 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.8046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.232 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 45.1200 0.0000 45.5000 0.7200 ;
    END
  END bot_N4END[6]
  PIN bot_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 28.8038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 143.213 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 43.7400 0.0000 44.1200 0.7200 ;
    END
  END bot_N4END[5]
  PIN bot_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.7073 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.1395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.3600 0.0000 42.7400 0.7200 ;
    END
  END bot_N4END[4]
  PIN bot_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.8808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 421.168 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 40.9800 0.0000 41.3600 0.7200 ;
    END
  END bot_N4END[3]
  PIN bot_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.48155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.5566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.576 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.6000 0.0000 39.9800 0.7200 ;
    END
  END bot_N4END[2]
  PIN bot_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.147 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 113.613 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 607.344 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 38.2200 0.0000 38.6000 0.7200 ;
    END
  END bot_N4END[1]
  PIN bot_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.19255 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.403 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.5268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 259.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.8400 0.0000 37.2200 0.7200 ;
    END
  END bot_N4END[0]
  PIN bot_NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.768 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.88391 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.0249 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 79.1600 0.0000 79.5400 0.7200 ;
    END
  END bot_NN4END[15]
  PIN bot_NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.9956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.86 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0314 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.7623 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.7800 0.0000 78.1600 0.7200 ;
    END
  END bot_NN4END[14]
  PIN bot_NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.0523 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.5734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 27.9438 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 140.069 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 76.4000 0.0000 76.7800 0.7200 ;
    END
  END bot_NN4END[13]
  PIN bot_NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26775 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.315 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.8413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.6815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.5062 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 8.84653 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.7906 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 75.0200 0.0000 75.4000 0.7200 ;
    END
  END bot_NN4END[12]
  PIN bot_NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 18.0041 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.1415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.0848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 25.968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.004 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 73.6400 0.0000 74.0200 0.7200 ;
    END
  END bot_NN4END[11]
  PIN bot_NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.9986 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 40.0949 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 203.942 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 72.2600 0.0000 72.6400 0.7200 ;
    END
  END bot_NN4END[10]
  PIN bot_NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15215 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.179 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 7.03535 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 35.9865 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 70.8800 0.0000 71.2600 0.7200 ;
    END
  END bot_NN4END[9]
  PIN bot_NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11815 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.139 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.4603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.0125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.2806 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.7437 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 105.246 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 69.5000 0.0000 69.8800 0.7200 ;
    END
  END bot_NN4END[8]
  PIN bot_NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61455 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.723 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.4182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.511 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 68.1200 0.0000 68.5000 0.7200 ;
    END
  END bot_NN4END[7]
  PIN bot_NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49895 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.587 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.0268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.78 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.7400 0.0000 67.1200 0.7200 ;
    END
  END bot_NN4END[6]
  PIN bot_NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.32555 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.383 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.7235 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 65.3600 0.0000 65.7400 0.7200 ;
    END
  END bot_NN4END[5]
  PIN bot_NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44115 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3467 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.2728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.592 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 63.9800 0.0000 64.3600 0.7200 ;
    END
  END bot_NN4END[4]
  PIN bot_NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55675 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.655 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.8598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 325.056 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.6000 0.0000 62.9800 0.7200 ;
    END
  END bot_NN4END[3]
  PIN bot_NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 116.078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 619.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.2200 0.0000 61.6000 0.7200 ;
    END
  END bot_NN4END[2]
  PIN bot_NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.5434 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 97.6395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 54.8384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 273.602 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 59.8400 0.0000 60.2200 0.7200 ;
    END
  END bot_NN4END[1]
  PIN bot_NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09435 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.111 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 97.2768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 519.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 58.4600 0.0000 58.8400 0.7200 ;
    END
  END bot_NN4END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.5904 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 8.86514 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 46.424 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 89.5100 0.0000 89.8900 0.7200 ;
    END
  END UserCLK
  PIN top_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.25603 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.5098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.70182 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.5158 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 71.3448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 382.368 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 92.8287 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 492.63 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.889308 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 439.2600 0.7200 439.6400 ;
    END
  END top_FrameData[31]
  PIN top_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.8984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 287.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 75.3841 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 400.273 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 121.422 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 651.328 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 139.966 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 729.092 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.13564 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 437.5600 0.7200 437.9400 ;
    END
  END top_FrameData[30]
  PIN top_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.4018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 291.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 76.9134 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 408.569 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 94.3218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 505.872 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 110.486 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 588.627 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 435.8600 0.7200 436.2400 ;
    END
  END top_FrameData[29]
  PIN top_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.6668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 31.8311 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 167.945 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 67.62 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 362.992 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 101.58 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 524.313 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 434.1600 0.7200 434.5400 ;
    END
  END top_FrameData[28]
  PIN top_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.7415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9825 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.0741 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.7071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 57.567 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.5948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.976 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 59.2038 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.332 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.735704 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 432.4600 0.7200 432.8400 ;
    END
  END top_FrameData[27]
  PIN top_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.8334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 282.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 74.3061 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 394.405 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 73.2648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 391.216 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 100.384 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 533.653 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.845767 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 430.7600 0.7200 431.1400 ;
    END
  END top_FrameData[26]
  PIN top_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 78.1407 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 419.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 118.192 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 605.087 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 428.7200 0.7200 429.1000 ;
    END
  END top_FrameData[25]
  PIN top_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 38.1282 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 200.799 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.261145 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 81.7992 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 438.144 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 114.34 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 592.17 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.88232 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 427.0200 0.7200 427.4000 ;
    END
  END top_FrameData[24]
  PIN top_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.9033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.0045 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 150.55 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 68.241 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 366.304 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 81.6378 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 419.895 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 425.3200 0.7200 425.7000 ;
    END
  END top_FrameData[23]
  PIN top_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 55.1794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 294.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 77.7071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 412.463 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 97.2738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 521.616 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 112.33 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 598.125 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 423.6200 0.7200 424.0000 ;
    END
  END top_FrameData[22]
  PIN top_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 70.7802 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 379.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 111.612 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 564.014 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.845767 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 421.9200 0.7200 422.3000 ;
    END
  END top_FrameData[21]
  PIN top_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.013 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 208.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 70.7823 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 378.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 111.087 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 561.012 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.927044 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 419.8800 0.7200 420.2600 ;
    END
  END top_FrameData[20]
  PIN top_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.0379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 109.449 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 30.089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 148.302 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 34.0661 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 170.142 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.6942 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.456 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 82.8961 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 438.682 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 418.1800 0.7200 418.5600 ;
    END
  END top_FrameData[19]
  PIN top_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.0716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 284.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 77.1122 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 409.495 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.6424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.504 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 93.002 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 494.743 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.02034 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 416.4800 0.7200 416.8600 ;
    END
  END top_FrameData[18]
  PIN top_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.56 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 107.284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 574.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 93.936 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 479.563 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.983979 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 94.5645 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 483.083 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.983979 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 414.7800 0.7200 415.1600 ;
    END
  END top_FrameData[17]
  PIN top_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.4162 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.3963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.032 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 35.2121 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 182.244 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 40.5325 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 198.876 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.987276 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 413.0800 0.7200 413.4600 ;
    END
  END top_FrameData[16]
  PIN top_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 101.73 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 513.061 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.642833 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 411.0400 0.7200 411.4200 ;
    END
  END top_FrameData[15]
  PIN top_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.8285 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 21.2125 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.37 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.4353 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.112 LAYER met3  ;
    ANTENNAGATEAREA 1.0605 LAYER met3  ;
    ANTENNAMAXAREACAR 45.1968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.717 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.612561 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.4636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.08 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 52.8104 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.699 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 409.3400 0.7200 409.7200 ;
    END
  END top_FrameData[14]
  PIN top_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.3874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 116.186 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met2  ;
    ANTENNAMAXAREACAR 27.3786 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 30.5012 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 149.926 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.412011 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.6946 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 79.312 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3195 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.422 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.763522 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 407.6400 0.7200 408.0200 ;
    END
  END top_FrameData[13]
  PIN top_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.2712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 263.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 68.4017 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 363.918 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 66.6276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 356.288 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 92.1169 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 490.733 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.594194 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 405.9400 0.7200 406.3200 ;
    END
  END top_FrameData[12]
  PIN top_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.3019 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 53.2603 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.728 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 404.2400 0.7200 404.6200 ;
    END
  END top_FrameData[11]
  PIN top_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.4636 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 64.2474 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 344.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 77.2302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.061 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.594194 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 402.2000 0.7200 402.5800 ;
    END
  END top_FrameData[10]
  PIN top_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.6556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 217.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 61.8042 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 331.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 80.1368 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 414.494 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 400.5000 0.7200 400.8800 ;
    END
  END top_FrameData[9]
  PIN top_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.9834 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 267.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 69.8622 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 370.87 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.104 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 89.2986 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 475.418 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 398.8000 0.7200 399.1800 ;
    END
  END top_FrameData[8]
  PIN top_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.549 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.011 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 58.3496 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 293.474 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.506709 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 397.1000 0.7200 397.4800 ;
    END
  END top_FrameData[7]
  PIN top_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.07 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.5665 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 75.5694 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 379.297 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.737317 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 395.4000 0.7200 395.7800 ;
    END
  END top_FrameData[6]
  PIN top_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.939 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.651 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.9474 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 72.3148 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 363.839 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.988889 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 393.3600 0.7200 393.7400 ;
    END
  END top_FrameData[5]
  PIN top_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 51.9386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.0312 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 60.5831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.726 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.699131 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 391.6600 0.7200 392.0400 ;
    END
  END top_FrameData[4]
  PIN top_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.8925 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 341.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 94.8314 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 503.886 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.892453 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 389.9600 0.7200 390.3400 ;
    END
  END top_FrameData[3]
  PIN top_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0611 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.9085 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.6119 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.3798 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.6586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.92 LAYER met3  ;
    ANTENNAGATEAREA 2.3325 LAYER met3  ;
    ANTENNAMAXAREACAR 52.779 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 262.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.582558 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 53.9467 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 268.429 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.582558 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 388.2600 0.7200 388.6400 ;
    END
  END top_FrameData[2]
  PIN top_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 58.501 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 314.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met3  ;
    ANTENNAMAXAREACAR 105.906 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 534.733 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.593246 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 106.365 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 537.359 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.05178 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 386.5600 0.7200 386.9400 ;
    END
  END top_FrameData[1]
  PIN top_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 102.501 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 56.0563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 275.278 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.9298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 293.896 LAYER met3  ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 95.9038 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 488.478 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.619583 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.3482 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.072 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 103.204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 528.12 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 384.8600 0.7200 385.2400 ;
    END
  END top_FrameData[0]
  PIN top_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.651 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 439.2600 210.2200 439.6400 ;
    END
  END top_FrameData_O[31]
  PIN top_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 437.5600 210.2200 437.9400 ;
    END
  END top_FrameData_O[30]
  PIN top_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 435.8600 210.2200 436.2400 ;
    END
  END top_FrameData_O[29]
  PIN top_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.96 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 434.1600 210.2200 434.5400 ;
    END
  END top_FrameData_O[28]
  PIN top_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.52 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 432.4600 210.2200 432.8400 ;
    END
  END top_FrameData_O[27]
  PIN top_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 430.7600 210.2200 431.1400 ;
    END
  END top_FrameData_O[26]
  PIN top_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 428.7200 210.2200 429.1000 ;
    END
  END top_FrameData_O[25]
  PIN top_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.56 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 427.0200 210.2200 427.4000 ;
    END
  END top_FrameData_O[24]
  PIN top_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 425.3200 210.2200 425.7000 ;
    END
  END top_FrameData_O[23]
  PIN top_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.687 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 423.6200 210.2200 424.0000 ;
    END
  END top_FrameData_O[22]
  PIN top_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.219 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 421.9200 210.2200 422.3000 ;
    END
  END top_FrameData_O[21]
  PIN top_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 419.8800 210.2200 420.2600 ;
    END
  END top_FrameData_O[20]
  PIN top_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.449 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 418.1800 210.2200 418.5600 ;
    END
  END top_FrameData_O[19]
  PIN top_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 416.4800 210.2200 416.8600 ;
    END
  END top_FrameData_O[18]
  PIN top_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.392 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 414.7800 210.2200 415.1600 ;
    END
  END top_FrameData_O[17]
  PIN top_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.174 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 413.0800 210.2200 413.4600 ;
    END
  END top_FrameData_O[16]
  PIN top_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 411.0400 210.2200 411.4200 ;
    END
  END top_FrameData_O[15]
  PIN top_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 409.3400 210.2200 409.7200 ;
    END
  END top_FrameData_O[14]
  PIN top_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 407.6400 210.2200 408.0200 ;
    END
  END top_FrameData_O[13]
  PIN top_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 405.9400 210.2200 406.3200 ;
    END
  END top_FrameData_O[12]
  PIN top_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.0508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 404.2400 210.2200 404.6200 ;
    END
  END top_FrameData_O[11]
  PIN top_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6128 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.946 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 402.2000 210.2200 402.5800 ;
    END
  END top_FrameData_O[10]
  PIN top_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 400.5000 210.2200 400.8800 ;
    END
  END top_FrameData_O[9]
  PIN top_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 398.8000 210.2200 399.1800 ;
    END
  END top_FrameData_O[8]
  PIN top_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.282 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 397.1000 210.2200 397.4800 ;
    END
  END top_FrameData_O[7]
  PIN top_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 395.4000 210.2200 395.7800 ;
    END
  END top_FrameData_O[6]
  PIN top_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 393.3600 210.2200 393.7400 ;
    END
  END top_FrameData_O[5]
  PIN top_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 391.6600 210.2200 392.0400 ;
    END
  END top_FrameData_O[4]
  PIN top_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.52 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 389.9600 210.2200 390.3400 ;
    END
  END top_FrameData_O[3]
  PIN top_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 388.2600 210.2200 388.6400 ;
    END
  END top_FrameData_O[2]
  PIN top_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.28 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 386.5600 210.2200 386.9400 ;
    END
  END top_FrameData_O[1]
  PIN top_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 384.8600 210.2200 385.2400 ;
    END
  END top_FrameData_O[0]
  PIN bot_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.0772 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 59.3175 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 293.499 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.858193 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 59.6203 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.281 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.858193 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 209.4200 0.7200 209.8000 ;
    END
  END bot_FrameData[31]
  PIN bot_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.2274 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 83.3967 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 425.732 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 207.7200 0.7200 208.1000 ;
    END
  END bot_FrameData[30]
  PIN bot_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.2275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 37.7272 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 183.282 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.669182 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 38.4646 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 187.949 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.732075 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.1042 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.104 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 58.5141 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 294.936 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.03353 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 206.0200 0.7200 206.4000 ;
    END
  END bot_FrameData[29]
  PIN bot_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.9658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 69.658 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.661 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.856376 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 204.3200 0.7200 204.7000 ;
    END
  END bot_FrameData[28]
  PIN bot_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.0768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 86.131 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 436.812 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.5426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.52 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 100.562 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 514.947 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.910273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 202.6200 0.7200 203.0000 ;
    END
  END bot_FrameData[27]
  PIN bot_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 44.7679 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 217.726 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.701 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 219.424 LAYER met3  ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 59.2548 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 295.827 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 200.9200 0.7200 201.3000 ;
    END
  END bot_FrameData[26]
  PIN bot_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.6332 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 97.9838 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 502.747 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 198.8800 0.7200 199.2600 ;
    END
  END bot_FrameData[25]
  PIN bot_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 58.1107 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 310.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 89.543 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 464.701 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.870786 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.9481 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.6 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 100.203 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 522.22 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 197.1800 0.7200 197.5600 ;
    END
  END bot_FrameData[24]
  PIN bot_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.0948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 42.1201 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 210.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.6627 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.352 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 66.2327 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 338.559 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 195.4800 0.7200 195.8600 ;
    END
  END bot_FrameData[23]
  PIN bot_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.9595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.7775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 39.4936 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 192.417 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.088 LAYER met3  ;
    ANTENNAGATEAREA 2.0145 LAYER met3  ;
    ANTENNAMAXAREACAR 55.2871 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 277.346 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.652351 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.3876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.008 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 62.2326 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.376 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 193.7800 0.7200 194.1600 ;
    END
  END bot_FrameData[22]
  PIN bot_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.1137 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 76.2447 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 392.633 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 192.0800 0.7200 192.4600 ;
    END
  END bot_FrameData[21]
  PIN bot_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.914 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met2  ;
    ANTENNAMAXAREACAR 47.1268 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 229.521 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.706918 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.765 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.68 LAYER met3  ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 80.7935 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 410.25 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.807547 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.4182 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.112 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 85.2135 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 434.494 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.807547 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 190.0400 0.7200 190.4200 ;
    END
  END bot_FrameData[20]
  PIN bot_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2765 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.501 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 88.2185 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 445.373 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 188.3400 0.7200 188.7200 ;
    END
  END bot_FrameData[19]
  PIN bot_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.3656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.7729 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 65.5678 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 347.014 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 186.6400 0.7200 187.0200 ;
    END
  END bot_FrameData[18]
  PIN bot_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.38 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.0406 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 75.1438 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 382.936 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.684157 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 184.9400 0.7200 185.3200 ;
    END
  END bot_FrameData[17]
  PIN bot_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 104.146 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 519.412 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.982162 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 183.2400 0.7200 183.6200 ;
    END
  END bot_FrameData[16]
  PIN bot_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.8857 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 203.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 114.243 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 587.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.1608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.68 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 123.911 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 640.005 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 181.2000 0.7200 181.5800 ;
    END
  END bot_FrameData[15]
  PIN bot_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.0525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.4408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 93.278 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 477.906 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.6006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.144 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 103.102 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 530.635 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 179.5000 0.7200 179.8800 ;
    END
  END bot_FrameData[14]
  PIN bot_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 84.3778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 451.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met3  ;
    ANTENNAMAXAREACAR 104.004 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 528.943 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.736208 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 104.372 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 531.073 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.736208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 177.8000 0.7200 178.1800 ;
    END
  END bot_FrameData[13]
  PIN bot_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.8538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 250.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 81.6425 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 427.514 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.261145 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.3719 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.664 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 92.8089 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 487.904 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 176.1000 0.7200 176.4800 ;
    END
  END bot_FrameData[12]
  PIN bot_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.5485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8555 LAYER met2  ;
    ANTENNAMAXAREACAR 32.5721 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 158.155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.486337 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.9069 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.632 LAYER met3  ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 38.8184 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 190.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.543728 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 39.0561 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 191.835 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 174.4000 0.7200 174.7800 ;
    END
  END bot_FrameData[11]
  PIN bot_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4633 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.97239 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.1051 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.696 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.6869 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.9088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.984 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 82.272 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 413.965 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.594194 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 172.3600 0.7200 172.7400 ;
    END
  END bot_FrameData[10]
  PIN bot_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.4818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 55.9542 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.908 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.604803 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 170.6600 0.7200 171.0400 ;
    END
  END bot_FrameData[9]
  PIN bot_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.013 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.829 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 69.5372 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 351.258 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04654 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 168.9600 0.7200 169.3400 ;
    END
  END bot_FrameData[8]
  PIN bot_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.563 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 58.3929 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 313.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 100.461 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 523.478 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 167.2600 0.7200 167.6400 ;
    END
  END bot_FrameData[7]
  PIN bot_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.4314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 45.1356 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 225.349 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.669514 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 46.1743 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 231.391 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.669514 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 165.5600 0.7200 165.9400 ;
    END
  END bot_FrameData[6]
  PIN bot_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.6305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.485 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.0802 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 122.037 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 631.952 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.34528 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 163.5200 0.7200 163.9000 ;
    END
  END bot_FrameData[5]
  PIN bot_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.5135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.8061 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 294.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 88.5848 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 444.56 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 161.8200 0.7200 162.2000 ;
    END
  END bot_FrameData[4]
  PIN bot_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.4536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 301.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.2794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 59.0684 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.749 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.987276 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 160.1200 0.7200 160.5000 ;
    END
  END bot_FrameData[3]
  PIN bot_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.7842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 87.7283 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 450.417 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.87673 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 158.4200 0.7200 158.8000 ;
    END
  END bot_FrameData[2]
  PIN bot_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.7539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 218.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 80.9948 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 424.274 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.2624 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.144 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 84.6476 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 444.257 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.00764 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 156.7200 0.7200 157.1000 ;
    END
  END bot_FrameData[1]
  PIN bot_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 62.589 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 335.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met3  ;
    ANTENNAMAXAREACAR 89.2537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 448.084 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 155.0200 0.7200 155.4000 ;
    END
  END bot_FrameData[0]
  PIN bot_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.633 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 209.4200 210.2200 209.8000 ;
    END
  END bot_FrameData_O[31]
  PIN bot_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.5348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.656 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 207.7200 210.2200 208.1000 ;
    END
  END bot_FrameData_O[30]
  PIN bot_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.064 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 206.0200 210.2200 206.4000 ;
    END
  END bot_FrameData_O[29]
  PIN bot_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 204.3200 210.2200 204.7000 ;
    END
  END bot_FrameData_O[28]
  PIN bot_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 202.6200 210.2200 203.0000 ;
    END
  END bot_FrameData_O[27]
  PIN bot_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 200.9200 210.2200 201.3000 ;
    END
  END bot_FrameData_O[26]
  PIN bot_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 198.8800 210.2200 199.2600 ;
    END
  END bot_FrameData_O[25]
  PIN bot_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 197.1800 210.2200 197.5600 ;
    END
  END bot_FrameData_O[24]
  PIN bot_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.0248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.936 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 195.4800 210.2200 195.8600 ;
    END
  END bot_FrameData_O[23]
  PIN bot_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 193.7800 210.2200 194.1600 ;
    END
  END bot_FrameData_O[22]
  PIN bot_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.0428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.032 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 192.0800 210.2200 192.4600 ;
    END
  END bot_FrameData_O[21]
  PIN bot_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.5148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.216 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 190.0400 210.2200 190.4200 ;
    END
  END bot_FrameData_O[20]
  PIN bot_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2765 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.824 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 188.3400 210.2200 188.7200 ;
    END
  END bot_FrameData_O[19]
  PIN bot_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.457 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 186.6400 210.2200 187.0200 ;
    END
  END bot_FrameData_O[18]
  PIN bot_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.904 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 184.9400 210.2200 185.3200 ;
    END
  END bot_FrameData_O[17]
  PIN bot_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 183.2400 210.2200 183.6200 ;
    END
  END bot_FrameData_O[16]
  PIN bot_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.6758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 181.2000 210.2200 181.5800 ;
    END
  END bot_FrameData_O[15]
  PIN bot_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.6308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.168 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 179.5000 210.2200 179.8800 ;
    END
  END bot_FrameData_O[14]
  PIN bot_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 177.8000 210.2200 178.1800 ;
    END
  END bot_FrameData_O[13]
  PIN bot_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.539 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 176.1000 210.2200 176.4800 ;
    END
  END bot_FrameData_O[12]
  PIN bot_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.3348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 306.256 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 174.4000 210.2200 174.7800 ;
    END
  END bot_FrameData_O[11]
  PIN bot_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.232 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 257.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 172.3600 210.2200 172.7400 ;
    END
  END bot_FrameData_O[10]
  PIN bot_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 170.6600 210.2200 171.0400 ;
    END
  END bot_FrameData_O[9]
  PIN bot_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 168.9600 210.2200 169.3400 ;
    END
  END bot_FrameData_O[8]
  PIN bot_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 167.2600 210.2200 167.6400 ;
    END
  END bot_FrameData_O[7]
  PIN bot_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 165.5600 210.2200 165.9400 ;
    END
  END bot_FrameData_O[6]
  PIN bot_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.015 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 163.5200 210.2200 163.9000 ;
    END
  END bot_FrameData_O[5]
  PIN bot_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 161.8200 210.2200 162.2000 ;
    END
  END bot_FrameData_O[4]
  PIN bot_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 160.1200 210.2200 160.5000 ;
    END
  END bot_FrameData_O[3]
  PIN bot_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.639 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 158.4200 210.2200 158.8000 ;
    END
  END bot_FrameData_O[2]
  PIN bot_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 156.7200 210.2200 157.1000 ;
    END
  END bot_FrameData_O[1]
  PIN bot_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.777 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.5000 155.0200 210.2200 155.4000 ;
    END
  END bot_FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.755 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.84094 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.8236 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 199.6800 0.0000 200.0600 0.7200 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.663 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.62168 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.7273 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 196.9200 0.0000 197.3000 0.7200 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.925 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.84606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8492 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 194.6200 0.0000 195.0000 0.7200 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.998 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 26.9754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.86 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 192.3200 0.0000 192.7000 0.7200 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.0168 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 190.0200 0.0000 190.4000 0.7200 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.9889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 208.604 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.9876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 17.4536 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.5529 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 187.2600 0.0000 187.6400 0.7200 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.139 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.97657 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.5926 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 185.4200 0.0000 185.8000 0.7200 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.5284 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 62.3714 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 310.741 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 183.1200 0.0000 183.5000 0.7200 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 76.7394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 410.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 48.6702 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.809 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.640709 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 180.3600 0.0000 180.7400 0.7200 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.2704 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 51.126 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 252.92 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.687444 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 178.5200 0.0000 178.9000 0.7200 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 72.9873 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 390.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 82.5836 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 435.411 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07583 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 175.7600 0.0000 176.1400 0.7200 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.8222 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 34.5529 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.384 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.547021 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 173.9200 0.0000 174.3000 0.7200 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.6248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 32.9342 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.22 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.66168 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 171.6200 0.0000 172.0000 0.7200 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 79.842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 428.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 47.4023 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.25 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.757449 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 169.3200 0.0000 169.7000 0.7200 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 60.1956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 324.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 44.1491 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219.901 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 167.0200 0.0000 167.4000 0.7200 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.319 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 75.0504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 404.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 79.1212 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 407.636 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.897005 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 164.2600 0.0000 164.6400 0.7200 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.5801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 157.042 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met2  ;
    ANTENNAMAXAREACAR 49.9013 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.076 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.512828 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 50.3818 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 242.199 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.560876 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.4578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.912 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 62.8947 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 314.592 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.976909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 162.4200 0.0000 162.8000 0.7200 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 62.6649 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 336.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 53.098 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 268.514 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.981971 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 160.1200 0.0000 160.5000 0.7200 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.8686 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 55.4722 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 277.517 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.730398 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.3600 0.0000 157.7400 0.7200 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.3296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 74.4417 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.014 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.790775 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 155.5200 0.0000 155.9000 0.7200 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.469 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 199.6800 449.1000 200.0600 449.8200 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 61.4214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 306.999 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 196.9200 449.1000 197.3000 449.8200 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.8241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.9595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.5116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 194.6200 449.1000 195.0000 449.8200 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.3200 449.1000 192.7000 449.8200 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.703 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.0200 449.1000 190.4000 449.8200 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.141 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 187.7200 449.1000 188.1000 449.8200 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.5888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 185.4200 449.1000 185.8000 449.8200 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.6666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 372.496 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 183.1200 449.1000 183.5000 449.8200 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.6378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 275.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 180.8200 449.1000 181.2000 449.8200 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.907 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.9456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 357.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 178.5200 449.1000 178.9000 449.8200 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.2200 449.1000 176.6000 449.8200 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.4728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 173.9200 449.1000 174.3000 449.8200 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.2718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 289.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 171.6200 449.1000 172.0000 449.8200 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.2998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 169.3200 449.1000 169.7000 449.8200 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.2228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 422.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 167.0200 449.1000 167.4000 449.8200 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.2286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 418.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 164.7200 449.1000 165.1000 449.8200 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 372.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 162.4200 449.1000 162.8000 449.8200 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 71.4018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 381.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 160.1200 449.1000 160.5000 449.8200 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2985 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 80.1858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 428.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 157.8200 449.1000 158.2000 449.8200 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.6158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 345.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 155.5200 449.1000 155.9000 449.8200 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 204.6600 7.4300 ;
        RECT 5.5600 442.2200 204.6600 444.2200 ;
        RECT 5.5600 224.5000 7.5600 224.9800 ;
        RECT 202.6600 224.5000 204.6600 224.9800 ;
        RECT 5.5600 55.8600 7.5600 56.3400 ;
        RECT 5.5600 12.3400 7.5600 12.8200 ;
        RECT 5.5600 17.7800 7.5600 18.2600 ;
        RECT 5.5600 23.2200 7.5600 23.7000 ;
        RECT 5.5600 28.6600 7.5600 29.1400 ;
        RECT 5.5600 34.1000 7.5600 34.5800 ;
        RECT 5.5600 39.5400 7.5600 40.0200 ;
        RECT 5.5600 44.9800 7.5600 45.4600 ;
        RECT 5.5600 50.4200 7.5600 50.9000 ;
        RECT 5.5600 61.3000 7.5600 61.7800 ;
        RECT 5.5600 66.7400 7.5600 67.2200 ;
        RECT 5.5600 72.1800 7.5600 72.6600 ;
        RECT 5.5600 77.6200 7.5600 78.1000 ;
        RECT 5.5600 83.0600 7.5600 83.5400 ;
        RECT 5.5600 88.5000 7.5600 88.9800 ;
        RECT 5.5600 93.9400 7.5600 94.4200 ;
        RECT 5.5600 99.3800 7.5600 99.8600 ;
        RECT 5.5600 104.8200 7.5600 105.3000 ;
        RECT 5.5600 110.2600 7.5600 110.7400 ;
        RECT 5.5600 115.7000 7.5600 116.1800 ;
        RECT 5.5600 121.1400 7.5600 121.6200 ;
        RECT 5.5600 126.5800 7.5600 127.0600 ;
        RECT 5.5600 132.0200 7.5600 132.5000 ;
        RECT 5.5600 137.4600 7.5600 137.9400 ;
        RECT 5.5600 142.9000 7.5600 143.3800 ;
        RECT 5.5600 148.3400 7.5600 148.8200 ;
        RECT 5.5600 153.7800 7.5600 154.2600 ;
        RECT 5.5600 159.2200 7.5600 159.7000 ;
        RECT 5.5600 164.6600 7.5600 165.1400 ;
        RECT 5.5600 170.1000 7.5600 170.5800 ;
        RECT 5.5600 175.5400 7.5600 176.0200 ;
        RECT 5.5600 180.9800 7.5600 181.4600 ;
        RECT 5.5600 186.4200 7.5600 186.9000 ;
        RECT 5.5600 191.8600 7.5600 192.3400 ;
        RECT 5.5600 197.3000 7.5600 197.7800 ;
        RECT 5.5600 202.7400 7.5600 203.2200 ;
        RECT 5.5600 208.1800 7.5600 208.6600 ;
        RECT 5.5600 213.6200 7.5600 214.1000 ;
        RECT 5.5600 219.0600 7.5600 219.5400 ;
        RECT 202.6600 55.8600 204.6600 56.3400 ;
        RECT 202.6600 12.3400 204.6600 12.8200 ;
        RECT 202.6600 17.7800 204.6600 18.2600 ;
        RECT 202.6600 23.2200 204.6600 23.7000 ;
        RECT 202.6600 28.6600 204.6600 29.1400 ;
        RECT 202.6600 34.1000 204.6600 34.5800 ;
        RECT 202.6600 39.5400 204.6600 40.0200 ;
        RECT 202.6600 44.9800 204.6600 45.4600 ;
        RECT 202.6600 50.4200 204.6600 50.9000 ;
        RECT 202.6600 61.3000 204.6600 61.7800 ;
        RECT 202.6600 66.7400 204.6600 67.2200 ;
        RECT 202.6600 72.1800 204.6600 72.6600 ;
        RECT 202.6600 77.6200 204.6600 78.1000 ;
        RECT 202.6600 83.0600 204.6600 83.5400 ;
        RECT 202.6600 88.5000 204.6600 88.9800 ;
        RECT 202.6600 93.9400 204.6600 94.4200 ;
        RECT 202.6600 99.3800 204.6600 99.8600 ;
        RECT 202.6600 104.8200 204.6600 105.3000 ;
        RECT 202.6600 110.2600 204.6600 110.7400 ;
        RECT 202.6600 115.7000 204.6600 116.1800 ;
        RECT 202.6600 121.1400 204.6600 121.6200 ;
        RECT 202.6600 126.5800 204.6600 127.0600 ;
        RECT 202.6600 132.0200 204.6600 132.5000 ;
        RECT 202.6600 137.4600 204.6600 137.9400 ;
        RECT 202.6600 142.9000 204.6600 143.3800 ;
        RECT 202.6600 148.3400 204.6600 148.8200 ;
        RECT 202.6600 153.7800 204.6600 154.2600 ;
        RECT 202.6600 159.2200 204.6600 159.7000 ;
        RECT 202.6600 164.6600 204.6600 165.1400 ;
        RECT 202.6600 170.1000 204.6600 170.5800 ;
        RECT 202.6600 175.5400 204.6600 176.0200 ;
        RECT 202.6600 180.9800 204.6600 181.4600 ;
        RECT 202.6600 186.4200 204.6600 186.9000 ;
        RECT 202.6600 191.8600 204.6600 192.3400 ;
        RECT 202.6600 197.3000 204.6600 197.7800 ;
        RECT 202.6600 202.7400 204.6600 203.2200 ;
        RECT 202.6600 208.1800 204.6600 208.6600 ;
        RECT 202.6600 213.6200 204.6600 214.1000 ;
        RECT 202.6600 219.0600 204.6600 219.5400 ;
        RECT 5.5600 229.9400 7.5600 230.4200 ;
        RECT 5.5600 235.3800 7.5600 235.8600 ;
        RECT 5.5600 240.8200 7.5600 241.3000 ;
        RECT 5.5600 246.2600 7.5600 246.7400 ;
        RECT 5.5600 251.7000 7.5600 252.1800 ;
        RECT 5.5600 257.1400 7.5600 257.6200 ;
        RECT 5.5600 262.5800 7.5600 263.0600 ;
        RECT 5.5600 268.0200 7.5600 268.5000 ;
        RECT 5.5600 273.4600 7.5600 273.9400 ;
        RECT 5.5600 278.9000 7.5600 279.3800 ;
        RECT 5.5600 284.3400 7.5600 284.8200 ;
        RECT 5.5600 289.7800 7.5600 290.2600 ;
        RECT 5.5600 295.2200 7.5600 295.7000 ;
        RECT 5.5600 300.6600 7.5600 301.1400 ;
        RECT 5.5600 306.1000 7.5600 306.5800 ;
        RECT 5.5600 311.5400 7.5600 312.0200 ;
        RECT 5.5600 316.9800 7.5600 317.4600 ;
        RECT 5.5600 322.4200 7.5600 322.9000 ;
        RECT 5.5600 327.8600 7.5600 328.3400 ;
        RECT 5.5600 333.3000 7.5600 333.7800 ;
        RECT 5.5600 393.1400 7.5600 393.6200 ;
        RECT 5.5600 338.7400 7.5600 339.2200 ;
        RECT 5.5600 344.1800 7.5600 344.6600 ;
        RECT 5.5600 349.6200 7.5600 350.1000 ;
        RECT 5.5600 355.0600 7.5600 355.5400 ;
        RECT 5.5600 360.5000 7.5600 360.9800 ;
        RECT 5.5600 365.9400 7.5600 366.4200 ;
        RECT 5.5600 371.3800 7.5600 371.8600 ;
        RECT 5.5600 376.8200 7.5600 377.3000 ;
        RECT 5.5600 382.2600 7.5600 382.7400 ;
        RECT 5.5600 387.7000 7.5600 388.1800 ;
        RECT 5.5600 398.5800 7.5600 399.0600 ;
        RECT 5.5600 404.0200 7.5600 404.5000 ;
        RECT 5.5600 409.4600 7.5600 409.9400 ;
        RECT 5.5600 414.9000 7.5600 415.3800 ;
        RECT 5.5600 420.3400 7.5600 420.8200 ;
        RECT 5.5600 425.7800 7.5600 426.2600 ;
        RECT 5.5600 431.2200 7.5600 431.7000 ;
        RECT 5.5600 436.6600 7.5600 437.1400 ;
        RECT 202.6600 229.9400 204.6600 230.4200 ;
        RECT 202.6600 235.3800 204.6600 235.8600 ;
        RECT 202.6600 240.8200 204.6600 241.3000 ;
        RECT 202.6600 246.2600 204.6600 246.7400 ;
        RECT 202.6600 251.7000 204.6600 252.1800 ;
        RECT 202.6600 257.1400 204.6600 257.6200 ;
        RECT 202.6600 262.5800 204.6600 263.0600 ;
        RECT 202.6600 268.0200 204.6600 268.5000 ;
        RECT 202.6600 273.4600 204.6600 273.9400 ;
        RECT 202.6600 278.9000 204.6600 279.3800 ;
        RECT 202.6600 284.3400 204.6600 284.8200 ;
        RECT 202.6600 289.7800 204.6600 290.2600 ;
        RECT 202.6600 295.2200 204.6600 295.7000 ;
        RECT 202.6600 300.6600 204.6600 301.1400 ;
        RECT 202.6600 306.1000 204.6600 306.5800 ;
        RECT 202.6600 311.5400 204.6600 312.0200 ;
        RECT 202.6600 316.9800 204.6600 317.4600 ;
        RECT 202.6600 322.4200 204.6600 322.9000 ;
        RECT 202.6600 327.8600 204.6600 328.3400 ;
        RECT 202.6600 333.3000 204.6600 333.7800 ;
        RECT 202.6600 393.1400 204.6600 393.6200 ;
        RECT 202.6600 338.7400 204.6600 339.2200 ;
        RECT 202.6600 344.1800 204.6600 344.6600 ;
        RECT 202.6600 349.6200 204.6600 350.1000 ;
        RECT 202.6600 355.0600 204.6600 355.5400 ;
        RECT 202.6600 360.5000 204.6600 360.9800 ;
        RECT 202.6600 365.9400 204.6600 366.4200 ;
        RECT 202.6600 371.3800 204.6600 371.8600 ;
        RECT 202.6600 376.8200 204.6600 377.3000 ;
        RECT 202.6600 382.2600 204.6600 382.7400 ;
        RECT 202.6600 387.7000 204.6600 388.1800 ;
        RECT 202.6600 398.5800 204.6600 399.0600 ;
        RECT 202.6600 404.0200 204.6600 404.5000 ;
        RECT 202.6600 409.4600 204.6600 409.9400 ;
        RECT 202.6600 414.9000 204.6600 415.3800 ;
        RECT 202.6600 420.3400 204.6600 420.8200 ;
        RECT 202.6600 425.7800 204.6600 426.2600 ;
        RECT 202.6600 431.2200 204.6600 431.7000 ;
        RECT 202.6600 436.6600 204.6600 437.1400 ;
      LAYER met4 ;
        RECT 190.1200 5.4300 191.7200 444.2200 ;
        RECT 145.1200 5.4300 146.7200 444.2200 ;
        RECT 100.1200 5.4300 101.7200 444.2200 ;
        RECT 55.1200 5.4300 56.7200 444.2200 ;
        RECT 10.1200 5.4300 11.7200 444.2200 ;
        RECT 202.6600 5.4300 204.6600 444.2200 ;
        RECT 5.5600 5.4300 7.5600 444.2200 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 2.4300 207.6600 4.4300 ;
        RECT 2.5600 445.2200 207.6600 447.2200 ;
        RECT 2.5600 9.6200 4.5600 10.1000 ;
        RECT 2.5600 15.0600 4.5600 15.5400 ;
        RECT 2.5600 20.5000 4.5600 20.9800 ;
        RECT 2.5600 25.9400 4.5600 26.4200 ;
        RECT 2.5600 31.3800 4.5600 31.8600 ;
        RECT 2.5600 36.8200 4.5600 37.3000 ;
        RECT 2.5600 42.2600 4.5600 42.7400 ;
        RECT 2.5600 47.7000 4.5600 48.1800 ;
        RECT 2.5600 53.1400 4.5600 53.6200 ;
        RECT 2.5600 58.5800 4.5600 59.0600 ;
        RECT 2.5600 64.0200 4.5600 64.5000 ;
        RECT 2.5600 69.4600 4.5600 69.9400 ;
        RECT 2.5600 74.9000 4.5600 75.3800 ;
        RECT 2.5600 80.3400 4.5600 80.8200 ;
        RECT 2.5600 85.7800 4.5600 86.2600 ;
        RECT 2.5600 91.2200 4.5600 91.7000 ;
        RECT 2.5600 96.6600 4.5600 97.1400 ;
        RECT 2.5600 102.1000 4.5600 102.5800 ;
        RECT 2.5600 107.5400 4.5600 108.0200 ;
        RECT 2.5600 140.1800 4.5600 140.6600 ;
        RECT 2.5600 112.9800 4.5600 113.4600 ;
        RECT 2.5600 118.4200 4.5600 118.9000 ;
        RECT 2.5600 123.8600 4.5600 124.3400 ;
        RECT 2.5600 129.3000 4.5600 129.7800 ;
        RECT 2.5600 134.7400 4.5600 135.2200 ;
        RECT 2.5600 145.6200 4.5600 146.1000 ;
        RECT 2.5600 151.0600 4.5600 151.5400 ;
        RECT 2.5600 156.5000 4.5600 156.9800 ;
        RECT 2.5600 161.9400 4.5600 162.4200 ;
        RECT 2.5600 167.3800 4.5600 167.8600 ;
        RECT 2.5600 172.8200 4.5600 173.3000 ;
        RECT 2.5600 178.2600 4.5600 178.7400 ;
        RECT 2.5600 183.7000 4.5600 184.1800 ;
        RECT 2.5600 189.1400 4.5600 189.6200 ;
        RECT 2.5600 194.5800 4.5600 195.0600 ;
        RECT 2.5600 200.0200 4.5600 200.5000 ;
        RECT 2.5600 205.4600 4.5600 205.9400 ;
        RECT 2.5600 210.9000 4.5600 211.3800 ;
        RECT 2.5600 216.3400 4.5600 216.8200 ;
        RECT 2.5600 221.7800 4.5600 222.2600 ;
        RECT 205.6600 9.6200 207.6600 10.1000 ;
        RECT 205.6600 15.0600 207.6600 15.5400 ;
        RECT 205.6600 20.5000 207.6600 20.9800 ;
        RECT 205.6600 25.9400 207.6600 26.4200 ;
        RECT 205.6600 31.3800 207.6600 31.8600 ;
        RECT 205.6600 36.8200 207.6600 37.3000 ;
        RECT 205.6600 42.2600 207.6600 42.7400 ;
        RECT 205.6600 47.7000 207.6600 48.1800 ;
        RECT 205.6600 53.1400 207.6600 53.6200 ;
        RECT 205.6600 58.5800 207.6600 59.0600 ;
        RECT 205.6600 64.0200 207.6600 64.5000 ;
        RECT 205.6600 69.4600 207.6600 69.9400 ;
        RECT 205.6600 74.9000 207.6600 75.3800 ;
        RECT 205.6600 80.3400 207.6600 80.8200 ;
        RECT 205.6600 85.7800 207.6600 86.2600 ;
        RECT 205.6600 91.2200 207.6600 91.7000 ;
        RECT 205.6600 96.6600 207.6600 97.1400 ;
        RECT 205.6600 102.1000 207.6600 102.5800 ;
        RECT 205.6600 107.5400 207.6600 108.0200 ;
        RECT 205.6600 140.1800 207.6600 140.6600 ;
        RECT 205.6600 112.9800 207.6600 113.4600 ;
        RECT 205.6600 118.4200 207.6600 118.9000 ;
        RECT 205.6600 123.8600 207.6600 124.3400 ;
        RECT 205.6600 129.3000 207.6600 129.7800 ;
        RECT 205.6600 134.7400 207.6600 135.2200 ;
        RECT 205.6600 145.6200 207.6600 146.1000 ;
        RECT 205.6600 151.0600 207.6600 151.5400 ;
        RECT 205.6600 156.5000 207.6600 156.9800 ;
        RECT 205.6600 161.9400 207.6600 162.4200 ;
        RECT 205.6600 167.3800 207.6600 167.8600 ;
        RECT 205.6600 172.8200 207.6600 173.3000 ;
        RECT 205.6600 178.2600 207.6600 178.7400 ;
        RECT 205.6600 183.7000 207.6600 184.1800 ;
        RECT 205.6600 189.1400 207.6600 189.6200 ;
        RECT 205.6600 194.5800 207.6600 195.0600 ;
        RECT 205.6600 200.0200 207.6600 200.5000 ;
        RECT 205.6600 205.4600 207.6600 205.9400 ;
        RECT 205.6600 210.9000 207.6600 211.3800 ;
        RECT 205.6600 216.3400 207.6600 216.8200 ;
        RECT 205.6600 221.7800 207.6600 222.2600 ;
        RECT 2.5600 227.2200 4.5600 227.7000 ;
        RECT 2.5600 232.6600 4.5600 233.1400 ;
        RECT 2.5600 238.1000 4.5600 238.5800 ;
        RECT 2.5600 243.5400 4.5600 244.0200 ;
        RECT 2.5600 248.9800 4.5600 249.4600 ;
        RECT 2.5600 254.4200 4.5600 254.9000 ;
        RECT 2.5600 259.8600 4.5600 260.3400 ;
        RECT 2.5600 265.3000 4.5600 265.7800 ;
        RECT 2.5600 270.7400 4.5600 271.2200 ;
        RECT 2.5600 276.1800 4.5600 276.6600 ;
        RECT 2.5600 308.8200 4.5600 309.3000 ;
        RECT 2.5600 281.6200 4.5600 282.1000 ;
        RECT 2.5600 287.0600 4.5600 287.5400 ;
        RECT 2.5600 292.5000 4.5600 292.9800 ;
        RECT 2.5600 297.9400 4.5600 298.4200 ;
        RECT 2.5600 303.3800 4.5600 303.8600 ;
        RECT 2.5600 314.2600 4.5600 314.7400 ;
        RECT 2.5600 319.7000 4.5600 320.1800 ;
        RECT 2.5600 325.1400 4.5600 325.6200 ;
        RECT 2.5600 330.5800 4.5600 331.0600 ;
        RECT 2.5600 336.0200 4.5600 336.5000 ;
        RECT 2.5600 341.4600 4.5600 341.9400 ;
        RECT 2.5600 346.9000 4.5600 347.3800 ;
        RECT 2.5600 352.3400 4.5600 352.8200 ;
        RECT 2.5600 357.7800 4.5600 358.2600 ;
        RECT 2.5600 363.2200 4.5600 363.7000 ;
        RECT 2.5600 368.6600 4.5600 369.1400 ;
        RECT 2.5600 374.1000 4.5600 374.5800 ;
        RECT 2.5600 379.5400 4.5600 380.0200 ;
        RECT 2.5600 384.9800 4.5600 385.4600 ;
        RECT 2.5600 390.4200 4.5600 390.9000 ;
        RECT 2.5600 395.8600 4.5600 396.3400 ;
        RECT 2.5600 401.3000 4.5600 401.7800 ;
        RECT 2.5600 406.7400 4.5600 407.2200 ;
        RECT 2.5600 412.1800 4.5600 412.6600 ;
        RECT 2.5600 417.6200 4.5600 418.1000 ;
        RECT 2.5600 423.0600 4.5600 423.5400 ;
        RECT 2.5600 428.5000 4.5600 428.9800 ;
        RECT 2.5600 433.9400 4.5600 434.4200 ;
        RECT 2.5600 439.3800 4.5600 439.8600 ;
        RECT 205.6600 227.2200 207.6600 227.7000 ;
        RECT 205.6600 232.6600 207.6600 233.1400 ;
        RECT 205.6600 238.1000 207.6600 238.5800 ;
        RECT 205.6600 243.5400 207.6600 244.0200 ;
        RECT 205.6600 248.9800 207.6600 249.4600 ;
        RECT 205.6600 254.4200 207.6600 254.9000 ;
        RECT 205.6600 259.8600 207.6600 260.3400 ;
        RECT 205.6600 265.3000 207.6600 265.7800 ;
        RECT 205.6600 270.7400 207.6600 271.2200 ;
        RECT 205.6600 276.1800 207.6600 276.6600 ;
        RECT 205.6600 308.8200 207.6600 309.3000 ;
        RECT 205.6600 281.6200 207.6600 282.1000 ;
        RECT 205.6600 287.0600 207.6600 287.5400 ;
        RECT 205.6600 292.5000 207.6600 292.9800 ;
        RECT 205.6600 297.9400 207.6600 298.4200 ;
        RECT 205.6600 303.3800 207.6600 303.8600 ;
        RECT 205.6600 314.2600 207.6600 314.7400 ;
        RECT 205.6600 319.7000 207.6600 320.1800 ;
        RECT 205.6600 325.1400 207.6600 325.6200 ;
        RECT 205.6600 330.5800 207.6600 331.0600 ;
        RECT 205.6600 336.0200 207.6600 336.5000 ;
        RECT 205.6600 341.4600 207.6600 341.9400 ;
        RECT 205.6600 346.9000 207.6600 347.3800 ;
        RECT 205.6600 352.3400 207.6600 352.8200 ;
        RECT 205.6600 357.7800 207.6600 358.2600 ;
        RECT 205.6600 363.2200 207.6600 363.7000 ;
        RECT 205.6600 368.6600 207.6600 369.1400 ;
        RECT 205.6600 374.1000 207.6600 374.5800 ;
        RECT 205.6600 379.5400 207.6600 380.0200 ;
        RECT 205.6600 384.9800 207.6600 385.4600 ;
        RECT 205.6600 390.4200 207.6600 390.9000 ;
        RECT 205.6600 395.8600 207.6600 396.3400 ;
        RECT 205.6600 401.3000 207.6600 401.7800 ;
        RECT 205.6600 406.7400 207.6600 407.2200 ;
        RECT 205.6600 412.1800 207.6600 412.6600 ;
        RECT 205.6600 417.6200 207.6600 418.1000 ;
        RECT 205.6600 423.0600 207.6600 423.5400 ;
        RECT 205.6600 428.5000 207.6600 428.9800 ;
        RECT 205.6600 433.9400 207.6600 434.4200 ;
        RECT 205.6600 439.3800 207.6600 439.8600 ;
      LAYER met4 ;
        RECT 193.3200 2.4300 194.9200 447.2200 ;
        RECT 148.3200 2.4300 149.9200 447.2200 ;
        RECT 103.3200 2.4300 104.9200 447.2200 ;
        RECT 58.3200 2.4300 59.9200 447.2200 ;
        RECT 13.3200 2.4300 14.9200 447.2200 ;
        RECT 205.6600 2.4300 207.6600 447.2200 ;
        RECT 2.5600 2.4300 4.5600 447.2200 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.6300 448.9300 210.2200 449.8200 ;
      RECT 148.7100 448.9300 148.9100 449.8200 ;
      RECT 147.3300 448.9300 147.9900 449.8200 ;
      RECT 145.9500 448.9300 146.6100 449.8200 ;
      RECT 144.5700 448.9300 145.2300 449.8200 ;
      RECT 143.1900 448.9300 143.8500 449.8200 ;
      RECT 141.8100 448.9300 142.4700 449.8200 ;
      RECT 140.4300 448.9300 141.0900 449.8200 ;
      RECT 139.0500 448.9300 139.7100 449.8200 ;
      RECT 137.6700 448.9300 138.3300 449.8200 ;
      RECT 136.2900 448.9300 136.9500 449.8200 ;
      RECT 134.9100 448.9300 135.5700 449.8200 ;
      RECT 133.5300 448.9300 134.1900 449.8200 ;
      RECT 132.1500 448.9300 132.8100 449.8200 ;
      RECT 130.7700 448.9300 131.4300 449.8200 ;
      RECT 129.3900 448.9300 130.0500 449.8200 ;
      RECT 128.0100 448.9300 128.6700 449.8200 ;
      RECT 126.6300 448.9300 127.2900 449.8200 ;
      RECT 125.7100 448.9300 125.9100 449.8200 ;
      RECT 124.3300 448.9300 124.9900 449.8200 ;
      RECT 122.9500 448.9300 123.6100 449.8200 ;
      RECT 121.5700 448.9300 122.2300 449.8200 ;
      RECT 120.1900 448.9300 120.8500 449.8200 ;
      RECT 118.8100 448.9300 119.4700 449.8200 ;
      RECT 117.4300 448.9300 118.0900 449.8200 ;
      RECT 116.0500 448.9300 116.7100 449.8200 ;
      RECT 114.6700 448.9300 115.3300 449.8200 ;
      RECT 113.2900 448.9300 113.9500 449.8200 ;
      RECT 111.9100 448.9300 112.5700 449.8200 ;
      RECT 110.5300 448.9300 111.1900 449.8200 ;
      RECT 109.1500 448.9300 109.8100 449.8200 ;
      RECT 107.7700 448.9300 108.4300 449.8200 ;
      RECT 106.3900 448.9300 107.0500 449.8200 ;
      RECT 105.0100 448.9300 105.6700 449.8200 ;
      RECT 103.6300 448.9300 104.2900 449.8200 ;
      RECT 102.7100 448.9300 102.9100 449.8200 ;
      RECT 101.3300 448.9300 101.9900 449.8200 ;
      RECT 99.9500 448.9300 100.6100 449.8200 ;
      RECT 98.5700 448.9300 99.2300 449.8200 ;
      RECT 97.1900 448.9300 97.8500 449.8200 ;
      RECT 95.8100 448.9300 96.4700 449.8200 ;
      RECT 94.4300 448.9300 95.0900 449.8200 ;
      RECT 93.0500 448.9300 93.7100 449.8200 ;
      RECT 91.6700 448.9300 92.3300 449.8200 ;
      RECT 90.2900 448.9300 90.9500 449.8200 ;
      RECT 88.9100 448.9300 89.5700 449.8200 ;
      RECT 87.5300 448.9300 88.1900 449.8200 ;
      RECT 86.1500 448.9300 86.8100 449.8200 ;
      RECT 84.7700 448.9300 85.4300 449.8200 ;
      RECT 83.3900 448.9300 84.0500 449.8200 ;
      RECT 82.0100 448.9300 82.6700 449.8200 ;
      RECT 80.6300 448.9300 81.2900 449.8200 ;
      RECT 79.7100 448.9300 79.9100 449.8200 ;
      RECT 78.3300 448.9300 78.9900 449.8200 ;
      RECT 76.9500 448.9300 77.6100 449.8200 ;
      RECT 75.5700 448.9300 76.2300 449.8200 ;
      RECT 74.1900 448.9300 74.8500 449.8200 ;
      RECT 72.8100 448.9300 73.4700 449.8200 ;
      RECT 71.4300 448.9300 72.0900 449.8200 ;
      RECT 70.0500 448.9300 70.7100 449.8200 ;
      RECT 68.6700 448.9300 69.3300 449.8200 ;
      RECT 67.2900 448.9300 67.9500 449.8200 ;
      RECT 65.9100 448.9300 66.5700 449.8200 ;
      RECT 64.5300 448.9300 65.1900 449.8200 ;
      RECT 63.1500 448.9300 63.8100 449.8200 ;
      RECT 61.7700 448.9300 62.4300 449.8200 ;
      RECT 60.3900 448.9300 61.0500 449.8200 ;
      RECT 59.0100 448.9300 59.6700 449.8200 ;
      RECT 57.6300 448.9300 58.2900 449.8200 ;
      RECT 56.7100 448.9300 56.9100 449.8200 ;
      RECT 55.3300 448.9300 55.9900 449.8200 ;
      RECT 53.9500 448.9300 54.6100 449.8200 ;
      RECT 52.5700 448.9300 53.2300 449.8200 ;
      RECT 51.1900 448.9300 51.8500 449.8200 ;
      RECT 49.8100 448.9300 50.4700 449.8200 ;
      RECT 48.4300 448.9300 49.0900 449.8200 ;
      RECT 47.0500 448.9300 47.7100 449.8200 ;
      RECT 45.6700 448.9300 46.3300 449.8200 ;
      RECT 44.2900 448.9300 44.9500 449.8200 ;
      RECT 42.9100 448.9300 43.5700 449.8200 ;
      RECT 41.5300 448.9300 42.1900 449.8200 ;
      RECT 40.1500 448.9300 40.8100 449.8200 ;
      RECT 38.7700 448.9300 39.4300 449.8200 ;
      RECT 37.3900 448.9300 38.0500 449.8200 ;
      RECT 36.0100 448.9300 36.6700 449.8200 ;
      RECT 34.6300 448.9300 35.2900 449.8200 ;
      RECT 33.7100 448.9300 33.9100 449.8200 ;
      RECT 32.3300 448.9300 32.9900 449.8200 ;
      RECT 30.9500 448.9300 31.6100 449.8200 ;
      RECT 29.5700 448.9300 30.2300 449.8200 ;
      RECT 28.1900 448.9300 28.8500 449.8200 ;
      RECT 26.8100 448.9300 27.4700 449.8200 ;
      RECT 25.4300 448.9300 26.0900 449.8200 ;
      RECT 24.0500 448.9300 24.7100 449.8200 ;
      RECT 22.6700 448.9300 23.3300 449.8200 ;
      RECT 21.2900 448.9300 21.9500 449.8200 ;
      RECT 19.9100 448.9300 20.5700 449.8200 ;
      RECT 18.5300 448.9300 19.1900 449.8200 ;
      RECT 17.1500 448.9300 17.8100 449.8200 ;
      RECT 15.7700 448.9300 16.4300 449.8200 ;
      RECT 14.3900 448.9300 15.0500 449.8200 ;
      RECT 13.0100 448.9300 13.6700 449.8200 ;
      RECT 11.6300 448.9300 12.2900 449.8200 ;
      RECT 10.7100 448.9300 10.9100 449.8200 ;
      RECT 0.0000 448.9300 9.9900 449.8200 ;
      RECT 0.0000 0.8900 210.2200 448.9300 ;
      RECT 149.6300 0.0000 210.2200 0.8900 ;
      RECT 148.7100 0.0000 148.9100 0.8900 ;
      RECT 147.3300 0.0000 147.9900 0.8900 ;
      RECT 145.9500 0.0000 146.6100 0.8900 ;
      RECT 144.5700 0.0000 145.2300 0.8900 ;
      RECT 143.1900 0.0000 143.8500 0.8900 ;
      RECT 141.8100 0.0000 142.4700 0.8900 ;
      RECT 140.4300 0.0000 141.0900 0.8900 ;
      RECT 139.0500 0.0000 139.7100 0.8900 ;
      RECT 137.6700 0.0000 138.3300 0.8900 ;
      RECT 136.2900 0.0000 136.9500 0.8900 ;
      RECT 134.9100 0.0000 135.5700 0.8900 ;
      RECT 133.5300 0.0000 134.1900 0.8900 ;
      RECT 132.1500 0.0000 132.8100 0.8900 ;
      RECT 130.7700 0.0000 131.4300 0.8900 ;
      RECT 129.3900 0.0000 130.0500 0.8900 ;
      RECT 128.0100 0.0000 128.6700 0.8900 ;
      RECT 126.6300 0.0000 127.2900 0.8900 ;
      RECT 125.7100 0.0000 125.9100 0.8900 ;
      RECT 124.3300 0.0000 124.9900 0.8900 ;
      RECT 122.9500 0.0000 123.6100 0.8900 ;
      RECT 121.5700 0.0000 122.2300 0.8900 ;
      RECT 120.1900 0.0000 120.8500 0.8900 ;
      RECT 118.8100 0.0000 119.4700 0.8900 ;
      RECT 117.4300 0.0000 118.0900 0.8900 ;
      RECT 116.0500 0.0000 116.7100 0.8900 ;
      RECT 114.6700 0.0000 115.3300 0.8900 ;
      RECT 113.2900 0.0000 113.9500 0.8900 ;
      RECT 111.9100 0.0000 112.5700 0.8900 ;
      RECT 110.5300 0.0000 111.1900 0.8900 ;
      RECT 109.1500 0.0000 109.8100 0.8900 ;
      RECT 107.7700 0.0000 108.4300 0.8900 ;
      RECT 106.3900 0.0000 107.0500 0.8900 ;
      RECT 105.0100 0.0000 105.6700 0.8900 ;
      RECT 103.6300 0.0000 104.2900 0.8900 ;
      RECT 102.7100 0.0000 102.9100 0.8900 ;
      RECT 101.3300 0.0000 101.9900 0.8900 ;
      RECT 99.9500 0.0000 100.6100 0.8900 ;
      RECT 98.5700 0.0000 99.2300 0.8900 ;
      RECT 97.1900 0.0000 97.8500 0.8900 ;
      RECT 95.8100 0.0000 96.4700 0.8900 ;
      RECT 94.4300 0.0000 95.0900 0.8900 ;
      RECT 93.0500 0.0000 93.7100 0.8900 ;
      RECT 91.6700 0.0000 92.3300 0.8900 ;
      RECT 90.2900 0.0000 90.9500 0.8900 ;
      RECT 88.9100 0.0000 89.5700 0.8900 ;
      RECT 87.5300 0.0000 88.1900 0.8900 ;
      RECT 86.1500 0.0000 86.8100 0.8900 ;
      RECT 84.7700 0.0000 85.4300 0.8900 ;
      RECT 83.3900 0.0000 84.0500 0.8900 ;
      RECT 82.0100 0.0000 82.6700 0.8900 ;
      RECT 80.6300 0.0000 81.2900 0.8900 ;
      RECT 79.7100 0.0000 79.9100 0.8900 ;
      RECT 78.3300 0.0000 78.9900 0.8900 ;
      RECT 76.9500 0.0000 77.6100 0.8900 ;
      RECT 75.5700 0.0000 76.2300 0.8900 ;
      RECT 74.1900 0.0000 74.8500 0.8900 ;
      RECT 72.8100 0.0000 73.4700 0.8900 ;
      RECT 71.4300 0.0000 72.0900 0.8900 ;
      RECT 70.0500 0.0000 70.7100 0.8900 ;
      RECT 68.6700 0.0000 69.3300 0.8900 ;
      RECT 67.2900 0.0000 67.9500 0.8900 ;
      RECT 65.9100 0.0000 66.5700 0.8900 ;
      RECT 64.5300 0.0000 65.1900 0.8900 ;
      RECT 63.1500 0.0000 63.8100 0.8900 ;
      RECT 61.7700 0.0000 62.4300 0.8900 ;
      RECT 60.3900 0.0000 61.0500 0.8900 ;
      RECT 59.0100 0.0000 59.6700 0.8900 ;
      RECT 57.6300 0.0000 58.2900 0.8900 ;
      RECT 56.7100 0.0000 56.9100 0.8900 ;
      RECT 55.3300 0.0000 55.9900 0.8900 ;
      RECT 53.9500 0.0000 54.6100 0.8900 ;
      RECT 52.5700 0.0000 53.2300 0.8900 ;
      RECT 51.1900 0.0000 51.8500 0.8900 ;
      RECT 49.8100 0.0000 50.4700 0.8900 ;
      RECT 48.4300 0.0000 49.0900 0.8900 ;
      RECT 47.0500 0.0000 47.7100 0.8900 ;
      RECT 45.6700 0.0000 46.3300 0.8900 ;
      RECT 44.2900 0.0000 44.9500 0.8900 ;
      RECT 42.9100 0.0000 43.5700 0.8900 ;
      RECT 41.5300 0.0000 42.1900 0.8900 ;
      RECT 40.1500 0.0000 40.8100 0.8900 ;
      RECT 38.7700 0.0000 39.4300 0.8900 ;
      RECT 37.3900 0.0000 38.0500 0.8900 ;
      RECT 36.0100 0.0000 36.6700 0.8900 ;
      RECT 34.6300 0.0000 35.2900 0.8900 ;
      RECT 33.7100 0.0000 33.9100 0.8900 ;
      RECT 32.3300 0.0000 32.9900 0.8900 ;
      RECT 30.9500 0.0000 31.6100 0.8900 ;
      RECT 29.5700 0.0000 30.2300 0.8900 ;
      RECT 28.1900 0.0000 28.8500 0.8900 ;
      RECT 26.8100 0.0000 27.4700 0.8900 ;
      RECT 25.4300 0.0000 26.0900 0.8900 ;
      RECT 24.0500 0.0000 24.7100 0.8900 ;
      RECT 22.6700 0.0000 23.3300 0.8900 ;
      RECT 21.2900 0.0000 21.9500 0.8900 ;
      RECT 19.9100 0.0000 20.5700 0.8900 ;
      RECT 18.5300 0.0000 19.1900 0.8900 ;
      RECT 17.1500 0.0000 17.8100 0.8900 ;
      RECT 15.7700 0.0000 16.4300 0.8900 ;
      RECT 14.3900 0.0000 15.0500 0.8900 ;
      RECT 13.0100 0.0000 13.6700 0.8900 ;
      RECT 11.6300 0.0000 12.2900 0.8900 ;
      RECT 10.7100 0.0000 10.9100 0.8900 ;
      RECT 0.0000 0.0000 9.9900 0.8900 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 210.2200 449.8200 ;
    LAYER met2 ;
      RECT 200.2000 448.9600 210.2200 449.8200 ;
      RECT 197.4400 448.9600 199.5400 449.8200 ;
      RECT 195.1400 448.9600 196.7800 449.8200 ;
      RECT 192.8400 448.9600 194.4800 449.8200 ;
      RECT 190.5400 448.9600 192.1800 449.8200 ;
      RECT 188.2400 448.9600 189.8800 449.8200 ;
      RECT 185.9400 448.9600 187.5800 449.8200 ;
      RECT 183.6400 448.9600 185.2800 449.8200 ;
      RECT 181.3400 448.9600 182.9800 449.8200 ;
      RECT 179.0400 448.9600 180.6800 449.8200 ;
      RECT 176.7400 448.9600 178.3800 449.8200 ;
      RECT 174.4400 448.9600 176.0800 449.8200 ;
      RECT 172.1400 448.9600 173.7800 449.8200 ;
      RECT 169.8400 448.9600 171.4800 449.8200 ;
      RECT 167.5400 448.9600 169.1800 449.8200 ;
      RECT 165.2400 448.9600 166.8800 449.8200 ;
      RECT 162.9400 448.9600 164.5800 449.8200 ;
      RECT 160.6400 448.9600 162.2800 449.8200 ;
      RECT 158.3400 448.9600 159.9800 449.8200 ;
      RECT 156.0400 448.9600 157.6800 449.8200 ;
      RECT 0.0000 448.9600 155.3800 449.8200 ;
      RECT 0.0000 439.7800 210.2200 448.9600 ;
      RECT 0.8600 439.1200 209.3600 439.7800 ;
      RECT 0.0000 438.0800 210.2200 439.1200 ;
      RECT 0.8600 437.4200 209.3600 438.0800 ;
      RECT 0.0000 436.3800 210.2200 437.4200 ;
      RECT 0.8600 435.7200 209.3600 436.3800 ;
      RECT 0.0000 434.6800 210.2200 435.7200 ;
      RECT 0.8600 434.0200 209.3600 434.6800 ;
      RECT 0.0000 432.9800 210.2200 434.0200 ;
      RECT 0.8600 432.3200 209.3600 432.9800 ;
      RECT 0.0000 431.2800 210.2200 432.3200 ;
      RECT 0.8600 430.6200 209.3600 431.2800 ;
      RECT 0.0000 429.2400 210.2200 430.6200 ;
      RECT 0.8600 428.5800 209.3600 429.2400 ;
      RECT 0.0000 427.5400 210.2200 428.5800 ;
      RECT 0.8600 426.8800 209.3600 427.5400 ;
      RECT 0.0000 425.8400 210.2200 426.8800 ;
      RECT 0.8600 425.1800 209.3600 425.8400 ;
      RECT 0.0000 424.1400 210.2200 425.1800 ;
      RECT 0.8600 423.4800 209.3600 424.1400 ;
      RECT 0.0000 422.4400 210.2200 423.4800 ;
      RECT 0.8600 421.7800 209.3600 422.4400 ;
      RECT 0.0000 420.4000 210.2200 421.7800 ;
      RECT 0.8600 419.7400 209.3600 420.4000 ;
      RECT 0.0000 418.7000 210.2200 419.7400 ;
      RECT 0.8600 418.0400 209.3600 418.7000 ;
      RECT 0.0000 417.0000 210.2200 418.0400 ;
      RECT 0.8600 416.3400 209.3600 417.0000 ;
      RECT 0.0000 415.3000 210.2200 416.3400 ;
      RECT 0.8600 414.6400 209.3600 415.3000 ;
      RECT 0.0000 413.6000 210.2200 414.6400 ;
      RECT 0.8600 412.9400 209.3600 413.6000 ;
      RECT 0.0000 411.5600 210.2200 412.9400 ;
      RECT 0.8600 410.9000 209.3600 411.5600 ;
      RECT 0.0000 409.8600 210.2200 410.9000 ;
      RECT 0.8600 409.2000 209.3600 409.8600 ;
      RECT 0.0000 408.1600 210.2200 409.2000 ;
      RECT 0.8600 407.5000 209.3600 408.1600 ;
      RECT 0.0000 406.4600 210.2200 407.5000 ;
      RECT 0.8600 405.8000 209.3600 406.4600 ;
      RECT 0.0000 404.7600 210.2200 405.8000 ;
      RECT 0.8600 404.1000 209.3600 404.7600 ;
      RECT 0.0000 402.7200 210.2200 404.1000 ;
      RECT 0.8600 402.0600 209.3600 402.7200 ;
      RECT 0.0000 401.0200 210.2200 402.0600 ;
      RECT 0.8600 400.3600 209.3600 401.0200 ;
      RECT 0.0000 399.3200 210.2200 400.3600 ;
      RECT 0.8600 398.6600 209.3600 399.3200 ;
      RECT 0.0000 397.6200 210.2200 398.6600 ;
      RECT 0.8600 396.9600 209.3600 397.6200 ;
      RECT 0.0000 395.9200 210.2200 396.9600 ;
      RECT 0.8600 395.2600 209.3600 395.9200 ;
      RECT 0.0000 393.8800 210.2200 395.2600 ;
      RECT 0.8600 393.2200 209.3600 393.8800 ;
      RECT 0.0000 392.1800 210.2200 393.2200 ;
      RECT 0.8600 391.5200 209.3600 392.1800 ;
      RECT 0.0000 390.4800 210.2200 391.5200 ;
      RECT 0.8600 389.8200 209.3600 390.4800 ;
      RECT 0.0000 388.7800 210.2200 389.8200 ;
      RECT 0.8600 388.1200 209.3600 388.7800 ;
      RECT 0.0000 387.0800 210.2200 388.1200 ;
      RECT 0.8600 386.4200 209.3600 387.0800 ;
      RECT 0.0000 385.3800 210.2200 386.4200 ;
      RECT 0.8600 384.7200 209.3600 385.3800 ;
      RECT 0.0000 380.2800 210.2200 384.7200 ;
      RECT 0.8600 379.6200 209.3600 380.2800 ;
      RECT 0.0000 378.5800 210.2200 379.6200 ;
      RECT 0.8600 377.9200 209.3600 378.5800 ;
      RECT 0.0000 377.2200 210.2200 377.9200 ;
      RECT 0.8600 376.5600 209.3600 377.2200 ;
      RECT 0.0000 375.8600 210.2200 376.5600 ;
      RECT 0.8600 375.2000 209.3600 375.8600 ;
      RECT 0.0000 374.1600 210.2200 375.2000 ;
      RECT 0.8600 373.5000 209.3600 374.1600 ;
      RECT 0.0000 372.8000 210.2200 373.5000 ;
      RECT 0.8600 372.1400 209.3600 372.8000 ;
      RECT 0.0000 371.4400 210.2200 372.1400 ;
      RECT 0.8600 370.7800 209.3600 371.4400 ;
      RECT 0.0000 369.7400 210.2200 370.7800 ;
      RECT 0.8600 369.0800 209.3600 369.7400 ;
      RECT 0.0000 368.3800 210.2200 369.0800 ;
      RECT 0.8600 367.7200 209.3600 368.3800 ;
      RECT 0.0000 367.0200 210.2200 367.7200 ;
      RECT 0.8600 366.3600 209.3600 367.0200 ;
      RECT 0.0000 365.3200 210.2200 366.3600 ;
      RECT 0.8600 364.6600 209.3600 365.3200 ;
      RECT 0.0000 363.9600 210.2200 364.6600 ;
      RECT 0.8600 363.3000 209.3600 363.9600 ;
      RECT 0.0000 362.6000 210.2200 363.3000 ;
      RECT 0.8600 361.9400 209.3600 362.6000 ;
      RECT 0.0000 360.9000 210.2200 361.9400 ;
      RECT 0.8600 360.2400 209.3600 360.9000 ;
      RECT 0.0000 359.5400 210.2200 360.2400 ;
      RECT 0.8600 358.8800 209.3600 359.5400 ;
      RECT 0.0000 358.1800 210.2200 358.8800 ;
      RECT 0.8600 357.5200 209.3600 358.1800 ;
      RECT 0.0000 356.4800 210.2200 357.5200 ;
      RECT 0.8600 355.8200 209.3600 356.4800 ;
      RECT 0.0000 355.1200 210.2200 355.8200 ;
      RECT 0.8600 354.4600 209.3600 355.1200 ;
      RECT 0.0000 353.7600 210.2200 354.4600 ;
      RECT 0.8600 353.1000 209.3600 353.7600 ;
      RECT 0.0000 352.0600 210.2200 353.1000 ;
      RECT 0.8600 351.4000 209.3600 352.0600 ;
      RECT 0.0000 350.7000 210.2200 351.4000 ;
      RECT 0.8600 350.0400 209.3600 350.7000 ;
      RECT 0.0000 349.3400 210.2200 350.0400 ;
      RECT 0.8600 348.6800 209.3600 349.3400 ;
      RECT 0.0000 347.6400 210.2200 348.6800 ;
      RECT 0.8600 346.9800 209.3600 347.6400 ;
      RECT 0.0000 346.2800 210.2200 346.9800 ;
      RECT 0.8600 345.6200 209.3600 346.2800 ;
      RECT 0.0000 344.9200 210.2200 345.6200 ;
      RECT 0.8600 344.2600 209.3600 344.9200 ;
      RECT 0.0000 343.2200 210.2200 344.2600 ;
      RECT 0.8600 342.5600 209.3600 343.2200 ;
      RECT 0.0000 341.8600 210.2200 342.5600 ;
      RECT 0.8600 341.2000 209.3600 341.8600 ;
      RECT 0.0000 340.5000 210.2200 341.2000 ;
      RECT 0.8600 339.8400 209.3600 340.5000 ;
      RECT 0.0000 338.8000 210.2200 339.8400 ;
      RECT 0.8600 338.1400 209.3600 338.8000 ;
      RECT 0.0000 337.4400 210.2200 338.1400 ;
      RECT 0.8600 336.7800 209.3600 337.4400 ;
      RECT 0.0000 336.0800 210.2200 336.7800 ;
      RECT 0.8600 335.4200 209.3600 336.0800 ;
      RECT 0.0000 334.3800 210.2200 335.4200 ;
      RECT 0.8600 333.7200 209.3600 334.3800 ;
      RECT 0.0000 333.0200 210.2200 333.7200 ;
      RECT 0.8600 332.3600 209.3600 333.0200 ;
      RECT 0.0000 331.6600 210.2200 332.3600 ;
      RECT 0.8600 331.0000 209.3600 331.6600 ;
      RECT 0.0000 329.9600 210.2200 331.0000 ;
      RECT 0.8600 329.3000 209.3600 329.9600 ;
      RECT 0.0000 328.6000 210.2200 329.3000 ;
      RECT 0.8600 327.9400 209.3600 328.6000 ;
      RECT 0.0000 327.2400 210.2200 327.9400 ;
      RECT 0.8600 326.5800 209.3600 327.2400 ;
      RECT 0.0000 325.5400 210.2200 326.5800 ;
      RECT 0.8600 324.8800 209.3600 325.5400 ;
      RECT 0.0000 324.1800 210.2200 324.8800 ;
      RECT 0.8600 323.5200 209.3600 324.1800 ;
      RECT 0.0000 322.8200 210.2200 323.5200 ;
      RECT 0.8600 322.1600 209.3600 322.8200 ;
      RECT 0.0000 321.1200 210.2200 322.1600 ;
      RECT 0.8600 320.4600 209.3600 321.1200 ;
      RECT 0.0000 319.7600 210.2200 320.4600 ;
      RECT 0.8600 319.1000 209.3600 319.7600 ;
      RECT 0.0000 318.4000 210.2200 319.1000 ;
      RECT 0.8600 317.7400 209.3600 318.4000 ;
      RECT 0.0000 316.7000 210.2200 317.7400 ;
      RECT 0.8600 316.0400 209.3600 316.7000 ;
      RECT 0.0000 315.3400 210.2200 316.0400 ;
      RECT 0.8600 314.6800 209.3600 315.3400 ;
      RECT 0.0000 313.9800 210.2200 314.6800 ;
      RECT 0.8600 313.3200 209.3600 313.9800 ;
      RECT 0.0000 312.2800 210.2200 313.3200 ;
      RECT 0.8600 311.6200 209.3600 312.2800 ;
      RECT 0.0000 310.9200 210.2200 311.6200 ;
      RECT 0.8600 310.2600 209.3600 310.9200 ;
      RECT 0.0000 309.5600 210.2200 310.2600 ;
      RECT 0.8600 308.9000 209.3600 309.5600 ;
      RECT 0.0000 308.2000 210.2200 308.9000 ;
      RECT 0.8600 307.5400 209.3600 308.2000 ;
      RECT 0.0000 306.5000 210.2200 307.5400 ;
      RECT 0.8600 305.8400 209.3600 306.5000 ;
      RECT 0.0000 305.1400 210.2200 305.8400 ;
      RECT 0.8600 304.4800 209.3600 305.1400 ;
      RECT 0.0000 303.7800 210.2200 304.4800 ;
      RECT 0.8600 303.1200 209.3600 303.7800 ;
      RECT 0.0000 302.0800 210.2200 303.1200 ;
      RECT 0.8600 301.4200 209.3600 302.0800 ;
      RECT 0.0000 300.7200 210.2200 301.4200 ;
      RECT 0.8600 300.0600 209.3600 300.7200 ;
      RECT 0.0000 299.3600 210.2200 300.0600 ;
      RECT 0.8600 298.7000 209.3600 299.3600 ;
      RECT 0.0000 297.6600 210.2200 298.7000 ;
      RECT 0.8600 297.0000 209.3600 297.6600 ;
      RECT 0.0000 296.3000 210.2200 297.0000 ;
      RECT 0.8600 295.6400 209.3600 296.3000 ;
      RECT 0.0000 294.9400 210.2200 295.6400 ;
      RECT 0.8600 294.2800 209.3600 294.9400 ;
      RECT 0.0000 293.2400 210.2200 294.2800 ;
      RECT 0.8600 292.5800 209.3600 293.2400 ;
      RECT 0.0000 291.8800 210.2200 292.5800 ;
      RECT 0.8600 291.2200 209.3600 291.8800 ;
      RECT 0.0000 290.5200 210.2200 291.2200 ;
      RECT 0.8600 289.8600 209.3600 290.5200 ;
      RECT 0.0000 288.8200 210.2200 289.8600 ;
      RECT 0.8600 288.1600 209.3600 288.8200 ;
      RECT 0.0000 287.4600 210.2200 288.1600 ;
      RECT 0.8600 286.8000 209.3600 287.4600 ;
      RECT 0.0000 286.1000 210.2200 286.8000 ;
      RECT 0.8600 285.4400 209.3600 286.1000 ;
      RECT 0.0000 284.4000 210.2200 285.4400 ;
      RECT 0.8600 283.7400 209.3600 284.4000 ;
      RECT 0.0000 283.0400 210.2200 283.7400 ;
      RECT 0.8600 282.3800 209.3600 283.0400 ;
      RECT 0.0000 281.6800 210.2200 282.3800 ;
      RECT 0.8600 281.0200 209.3600 281.6800 ;
      RECT 0.0000 279.9800 210.2200 281.0200 ;
      RECT 0.8600 279.3200 209.3600 279.9800 ;
      RECT 0.0000 278.6200 210.2200 279.3200 ;
      RECT 0.8600 277.9600 209.3600 278.6200 ;
      RECT 0.0000 277.2600 210.2200 277.9600 ;
      RECT 0.8600 276.6000 209.3600 277.2600 ;
      RECT 0.0000 275.5600 210.2200 276.6000 ;
      RECT 0.8600 274.9000 209.3600 275.5600 ;
      RECT 0.0000 274.2000 210.2200 274.9000 ;
      RECT 0.8600 273.5400 209.3600 274.2000 ;
      RECT 0.0000 272.8400 210.2200 273.5400 ;
      RECT 0.8600 272.1800 209.3600 272.8400 ;
      RECT 0.0000 271.1400 210.2200 272.1800 ;
      RECT 0.8600 270.4800 209.3600 271.1400 ;
      RECT 0.0000 269.7800 210.2200 270.4800 ;
      RECT 0.8600 269.1200 209.3600 269.7800 ;
      RECT 0.0000 268.4200 210.2200 269.1200 ;
      RECT 0.8600 267.7600 209.3600 268.4200 ;
      RECT 0.0000 266.7200 210.2200 267.7600 ;
      RECT 0.8600 266.0600 209.3600 266.7200 ;
      RECT 0.0000 265.3600 210.2200 266.0600 ;
      RECT 0.8600 264.7000 209.3600 265.3600 ;
      RECT 0.0000 264.0000 210.2200 264.7000 ;
      RECT 0.8600 263.3400 209.3600 264.0000 ;
      RECT 0.0000 262.3000 210.2200 263.3400 ;
      RECT 0.8600 261.6400 209.3600 262.3000 ;
      RECT 0.0000 260.9400 210.2200 261.6400 ;
      RECT 0.8600 260.2800 209.3600 260.9400 ;
      RECT 0.0000 259.5800 210.2200 260.2800 ;
      RECT 0.8600 258.9200 209.3600 259.5800 ;
      RECT 0.0000 257.8800 210.2200 258.9200 ;
      RECT 0.8600 257.2200 209.3600 257.8800 ;
      RECT 0.0000 256.5200 210.2200 257.2200 ;
      RECT 0.8600 255.8600 209.3600 256.5200 ;
      RECT 0.0000 255.1600 210.2200 255.8600 ;
      RECT 0.8600 254.5000 209.3600 255.1600 ;
      RECT 0.0000 253.4600 210.2200 254.5000 ;
      RECT 0.8600 252.8000 209.3600 253.4600 ;
      RECT 0.0000 252.1000 210.2200 252.8000 ;
      RECT 0.8600 251.4400 209.3600 252.1000 ;
      RECT 0.0000 250.7400 210.2200 251.4400 ;
      RECT 0.8600 250.0800 209.3600 250.7400 ;
      RECT 0.0000 249.0400 210.2200 250.0800 ;
      RECT 0.8600 248.3800 209.3600 249.0400 ;
      RECT 0.0000 247.6800 210.2200 248.3800 ;
      RECT 0.8600 247.0200 209.3600 247.6800 ;
      RECT 0.0000 246.3200 210.2200 247.0200 ;
      RECT 0.8600 245.6600 209.3600 246.3200 ;
      RECT 0.0000 244.6200 210.2200 245.6600 ;
      RECT 0.8600 243.9600 209.3600 244.6200 ;
      RECT 0.0000 243.2600 210.2200 243.9600 ;
      RECT 0.8600 242.6000 209.3600 243.2600 ;
      RECT 0.0000 241.9000 210.2200 242.6000 ;
      RECT 0.8600 241.2400 209.3600 241.9000 ;
      RECT 0.0000 240.5400 210.2200 241.2400 ;
      RECT 0.8600 239.8800 209.3600 240.5400 ;
      RECT 0.0000 209.9400 210.2200 239.8800 ;
      RECT 0.8600 209.2800 209.3600 209.9400 ;
      RECT 0.0000 208.2400 210.2200 209.2800 ;
      RECT 0.8600 207.5800 209.3600 208.2400 ;
      RECT 0.0000 206.5400 210.2200 207.5800 ;
      RECT 0.8600 205.8800 209.3600 206.5400 ;
      RECT 0.0000 204.8400 210.2200 205.8800 ;
      RECT 0.8600 204.1800 209.3600 204.8400 ;
      RECT 0.0000 203.1400 210.2200 204.1800 ;
      RECT 0.8600 202.4800 209.3600 203.1400 ;
      RECT 0.0000 201.4400 210.2200 202.4800 ;
      RECT 0.8600 200.7800 209.3600 201.4400 ;
      RECT 0.0000 199.4000 210.2200 200.7800 ;
      RECT 0.8600 198.7400 209.3600 199.4000 ;
      RECT 0.0000 197.7000 210.2200 198.7400 ;
      RECT 0.8600 197.0400 209.3600 197.7000 ;
      RECT 0.0000 196.0000 210.2200 197.0400 ;
      RECT 0.8600 195.3400 209.3600 196.0000 ;
      RECT 0.0000 194.3000 210.2200 195.3400 ;
      RECT 0.8600 193.6400 209.3600 194.3000 ;
      RECT 0.0000 192.6000 210.2200 193.6400 ;
      RECT 0.8600 191.9400 209.3600 192.6000 ;
      RECT 0.0000 190.5600 210.2200 191.9400 ;
      RECT 0.8600 189.9000 209.3600 190.5600 ;
      RECT 0.0000 188.8600 210.2200 189.9000 ;
      RECT 0.8600 188.2000 209.3600 188.8600 ;
      RECT 0.0000 187.1600 210.2200 188.2000 ;
      RECT 0.8600 186.5000 209.3600 187.1600 ;
      RECT 0.0000 185.4600 210.2200 186.5000 ;
      RECT 0.8600 184.8000 209.3600 185.4600 ;
      RECT 0.0000 183.7600 210.2200 184.8000 ;
      RECT 0.8600 183.1000 209.3600 183.7600 ;
      RECT 0.0000 181.7200 210.2200 183.1000 ;
      RECT 0.8600 181.0600 209.3600 181.7200 ;
      RECT 0.0000 180.0200 210.2200 181.0600 ;
      RECT 0.8600 179.3600 209.3600 180.0200 ;
      RECT 0.0000 178.3200 210.2200 179.3600 ;
      RECT 0.8600 177.6600 209.3600 178.3200 ;
      RECT 0.0000 176.6200 210.2200 177.6600 ;
      RECT 0.8600 175.9600 209.3600 176.6200 ;
      RECT 0.0000 174.9200 210.2200 175.9600 ;
      RECT 0.8600 174.2600 209.3600 174.9200 ;
      RECT 0.0000 172.8800 210.2200 174.2600 ;
      RECT 0.8600 172.2200 209.3600 172.8800 ;
      RECT 0.0000 171.1800 210.2200 172.2200 ;
      RECT 0.8600 170.5200 209.3600 171.1800 ;
      RECT 0.0000 169.4800 210.2200 170.5200 ;
      RECT 0.8600 168.8200 209.3600 169.4800 ;
      RECT 0.0000 167.7800 210.2200 168.8200 ;
      RECT 0.8600 167.1200 209.3600 167.7800 ;
      RECT 0.0000 166.0800 210.2200 167.1200 ;
      RECT 0.8600 165.4200 209.3600 166.0800 ;
      RECT 0.0000 164.0400 210.2200 165.4200 ;
      RECT 0.8600 163.3800 209.3600 164.0400 ;
      RECT 0.0000 162.3400 210.2200 163.3800 ;
      RECT 0.8600 161.6800 209.3600 162.3400 ;
      RECT 0.0000 160.6400 210.2200 161.6800 ;
      RECT 0.8600 159.9800 209.3600 160.6400 ;
      RECT 0.0000 158.9400 210.2200 159.9800 ;
      RECT 0.8600 158.2800 209.3600 158.9400 ;
      RECT 0.0000 157.2400 210.2200 158.2800 ;
      RECT 0.8600 156.5800 209.3600 157.2400 ;
      RECT 0.0000 155.5400 210.2200 156.5800 ;
      RECT 0.8600 154.8800 209.3600 155.5400 ;
      RECT 0.0000 150.1000 210.2200 154.8800 ;
      RECT 0.8600 149.4400 209.3600 150.1000 ;
      RECT 0.0000 148.4000 210.2200 149.4400 ;
      RECT 0.8600 147.7400 209.3600 148.4000 ;
      RECT 0.0000 147.0400 210.2200 147.7400 ;
      RECT 0.8600 146.3800 209.3600 147.0400 ;
      RECT 0.0000 145.6800 210.2200 146.3800 ;
      RECT 0.8600 145.0200 209.3600 145.6800 ;
      RECT 0.0000 143.9800 210.2200 145.0200 ;
      RECT 0.8600 143.3200 209.3600 143.9800 ;
      RECT 0.0000 142.6200 210.2200 143.3200 ;
      RECT 0.8600 141.9600 209.3600 142.6200 ;
      RECT 0.0000 141.2600 210.2200 141.9600 ;
      RECT 0.8600 140.6000 209.3600 141.2600 ;
      RECT 0.0000 139.5600 210.2200 140.6000 ;
      RECT 0.8600 138.9000 209.3600 139.5600 ;
      RECT 0.0000 138.2000 210.2200 138.9000 ;
      RECT 0.8600 137.5400 209.3600 138.2000 ;
      RECT 0.0000 136.8400 210.2200 137.5400 ;
      RECT 0.8600 136.1800 209.3600 136.8400 ;
      RECT 0.0000 135.1400 210.2200 136.1800 ;
      RECT 0.8600 134.4800 209.3600 135.1400 ;
      RECT 0.0000 133.7800 210.2200 134.4800 ;
      RECT 0.8600 133.1200 209.3600 133.7800 ;
      RECT 0.0000 132.4200 210.2200 133.1200 ;
      RECT 0.8600 131.7600 209.3600 132.4200 ;
      RECT 0.0000 130.7200 210.2200 131.7600 ;
      RECT 0.8600 130.0600 209.3600 130.7200 ;
      RECT 0.0000 129.3600 210.2200 130.0600 ;
      RECT 0.8600 128.7000 209.3600 129.3600 ;
      RECT 0.0000 128.0000 210.2200 128.7000 ;
      RECT 0.8600 127.3400 209.3600 128.0000 ;
      RECT 0.0000 126.3000 210.2200 127.3400 ;
      RECT 0.8600 125.6400 209.3600 126.3000 ;
      RECT 0.0000 124.9400 210.2200 125.6400 ;
      RECT 0.8600 124.2800 209.3600 124.9400 ;
      RECT 0.0000 123.5800 210.2200 124.2800 ;
      RECT 0.8600 122.9200 209.3600 123.5800 ;
      RECT 0.0000 121.8800 210.2200 122.9200 ;
      RECT 0.8600 121.2200 209.3600 121.8800 ;
      RECT 0.0000 120.5200 210.2200 121.2200 ;
      RECT 0.8600 119.8600 209.3600 120.5200 ;
      RECT 0.0000 119.1600 210.2200 119.8600 ;
      RECT 0.8600 118.5000 209.3600 119.1600 ;
      RECT 0.0000 117.4600 210.2200 118.5000 ;
      RECT 0.8600 116.8000 209.3600 117.4600 ;
      RECT 0.0000 116.1000 210.2200 116.8000 ;
      RECT 0.8600 115.4400 209.3600 116.1000 ;
      RECT 0.0000 114.7400 210.2200 115.4400 ;
      RECT 0.8600 114.0800 209.3600 114.7400 ;
      RECT 0.0000 113.0400 210.2200 114.0800 ;
      RECT 0.8600 112.3800 209.3600 113.0400 ;
      RECT 0.0000 111.6800 210.2200 112.3800 ;
      RECT 0.8600 111.0200 209.3600 111.6800 ;
      RECT 0.0000 110.3200 210.2200 111.0200 ;
      RECT 0.8600 109.6600 209.3600 110.3200 ;
      RECT 0.0000 108.6200 210.2200 109.6600 ;
      RECT 0.8600 107.9600 209.3600 108.6200 ;
      RECT 0.0000 107.2600 210.2200 107.9600 ;
      RECT 0.8600 106.6000 209.3600 107.2600 ;
      RECT 0.0000 105.9000 210.2200 106.6000 ;
      RECT 0.8600 105.2400 209.3600 105.9000 ;
      RECT 0.0000 104.2000 210.2200 105.2400 ;
      RECT 0.8600 103.5400 209.3600 104.2000 ;
      RECT 0.0000 102.8400 210.2200 103.5400 ;
      RECT 0.8600 102.1800 209.3600 102.8400 ;
      RECT 0.0000 101.4800 210.2200 102.1800 ;
      RECT 0.8600 100.8200 209.3600 101.4800 ;
      RECT 0.0000 99.7800 210.2200 100.8200 ;
      RECT 0.8600 99.1200 209.3600 99.7800 ;
      RECT 0.0000 98.4200 210.2200 99.1200 ;
      RECT 0.8600 97.7600 209.3600 98.4200 ;
      RECT 0.0000 97.0600 210.2200 97.7600 ;
      RECT 0.8600 96.4000 209.3600 97.0600 ;
      RECT 0.0000 95.3600 210.2200 96.4000 ;
      RECT 0.8600 94.7000 209.3600 95.3600 ;
      RECT 0.0000 94.0000 210.2200 94.7000 ;
      RECT 0.8600 93.3400 209.3600 94.0000 ;
      RECT 0.0000 92.6400 210.2200 93.3400 ;
      RECT 0.8600 91.9800 209.3600 92.6400 ;
      RECT 0.0000 90.9400 210.2200 91.9800 ;
      RECT 0.8600 90.2800 209.3600 90.9400 ;
      RECT 0.0000 89.5800 210.2200 90.2800 ;
      RECT 0.8600 88.9200 209.3600 89.5800 ;
      RECT 0.0000 88.2200 210.2200 88.9200 ;
      RECT 0.8600 87.5600 209.3600 88.2200 ;
      RECT 0.0000 86.5200 210.2200 87.5600 ;
      RECT 0.8600 85.8600 209.3600 86.5200 ;
      RECT 0.0000 85.1600 210.2200 85.8600 ;
      RECT 0.8600 84.5000 209.3600 85.1600 ;
      RECT 0.0000 83.8000 210.2200 84.5000 ;
      RECT 0.8600 83.1400 209.3600 83.8000 ;
      RECT 0.0000 82.1000 210.2200 83.1400 ;
      RECT 0.8600 81.4400 209.3600 82.1000 ;
      RECT 0.0000 80.7400 210.2200 81.4400 ;
      RECT 0.8600 80.0800 209.3600 80.7400 ;
      RECT 0.0000 79.3800 210.2200 80.0800 ;
      RECT 0.8600 78.7200 209.3600 79.3800 ;
      RECT 0.0000 78.0200 210.2200 78.7200 ;
      RECT 0.8600 77.3600 209.3600 78.0200 ;
      RECT 0.0000 76.3200 210.2200 77.3600 ;
      RECT 0.8600 75.6600 209.3600 76.3200 ;
      RECT 0.0000 74.9600 210.2200 75.6600 ;
      RECT 0.8600 74.3000 209.3600 74.9600 ;
      RECT 0.0000 73.6000 210.2200 74.3000 ;
      RECT 0.8600 72.9400 209.3600 73.6000 ;
      RECT 0.0000 71.9000 210.2200 72.9400 ;
      RECT 0.8600 71.2400 209.3600 71.9000 ;
      RECT 0.0000 70.5400 210.2200 71.2400 ;
      RECT 0.8600 69.8800 209.3600 70.5400 ;
      RECT 0.0000 69.1800 210.2200 69.8800 ;
      RECT 0.8600 68.5200 209.3600 69.1800 ;
      RECT 0.0000 67.4800 210.2200 68.5200 ;
      RECT 0.8600 66.8200 209.3600 67.4800 ;
      RECT 0.0000 66.1200 210.2200 66.8200 ;
      RECT 0.8600 65.4600 209.3600 66.1200 ;
      RECT 0.0000 64.7600 210.2200 65.4600 ;
      RECT 0.8600 64.1000 209.3600 64.7600 ;
      RECT 0.0000 63.0600 210.2200 64.1000 ;
      RECT 0.8600 62.4000 209.3600 63.0600 ;
      RECT 0.0000 61.7000 210.2200 62.4000 ;
      RECT 0.8600 61.0400 209.3600 61.7000 ;
      RECT 0.0000 60.3400 210.2200 61.0400 ;
      RECT 0.8600 59.6800 209.3600 60.3400 ;
      RECT 0.0000 58.6400 210.2200 59.6800 ;
      RECT 0.8600 57.9800 209.3600 58.6400 ;
      RECT 0.0000 57.2800 210.2200 57.9800 ;
      RECT 0.8600 56.6200 209.3600 57.2800 ;
      RECT 0.0000 55.9200 210.2200 56.6200 ;
      RECT 0.8600 55.2600 209.3600 55.9200 ;
      RECT 0.0000 54.2200 210.2200 55.2600 ;
      RECT 0.8600 53.5600 209.3600 54.2200 ;
      RECT 0.0000 52.8600 210.2200 53.5600 ;
      RECT 0.8600 52.2000 209.3600 52.8600 ;
      RECT 0.0000 51.5000 210.2200 52.2000 ;
      RECT 0.8600 50.8400 209.3600 51.5000 ;
      RECT 0.0000 49.8000 210.2200 50.8400 ;
      RECT 0.8600 49.1400 209.3600 49.8000 ;
      RECT 0.0000 48.4400 210.2200 49.1400 ;
      RECT 0.8600 47.7800 209.3600 48.4400 ;
      RECT 0.0000 47.0800 210.2200 47.7800 ;
      RECT 0.8600 46.4200 209.3600 47.0800 ;
      RECT 0.0000 45.3800 210.2200 46.4200 ;
      RECT 0.8600 44.7200 209.3600 45.3800 ;
      RECT 0.0000 44.0200 210.2200 44.7200 ;
      RECT 0.8600 43.3600 209.3600 44.0200 ;
      RECT 0.0000 42.6600 210.2200 43.3600 ;
      RECT 0.8600 42.0000 209.3600 42.6600 ;
      RECT 0.0000 40.9600 210.2200 42.0000 ;
      RECT 0.8600 40.3000 209.3600 40.9600 ;
      RECT 0.0000 39.6000 210.2200 40.3000 ;
      RECT 0.8600 38.9400 209.3600 39.6000 ;
      RECT 0.0000 38.2400 210.2200 38.9400 ;
      RECT 0.8600 37.5800 209.3600 38.2400 ;
      RECT 0.0000 36.5400 210.2200 37.5800 ;
      RECT 0.8600 35.8800 209.3600 36.5400 ;
      RECT 0.0000 35.1800 210.2200 35.8800 ;
      RECT 0.8600 34.5200 209.3600 35.1800 ;
      RECT 0.0000 33.8200 210.2200 34.5200 ;
      RECT 0.8600 33.1600 209.3600 33.8200 ;
      RECT 0.0000 32.1200 210.2200 33.1600 ;
      RECT 0.8600 31.4600 209.3600 32.1200 ;
      RECT 0.0000 30.7600 210.2200 31.4600 ;
      RECT 0.8600 30.1000 209.3600 30.7600 ;
      RECT 0.0000 29.4000 210.2200 30.1000 ;
      RECT 0.8600 28.7400 209.3600 29.4000 ;
      RECT 0.0000 27.7000 210.2200 28.7400 ;
      RECT 0.8600 27.0400 209.3600 27.7000 ;
      RECT 0.0000 26.3400 210.2200 27.0400 ;
      RECT 0.8600 25.6800 209.3600 26.3400 ;
      RECT 0.0000 24.9800 210.2200 25.6800 ;
      RECT 0.8600 24.3200 209.3600 24.9800 ;
      RECT 0.0000 23.2800 210.2200 24.3200 ;
      RECT 0.8600 22.6200 209.3600 23.2800 ;
      RECT 0.0000 21.9200 210.2200 22.6200 ;
      RECT 0.8600 21.2600 209.3600 21.9200 ;
      RECT 0.0000 20.5600 210.2200 21.2600 ;
      RECT 0.8600 19.9000 209.3600 20.5600 ;
      RECT 0.0000 18.8600 210.2200 19.9000 ;
      RECT 0.8600 18.2000 209.3600 18.8600 ;
      RECT 0.0000 17.5000 210.2200 18.2000 ;
      RECT 0.8600 16.8400 209.3600 17.5000 ;
      RECT 0.0000 16.1400 210.2200 16.8400 ;
      RECT 0.8600 15.4800 209.3600 16.1400 ;
      RECT 0.0000 14.4400 210.2200 15.4800 ;
      RECT 0.8600 13.7800 209.3600 14.4400 ;
      RECT 0.0000 13.0800 210.2200 13.7800 ;
      RECT 0.8600 12.4200 209.3600 13.0800 ;
      RECT 0.0000 11.7200 210.2200 12.4200 ;
      RECT 0.8600 11.0600 209.3600 11.7200 ;
      RECT 0.0000 10.3600 210.2200 11.0600 ;
      RECT 0.8600 9.7000 209.3600 10.3600 ;
      RECT 0.0000 0.8600 210.2200 9.7000 ;
      RECT 200.2000 0.0000 210.2200 0.8600 ;
      RECT 197.4400 0.0000 199.5400 0.8600 ;
      RECT 195.1400 0.0000 196.7800 0.8600 ;
      RECT 192.8400 0.0000 194.4800 0.8600 ;
      RECT 190.5400 0.0000 192.1800 0.8600 ;
      RECT 187.7800 0.0000 189.8800 0.8600 ;
      RECT 185.9400 0.0000 187.1200 0.8600 ;
      RECT 183.6400 0.0000 185.2800 0.8600 ;
      RECT 180.8800 0.0000 182.9800 0.8600 ;
      RECT 179.0400 0.0000 180.2200 0.8600 ;
      RECT 176.2800 0.0000 178.3800 0.8600 ;
      RECT 174.4400 0.0000 175.6200 0.8600 ;
      RECT 172.1400 0.0000 173.7800 0.8600 ;
      RECT 169.8400 0.0000 171.4800 0.8600 ;
      RECT 167.5400 0.0000 169.1800 0.8600 ;
      RECT 164.7800 0.0000 166.8800 0.8600 ;
      RECT 162.9400 0.0000 164.1200 0.8600 ;
      RECT 160.6400 0.0000 162.2800 0.8600 ;
      RECT 157.8800 0.0000 159.9800 0.8600 ;
      RECT 156.0400 0.0000 157.2200 0.8600 ;
      RECT 0.0000 0.0000 155.3800 0.8600 ;
    LAYER met3 ;
      RECT 0.0000 447.5200 210.2200 449.8200 ;
      RECT 207.9600 444.9200 210.2200 447.5200 ;
      RECT 0.0000 444.9200 2.2600 447.5200 ;
      RECT 0.0000 444.5200 210.2200 444.9200 ;
      RECT 204.9600 441.9200 210.2200 444.5200 ;
      RECT 0.0000 441.9200 5.2600 444.5200 ;
      RECT 0.0000 440.1600 210.2200 441.9200 ;
      RECT 207.9600 439.0800 210.2200 440.1600 ;
      RECT 4.8600 439.0800 205.3600 440.1600 ;
      RECT 0.0000 439.0800 2.2600 440.1600 ;
      RECT 0.0000 437.4400 210.2200 439.0800 ;
      RECT 204.9600 436.3600 210.2200 437.4400 ;
      RECT 7.8600 436.3600 202.3600 437.4400 ;
      RECT 0.0000 436.3600 5.2600 437.4400 ;
      RECT 0.0000 434.7200 210.2200 436.3600 ;
      RECT 207.9600 433.6400 210.2200 434.7200 ;
      RECT 4.8600 433.6400 205.3600 434.7200 ;
      RECT 0.0000 433.6400 2.2600 434.7200 ;
      RECT 0.0000 432.0000 210.2200 433.6400 ;
      RECT 204.9600 430.9200 210.2200 432.0000 ;
      RECT 7.8600 430.9200 202.3600 432.0000 ;
      RECT 0.0000 430.9200 5.2600 432.0000 ;
      RECT 0.0000 429.2800 210.2200 430.9200 ;
      RECT 207.9600 428.2000 210.2200 429.2800 ;
      RECT 4.8600 428.2000 205.3600 429.2800 ;
      RECT 0.0000 428.2000 2.2600 429.2800 ;
      RECT 0.0000 426.5600 210.2200 428.2000 ;
      RECT 204.9600 425.4800 210.2200 426.5600 ;
      RECT 7.8600 425.4800 202.3600 426.5600 ;
      RECT 0.0000 425.4800 5.2600 426.5600 ;
      RECT 0.0000 423.8400 210.2200 425.4800 ;
      RECT 207.9600 422.7600 210.2200 423.8400 ;
      RECT 4.8600 422.7600 205.3600 423.8400 ;
      RECT 0.0000 422.7600 2.2600 423.8400 ;
      RECT 0.0000 421.1200 210.2200 422.7600 ;
      RECT 204.9600 420.0400 210.2200 421.1200 ;
      RECT 7.8600 420.0400 202.3600 421.1200 ;
      RECT 0.0000 420.0400 5.2600 421.1200 ;
      RECT 0.0000 418.4000 210.2200 420.0400 ;
      RECT 207.9600 417.3200 210.2200 418.4000 ;
      RECT 4.8600 417.3200 205.3600 418.4000 ;
      RECT 0.0000 417.3200 2.2600 418.4000 ;
      RECT 0.0000 415.6800 210.2200 417.3200 ;
      RECT 204.9600 414.6000 210.2200 415.6800 ;
      RECT 7.8600 414.6000 202.3600 415.6800 ;
      RECT 0.0000 414.6000 5.2600 415.6800 ;
      RECT 0.0000 412.9600 210.2200 414.6000 ;
      RECT 207.9600 411.8800 210.2200 412.9600 ;
      RECT 4.8600 411.8800 205.3600 412.9600 ;
      RECT 0.0000 411.8800 2.2600 412.9600 ;
      RECT 0.0000 410.2400 210.2200 411.8800 ;
      RECT 204.9600 409.1600 210.2200 410.2400 ;
      RECT 7.8600 409.1600 202.3600 410.2400 ;
      RECT 0.0000 409.1600 5.2600 410.2400 ;
      RECT 0.0000 407.5200 210.2200 409.1600 ;
      RECT 207.9600 406.4400 210.2200 407.5200 ;
      RECT 4.8600 406.4400 205.3600 407.5200 ;
      RECT 0.0000 406.4400 2.2600 407.5200 ;
      RECT 0.0000 404.8000 210.2200 406.4400 ;
      RECT 204.9600 403.7200 210.2200 404.8000 ;
      RECT 7.8600 403.7200 202.3600 404.8000 ;
      RECT 0.0000 403.7200 5.2600 404.8000 ;
      RECT 0.0000 402.0800 210.2200 403.7200 ;
      RECT 207.9600 401.0000 210.2200 402.0800 ;
      RECT 4.8600 401.0000 205.3600 402.0800 ;
      RECT 0.0000 401.0000 2.2600 402.0800 ;
      RECT 0.0000 399.3600 210.2200 401.0000 ;
      RECT 204.9600 398.2800 210.2200 399.3600 ;
      RECT 7.8600 398.2800 202.3600 399.3600 ;
      RECT 0.0000 398.2800 5.2600 399.3600 ;
      RECT 0.0000 396.6400 210.2200 398.2800 ;
      RECT 207.9600 395.5600 210.2200 396.6400 ;
      RECT 4.8600 395.5600 205.3600 396.6400 ;
      RECT 0.0000 395.5600 2.2600 396.6400 ;
      RECT 0.0000 393.9200 210.2200 395.5600 ;
      RECT 204.9600 392.8400 210.2200 393.9200 ;
      RECT 7.8600 392.8400 202.3600 393.9200 ;
      RECT 0.0000 392.8400 5.2600 393.9200 ;
      RECT 0.0000 391.2000 210.2200 392.8400 ;
      RECT 207.9600 390.1200 210.2200 391.2000 ;
      RECT 4.8600 390.1200 205.3600 391.2000 ;
      RECT 0.0000 390.1200 2.2600 391.2000 ;
      RECT 0.0000 388.4800 210.2200 390.1200 ;
      RECT 204.9600 387.4000 210.2200 388.4800 ;
      RECT 7.8600 387.4000 202.3600 388.4800 ;
      RECT 0.0000 387.4000 5.2600 388.4800 ;
      RECT 0.0000 385.7600 210.2200 387.4000 ;
      RECT 207.9600 384.6800 210.2200 385.7600 ;
      RECT 4.8600 384.6800 205.3600 385.7600 ;
      RECT 0.0000 384.6800 2.2600 385.7600 ;
      RECT 0.0000 383.0400 210.2200 384.6800 ;
      RECT 204.9600 381.9600 210.2200 383.0400 ;
      RECT 7.8600 381.9600 202.3600 383.0400 ;
      RECT 0.0000 381.9600 5.2600 383.0400 ;
      RECT 0.0000 380.3200 210.2200 381.9600 ;
      RECT 207.9600 379.2400 210.2200 380.3200 ;
      RECT 4.8600 379.2400 205.3600 380.3200 ;
      RECT 0.0000 379.2400 2.2600 380.3200 ;
      RECT 0.0000 377.6000 210.2200 379.2400 ;
      RECT 204.9600 376.5200 210.2200 377.6000 ;
      RECT 7.8600 376.5200 202.3600 377.6000 ;
      RECT 0.0000 376.5200 5.2600 377.6000 ;
      RECT 0.0000 374.8800 210.2200 376.5200 ;
      RECT 207.9600 373.8000 210.2200 374.8800 ;
      RECT 4.8600 373.8000 205.3600 374.8800 ;
      RECT 0.0000 373.8000 2.2600 374.8800 ;
      RECT 0.0000 372.1600 210.2200 373.8000 ;
      RECT 204.9600 371.0800 210.2200 372.1600 ;
      RECT 7.8600 371.0800 202.3600 372.1600 ;
      RECT 0.0000 371.0800 5.2600 372.1600 ;
      RECT 0.0000 369.4400 210.2200 371.0800 ;
      RECT 207.9600 368.3600 210.2200 369.4400 ;
      RECT 4.8600 368.3600 205.3600 369.4400 ;
      RECT 0.0000 368.3600 2.2600 369.4400 ;
      RECT 0.0000 366.7200 210.2200 368.3600 ;
      RECT 204.9600 365.6400 210.2200 366.7200 ;
      RECT 7.8600 365.6400 202.3600 366.7200 ;
      RECT 0.0000 365.6400 5.2600 366.7200 ;
      RECT 0.0000 364.0000 210.2200 365.6400 ;
      RECT 207.9600 362.9200 210.2200 364.0000 ;
      RECT 4.8600 362.9200 205.3600 364.0000 ;
      RECT 0.0000 362.9200 2.2600 364.0000 ;
      RECT 0.0000 361.2800 210.2200 362.9200 ;
      RECT 204.9600 360.2000 210.2200 361.2800 ;
      RECT 7.8600 360.2000 202.3600 361.2800 ;
      RECT 0.0000 360.2000 5.2600 361.2800 ;
      RECT 0.0000 358.5600 210.2200 360.2000 ;
      RECT 207.9600 357.4800 210.2200 358.5600 ;
      RECT 4.8600 357.4800 205.3600 358.5600 ;
      RECT 0.0000 357.4800 2.2600 358.5600 ;
      RECT 0.0000 355.8400 210.2200 357.4800 ;
      RECT 204.9600 354.7600 210.2200 355.8400 ;
      RECT 7.8600 354.7600 202.3600 355.8400 ;
      RECT 0.0000 354.7600 5.2600 355.8400 ;
      RECT 0.0000 353.1200 210.2200 354.7600 ;
      RECT 207.9600 352.0400 210.2200 353.1200 ;
      RECT 4.8600 352.0400 205.3600 353.1200 ;
      RECT 0.0000 352.0400 2.2600 353.1200 ;
      RECT 0.0000 350.4000 210.2200 352.0400 ;
      RECT 204.9600 349.3200 210.2200 350.4000 ;
      RECT 7.8600 349.3200 202.3600 350.4000 ;
      RECT 0.0000 349.3200 5.2600 350.4000 ;
      RECT 0.0000 347.6800 210.2200 349.3200 ;
      RECT 207.9600 346.6000 210.2200 347.6800 ;
      RECT 4.8600 346.6000 205.3600 347.6800 ;
      RECT 0.0000 346.6000 2.2600 347.6800 ;
      RECT 0.0000 344.9600 210.2200 346.6000 ;
      RECT 204.9600 343.8800 210.2200 344.9600 ;
      RECT 7.8600 343.8800 202.3600 344.9600 ;
      RECT 0.0000 343.8800 5.2600 344.9600 ;
      RECT 0.0000 342.2400 210.2200 343.8800 ;
      RECT 207.9600 341.1600 210.2200 342.2400 ;
      RECT 4.8600 341.1600 205.3600 342.2400 ;
      RECT 0.0000 341.1600 2.2600 342.2400 ;
      RECT 0.0000 339.5200 210.2200 341.1600 ;
      RECT 204.9600 338.4400 210.2200 339.5200 ;
      RECT 7.8600 338.4400 202.3600 339.5200 ;
      RECT 0.0000 338.4400 5.2600 339.5200 ;
      RECT 0.0000 336.8000 210.2200 338.4400 ;
      RECT 207.9600 335.7200 210.2200 336.8000 ;
      RECT 4.8600 335.7200 205.3600 336.8000 ;
      RECT 0.0000 335.7200 2.2600 336.8000 ;
      RECT 0.0000 334.0800 210.2200 335.7200 ;
      RECT 204.9600 333.0000 210.2200 334.0800 ;
      RECT 7.8600 333.0000 202.3600 334.0800 ;
      RECT 0.0000 333.0000 5.2600 334.0800 ;
      RECT 0.0000 331.3600 210.2200 333.0000 ;
      RECT 207.9600 330.2800 210.2200 331.3600 ;
      RECT 4.8600 330.2800 205.3600 331.3600 ;
      RECT 0.0000 330.2800 2.2600 331.3600 ;
      RECT 0.0000 328.6400 210.2200 330.2800 ;
      RECT 204.9600 327.5600 210.2200 328.6400 ;
      RECT 7.8600 327.5600 202.3600 328.6400 ;
      RECT 0.0000 327.5600 5.2600 328.6400 ;
      RECT 0.0000 325.9200 210.2200 327.5600 ;
      RECT 207.9600 324.8400 210.2200 325.9200 ;
      RECT 4.8600 324.8400 205.3600 325.9200 ;
      RECT 0.0000 324.8400 2.2600 325.9200 ;
      RECT 0.0000 323.2000 210.2200 324.8400 ;
      RECT 204.9600 322.1200 210.2200 323.2000 ;
      RECT 7.8600 322.1200 202.3600 323.2000 ;
      RECT 0.0000 322.1200 5.2600 323.2000 ;
      RECT 0.0000 320.4800 210.2200 322.1200 ;
      RECT 207.9600 319.4000 210.2200 320.4800 ;
      RECT 4.8600 319.4000 205.3600 320.4800 ;
      RECT 0.0000 319.4000 2.2600 320.4800 ;
      RECT 0.0000 317.7600 210.2200 319.4000 ;
      RECT 204.9600 316.6800 210.2200 317.7600 ;
      RECT 7.8600 316.6800 202.3600 317.7600 ;
      RECT 0.0000 316.6800 5.2600 317.7600 ;
      RECT 0.0000 315.0400 210.2200 316.6800 ;
      RECT 207.9600 313.9600 210.2200 315.0400 ;
      RECT 4.8600 313.9600 205.3600 315.0400 ;
      RECT 0.0000 313.9600 2.2600 315.0400 ;
      RECT 0.0000 312.3200 210.2200 313.9600 ;
      RECT 204.9600 311.2400 210.2200 312.3200 ;
      RECT 7.8600 311.2400 202.3600 312.3200 ;
      RECT 0.0000 311.2400 5.2600 312.3200 ;
      RECT 0.0000 309.6000 210.2200 311.2400 ;
      RECT 207.9600 308.5200 210.2200 309.6000 ;
      RECT 4.8600 308.5200 205.3600 309.6000 ;
      RECT 0.0000 308.5200 2.2600 309.6000 ;
      RECT 0.0000 306.8800 210.2200 308.5200 ;
      RECT 204.9600 305.8000 210.2200 306.8800 ;
      RECT 7.8600 305.8000 202.3600 306.8800 ;
      RECT 0.0000 305.8000 5.2600 306.8800 ;
      RECT 0.0000 304.1600 210.2200 305.8000 ;
      RECT 207.9600 303.0800 210.2200 304.1600 ;
      RECT 4.8600 303.0800 205.3600 304.1600 ;
      RECT 0.0000 303.0800 2.2600 304.1600 ;
      RECT 0.0000 301.4400 210.2200 303.0800 ;
      RECT 204.9600 300.3600 210.2200 301.4400 ;
      RECT 7.8600 300.3600 202.3600 301.4400 ;
      RECT 0.0000 300.3600 5.2600 301.4400 ;
      RECT 0.0000 298.7200 210.2200 300.3600 ;
      RECT 207.9600 297.6400 210.2200 298.7200 ;
      RECT 4.8600 297.6400 205.3600 298.7200 ;
      RECT 0.0000 297.6400 2.2600 298.7200 ;
      RECT 0.0000 296.0000 210.2200 297.6400 ;
      RECT 204.9600 294.9200 210.2200 296.0000 ;
      RECT 7.8600 294.9200 202.3600 296.0000 ;
      RECT 0.0000 294.9200 5.2600 296.0000 ;
      RECT 0.0000 293.2800 210.2200 294.9200 ;
      RECT 207.9600 292.2000 210.2200 293.2800 ;
      RECT 4.8600 292.2000 205.3600 293.2800 ;
      RECT 0.0000 292.2000 2.2600 293.2800 ;
      RECT 0.0000 290.5600 210.2200 292.2000 ;
      RECT 204.9600 289.4800 210.2200 290.5600 ;
      RECT 7.8600 289.4800 202.3600 290.5600 ;
      RECT 0.0000 289.4800 5.2600 290.5600 ;
      RECT 0.0000 287.8400 210.2200 289.4800 ;
      RECT 207.9600 286.7600 210.2200 287.8400 ;
      RECT 4.8600 286.7600 205.3600 287.8400 ;
      RECT 0.0000 286.7600 2.2600 287.8400 ;
      RECT 0.0000 285.1200 210.2200 286.7600 ;
      RECT 204.9600 284.0400 210.2200 285.1200 ;
      RECT 7.8600 284.0400 202.3600 285.1200 ;
      RECT 0.0000 284.0400 5.2600 285.1200 ;
      RECT 0.0000 282.4000 210.2200 284.0400 ;
      RECT 207.9600 281.3200 210.2200 282.4000 ;
      RECT 4.8600 281.3200 205.3600 282.4000 ;
      RECT 0.0000 281.3200 2.2600 282.4000 ;
      RECT 0.0000 279.6800 210.2200 281.3200 ;
      RECT 204.9600 278.6000 210.2200 279.6800 ;
      RECT 7.8600 278.6000 202.3600 279.6800 ;
      RECT 0.0000 278.6000 5.2600 279.6800 ;
      RECT 0.0000 276.9600 210.2200 278.6000 ;
      RECT 207.9600 275.8800 210.2200 276.9600 ;
      RECT 4.8600 275.8800 205.3600 276.9600 ;
      RECT 0.0000 275.8800 2.2600 276.9600 ;
      RECT 0.0000 274.2400 210.2200 275.8800 ;
      RECT 204.9600 273.1600 210.2200 274.2400 ;
      RECT 7.8600 273.1600 202.3600 274.2400 ;
      RECT 0.0000 273.1600 5.2600 274.2400 ;
      RECT 0.0000 271.5200 210.2200 273.1600 ;
      RECT 207.9600 270.4400 210.2200 271.5200 ;
      RECT 4.8600 270.4400 205.3600 271.5200 ;
      RECT 0.0000 270.4400 2.2600 271.5200 ;
      RECT 0.0000 268.8000 210.2200 270.4400 ;
      RECT 204.9600 267.7200 210.2200 268.8000 ;
      RECT 7.8600 267.7200 202.3600 268.8000 ;
      RECT 0.0000 267.7200 5.2600 268.8000 ;
      RECT 0.0000 266.0800 210.2200 267.7200 ;
      RECT 207.9600 265.0000 210.2200 266.0800 ;
      RECT 4.8600 265.0000 205.3600 266.0800 ;
      RECT 0.0000 265.0000 2.2600 266.0800 ;
      RECT 0.0000 263.3600 210.2200 265.0000 ;
      RECT 204.9600 262.2800 210.2200 263.3600 ;
      RECT 7.8600 262.2800 202.3600 263.3600 ;
      RECT 0.0000 262.2800 5.2600 263.3600 ;
      RECT 0.0000 260.6400 210.2200 262.2800 ;
      RECT 207.9600 259.5600 210.2200 260.6400 ;
      RECT 4.8600 259.5600 205.3600 260.6400 ;
      RECT 0.0000 259.5600 2.2600 260.6400 ;
      RECT 0.0000 257.9200 210.2200 259.5600 ;
      RECT 204.9600 256.8400 210.2200 257.9200 ;
      RECT 7.8600 256.8400 202.3600 257.9200 ;
      RECT 0.0000 256.8400 5.2600 257.9200 ;
      RECT 0.0000 255.2000 210.2200 256.8400 ;
      RECT 207.9600 254.1200 210.2200 255.2000 ;
      RECT 4.8600 254.1200 205.3600 255.2000 ;
      RECT 0.0000 254.1200 2.2600 255.2000 ;
      RECT 0.0000 252.4800 210.2200 254.1200 ;
      RECT 204.9600 251.4000 210.2200 252.4800 ;
      RECT 7.8600 251.4000 202.3600 252.4800 ;
      RECT 0.0000 251.4000 5.2600 252.4800 ;
      RECT 0.0000 249.7600 210.2200 251.4000 ;
      RECT 207.9600 248.6800 210.2200 249.7600 ;
      RECT 4.8600 248.6800 205.3600 249.7600 ;
      RECT 0.0000 248.6800 2.2600 249.7600 ;
      RECT 0.0000 247.0400 210.2200 248.6800 ;
      RECT 204.9600 245.9600 210.2200 247.0400 ;
      RECT 7.8600 245.9600 202.3600 247.0400 ;
      RECT 0.0000 245.9600 5.2600 247.0400 ;
      RECT 0.0000 244.3200 210.2200 245.9600 ;
      RECT 207.9600 243.2400 210.2200 244.3200 ;
      RECT 4.8600 243.2400 205.3600 244.3200 ;
      RECT 0.0000 243.2400 2.2600 244.3200 ;
      RECT 0.0000 241.6000 210.2200 243.2400 ;
      RECT 204.9600 240.5200 210.2200 241.6000 ;
      RECT 7.8600 240.5200 202.3600 241.6000 ;
      RECT 0.0000 240.5200 5.2600 241.6000 ;
      RECT 0.0000 238.8800 210.2200 240.5200 ;
      RECT 207.9600 237.8000 210.2200 238.8800 ;
      RECT 4.8600 237.8000 205.3600 238.8800 ;
      RECT 0.0000 237.8000 2.2600 238.8800 ;
      RECT 0.0000 236.1600 210.2200 237.8000 ;
      RECT 204.9600 235.0800 210.2200 236.1600 ;
      RECT 7.8600 235.0800 202.3600 236.1600 ;
      RECT 0.0000 235.0800 5.2600 236.1600 ;
      RECT 0.0000 233.4400 210.2200 235.0800 ;
      RECT 207.9600 232.3600 210.2200 233.4400 ;
      RECT 4.8600 232.3600 205.3600 233.4400 ;
      RECT 0.0000 232.3600 2.2600 233.4400 ;
      RECT 0.0000 230.7200 210.2200 232.3600 ;
      RECT 204.9600 229.6400 210.2200 230.7200 ;
      RECT 7.8600 229.6400 202.3600 230.7200 ;
      RECT 0.0000 229.6400 5.2600 230.7200 ;
      RECT 0.0000 228.0000 210.2200 229.6400 ;
      RECT 207.9600 226.9200 210.2200 228.0000 ;
      RECT 4.8600 226.9200 205.3600 228.0000 ;
      RECT 0.0000 226.9200 2.2600 228.0000 ;
      RECT 0.0000 225.2800 210.2200 226.9200 ;
      RECT 204.9600 224.2000 210.2200 225.2800 ;
      RECT 7.8600 224.2000 202.3600 225.2800 ;
      RECT 0.0000 224.2000 5.2600 225.2800 ;
      RECT 0.0000 222.5600 210.2200 224.2000 ;
      RECT 207.9600 221.4800 210.2200 222.5600 ;
      RECT 4.8600 221.4800 205.3600 222.5600 ;
      RECT 0.0000 221.4800 2.2600 222.5600 ;
      RECT 0.0000 219.8400 210.2200 221.4800 ;
      RECT 204.9600 218.7600 210.2200 219.8400 ;
      RECT 7.8600 218.7600 202.3600 219.8400 ;
      RECT 0.0000 218.7600 5.2600 219.8400 ;
      RECT 0.0000 217.1200 210.2200 218.7600 ;
      RECT 207.9600 216.0400 210.2200 217.1200 ;
      RECT 4.8600 216.0400 205.3600 217.1200 ;
      RECT 0.0000 216.0400 2.2600 217.1200 ;
      RECT 0.0000 214.4000 210.2200 216.0400 ;
      RECT 204.9600 213.3200 210.2200 214.4000 ;
      RECT 7.8600 213.3200 202.3600 214.4000 ;
      RECT 0.0000 213.3200 5.2600 214.4000 ;
      RECT 0.0000 211.6800 210.2200 213.3200 ;
      RECT 207.9600 210.6000 210.2200 211.6800 ;
      RECT 4.8600 210.6000 205.3600 211.6800 ;
      RECT 0.0000 210.6000 2.2600 211.6800 ;
      RECT 0.0000 208.9600 210.2200 210.6000 ;
      RECT 204.9600 207.8800 210.2200 208.9600 ;
      RECT 7.8600 207.8800 202.3600 208.9600 ;
      RECT 0.0000 207.8800 5.2600 208.9600 ;
      RECT 0.0000 206.2400 210.2200 207.8800 ;
      RECT 207.9600 205.1600 210.2200 206.2400 ;
      RECT 4.8600 205.1600 205.3600 206.2400 ;
      RECT 0.0000 205.1600 2.2600 206.2400 ;
      RECT 0.0000 203.5200 210.2200 205.1600 ;
      RECT 204.9600 202.4400 210.2200 203.5200 ;
      RECT 7.8600 202.4400 202.3600 203.5200 ;
      RECT 0.0000 202.4400 5.2600 203.5200 ;
      RECT 0.0000 200.8000 210.2200 202.4400 ;
      RECT 207.9600 199.7200 210.2200 200.8000 ;
      RECT 4.8600 199.7200 205.3600 200.8000 ;
      RECT 0.0000 199.7200 2.2600 200.8000 ;
      RECT 0.0000 198.0800 210.2200 199.7200 ;
      RECT 204.9600 197.0000 210.2200 198.0800 ;
      RECT 7.8600 197.0000 202.3600 198.0800 ;
      RECT 0.0000 197.0000 5.2600 198.0800 ;
      RECT 0.0000 195.3600 210.2200 197.0000 ;
      RECT 207.9600 194.2800 210.2200 195.3600 ;
      RECT 4.8600 194.2800 205.3600 195.3600 ;
      RECT 0.0000 194.2800 2.2600 195.3600 ;
      RECT 0.0000 192.6400 210.2200 194.2800 ;
      RECT 204.9600 191.5600 210.2200 192.6400 ;
      RECT 7.8600 191.5600 202.3600 192.6400 ;
      RECT 0.0000 191.5600 5.2600 192.6400 ;
      RECT 0.0000 189.9200 210.2200 191.5600 ;
      RECT 207.9600 188.8400 210.2200 189.9200 ;
      RECT 4.8600 188.8400 205.3600 189.9200 ;
      RECT 0.0000 188.8400 2.2600 189.9200 ;
      RECT 0.0000 187.2000 210.2200 188.8400 ;
      RECT 204.9600 186.1200 210.2200 187.2000 ;
      RECT 7.8600 186.1200 202.3600 187.2000 ;
      RECT 0.0000 186.1200 5.2600 187.2000 ;
      RECT 0.0000 184.4800 210.2200 186.1200 ;
      RECT 207.9600 183.4000 210.2200 184.4800 ;
      RECT 4.8600 183.4000 205.3600 184.4800 ;
      RECT 0.0000 183.4000 2.2600 184.4800 ;
      RECT 0.0000 181.7600 210.2200 183.4000 ;
      RECT 204.9600 180.6800 210.2200 181.7600 ;
      RECT 7.8600 180.6800 202.3600 181.7600 ;
      RECT 0.0000 180.6800 5.2600 181.7600 ;
      RECT 0.0000 179.0400 210.2200 180.6800 ;
      RECT 207.9600 177.9600 210.2200 179.0400 ;
      RECT 4.8600 177.9600 205.3600 179.0400 ;
      RECT 0.0000 177.9600 2.2600 179.0400 ;
      RECT 0.0000 176.3200 210.2200 177.9600 ;
      RECT 204.9600 175.2400 210.2200 176.3200 ;
      RECT 7.8600 175.2400 202.3600 176.3200 ;
      RECT 0.0000 175.2400 5.2600 176.3200 ;
      RECT 0.0000 173.6000 210.2200 175.2400 ;
      RECT 207.9600 172.5200 210.2200 173.6000 ;
      RECT 4.8600 172.5200 205.3600 173.6000 ;
      RECT 0.0000 172.5200 2.2600 173.6000 ;
      RECT 0.0000 170.8800 210.2200 172.5200 ;
      RECT 204.9600 169.8000 210.2200 170.8800 ;
      RECT 7.8600 169.8000 202.3600 170.8800 ;
      RECT 0.0000 169.8000 5.2600 170.8800 ;
      RECT 0.0000 168.1600 210.2200 169.8000 ;
      RECT 207.9600 167.0800 210.2200 168.1600 ;
      RECT 4.8600 167.0800 205.3600 168.1600 ;
      RECT 0.0000 167.0800 2.2600 168.1600 ;
      RECT 0.0000 165.4400 210.2200 167.0800 ;
      RECT 204.9600 164.3600 210.2200 165.4400 ;
      RECT 7.8600 164.3600 202.3600 165.4400 ;
      RECT 0.0000 164.3600 5.2600 165.4400 ;
      RECT 0.0000 162.7200 210.2200 164.3600 ;
      RECT 207.9600 161.6400 210.2200 162.7200 ;
      RECT 4.8600 161.6400 205.3600 162.7200 ;
      RECT 0.0000 161.6400 2.2600 162.7200 ;
      RECT 0.0000 160.0000 210.2200 161.6400 ;
      RECT 204.9600 158.9200 210.2200 160.0000 ;
      RECT 7.8600 158.9200 202.3600 160.0000 ;
      RECT 0.0000 158.9200 5.2600 160.0000 ;
      RECT 0.0000 157.2800 210.2200 158.9200 ;
      RECT 207.9600 156.2000 210.2200 157.2800 ;
      RECT 4.8600 156.2000 205.3600 157.2800 ;
      RECT 0.0000 156.2000 2.2600 157.2800 ;
      RECT 0.0000 154.5600 210.2200 156.2000 ;
      RECT 204.9600 153.4800 210.2200 154.5600 ;
      RECT 7.8600 153.4800 202.3600 154.5600 ;
      RECT 0.0000 153.4800 5.2600 154.5600 ;
      RECT 0.0000 151.8400 210.2200 153.4800 ;
      RECT 207.9600 150.7600 210.2200 151.8400 ;
      RECT 4.8600 150.7600 205.3600 151.8400 ;
      RECT 0.0000 150.7600 2.2600 151.8400 ;
      RECT 0.0000 149.1200 210.2200 150.7600 ;
      RECT 204.9600 148.0400 210.2200 149.1200 ;
      RECT 7.8600 148.0400 202.3600 149.1200 ;
      RECT 0.0000 148.0400 5.2600 149.1200 ;
      RECT 0.0000 146.4000 210.2200 148.0400 ;
      RECT 207.9600 145.3200 210.2200 146.4000 ;
      RECT 4.8600 145.3200 205.3600 146.4000 ;
      RECT 0.0000 145.3200 2.2600 146.4000 ;
      RECT 0.0000 143.6800 210.2200 145.3200 ;
      RECT 204.9600 142.6000 210.2200 143.6800 ;
      RECT 7.8600 142.6000 202.3600 143.6800 ;
      RECT 0.0000 142.6000 5.2600 143.6800 ;
      RECT 0.0000 140.9600 210.2200 142.6000 ;
      RECT 207.9600 139.8800 210.2200 140.9600 ;
      RECT 4.8600 139.8800 205.3600 140.9600 ;
      RECT 0.0000 139.8800 2.2600 140.9600 ;
      RECT 0.0000 138.2400 210.2200 139.8800 ;
      RECT 204.9600 137.1600 210.2200 138.2400 ;
      RECT 7.8600 137.1600 202.3600 138.2400 ;
      RECT 0.0000 137.1600 5.2600 138.2400 ;
      RECT 0.0000 135.5200 210.2200 137.1600 ;
      RECT 207.9600 134.4400 210.2200 135.5200 ;
      RECT 4.8600 134.4400 205.3600 135.5200 ;
      RECT 0.0000 134.4400 2.2600 135.5200 ;
      RECT 0.0000 132.8000 210.2200 134.4400 ;
      RECT 204.9600 131.7200 210.2200 132.8000 ;
      RECT 7.8600 131.7200 202.3600 132.8000 ;
      RECT 0.0000 131.7200 5.2600 132.8000 ;
      RECT 0.0000 130.0800 210.2200 131.7200 ;
      RECT 207.9600 129.0000 210.2200 130.0800 ;
      RECT 4.8600 129.0000 205.3600 130.0800 ;
      RECT 0.0000 129.0000 2.2600 130.0800 ;
      RECT 0.0000 127.3600 210.2200 129.0000 ;
      RECT 204.9600 126.2800 210.2200 127.3600 ;
      RECT 7.8600 126.2800 202.3600 127.3600 ;
      RECT 0.0000 126.2800 5.2600 127.3600 ;
      RECT 0.0000 124.6400 210.2200 126.2800 ;
      RECT 207.9600 123.5600 210.2200 124.6400 ;
      RECT 4.8600 123.5600 205.3600 124.6400 ;
      RECT 0.0000 123.5600 2.2600 124.6400 ;
      RECT 0.0000 121.9200 210.2200 123.5600 ;
      RECT 204.9600 120.8400 210.2200 121.9200 ;
      RECT 7.8600 120.8400 202.3600 121.9200 ;
      RECT 0.0000 120.8400 5.2600 121.9200 ;
      RECT 0.0000 119.2000 210.2200 120.8400 ;
      RECT 207.9600 118.1200 210.2200 119.2000 ;
      RECT 4.8600 118.1200 205.3600 119.2000 ;
      RECT 0.0000 118.1200 2.2600 119.2000 ;
      RECT 0.0000 116.4800 210.2200 118.1200 ;
      RECT 204.9600 115.4000 210.2200 116.4800 ;
      RECT 7.8600 115.4000 202.3600 116.4800 ;
      RECT 0.0000 115.4000 5.2600 116.4800 ;
      RECT 0.0000 113.7600 210.2200 115.4000 ;
      RECT 207.9600 112.6800 210.2200 113.7600 ;
      RECT 4.8600 112.6800 205.3600 113.7600 ;
      RECT 0.0000 112.6800 2.2600 113.7600 ;
      RECT 0.0000 111.0400 210.2200 112.6800 ;
      RECT 204.9600 109.9600 210.2200 111.0400 ;
      RECT 7.8600 109.9600 202.3600 111.0400 ;
      RECT 0.0000 109.9600 5.2600 111.0400 ;
      RECT 0.0000 108.3200 210.2200 109.9600 ;
      RECT 207.9600 107.2400 210.2200 108.3200 ;
      RECT 4.8600 107.2400 205.3600 108.3200 ;
      RECT 0.0000 107.2400 2.2600 108.3200 ;
      RECT 0.0000 105.6000 210.2200 107.2400 ;
      RECT 204.9600 104.5200 210.2200 105.6000 ;
      RECT 7.8600 104.5200 202.3600 105.6000 ;
      RECT 0.0000 104.5200 5.2600 105.6000 ;
      RECT 0.0000 102.8800 210.2200 104.5200 ;
      RECT 207.9600 101.8000 210.2200 102.8800 ;
      RECT 4.8600 101.8000 205.3600 102.8800 ;
      RECT 0.0000 101.8000 2.2600 102.8800 ;
      RECT 0.0000 100.1600 210.2200 101.8000 ;
      RECT 204.9600 99.0800 210.2200 100.1600 ;
      RECT 7.8600 99.0800 202.3600 100.1600 ;
      RECT 0.0000 99.0800 5.2600 100.1600 ;
      RECT 0.0000 97.4400 210.2200 99.0800 ;
      RECT 207.9600 96.3600 210.2200 97.4400 ;
      RECT 4.8600 96.3600 205.3600 97.4400 ;
      RECT 0.0000 96.3600 2.2600 97.4400 ;
      RECT 0.0000 94.7200 210.2200 96.3600 ;
      RECT 204.9600 93.6400 210.2200 94.7200 ;
      RECT 7.8600 93.6400 202.3600 94.7200 ;
      RECT 0.0000 93.6400 5.2600 94.7200 ;
      RECT 0.0000 92.0000 210.2200 93.6400 ;
      RECT 207.9600 90.9200 210.2200 92.0000 ;
      RECT 4.8600 90.9200 205.3600 92.0000 ;
      RECT 0.0000 90.9200 2.2600 92.0000 ;
      RECT 0.0000 89.2800 210.2200 90.9200 ;
      RECT 204.9600 88.2000 210.2200 89.2800 ;
      RECT 7.8600 88.2000 202.3600 89.2800 ;
      RECT 0.0000 88.2000 5.2600 89.2800 ;
      RECT 0.0000 86.5600 210.2200 88.2000 ;
      RECT 207.9600 85.4800 210.2200 86.5600 ;
      RECT 4.8600 85.4800 205.3600 86.5600 ;
      RECT 0.0000 85.4800 2.2600 86.5600 ;
      RECT 0.0000 83.8400 210.2200 85.4800 ;
      RECT 204.9600 82.7600 210.2200 83.8400 ;
      RECT 7.8600 82.7600 202.3600 83.8400 ;
      RECT 0.0000 82.7600 5.2600 83.8400 ;
      RECT 0.0000 81.1200 210.2200 82.7600 ;
      RECT 207.9600 80.0400 210.2200 81.1200 ;
      RECT 4.8600 80.0400 205.3600 81.1200 ;
      RECT 0.0000 80.0400 2.2600 81.1200 ;
      RECT 0.0000 78.4000 210.2200 80.0400 ;
      RECT 204.9600 77.3200 210.2200 78.4000 ;
      RECT 7.8600 77.3200 202.3600 78.4000 ;
      RECT 0.0000 77.3200 5.2600 78.4000 ;
      RECT 0.0000 75.6800 210.2200 77.3200 ;
      RECT 207.9600 74.6000 210.2200 75.6800 ;
      RECT 4.8600 74.6000 205.3600 75.6800 ;
      RECT 0.0000 74.6000 2.2600 75.6800 ;
      RECT 0.0000 72.9600 210.2200 74.6000 ;
      RECT 204.9600 71.8800 210.2200 72.9600 ;
      RECT 7.8600 71.8800 202.3600 72.9600 ;
      RECT 0.0000 71.8800 5.2600 72.9600 ;
      RECT 0.0000 70.2400 210.2200 71.8800 ;
      RECT 207.9600 69.1600 210.2200 70.2400 ;
      RECT 4.8600 69.1600 205.3600 70.2400 ;
      RECT 0.0000 69.1600 2.2600 70.2400 ;
      RECT 0.0000 67.5200 210.2200 69.1600 ;
      RECT 204.9600 66.4400 210.2200 67.5200 ;
      RECT 7.8600 66.4400 202.3600 67.5200 ;
      RECT 0.0000 66.4400 5.2600 67.5200 ;
      RECT 0.0000 64.8000 210.2200 66.4400 ;
      RECT 207.9600 63.7200 210.2200 64.8000 ;
      RECT 4.8600 63.7200 205.3600 64.8000 ;
      RECT 0.0000 63.7200 2.2600 64.8000 ;
      RECT 0.0000 62.0800 210.2200 63.7200 ;
      RECT 204.9600 61.0000 210.2200 62.0800 ;
      RECT 7.8600 61.0000 202.3600 62.0800 ;
      RECT 0.0000 61.0000 5.2600 62.0800 ;
      RECT 0.0000 59.3600 210.2200 61.0000 ;
      RECT 207.9600 58.2800 210.2200 59.3600 ;
      RECT 4.8600 58.2800 205.3600 59.3600 ;
      RECT 0.0000 58.2800 2.2600 59.3600 ;
      RECT 0.0000 56.6400 210.2200 58.2800 ;
      RECT 204.9600 55.5600 210.2200 56.6400 ;
      RECT 7.8600 55.5600 202.3600 56.6400 ;
      RECT 0.0000 55.5600 5.2600 56.6400 ;
      RECT 0.0000 53.9200 210.2200 55.5600 ;
      RECT 207.9600 52.8400 210.2200 53.9200 ;
      RECT 4.8600 52.8400 205.3600 53.9200 ;
      RECT 0.0000 52.8400 2.2600 53.9200 ;
      RECT 0.0000 51.2000 210.2200 52.8400 ;
      RECT 204.9600 50.1200 210.2200 51.2000 ;
      RECT 7.8600 50.1200 202.3600 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 210.2200 50.1200 ;
      RECT 207.9600 47.4000 210.2200 48.4800 ;
      RECT 4.8600 47.4000 205.3600 48.4800 ;
      RECT 0.0000 47.4000 2.2600 48.4800 ;
      RECT 0.0000 45.7600 210.2200 47.4000 ;
      RECT 204.9600 44.6800 210.2200 45.7600 ;
      RECT 7.8600 44.6800 202.3600 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 210.2200 44.6800 ;
      RECT 207.9600 41.9600 210.2200 43.0400 ;
      RECT 4.8600 41.9600 205.3600 43.0400 ;
      RECT 0.0000 41.9600 2.2600 43.0400 ;
      RECT 0.0000 40.3200 210.2200 41.9600 ;
      RECT 204.9600 39.2400 210.2200 40.3200 ;
      RECT 7.8600 39.2400 202.3600 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 210.2200 39.2400 ;
      RECT 207.9600 36.5200 210.2200 37.6000 ;
      RECT 4.8600 36.5200 205.3600 37.6000 ;
      RECT 0.0000 36.5200 2.2600 37.6000 ;
      RECT 0.0000 34.8800 210.2200 36.5200 ;
      RECT 204.9600 33.8000 210.2200 34.8800 ;
      RECT 7.8600 33.8000 202.3600 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 210.2200 33.8000 ;
      RECT 207.9600 31.0800 210.2200 32.1600 ;
      RECT 4.8600 31.0800 205.3600 32.1600 ;
      RECT 0.0000 31.0800 2.2600 32.1600 ;
      RECT 0.0000 29.4400 210.2200 31.0800 ;
      RECT 204.9600 28.3600 210.2200 29.4400 ;
      RECT 7.8600 28.3600 202.3600 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 210.2200 28.3600 ;
      RECT 207.9600 25.6400 210.2200 26.7200 ;
      RECT 4.8600 25.6400 205.3600 26.7200 ;
      RECT 0.0000 25.6400 2.2600 26.7200 ;
      RECT 0.0000 24.0000 210.2200 25.6400 ;
      RECT 204.9600 22.9200 210.2200 24.0000 ;
      RECT 7.8600 22.9200 202.3600 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 210.2200 22.9200 ;
      RECT 207.9600 20.2000 210.2200 21.2800 ;
      RECT 4.8600 20.2000 205.3600 21.2800 ;
      RECT 0.0000 20.2000 2.2600 21.2800 ;
      RECT 0.0000 18.5600 210.2200 20.2000 ;
      RECT 204.9600 17.4800 210.2200 18.5600 ;
      RECT 7.8600 17.4800 202.3600 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 210.2200 17.4800 ;
      RECT 207.9600 14.7600 210.2200 15.8400 ;
      RECT 4.8600 14.7600 205.3600 15.8400 ;
      RECT 0.0000 14.7600 2.2600 15.8400 ;
      RECT 0.0000 13.1200 210.2200 14.7600 ;
      RECT 204.9600 12.0400 210.2200 13.1200 ;
      RECT 7.8600 12.0400 202.3600 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 210.2200 12.0400 ;
      RECT 207.9600 9.3200 210.2200 10.4000 ;
      RECT 4.8600 9.3200 205.3600 10.4000 ;
      RECT 0.0000 9.3200 2.2600 10.4000 ;
      RECT 0.0000 7.7300 210.2200 9.3200 ;
      RECT 204.9600 5.1300 210.2200 7.7300 ;
      RECT 0.0000 5.1300 5.2600 7.7300 ;
      RECT 0.0000 4.7300 210.2200 5.1300 ;
      RECT 207.9600 2.1300 210.2200 4.7300 ;
      RECT 0.0000 2.1300 2.2600 4.7300 ;
      RECT 0.0000 0.0000 210.2200 2.1300 ;
    LAYER met4 ;
      RECT 0.0000 447.5200 210.2200 449.8200 ;
      RECT 195.2200 444.5200 205.3600 447.5200 ;
      RECT 150.2200 444.5200 193.0200 447.5200 ;
      RECT 105.2200 444.5200 148.0200 447.5200 ;
      RECT 60.2200 444.5200 103.0200 447.5200 ;
      RECT 15.2200 444.5200 58.0200 447.5200 ;
      RECT 4.8600 444.5200 13.0200 447.5200 ;
      RECT 204.9600 5.1300 205.3600 444.5200 ;
      RECT 195.2200 5.1300 202.3600 444.5200 ;
      RECT 192.0200 5.1300 193.0200 444.5200 ;
      RECT 150.2200 5.1300 189.8200 444.5200 ;
      RECT 147.0200 5.1300 148.0200 444.5200 ;
      RECT 105.2200 5.1300 144.8200 444.5200 ;
      RECT 102.0200 5.1300 103.0200 444.5200 ;
      RECT 60.2200 5.1300 99.8200 444.5200 ;
      RECT 57.0200 5.1300 58.0200 444.5200 ;
      RECT 15.2200 5.1300 54.8200 444.5200 ;
      RECT 12.0200 5.1300 13.0200 444.5200 ;
      RECT 7.8600 5.1300 9.8200 444.5200 ;
      RECT 4.8600 5.1300 5.2600 444.5200 ;
      RECT 207.9600 2.1300 210.2200 447.5200 ;
      RECT 195.2200 2.1300 205.3600 5.1300 ;
      RECT 150.2200 2.1300 193.0200 5.1300 ;
      RECT 105.2200 2.1300 148.0200 5.1300 ;
      RECT 60.2200 2.1300 103.0200 5.1300 ;
      RECT 15.2200 2.1300 58.0200 5.1300 ;
      RECT 4.8600 2.1300 13.0200 5.1300 ;
      RECT 0.0000 2.1300 2.2600 447.5200 ;
      RECT 0.0000 1.0200 210.2200 2.1300 ;
      RECT 90.1900 0.0000 210.2200 1.0200 ;
      RECT 0.0000 0.0000 89.2100 1.0200 ;
  END
END DSP

END LIBRARY
