##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Wed Jun 30 15:39:28 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO eFPGA_top
  CLASS BLOCK ;
  SIZE 3390.2000 BY 2889.6600 ;
  FOREIGN eFPGA_top 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.4656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 56.5486 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 298.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.6587 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 94.4265 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 506.896 LAYER met4  ;
    ANTENNAGATEAREA 7.917 LAYER met4  ;
    ANTENNAMAXAREACAR 78.6355 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 395.707 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2799.4100 0.8000 2799.7100 ;
    END
  END wb_clk_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2774.4000 0.8000 2774.7000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2749.3900 0.8000 2749.6900 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2723.7700 0.8000 2724.0700 ;
    END
  END wbs_we_i
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2698.7600 0.8000 2699.0600 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2673.7500 0.8000 2674.0500 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2648.1300 0.8000 2648.4300 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2623.1200 0.8000 2623.4200 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2598.1100 0.8000 2598.4100 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2572.4900 0.8000 2572.7900 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2547.4800 0.8000 2547.7800 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2522.4700 0.8000 2522.7700 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2496.8500 0.8000 2497.1500 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2471.8400 0.8000 2472.1400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2446.8300 0.8000 2447.1300 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2421.2100 0.8000 2421.5100 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2396.2000 0.8000 2396.5000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2370.5800 0.8000 2370.8800 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2345.5700 0.8000 2345.8700 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2320.5600 0.8000 2320.8600 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2294.9400 0.8000 2295.2400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2269.9300 0.8000 2270.2300 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2244.9200 0.8000 2245.2200 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2219.3000 0.8000 2219.6000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2194.2900 0.8000 2194.5900 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2169.2800 0.8000 2169.5800 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2143.6600 0.8000 2143.9600 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2118.6500 0.8000 2118.9500 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2093.6400 0.8000 2093.9400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2068.0200 0.8000 2068.3200 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2043.0100 0.8000 2043.3100 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2017.3900 0.8000 2017.6900 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1992.3800 0.8000 1992.6800 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1967.3700 0.8000 1967.6700 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1941.7500 0.8000 1942.0500 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1916.7400 0.8000 1917.0400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1891.7300 0.8000 1892.0300 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1866.1100 0.8000 1866.4100 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1841.1000 0.8000 1841.4000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1816.0900 0.8000 1816.3900 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1790.4700 0.8000 1790.7700 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1765.4600 0.8000 1765.7600 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1740.4500 0.8000 1740.7500 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1714.8300 0.8000 1715.1300 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1689.8200 0.8000 1690.1200 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1664.8100 0.8000 1665.1100 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1639.1900 0.8000 1639.4900 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1614.1800 0.8000 1614.4800 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1588.5600 0.8000 1588.8600 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1563.5500 0.8000 1563.8500 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1538.5400 0.8000 1538.8400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1512.9200 0.8000 1513.2200 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1487.9100 0.8000 1488.2100 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1462.9000 0.8000 1463.2000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1437.2800 0.8000 1437.5800 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1412.2700 0.8000 1412.5700 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1387.2600 0.8000 1387.5600 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1361.6400 0.8000 1361.9400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1336.6300 0.8000 1336.9300 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1311.6200 0.8000 1311.9200 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1286.0000 0.8000 1286.3000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1260.9900 0.8000 1261.2900 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1235.3700 0.8000 1235.6700 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1210.3600 0.8000 1210.6600 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1185.3500 0.8000 1185.6500 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1159.7300 0.8000 1160.0300 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1134.7200 0.8000 1135.0200 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1109.7100 0.8000 1110.0100 ;
    END
  END wbs_adr_i[0]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2155 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1084.0900 0.8000 1084.3900 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1059.0800 0.8000 1059.3800 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.8032 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1034.0700 0.8000 1034.3700 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.8064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1008.4500 0.8000 1008.7500 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 93.3138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 498.144 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 983.4400 0.8000 983.7400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 958.4300 0.8000 958.7300 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 932.8100 0.8000 933.1100 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.8758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.808 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 907.8000 0.8000 908.1000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5983 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.9038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.624 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 882.7900 0.8000 883.0900 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.5844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 857.1700 0.8000 857.4700 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 832.1600 0.8000 832.4600 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 806.5400 0.8000 806.8400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 781.5300 0.8000 781.8300 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.3969 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.8168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 202.16 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 756.5200 0.8000 756.8200 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 240.605 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1283.7 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 730.9000 0.8000 731.2000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 262.781 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1401.97 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 705.8900 0.8000 706.1900 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.431 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 594.768 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 680.8800 0.8000 681.1800 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 120.263 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 641.872 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 655.2600 0.8000 655.5600 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 93.1068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 497.04 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 630.2500 0.8000 630.5500 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 102.05 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 544.736 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 605.2400 0.8000 605.5400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.0304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.824 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 579.6200 0.8000 579.9200 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7232 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 554.6100 0.8000 554.9100 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.6188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 489.104 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 529.6000 0.8000 529.9000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.888 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 503.9800 0.8000 504.2800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 148.166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 790.688 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 478.9700 0.8000 479.2700 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.8418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 372.96 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 453.3500 0.8000 453.6500 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.5188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 477.904 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 428.3400 0.8000 428.6400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.3974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 340.865 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1818.42 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 403.3300 0.8000 403.6300 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 313.598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1672.99 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 377.7100 0.8000 378.0100 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.902 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1376.42 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 352.7000 0.8000 353.0000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 213.434 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1138.78 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 327.6900 0.8000 327.9900 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 203.846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1087.65 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 302.0700 0.8000 302.3700 ;
    END
  END wbs_dat_o[0]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.0944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 277.0600 0.8000 277.3600 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 252.0500 0.8000 252.3500 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.1608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 237.608 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1260.53 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521429 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 226.4300 0.8000 226.7300 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.1232 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 198.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.064 LAYER met3  ;
    ANTENNAMAXAREACAR 87.47 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 425.613 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.328572 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 201.4200 0.8000 201.7200 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 176.4100 0.8000 176.7100 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4199 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 35.3706 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.131 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 150.7900 0.8000 151.0900 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 125.7800 0.8000 126.0800 ;
    END
  END la_data_out[0]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.3274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 141.358 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.8485 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 14.318 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 77.877 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.9800 2889.1750 100.1200 2889.6600 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.6268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 142.737 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.4474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met3  ;
    ANTENNAMAXAREACAR 29.8502 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 161.476 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0647249 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 32.4113 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.896 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0647249 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 580.2200 2889.1750 580.3600 2889.6600 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.616 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 253.794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1354.5 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.8485 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 14.318 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 77.877 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1060.0000 2889.1750 1060.1400 2889.6600 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.651 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.4474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met3  ;
    ANTENNAMAXAREACAR 29.8502 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 161.476 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0647249 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 32.4113 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.896 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0647249 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1540.2400 2889.1750 1540.3800 2889.6600 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.8778 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.992 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.8485 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 14.318 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 77.877 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2020.0200 2889.1750 2020.1600 2889.6600 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 77.0673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 384.822 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.4474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met3  ;
    ANTENNAMAXAREACAR 29.8502 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 161.476 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0647249 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 32.4113 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.896 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0647249 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2499.8000 2889.1750 2499.9400 2889.6600 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 105.24 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 525.819 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.8628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 10.8687 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 49.373 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2980.0400 2889.1750 2980.1800 2889.6600 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 10.5052 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 49.1032 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 2592.0100 3390.2000 2592.3100 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5219 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 57.9083 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.246 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 2280.9100 3390.2000 2281.2100 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 40.2837 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 205.044 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1969.2000 3390.2000 1969.5000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.9494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 9.97897 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 48.25 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1657.4900 3390.2000 1657.7900 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 9.51468 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 45.3532 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1346.3900 3390.2000 1346.6900 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5432 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 40.0782 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 205.119 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1034.6800 3390.2000 1034.9800 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 9.51468 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 45.3532 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 723.5800 3390.2000 723.8800 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 56.9139 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.615 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 411.8700 3390.2000 412.1700 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 8.67937 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 40.4722 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 100.7700 3390.2000 101.0700 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 115.853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 578.75 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 36.2036 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.492 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 3154.3800 0.0000 3154.5200 0.4850 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 74.4882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 372.162 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 76.8268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 410.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 58.5131 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 303 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2936.3400 0.0000 2936.4800 0.4850 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.3404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 291.305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.0678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 9.59722 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 45.5754 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2718.3000 0.0000 2718.4400 0.4850 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.5035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 45.7091 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 215.73 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 2500.2600 0.0000 2500.4000 0.4850 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.782 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.1116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 78.0591 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 410.345 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2281.7600 0.0000 2281.9000 0.4850 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 212.093 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 6.05913 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 23.7222 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2063.7200 0.0000 2063.8600 0.4850 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1663 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.6605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 7.15437 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 29.5635 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1845.6800 0.0000 1845.8200 0.4850 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 93.9131 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 484.992 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1627.1800 0.0000 1627.3200 0.4850 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.1400 0.0000 1409.2800 0.4850 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 192.903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 963.956 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.5399 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 24.181 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.698 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1191.1000 0.0000 1191.2400 0.4850 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 169.554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 847.371 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.5618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 42.5 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 217.813 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 973.0600 0.0000 973.2000 0.4850 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 211.365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1056.55 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.77 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 64.9873 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 328.131 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 754.5600 0.0000 754.7000 0.4850 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 196.21 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 980.574 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.9888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 7.95833 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.1468 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.362698 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 536.5200 0.0000 536.6600 0.4850 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 188.303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 941.234 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.2248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 61.8071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 304.298 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.362698 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 318.4800 0.0000 318.6200 0.4850 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 197.034 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 984.774 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 7.27183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 29.25 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 100.4400 0.0000 100.5800 0.4850 ;
    END
  END io_in[0]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.2006 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 165.606 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 260.0600 2889.1750 260.2000 2889.6600 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 29.6039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 147.676 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 740.3000 2889.1750 740.4400 2889.6600 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.7976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 234.528 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1220.0800 2889.1750 1220.2200 2889.6600 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1554 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.616 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 66.5418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 355.36 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1699.8600 2889.1750 1700.0000 2889.6600 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.566 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2180.1000 2889.1750 2180.2400 2889.6600 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 94.0331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 469.703 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2659.8800 2889.1750 2660.0200 2889.6600 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 112.277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 560.868 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 3140.1200 2889.1750 3140.2600 2889.6600 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.1364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 2695.7100 3390.2000 2696.0100 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0282 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 2384.6100 3390.2000 2384.9100 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 2072.9000 3390.2000 2073.2000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.2942 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1761.8000 3390.2000 1762.1000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.52 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1450.0900 3390.2000 1450.3900 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 176.171 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 940.984 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1138.3800 3390.2000 1138.6800 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.912 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 827.2800 3390.2000 827.5800 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.3692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 515.5700 3390.2000 515.8700 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 204.4700 3390.2000 204.7700 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 127.576 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 637.364 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 3227.0600 0.0000 3227.2000 0.4850 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 54.7997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 273.655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 3009.0200 0.0000 3009.1600 0.4850 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.876 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.4188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2790.9800 0.0000 2791.1200 0.4850 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.4335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2572.9400 0.0000 2573.0800 0.4850 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.146 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2354.4400 0.0000 2354.5800 0.4850 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 55.1411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 275.243 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2136.4000 0.0000 2136.5400 0.4850 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.937 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1918.3600 0.0000 1918.5000 0.4850 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.3855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1700.3200 0.0000 1700.4600 0.4850 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4464 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 120.385 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 642.992 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1481.8200 0.0000 1481.9600 0.4850 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3955 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1263.7800 0.0000 1263.9200 0.4850 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.0723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.1355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1045.7400 0.0000 1045.8800 0.4850 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 827.2400 0.0000 827.3800 0.4850 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.8275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.7935 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 609.2000 0.0000 609.3400 0.4850 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.1437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.5418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 275.36 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 391.1600 0.0000 391.3000 0.4850 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 199.713 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 998.284 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.1828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 173.1200 0.0000 173.2600 0.4850 ;
    END
  END io_out[0]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.1029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 170.118 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 420.1400 2889.1750 420.2800 2889.6600 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 189.378 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 899.9200 2889.1750 900.0600 2889.6600 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.8176 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 243.691 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1380.1600 2889.1750 1380.3000 2889.6600 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.7054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.13 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1859.9400 2889.1750 1860.0800 2889.6600 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 80.2784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 400.995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2340.1800 2889.1750 2340.3200 2889.6600 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 72.9524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 364.483 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.8996 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.072 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2819.9600 2889.1750 2820.1000 2889.6600 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 130.847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 653.604 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 3299.7400 2889.1750 3299.8800 2889.6600 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.6632 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 2799.4100 3390.2000 2799.7100 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3772 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 2488.3100 3390.2000 2488.6100 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.2452 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 2176.6000 3390.2000 2176.9000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.6712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1865.5000 3390.2000 1865.8000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.1452 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1553.7900 3390.2000 1554.0900 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.1892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 1242.6900 3390.2000 1242.9900 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.54 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 930.9800 3390.2000 931.2800 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.0602 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 619.2700 3390.2000 619.5700 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.9372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.464 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 3389.4000 308.1700 3390.2000 308.4700 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 91.8744 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 458.857 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 3299.7400 0.0000 3299.8800 0.4850 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 127.04 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 634.683 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 3081.7000 0.0000 3081.8400 0.4850 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 81.5594 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 407.4 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2863.6600 0.0000 2863.8000 0.4850 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.0348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 294.777 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 83.9946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 448.912 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2645.6200 0.0000 2645.7600 0.4850 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.763 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2427.1200 0.0000 2427.2600 0.4850 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 268.555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2209.0800 0.0000 2209.2200 0.4850 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.6144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1991.0400 0.0000 1991.1800 0.4850 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.742 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1773.0000 0.0000 1773.1400 0.4850 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.8607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.9595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1554.5000 0.0000 1554.6400 0.4850 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4884 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.281 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 58.3548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 311.696 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1336.4600 0.0000 1336.6000 0.4850 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1118.4200 0.0000 1118.5600 0.4850 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.6815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.0635 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 900.3800 0.0000 900.5200 0.4850 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 57.6389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 287.85 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 681.8800 0.0000 682.0200 0.4850 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.704 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 463.8400 0.0000 463.9800 0.4850 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 403.086 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2015.21 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 245.8000 0.0000 245.9400 0.4850 ;
    END
  END io_oeb[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 28.604 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.46 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 100.7700 0.8000 101.0700 ;
    END
  END user_clock2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.0000 2.0000 3388.2000 5.0000 ;
        RECT 2.0000 2884.6600 3388.2000 2887.6600 ;
        RECT 2.0000 12.3400 5.0000 12.8200 ;
        RECT 2.0000 23.2200 5.0000 23.7000 ;
        RECT 2.0000 17.7800 5.0000 18.2600 ;
        RECT 2.0000 39.5400 5.0000 40.0200 ;
        RECT 2.0000 34.1000 5.0000 34.5800 ;
        RECT 2.0000 28.6600 5.0000 29.1400 ;
        RECT 2.0000 50.4200 5.0000 50.9000 ;
        RECT 2.0000 44.9800 5.0000 45.4600 ;
        RECT 2.0000 66.7400 5.0000 67.2200 ;
        RECT 2.0000 61.3000 5.0000 61.7800 ;
        RECT 2.0000 55.8600 5.0000 56.3400 ;
        RECT 2.0000 93.9400 5.0000 94.4200 ;
        RECT 2.0000 77.6200 5.0000 78.1000 ;
        RECT 2.0000 72.1800 5.0000 72.6600 ;
        RECT 2.0000 88.5000 5.0000 88.9800 ;
        RECT 2.0000 83.0600 5.0000 83.5400 ;
        RECT 2.0000 104.8200 5.0000 105.3000 ;
        RECT 2.0000 99.3800 5.0000 99.8600 ;
        RECT 2.0000 115.7000 5.0000 116.1800 ;
        RECT 2.0000 110.2600 5.0000 110.7400 ;
        RECT 2.0000 132.0200 5.0000 132.5000 ;
        RECT 2.0000 126.5800 5.0000 127.0600 ;
        RECT 2.0000 121.1400 5.0000 121.6200 ;
        RECT 2.0000 142.9000 5.0000 143.3800 ;
        RECT 2.0000 137.4600 5.0000 137.9400 ;
        RECT 2.0000 159.2200 5.0000 159.7000 ;
        RECT 2.0000 153.7800 5.0000 154.2600 ;
        RECT 2.0000 148.3400 5.0000 148.8200 ;
        RECT 2.0000 170.1000 5.0000 170.5800 ;
        RECT 2.0000 164.6600 5.0000 165.1400 ;
        RECT 2.0000 186.4200 5.0000 186.9000 ;
        RECT 2.0000 180.9800 5.0000 181.4600 ;
        RECT 2.0000 175.5400 5.0000 176.0200 ;
        RECT 2.0000 197.3000 5.0000 197.7800 ;
        RECT 2.0000 191.8600 5.0000 192.3400 ;
        RECT 2.0000 208.1800 5.0000 208.6600 ;
        RECT 2.0000 202.7400 5.0000 203.2200 ;
        RECT 2.0000 224.5000 5.0000 224.9800 ;
        RECT 2.0000 219.0600 5.0000 219.5400 ;
        RECT 2.0000 213.6200 5.0000 214.1000 ;
        RECT 2.0000 235.3800 5.0000 235.8600 ;
        RECT 2.0000 229.9400 5.0000 230.4200 ;
        RECT 2.0000 251.7000 5.0000 252.1800 ;
        RECT 2.0000 246.2600 5.0000 246.7400 ;
        RECT 2.0000 240.8200 5.0000 241.3000 ;
        RECT 2.0000 262.5800 5.0000 263.0600 ;
        RECT 2.0000 257.1400 5.0000 257.6200 ;
        RECT 2.0000 278.9000 5.0000 279.3800 ;
        RECT 2.0000 273.4600 5.0000 273.9400 ;
        RECT 2.0000 268.0200 5.0000 268.5000 ;
        RECT 2.0000 289.7800 5.0000 290.2600 ;
        RECT 2.0000 284.3400 5.0000 284.8200 ;
        RECT 2.0000 300.6600 5.0000 301.1400 ;
        RECT 2.0000 295.2200 5.0000 295.7000 ;
        RECT 2.0000 316.9800 5.0000 317.4600 ;
        RECT 2.0000 311.5400 5.0000 312.0200 ;
        RECT 2.0000 306.1000 5.0000 306.5800 ;
        RECT 2.0000 327.8600 5.0000 328.3400 ;
        RECT 2.0000 322.4200 5.0000 322.9000 ;
        RECT 2.0000 344.1800 5.0000 344.6600 ;
        RECT 2.0000 338.7400 5.0000 339.2200 ;
        RECT 2.0000 333.3000 5.0000 333.7800 ;
        RECT 2.0000 355.0600 5.0000 355.5400 ;
        RECT 2.0000 349.6200 5.0000 350.1000 ;
        RECT 2.0000 371.3800 5.0000 371.8600 ;
        RECT 2.0000 365.9400 5.0000 366.4200 ;
        RECT 2.0000 360.5000 5.0000 360.9800 ;
        RECT 2.0000 382.2600 5.0000 382.7400 ;
        RECT 2.0000 376.8200 5.0000 377.3000 ;
        RECT 2.0000 491.0600 5.0000 491.5400 ;
        RECT 2.0000 398.5800 5.0000 399.0600 ;
        RECT 2.0000 393.1400 5.0000 393.6200 ;
        RECT 2.0000 387.7000 5.0000 388.1800 ;
        RECT 2.0000 409.4600 5.0000 409.9400 ;
        RECT 2.0000 404.0200 5.0000 404.5000 ;
        RECT 2.0000 420.3400 5.0000 420.8200 ;
        RECT 2.0000 414.9000 5.0000 415.3800 ;
        RECT 2.0000 436.6600 5.0000 437.1400 ;
        RECT 2.0000 431.2200 5.0000 431.7000 ;
        RECT 2.0000 425.7800 5.0000 426.2600 ;
        RECT 2.0000 447.5400 5.0000 448.0200 ;
        RECT 2.0000 442.1000 5.0000 442.5800 ;
        RECT 2.0000 463.8600 5.0000 464.3400 ;
        RECT 2.0000 458.4200 5.0000 458.9000 ;
        RECT 2.0000 452.9800 5.0000 453.4600 ;
        RECT 2.0000 474.7400 5.0000 475.2200 ;
        RECT 2.0000 469.3000 5.0000 469.7800 ;
        RECT 2.0000 485.6200 5.0000 486.1000 ;
        RECT 2.0000 480.1800 5.0000 480.6600 ;
        RECT 2.0000 501.9400 5.0000 502.4200 ;
        RECT 2.0000 496.5000 5.0000 496.9800 ;
        RECT 2.0000 512.8200 5.0000 513.3000 ;
        RECT 2.0000 507.3800 5.0000 507.8600 ;
        RECT 2.0000 529.1400 5.0000 529.6200 ;
        RECT 2.0000 523.7000 5.0000 524.1800 ;
        RECT 2.0000 518.2600 5.0000 518.7400 ;
        RECT 2.0000 540.0200 5.0000 540.5000 ;
        RECT 2.0000 534.5800 5.0000 535.0600 ;
        RECT 2.0000 556.3400 5.0000 556.8200 ;
        RECT 2.0000 550.9000 5.0000 551.3800 ;
        RECT 2.0000 545.4600 5.0000 545.9400 ;
        RECT 2.0000 567.2200 5.0000 567.7000 ;
        RECT 2.0000 561.7800 5.0000 562.2600 ;
        RECT 2.0000 583.5400 5.0000 584.0200 ;
        RECT 2.0000 578.1000 5.0000 578.5800 ;
        RECT 2.0000 572.6600 5.0000 573.1400 ;
        RECT 2.0000 594.4200 5.0000 594.9000 ;
        RECT 2.0000 588.9800 5.0000 589.4600 ;
        RECT 2.0000 703.2200 5.0000 703.7000 ;
        RECT 2.0000 605.3000 5.0000 605.7800 ;
        RECT 2.0000 599.8600 5.0000 600.3400 ;
        RECT 2.0000 621.6200 5.0000 622.1000 ;
        RECT 2.0000 616.1800 5.0000 616.6600 ;
        RECT 2.0000 610.7400 5.0000 611.2200 ;
        RECT 2.0000 632.5000 5.0000 632.9800 ;
        RECT 2.0000 627.0600 5.0000 627.5400 ;
        RECT 2.0000 648.8200 5.0000 649.3000 ;
        RECT 2.0000 643.3800 5.0000 643.8600 ;
        RECT 2.0000 637.9400 5.0000 638.4200 ;
        RECT 2.0000 659.7000 5.0000 660.1800 ;
        RECT 2.0000 654.2600 5.0000 654.7400 ;
        RECT 2.0000 676.0200 5.0000 676.5000 ;
        RECT 2.0000 670.5800 5.0000 671.0600 ;
        RECT 2.0000 665.1400 5.0000 665.6200 ;
        RECT 2.0000 686.9000 5.0000 687.3800 ;
        RECT 2.0000 681.4600 5.0000 681.9400 ;
        RECT 2.0000 697.7800 5.0000 698.2600 ;
        RECT 2.0000 692.3400 5.0000 692.8200 ;
        RECT 2.0000 714.1000 5.0000 714.5800 ;
        RECT 2.0000 708.6600 5.0000 709.1400 ;
        RECT 2.0000 724.9800 5.0000 725.4600 ;
        RECT 2.0000 719.5400 5.0000 720.0200 ;
        RECT 2.0000 741.3000 5.0000 741.7800 ;
        RECT 2.0000 735.8600 5.0000 736.3400 ;
        RECT 2.0000 730.4200 5.0000 730.9000 ;
        RECT 2.0000 752.1800 5.0000 752.6600 ;
        RECT 2.0000 746.7400 5.0000 747.2200 ;
        RECT 2.0000 768.5000 5.0000 768.9800 ;
        RECT 2.0000 763.0600 5.0000 763.5400 ;
        RECT 2.0000 757.6200 5.0000 758.1000 ;
        RECT 2.0000 779.3800 5.0000 779.8600 ;
        RECT 2.0000 773.9400 5.0000 774.4200 ;
        RECT 2.0000 795.7000 5.0000 796.1800 ;
        RECT 2.0000 790.2600 5.0000 790.7400 ;
        RECT 2.0000 784.8200 5.0000 785.3000 ;
        RECT 2.0000 806.5800 5.0000 807.0600 ;
        RECT 2.0000 801.1400 5.0000 801.6200 ;
        RECT 2.0000 817.4600 5.0000 817.9400 ;
        RECT 2.0000 812.0200 5.0000 812.5000 ;
        RECT 2.0000 833.7800 5.0000 834.2600 ;
        RECT 2.0000 828.3400 5.0000 828.8200 ;
        RECT 2.0000 822.9000 5.0000 823.3800 ;
        RECT 2.0000 844.6600 5.0000 845.1400 ;
        RECT 2.0000 839.2200 5.0000 839.7000 ;
        RECT 2.0000 860.9800 5.0000 861.4600 ;
        RECT 2.0000 855.5400 5.0000 856.0200 ;
        RECT 2.0000 850.1000 5.0000 850.5800 ;
        RECT 2.0000 888.1800 5.0000 888.6600 ;
        RECT 2.0000 871.8600 5.0000 872.3400 ;
        RECT 2.0000 866.4200 5.0000 866.9000 ;
        RECT 2.0000 882.7400 5.0000 883.2200 ;
        RECT 2.0000 877.3000 5.0000 877.7800 ;
        RECT 2.0000 899.0600 5.0000 899.5400 ;
        RECT 2.0000 893.6200 5.0000 894.1000 ;
        RECT 2.0000 909.9400 5.0000 910.4200 ;
        RECT 2.0000 904.5000 5.0000 904.9800 ;
        RECT 2.0000 926.2600 5.0000 926.7400 ;
        RECT 2.0000 920.8200 5.0000 921.3000 ;
        RECT 2.0000 915.3800 5.0000 915.8600 ;
        RECT 2.0000 937.1400 5.0000 937.6200 ;
        RECT 2.0000 931.7000 5.0000 932.1800 ;
        RECT 2.0000 953.4600 5.0000 953.9400 ;
        RECT 2.0000 948.0200 5.0000 948.5000 ;
        RECT 2.0000 942.5800 5.0000 943.0600 ;
        RECT 2.0000 964.3400 5.0000 964.8200 ;
        RECT 2.0000 958.9000 5.0000 959.3800 ;
        RECT 2.0000 980.6600 5.0000 981.1400 ;
        RECT 2.0000 975.2200 5.0000 975.7000 ;
        RECT 2.0000 969.7800 5.0000 970.2600 ;
        RECT 2.0000 991.5400 5.0000 992.0200 ;
        RECT 2.0000 986.1000 5.0000 986.5800 ;
        RECT 2.0000 1002.4200 5.0000 1002.9000 ;
        RECT 2.0000 996.9800 5.0000 997.4600 ;
        RECT 2.0000 1018.7400 5.0000 1019.2200 ;
        RECT 2.0000 1013.3000 5.0000 1013.7800 ;
        RECT 2.0000 1007.8600 5.0000 1008.3400 ;
        RECT 2.0000 1029.6200 5.0000 1030.1000 ;
        RECT 2.0000 1024.1800 5.0000 1024.6600 ;
        RECT 2.0000 1045.9400 5.0000 1046.4200 ;
        RECT 2.0000 1040.5000 5.0000 1040.9800 ;
        RECT 2.0000 1035.0600 5.0000 1035.5400 ;
        RECT 2.0000 1056.8200 5.0000 1057.3000 ;
        RECT 2.0000 1051.3800 5.0000 1051.8600 ;
        RECT 2.0000 1073.1400 5.0000 1073.6200 ;
        RECT 2.0000 1067.7000 5.0000 1068.1800 ;
        RECT 2.0000 1062.2600 5.0000 1062.7400 ;
        RECT 2.0000 1100.3400 5.0000 1100.8200 ;
        RECT 2.0000 1084.0200 5.0000 1084.5000 ;
        RECT 2.0000 1078.5800 5.0000 1079.0600 ;
        RECT 2.0000 1094.9000 5.0000 1095.3800 ;
        RECT 2.0000 1089.4600 5.0000 1089.9400 ;
        RECT 2.0000 1111.2200 5.0000 1111.7000 ;
        RECT 2.0000 1105.7800 5.0000 1106.2600 ;
        RECT 2.0000 1122.1000 5.0000 1122.5800 ;
        RECT 2.0000 1116.6600 5.0000 1117.1400 ;
        RECT 2.0000 1138.4200 5.0000 1138.9000 ;
        RECT 2.0000 1132.9800 5.0000 1133.4600 ;
        RECT 2.0000 1127.5400 5.0000 1128.0200 ;
        RECT 2.0000 1149.3000 5.0000 1149.7800 ;
        RECT 2.0000 1143.8600 5.0000 1144.3400 ;
        RECT 2.0000 1165.6200 5.0000 1166.1000 ;
        RECT 2.0000 1160.1800 5.0000 1160.6600 ;
        RECT 2.0000 1154.7400 5.0000 1155.2200 ;
        RECT 2.0000 1176.5000 5.0000 1176.9800 ;
        RECT 2.0000 1171.0600 5.0000 1171.5400 ;
        RECT 2.0000 1192.8200 5.0000 1193.3000 ;
        RECT 2.0000 1187.3800 5.0000 1187.8600 ;
        RECT 2.0000 1181.9400 5.0000 1182.4200 ;
        RECT 2.0000 1203.7000 5.0000 1204.1800 ;
        RECT 2.0000 1198.2600 5.0000 1198.7400 ;
        RECT 2.0000 1214.5800 5.0000 1215.0600 ;
        RECT 2.0000 1209.1400 5.0000 1209.6200 ;
        RECT 2.0000 1230.9000 5.0000 1231.3800 ;
        RECT 2.0000 1225.4600 5.0000 1225.9400 ;
        RECT 2.0000 1220.0200 5.0000 1220.5000 ;
        RECT 2.0000 1241.7800 5.0000 1242.2600 ;
        RECT 2.0000 1236.3400 5.0000 1236.8200 ;
        RECT 2.0000 1258.1000 5.0000 1258.5800 ;
        RECT 2.0000 1252.6600 5.0000 1253.1400 ;
        RECT 2.0000 1247.2200 5.0000 1247.7000 ;
        RECT 2.0000 1268.9800 5.0000 1269.4600 ;
        RECT 2.0000 1263.5400 5.0000 1264.0200 ;
        RECT 2.0000 1285.3000 5.0000 1285.7800 ;
        RECT 2.0000 1279.8600 5.0000 1280.3400 ;
        RECT 2.0000 1274.4200 5.0000 1274.9000 ;
        RECT 2.0000 1296.1800 5.0000 1296.6600 ;
        RECT 2.0000 1290.7400 5.0000 1291.2200 ;
        RECT 2.0000 1307.0600 5.0000 1307.5400 ;
        RECT 2.0000 1301.6200 5.0000 1302.1000 ;
        RECT 2.0000 1323.3800 5.0000 1323.8600 ;
        RECT 2.0000 1317.9400 5.0000 1318.4200 ;
        RECT 2.0000 1312.5000 5.0000 1312.9800 ;
        RECT 2.0000 1334.2600 5.0000 1334.7400 ;
        RECT 2.0000 1328.8200 5.0000 1329.3000 ;
        RECT 2.0000 1350.5800 5.0000 1351.0600 ;
        RECT 2.0000 1345.1400 5.0000 1345.6200 ;
        RECT 2.0000 1339.7000 5.0000 1340.1800 ;
        RECT 2.0000 1361.4600 5.0000 1361.9400 ;
        RECT 2.0000 1356.0200 5.0000 1356.5000 ;
        RECT 2.0000 1377.7800 5.0000 1378.2600 ;
        RECT 2.0000 1372.3400 5.0000 1372.8200 ;
        RECT 2.0000 1366.9000 5.0000 1367.3800 ;
        RECT 2.0000 1388.6600 5.0000 1389.1400 ;
        RECT 2.0000 1383.2200 5.0000 1383.7000 ;
        RECT 2.0000 1404.9800 5.0000 1405.4600 ;
        RECT 2.0000 1399.5400 5.0000 1400.0200 ;
        RECT 2.0000 1394.1000 5.0000 1394.5800 ;
        RECT 2.0000 1415.8600 5.0000 1416.3400 ;
        RECT 2.0000 1410.4200 5.0000 1410.9000 ;
        RECT 2.0000 1426.7400 5.0000 1427.2200 ;
        RECT 2.0000 1421.3000 5.0000 1421.7800 ;
        RECT 2.0000 1443.0600 5.0000 1443.5400 ;
        RECT 2.0000 1437.6200 5.0000 1438.1000 ;
        RECT 2.0000 1432.1800 5.0000 1432.6600 ;
        RECT 3385.2000 12.3400 3388.2000 12.8200 ;
        RECT 3385.2000 23.2200 3388.2000 23.7000 ;
        RECT 3385.2000 17.7800 3388.2000 18.2600 ;
        RECT 3385.2000 39.5400 3388.2000 40.0200 ;
        RECT 3385.2000 34.1000 3388.2000 34.5800 ;
        RECT 3385.2000 28.6600 3388.2000 29.1400 ;
        RECT 3385.2000 50.4200 3388.2000 50.9000 ;
        RECT 3385.2000 44.9800 3388.2000 45.4600 ;
        RECT 3385.2000 66.7400 3388.2000 67.2200 ;
        RECT 3385.2000 61.3000 3388.2000 61.7800 ;
        RECT 3385.2000 55.8600 3388.2000 56.3400 ;
        RECT 3385.2000 93.9400 3388.2000 94.4200 ;
        RECT 3385.2000 77.6200 3388.2000 78.1000 ;
        RECT 3385.2000 72.1800 3388.2000 72.6600 ;
        RECT 3385.2000 88.5000 3388.2000 88.9800 ;
        RECT 3385.2000 83.0600 3388.2000 83.5400 ;
        RECT 3385.2000 104.8200 3388.2000 105.3000 ;
        RECT 3385.2000 99.3800 3388.2000 99.8600 ;
        RECT 3385.2000 115.7000 3388.2000 116.1800 ;
        RECT 3385.2000 110.2600 3388.2000 110.7400 ;
        RECT 3385.2000 132.0200 3388.2000 132.5000 ;
        RECT 3385.2000 126.5800 3388.2000 127.0600 ;
        RECT 3385.2000 121.1400 3388.2000 121.6200 ;
        RECT 3385.2000 142.9000 3388.2000 143.3800 ;
        RECT 3385.2000 137.4600 3388.2000 137.9400 ;
        RECT 3385.2000 159.2200 3388.2000 159.7000 ;
        RECT 3385.2000 153.7800 3388.2000 154.2600 ;
        RECT 3385.2000 148.3400 3388.2000 148.8200 ;
        RECT 3385.2000 170.1000 3388.2000 170.5800 ;
        RECT 3385.2000 164.6600 3388.2000 165.1400 ;
        RECT 3385.2000 186.4200 3388.2000 186.9000 ;
        RECT 3385.2000 180.9800 3388.2000 181.4600 ;
        RECT 3385.2000 175.5400 3388.2000 176.0200 ;
        RECT 3385.2000 197.3000 3388.2000 197.7800 ;
        RECT 3385.2000 191.8600 3388.2000 192.3400 ;
        RECT 3385.2000 208.1800 3388.2000 208.6600 ;
        RECT 3385.2000 202.7400 3388.2000 203.2200 ;
        RECT 3385.2000 224.5000 3388.2000 224.9800 ;
        RECT 3385.2000 219.0600 3388.2000 219.5400 ;
        RECT 3385.2000 213.6200 3388.2000 214.1000 ;
        RECT 3385.2000 235.3800 3388.2000 235.8600 ;
        RECT 3385.2000 229.9400 3388.2000 230.4200 ;
        RECT 3385.2000 251.7000 3388.2000 252.1800 ;
        RECT 3385.2000 246.2600 3388.2000 246.7400 ;
        RECT 3385.2000 240.8200 3388.2000 241.3000 ;
        RECT 3385.2000 262.5800 3388.2000 263.0600 ;
        RECT 3385.2000 257.1400 3388.2000 257.6200 ;
        RECT 3385.2000 278.9000 3388.2000 279.3800 ;
        RECT 3385.2000 273.4600 3388.2000 273.9400 ;
        RECT 3385.2000 268.0200 3388.2000 268.5000 ;
        RECT 3385.2000 289.7800 3388.2000 290.2600 ;
        RECT 3385.2000 284.3400 3388.2000 284.8200 ;
        RECT 3385.2000 300.6600 3388.2000 301.1400 ;
        RECT 3385.2000 295.2200 3388.2000 295.7000 ;
        RECT 3385.2000 316.9800 3388.2000 317.4600 ;
        RECT 3385.2000 311.5400 3388.2000 312.0200 ;
        RECT 3385.2000 306.1000 3388.2000 306.5800 ;
        RECT 3385.2000 327.8600 3388.2000 328.3400 ;
        RECT 3385.2000 322.4200 3388.2000 322.9000 ;
        RECT 3385.2000 344.1800 3388.2000 344.6600 ;
        RECT 3385.2000 338.7400 3388.2000 339.2200 ;
        RECT 3385.2000 333.3000 3388.2000 333.7800 ;
        RECT 3385.2000 355.0600 3388.2000 355.5400 ;
        RECT 3385.2000 349.6200 3388.2000 350.1000 ;
        RECT 3385.2000 371.3800 3388.2000 371.8600 ;
        RECT 3385.2000 365.9400 3388.2000 366.4200 ;
        RECT 3385.2000 360.5000 3388.2000 360.9800 ;
        RECT 3385.2000 382.2600 3388.2000 382.7400 ;
        RECT 3385.2000 376.8200 3388.2000 377.3000 ;
        RECT 3385.2000 491.0600 3388.2000 491.5400 ;
        RECT 3385.2000 398.5800 3388.2000 399.0600 ;
        RECT 3385.2000 393.1400 3388.2000 393.6200 ;
        RECT 3385.2000 387.7000 3388.2000 388.1800 ;
        RECT 3385.2000 409.4600 3388.2000 409.9400 ;
        RECT 3385.2000 404.0200 3388.2000 404.5000 ;
        RECT 3385.2000 420.3400 3388.2000 420.8200 ;
        RECT 3385.2000 414.9000 3388.2000 415.3800 ;
        RECT 3385.2000 436.6600 3388.2000 437.1400 ;
        RECT 3385.2000 431.2200 3388.2000 431.7000 ;
        RECT 3385.2000 425.7800 3388.2000 426.2600 ;
        RECT 3385.2000 447.5400 3388.2000 448.0200 ;
        RECT 3385.2000 442.1000 3388.2000 442.5800 ;
        RECT 3385.2000 463.8600 3388.2000 464.3400 ;
        RECT 3385.2000 458.4200 3388.2000 458.9000 ;
        RECT 3385.2000 452.9800 3388.2000 453.4600 ;
        RECT 3385.2000 474.7400 3388.2000 475.2200 ;
        RECT 3385.2000 469.3000 3388.2000 469.7800 ;
        RECT 3385.2000 485.6200 3388.2000 486.1000 ;
        RECT 3385.2000 480.1800 3388.2000 480.6600 ;
        RECT 3385.2000 501.9400 3388.2000 502.4200 ;
        RECT 3385.2000 496.5000 3388.2000 496.9800 ;
        RECT 3385.2000 512.8200 3388.2000 513.3000 ;
        RECT 3385.2000 507.3800 3388.2000 507.8600 ;
        RECT 3385.2000 529.1400 3388.2000 529.6200 ;
        RECT 3385.2000 523.7000 3388.2000 524.1800 ;
        RECT 3385.2000 518.2600 3388.2000 518.7400 ;
        RECT 3385.2000 540.0200 3388.2000 540.5000 ;
        RECT 3385.2000 534.5800 3388.2000 535.0600 ;
        RECT 3385.2000 556.3400 3388.2000 556.8200 ;
        RECT 3385.2000 550.9000 3388.2000 551.3800 ;
        RECT 3385.2000 545.4600 3388.2000 545.9400 ;
        RECT 3385.2000 567.2200 3388.2000 567.7000 ;
        RECT 3385.2000 561.7800 3388.2000 562.2600 ;
        RECT 3385.2000 583.5400 3388.2000 584.0200 ;
        RECT 3385.2000 578.1000 3388.2000 578.5800 ;
        RECT 3385.2000 572.6600 3388.2000 573.1400 ;
        RECT 3385.2000 594.4200 3388.2000 594.9000 ;
        RECT 3385.2000 588.9800 3388.2000 589.4600 ;
        RECT 3385.2000 703.2200 3388.2000 703.7000 ;
        RECT 3385.2000 605.3000 3388.2000 605.7800 ;
        RECT 3385.2000 599.8600 3388.2000 600.3400 ;
        RECT 3385.2000 621.6200 3388.2000 622.1000 ;
        RECT 3385.2000 616.1800 3388.2000 616.6600 ;
        RECT 3385.2000 610.7400 3388.2000 611.2200 ;
        RECT 3385.2000 632.5000 3388.2000 632.9800 ;
        RECT 3385.2000 627.0600 3388.2000 627.5400 ;
        RECT 3385.2000 648.8200 3388.2000 649.3000 ;
        RECT 3385.2000 643.3800 3388.2000 643.8600 ;
        RECT 3385.2000 637.9400 3388.2000 638.4200 ;
        RECT 3385.2000 659.7000 3388.2000 660.1800 ;
        RECT 3385.2000 654.2600 3388.2000 654.7400 ;
        RECT 3385.2000 676.0200 3388.2000 676.5000 ;
        RECT 3385.2000 670.5800 3388.2000 671.0600 ;
        RECT 3385.2000 665.1400 3388.2000 665.6200 ;
        RECT 3385.2000 686.9000 3388.2000 687.3800 ;
        RECT 3385.2000 681.4600 3388.2000 681.9400 ;
        RECT 3385.2000 697.7800 3388.2000 698.2600 ;
        RECT 3385.2000 692.3400 3388.2000 692.8200 ;
        RECT 3385.2000 714.1000 3388.2000 714.5800 ;
        RECT 3385.2000 708.6600 3388.2000 709.1400 ;
        RECT 3385.2000 724.9800 3388.2000 725.4600 ;
        RECT 3385.2000 719.5400 3388.2000 720.0200 ;
        RECT 3385.2000 741.3000 3388.2000 741.7800 ;
        RECT 3385.2000 735.8600 3388.2000 736.3400 ;
        RECT 3385.2000 730.4200 3388.2000 730.9000 ;
        RECT 3385.2000 752.1800 3388.2000 752.6600 ;
        RECT 3385.2000 746.7400 3388.2000 747.2200 ;
        RECT 3385.2000 768.5000 3388.2000 768.9800 ;
        RECT 3385.2000 763.0600 3388.2000 763.5400 ;
        RECT 3385.2000 757.6200 3388.2000 758.1000 ;
        RECT 3385.2000 779.3800 3388.2000 779.8600 ;
        RECT 3385.2000 773.9400 3388.2000 774.4200 ;
        RECT 3385.2000 795.7000 3388.2000 796.1800 ;
        RECT 3385.2000 790.2600 3388.2000 790.7400 ;
        RECT 3385.2000 784.8200 3388.2000 785.3000 ;
        RECT 3385.2000 806.5800 3388.2000 807.0600 ;
        RECT 3385.2000 801.1400 3388.2000 801.6200 ;
        RECT 3385.2000 817.4600 3388.2000 817.9400 ;
        RECT 3385.2000 812.0200 3388.2000 812.5000 ;
        RECT 3385.2000 833.7800 3388.2000 834.2600 ;
        RECT 3385.2000 828.3400 3388.2000 828.8200 ;
        RECT 3385.2000 822.9000 3388.2000 823.3800 ;
        RECT 3385.2000 844.6600 3388.2000 845.1400 ;
        RECT 3385.2000 839.2200 3388.2000 839.7000 ;
        RECT 3385.2000 860.9800 3388.2000 861.4600 ;
        RECT 3385.2000 855.5400 3388.2000 856.0200 ;
        RECT 3385.2000 850.1000 3388.2000 850.5800 ;
        RECT 3385.2000 888.1800 3388.2000 888.6600 ;
        RECT 3385.2000 871.8600 3388.2000 872.3400 ;
        RECT 3385.2000 866.4200 3388.2000 866.9000 ;
        RECT 3385.2000 882.7400 3388.2000 883.2200 ;
        RECT 3385.2000 877.3000 3388.2000 877.7800 ;
        RECT 3385.2000 899.0600 3388.2000 899.5400 ;
        RECT 3385.2000 893.6200 3388.2000 894.1000 ;
        RECT 3385.2000 909.9400 3388.2000 910.4200 ;
        RECT 3385.2000 904.5000 3388.2000 904.9800 ;
        RECT 3385.2000 926.2600 3388.2000 926.7400 ;
        RECT 3385.2000 920.8200 3388.2000 921.3000 ;
        RECT 3385.2000 915.3800 3388.2000 915.8600 ;
        RECT 3385.2000 937.1400 3388.2000 937.6200 ;
        RECT 3385.2000 931.7000 3388.2000 932.1800 ;
        RECT 3385.2000 953.4600 3388.2000 953.9400 ;
        RECT 3385.2000 948.0200 3388.2000 948.5000 ;
        RECT 3385.2000 942.5800 3388.2000 943.0600 ;
        RECT 3385.2000 964.3400 3388.2000 964.8200 ;
        RECT 3385.2000 958.9000 3388.2000 959.3800 ;
        RECT 3385.2000 980.6600 3388.2000 981.1400 ;
        RECT 3385.2000 975.2200 3388.2000 975.7000 ;
        RECT 3385.2000 969.7800 3388.2000 970.2600 ;
        RECT 3385.2000 991.5400 3388.2000 992.0200 ;
        RECT 3385.2000 986.1000 3388.2000 986.5800 ;
        RECT 3385.2000 1002.4200 3388.2000 1002.9000 ;
        RECT 3385.2000 996.9800 3388.2000 997.4600 ;
        RECT 3385.2000 1018.7400 3388.2000 1019.2200 ;
        RECT 3385.2000 1013.3000 3388.2000 1013.7800 ;
        RECT 3385.2000 1007.8600 3388.2000 1008.3400 ;
        RECT 3385.2000 1029.6200 3388.2000 1030.1000 ;
        RECT 3385.2000 1024.1800 3388.2000 1024.6600 ;
        RECT 3385.2000 1045.9400 3388.2000 1046.4200 ;
        RECT 3385.2000 1040.5000 3388.2000 1040.9800 ;
        RECT 3385.2000 1035.0600 3388.2000 1035.5400 ;
        RECT 3385.2000 1056.8200 3388.2000 1057.3000 ;
        RECT 3385.2000 1051.3800 3388.2000 1051.8600 ;
        RECT 3385.2000 1073.1400 3388.2000 1073.6200 ;
        RECT 3385.2000 1067.7000 3388.2000 1068.1800 ;
        RECT 3385.2000 1062.2600 3388.2000 1062.7400 ;
        RECT 3385.2000 1100.3400 3388.2000 1100.8200 ;
        RECT 3385.2000 1084.0200 3388.2000 1084.5000 ;
        RECT 3385.2000 1078.5800 3388.2000 1079.0600 ;
        RECT 3385.2000 1094.9000 3388.2000 1095.3800 ;
        RECT 3385.2000 1089.4600 3388.2000 1089.9400 ;
        RECT 3385.2000 1111.2200 3388.2000 1111.7000 ;
        RECT 3385.2000 1105.7800 3388.2000 1106.2600 ;
        RECT 3385.2000 1122.1000 3388.2000 1122.5800 ;
        RECT 3385.2000 1116.6600 3388.2000 1117.1400 ;
        RECT 3385.2000 1138.4200 3388.2000 1138.9000 ;
        RECT 3385.2000 1132.9800 3388.2000 1133.4600 ;
        RECT 3385.2000 1127.5400 3388.2000 1128.0200 ;
        RECT 3385.2000 1149.3000 3388.2000 1149.7800 ;
        RECT 3385.2000 1143.8600 3388.2000 1144.3400 ;
        RECT 3385.2000 1165.6200 3388.2000 1166.1000 ;
        RECT 3385.2000 1160.1800 3388.2000 1160.6600 ;
        RECT 3385.2000 1154.7400 3388.2000 1155.2200 ;
        RECT 3385.2000 1176.5000 3388.2000 1176.9800 ;
        RECT 3385.2000 1171.0600 3388.2000 1171.5400 ;
        RECT 3385.2000 1192.8200 3388.2000 1193.3000 ;
        RECT 3385.2000 1187.3800 3388.2000 1187.8600 ;
        RECT 3385.2000 1181.9400 3388.2000 1182.4200 ;
        RECT 3385.2000 1203.7000 3388.2000 1204.1800 ;
        RECT 3385.2000 1198.2600 3388.2000 1198.7400 ;
        RECT 3385.2000 1214.5800 3388.2000 1215.0600 ;
        RECT 3385.2000 1209.1400 3388.2000 1209.6200 ;
        RECT 3385.2000 1230.9000 3388.2000 1231.3800 ;
        RECT 3385.2000 1225.4600 3388.2000 1225.9400 ;
        RECT 3385.2000 1220.0200 3388.2000 1220.5000 ;
        RECT 3385.2000 1241.7800 3388.2000 1242.2600 ;
        RECT 3385.2000 1236.3400 3388.2000 1236.8200 ;
        RECT 3385.2000 1258.1000 3388.2000 1258.5800 ;
        RECT 3385.2000 1252.6600 3388.2000 1253.1400 ;
        RECT 3385.2000 1247.2200 3388.2000 1247.7000 ;
        RECT 3385.2000 1268.9800 3388.2000 1269.4600 ;
        RECT 3385.2000 1263.5400 3388.2000 1264.0200 ;
        RECT 3385.2000 1285.3000 3388.2000 1285.7800 ;
        RECT 3385.2000 1279.8600 3388.2000 1280.3400 ;
        RECT 3385.2000 1274.4200 3388.2000 1274.9000 ;
        RECT 3385.2000 1296.1800 3388.2000 1296.6600 ;
        RECT 3385.2000 1290.7400 3388.2000 1291.2200 ;
        RECT 3385.2000 1307.0600 3388.2000 1307.5400 ;
        RECT 3385.2000 1301.6200 3388.2000 1302.1000 ;
        RECT 3385.2000 1323.3800 3388.2000 1323.8600 ;
        RECT 3385.2000 1317.9400 3388.2000 1318.4200 ;
        RECT 3385.2000 1312.5000 3388.2000 1312.9800 ;
        RECT 3385.2000 1334.2600 3388.2000 1334.7400 ;
        RECT 3385.2000 1328.8200 3388.2000 1329.3000 ;
        RECT 3385.2000 1350.5800 3388.2000 1351.0600 ;
        RECT 3385.2000 1345.1400 3388.2000 1345.6200 ;
        RECT 3385.2000 1339.7000 3388.2000 1340.1800 ;
        RECT 3385.2000 1361.4600 3388.2000 1361.9400 ;
        RECT 3385.2000 1356.0200 3388.2000 1356.5000 ;
        RECT 3385.2000 1377.7800 3388.2000 1378.2600 ;
        RECT 3385.2000 1372.3400 3388.2000 1372.8200 ;
        RECT 3385.2000 1366.9000 3388.2000 1367.3800 ;
        RECT 3385.2000 1388.6600 3388.2000 1389.1400 ;
        RECT 3385.2000 1383.2200 3388.2000 1383.7000 ;
        RECT 3385.2000 1404.9800 3388.2000 1405.4600 ;
        RECT 3385.2000 1399.5400 3388.2000 1400.0200 ;
        RECT 3385.2000 1394.1000 3388.2000 1394.5800 ;
        RECT 3385.2000 1415.8600 3388.2000 1416.3400 ;
        RECT 3385.2000 1410.4200 3388.2000 1410.9000 ;
        RECT 3385.2000 1426.7400 3388.2000 1427.2200 ;
        RECT 3385.2000 1421.3000 3388.2000 1421.7800 ;
        RECT 3385.2000 1443.0600 3388.2000 1443.5400 ;
        RECT 3385.2000 1437.6200 3388.2000 1438.1000 ;
        RECT 3385.2000 1432.1800 3388.2000 1432.6600 ;
        RECT 2.0000 1497.4600 5.0000 1497.9400 ;
        RECT 2.0000 1453.9400 5.0000 1454.4200 ;
        RECT 2.0000 1448.5000 5.0000 1448.9800 ;
        RECT 2.0000 1470.2600 5.0000 1470.7400 ;
        RECT 2.0000 1464.8200 5.0000 1465.3000 ;
        RECT 2.0000 1459.3800 5.0000 1459.8600 ;
        RECT 2.0000 1481.1400 5.0000 1481.6200 ;
        RECT 2.0000 1475.7000 5.0000 1476.1800 ;
        RECT 2.0000 1492.0200 5.0000 1492.5000 ;
        RECT 2.0000 1486.5800 5.0000 1487.0600 ;
        RECT 2.0000 1508.3400 5.0000 1508.8200 ;
        RECT 2.0000 1502.9000 5.0000 1503.3800 ;
        RECT 2.0000 1519.2200 5.0000 1519.7000 ;
        RECT 2.0000 1513.7800 5.0000 1514.2600 ;
        RECT 2.0000 1535.5400 5.0000 1536.0200 ;
        RECT 2.0000 1530.1000 5.0000 1530.5800 ;
        RECT 2.0000 1524.6600 5.0000 1525.1400 ;
        RECT 2.0000 1546.4200 5.0000 1546.9000 ;
        RECT 2.0000 1540.9800 5.0000 1541.4600 ;
        RECT 2.0000 1562.7400 5.0000 1563.2200 ;
        RECT 2.0000 1557.3000 5.0000 1557.7800 ;
        RECT 2.0000 1551.8600 5.0000 1552.3400 ;
        RECT 2.0000 1573.6200 5.0000 1574.1000 ;
        RECT 2.0000 1568.1800 5.0000 1568.6600 ;
        RECT 2.0000 1589.9400 5.0000 1590.4200 ;
        RECT 2.0000 1584.5000 5.0000 1584.9800 ;
        RECT 2.0000 1579.0600 5.0000 1579.5400 ;
        RECT 2.0000 1600.8200 5.0000 1601.3000 ;
        RECT 2.0000 1595.3800 5.0000 1595.8600 ;
        RECT 2.0000 1611.7000 5.0000 1612.1800 ;
        RECT 2.0000 1606.2600 5.0000 1606.7400 ;
        RECT 2.0000 1628.0200 5.0000 1628.5000 ;
        RECT 2.0000 1622.5800 5.0000 1623.0600 ;
        RECT 2.0000 1617.1400 5.0000 1617.6200 ;
        RECT 2.0000 1638.9000 5.0000 1639.3800 ;
        RECT 2.0000 1633.4600 5.0000 1633.9400 ;
        RECT 2.0000 1655.2200 5.0000 1655.7000 ;
        RECT 2.0000 1649.7800 5.0000 1650.2600 ;
        RECT 2.0000 1644.3400 5.0000 1644.8200 ;
        RECT 2.0000 1709.6200 5.0000 1710.1000 ;
        RECT 2.0000 1666.1000 5.0000 1666.5800 ;
        RECT 2.0000 1660.6600 5.0000 1661.1400 ;
        RECT 2.0000 1682.4200 5.0000 1682.9000 ;
        RECT 2.0000 1676.9800 5.0000 1677.4600 ;
        RECT 2.0000 1671.5400 5.0000 1672.0200 ;
        RECT 2.0000 1693.3000 5.0000 1693.7800 ;
        RECT 2.0000 1687.8600 5.0000 1688.3400 ;
        RECT 2.0000 1704.1800 5.0000 1704.6600 ;
        RECT 2.0000 1698.7400 5.0000 1699.2200 ;
        RECT 2.0000 1720.5000 5.0000 1720.9800 ;
        RECT 2.0000 1715.0600 5.0000 1715.5400 ;
        RECT 2.0000 1731.3800 5.0000 1731.8600 ;
        RECT 2.0000 1725.9400 5.0000 1726.4200 ;
        RECT 2.0000 1747.7000 5.0000 1748.1800 ;
        RECT 2.0000 1742.2600 5.0000 1742.7400 ;
        RECT 2.0000 1736.8200 5.0000 1737.3000 ;
        RECT 2.0000 1758.5800 5.0000 1759.0600 ;
        RECT 2.0000 1753.1400 5.0000 1753.6200 ;
        RECT 2.0000 1774.9000 5.0000 1775.3800 ;
        RECT 2.0000 1769.4600 5.0000 1769.9400 ;
        RECT 2.0000 1764.0200 5.0000 1764.5000 ;
        RECT 2.0000 1785.7800 5.0000 1786.2600 ;
        RECT 2.0000 1780.3400 5.0000 1780.8200 ;
        RECT 2.0000 1802.1000 5.0000 1802.5800 ;
        RECT 2.0000 1796.6600 5.0000 1797.1400 ;
        RECT 2.0000 1791.2200 5.0000 1791.7000 ;
        RECT 2.0000 1812.9800 5.0000 1813.4600 ;
        RECT 2.0000 1807.5400 5.0000 1808.0200 ;
        RECT 2.0000 1823.8600 5.0000 1824.3400 ;
        RECT 2.0000 1818.4200 5.0000 1818.9000 ;
        RECT 2.0000 1840.1800 5.0000 1840.6600 ;
        RECT 2.0000 1834.7400 5.0000 1835.2200 ;
        RECT 2.0000 1829.3000 5.0000 1829.7800 ;
        RECT 2.0000 1851.0600 5.0000 1851.5400 ;
        RECT 2.0000 1845.6200 5.0000 1846.1000 ;
        RECT 2.0000 1867.3800 5.0000 1867.8600 ;
        RECT 2.0000 1861.9400 5.0000 1862.4200 ;
        RECT 2.0000 1856.5000 5.0000 1856.9800 ;
        RECT 2.0000 1878.2600 5.0000 1878.7400 ;
        RECT 2.0000 1872.8200 5.0000 1873.3000 ;
        RECT 2.0000 1894.5800 5.0000 1895.0600 ;
        RECT 2.0000 1889.1400 5.0000 1889.6200 ;
        RECT 2.0000 1883.7000 5.0000 1884.1800 ;
        RECT 2.0000 1905.4600 5.0000 1905.9400 ;
        RECT 2.0000 1900.0200 5.0000 1900.5000 ;
        RECT 2.0000 1916.3400 5.0000 1916.8200 ;
        RECT 2.0000 1910.9000 5.0000 1911.3800 ;
        RECT 2.0000 1932.6600 5.0000 1933.1400 ;
        RECT 2.0000 1927.2200 5.0000 1927.7000 ;
        RECT 2.0000 1921.7800 5.0000 1922.2600 ;
        RECT 2.0000 1943.5400 5.0000 1944.0200 ;
        RECT 2.0000 1938.1000 5.0000 1938.5800 ;
        RECT 2.0000 1959.8600 5.0000 1960.3400 ;
        RECT 2.0000 1954.4200 5.0000 1954.9000 ;
        RECT 2.0000 1948.9800 5.0000 1949.4600 ;
        RECT 2.0000 1970.7400 5.0000 1971.2200 ;
        RECT 2.0000 1965.3000 5.0000 1965.7800 ;
        RECT 2.0000 1987.0600 5.0000 1987.5400 ;
        RECT 2.0000 1981.6200 5.0000 1982.1000 ;
        RECT 2.0000 1976.1800 5.0000 1976.6600 ;
        RECT 2.0000 1997.9400 5.0000 1998.4200 ;
        RECT 2.0000 1992.5000 5.0000 1992.9800 ;
        RECT 2.0000 2014.2600 5.0000 2014.7400 ;
        RECT 2.0000 2008.8200 5.0000 2009.3000 ;
        RECT 2.0000 2003.3800 5.0000 2003.8600 ;
        RECT 2.0000 2025.1400 5.0000 2025.6200 ;
        RECT 2.0000 2019.7000 5.0000 2020.1800 ;
        RECT 2.0000 2036.0200 5.0000 2036.5000 ;
        RECT 2.0000 2030.5800 5.0000 2031.0600 ;
        RECT 2.0000 2052.3400 5.0000 2052.8200 ;
        RECT 2.0000 2046.9000 5.0000 2047.3800 ;
        RECT 2.0000 2041.4600 5.0000 2041.9400 ;
        RECT 2.0000 2063.2200 5.0000 2063.7000 ;
        RECT 2.0000 2057.7800 5.0000 2058.2600 ;
        RECT 2.0000 2079.5400 5.0000 2080.0200 ;
        RECT 2.0000 2074.1000 5.0000 2074.5800 ;
        RECT 2.0000 2068.6600 5.0000 2069.1400 ;
        RECT 2.0000 2106.7400 5.0000 2107.2200 ;
        RECT 2.0000 2090.4200 5.0000 2090.9000 ;
        RECT 2.0000 2084.9800 5.0000 2085.4600 ;
        RECT 2.0000 2101.3000 5.0000 2101.7800 ;
        RECT 2.0000 2095.8600 5.0000 2096.3400 ;
        RECT 2.0000 2117.6200 5.0000 2118.1000 ;
        RECT 2.0000 2112.1800 5.0000 2112.6600 ;
        RECT 2.0000 2128.5000 5.0000 2128.9800 ;
        RECT 2.0000 2123.0600 5.0000 2123.5400 ;
        RECT 2.0000 2144.8200 5.0000 2145.3000 ;
        RECT 2.0000 2139.3800 5.0000 2139.8600 ;
        RECT 2.0000 2133.9400 5.0000 2134.4200 ;
        RECT 2.0000 2155.7000 5.0000 2156.1800 ;
        RECT 2.0000 2150.2600 5.0000 2150.7400 ;
        RECT 2.0000 2172.0200 5.0000 2172.5000 ;
        RECT 2.0000 2166.5800 5.0000 2167.0600 ;
        RECT 2.0000 2161.1400 5.0000 2161.6200 ;
        RECT 2.0000 2182.9000 5.0000 2183.3800 ;
        RECT 2.0000 2177.4600 5.0000 2177.9400 ;
        RECT 2.0000 2199.2200 5.0000 2199.7000 ;
        RECT 2.0000 2193.7800 5.0000 2194.2600 ;
        RECT 2.0000 2188.3400 5.0000 2188.8200 ;
        RECT 2.0000 2210.1000 5.0000 2210.5800 ;
        RECT 2.0000 2204.6600 5.0000 2205.1400 ;
        RECT 2.0000 2220.9800 5.0000 2221.4600 ;
        RECT 2.0000 2215.5400 5.0000 2216.0200 ;
        RECT 2.0000 2237.3000 5.0000 2237.7800 ;
        RECT 2.0000 2231.8600 5.0000 2232.3400 ;
        RECT 2.0000 2226.4200 5.0000 2226.9000 ;
        RECT 2.0000 2248.1800 5.0000 2248.6600 ;
        RECT 2.0000 2242.7400 5.0000 2243.2200 ;
        RECT 2.0000 2264.5000 5.0000 2264.9800 ;
        RECT 2.0000 2259.0600 5.0000 2259.5400 ;
        RECT 2.0000 2253.6200 5.0000 2254.1000 ;
        RECT 2.0000 2275.3800 5.0000 2275.8600 ;
        RECT 2.0000 2269.9400 5.0000 2270.4200 ;
        RECT 2.0000 2291.7000 5.0000 2292.1800 ;
        RECT 2.0000 2286.2600 5.0000 2286.7400 ;
        RECT 2.0000 2280.8200 5.0000 2281.3000 ;
        RECT 2.0000 2716.0200 5.0000 2716.5000 ;
        RECT 2.0000 2503.8600 5.0000 2504.3400 ;
        RECT 2.0000 2302.5800 5.0000 2303.0600 ;
        RECT 2.0000 2297.1400 5.0000 2297.6200 ;
        RECT 2.0000 2313.4600 5.0000 2313.9400 ;
        RECT 2.0000 2308.0200 5.0000 2308.5000 ;
        RECT 2.0000 2329.7800 5.0000 2330.2600 ;
        RECT 2.0000 2324.3400 5.0000 2324.8200 ;
        RECT 2.0000 2318.9000 5.0000 2319.3800 ;
        RECT 2.0000 2340.6600 5.0000 2341.1400 ;
        RECT 2.0000 2335.2200 5.0000 2335.7000 ;
        RECT 2.0000 2356.9800 5.0000 2357.4600 ;
        RECT 2.0000 2351.5400 5.0000 2352.0200 ;
        RECT 2.0000 2346.1000 5.0000 2346.5800 ;
        RECT 2.0000 2367.8600 5.0000 2368.3400 ;
        RECT 2.0000 2362.4200 5.0000 2362.9000 ;
        RECT 2.0000 2384.1800 5.0000 2384.6600 ;
        RECT 2.0000 2378.7400 5.0000 2379.2200 ;
        RECT 2.0000 2373.3000 5.0000 2373.7800 ;
        RECT 2.0000 2395.0600 5.0000 2395.5400 ;
        RECT 2.0000 2389.6200 5.0000 2390.1000 ;
        RECT 2.0000 2411.3800 5.0000 2411.8600 ;
        RECT 2.0000 2405.9400 5.0000 2406.4200 ;
        RECT 2.0000 2400.5000 5.0000 2400.9800 ;
        RECT 2.0000 2422.2600 5.0000 2422.7400 ;
        RECT 2.0000 2416.8200 5.0000 2417.3000 ;
        RECT 2.0000 2433.1400 5.0000 2433.6200 ;
        RECT 2.0000 2427.7000 5.0000 2428.1800 ;
        RECT 2.0000 2449.4600 5.0000 2449.9400 ;
        RECT 2.0000 2444.0200 5.0000 2444.5000 ;
        RECT 2.0000 2438.5800 5.0000 2439.0600 ;
        RECT 2.0000 2460.3400 5.0000 2460.8200 ;
        RECT 2.0000 2454.9000 5.0000 2455.3800 ;
        RECT 2.0000 2476.6600 5.0000 2477.1400 ;
        RECT 2.0000 2471.2200 5.0000 2471.7000 ;
        RECT 2.0000 2465.7800 5.0000 2466.2600 ;
        RECT 2.0000 2487.5400 5.0000 2488.0200 ;
        RECT 2.0000 2482.1000 5.0000 2482.5800 ;
        RECT 2.0000 2498.4200 5.0000 2498.9000 ;
        RECT 2.0000 2492.9800 5.0000 2493.4600 ;
        RECT 2.0000 2514.7400 5.0000 2515.2200 ;
        RECT 2.0000 2509.3000 5.0000 2509.7800 ;
        RECT 2.0000 2525.6200 5.0000 2526.1000 ;
        RECT 2.0000 2520.1800 5.0000 2520.6600 ;
        RECT 2.0000 2541.9400 5.0000 2542.4200 ;
        RECT 2.0000 2536.5000 5.0000 2536.9800 ;
        RECT 2.0000 2531.0600 5.0000 2531.5400 ;
        RECT 2.0000 2552.8200 5.0000 2553.3000 ;
        RECT 2.0000 2547.3800 5.0000 2547.8600 ;
        RECT 2.0000 2569.1400 5.0000 2569.6200 ;
        RECT 2.0000 2563.7000 5.0000 2564.1800 ;
        RECT 2.0000 2558.2600 5.0000 2558.7400 ;
        RECT 2.0000 2580.0200 5.0000 2580.5000 ;
        RECT 2.0000 2574.5800 5.0000 2575.0600 ;
        RECT 2.0000 2596.3400 5.0000 2596.8200 ;
        RECT 2.0000 2590.9000 5.0000 2591.3800 ;
        RECT 2.0000 2585.4600 5.0000 2585.9400 ;
        RECT 2.0000 2607.2200 5.0000 2607.7000 ;
        RECT 2.0000 2601.7800 5.0000 2602.2600 ;
        RECT 2.0000 2618.1000 5.0000 2618.5800 ;
        RECT 2.0000 2612.6600 5.0000 2613.1400 ;
        RECT 2.0000 2634.4200 5.0000 2634.9000 ;
        RECT 2.0000 2628.9800 5.0000 2629.4600 ;
        RECT 2.0000 2623.5400 5.0000 2624.0200 ;
        RECT 2.0000 2645.3000 5.0000 2645.7800 ;
        RECT 2.0000 2639.8600 5.0000 2640.3400 ;
        RECT 2.0000 2661.6200 5.0000 2662.1000 ;
        RECT 2.0000 2656.1800 5.0000 2656.6600 ;
        RECT 2.0000 2650.7400 5.0000 2651.2200 ;
        RECT 2.0000 2672.5000 5.0000 2672.9800 ;
        RECT 2.0000 2667.0600 5.0000 2667.5400 ;
        RECT 2.0000 2688.8200 5.0000 2689.3000 ;
        RECT 2.0000 2683.3800 5.0000 2683.8600 ;
        RECT 2.0000 2677.9400 5.0000 2678.4200 ;
        RECT 2.0000 2699.7000 5.0000 2700.1800 ;
        RECT 2.0000 2694.2600 5.0000 2694.7400 ;
        RECT 2.0000 2710.5800 5.0000 2711.0600 ;
        RECT 2.0000 2705.1400 5.0000 2705.6200 ;
        RECT 2.0000 2726.9000 5.0000 2727.3800 ;
        RECT 2.0000 2721.4600 5.0000 2721.9400 ;
        RECT 2.0000 2737.7800 5.0000 2738.2600 ;
        RECT 2.0000 2732.3400 5.0000 2732.8200 ;
        RECT 2.0000 2754.1000 5.0000 2754.5800 ;
        RECT 2.0000 2748.6600 5.0000 2749.1400 ;
        RECT 2.0000 2743.2200 5.0000 2743.7000 ;
        RECT 2.0000 2764.9800 5.0000 2765.4600 ;
        RECT 2.0000 2759.5400 5.0000 2760.0200 ;
        RECT 2.0000 2781.3000 5.0000 2781.7800 ;
        RECT 2.0000 2775.8600 5.0000 2776.3400 ;
        RECT 2.0000 2770.4200 5.0000 2770.9000 ;
        RECT 2.0000 2792.1800 5.0000 2792.6600 ;
        RECT 2.0000 2786.7400 5.0000 2787.2200 ;
        RECT 2.0000 2808.5000 5.0000 2808.9800 ;
        RECT 2.0000 2803.0600 5.0000 2803.5400 ;
        RECT 2.0000 2797.6200 5.0000 2798.1000 ;
        RECT 2.0000 2819.3800 5.0000 2819.8600 ;
        RECT 2.0000 2813.9400 5.0000 2814.4200 ;
        RECT 2.0000 2830.2600 5.0000 2830.7400 ;
        RECT 2.0000 2824.8200 5.0000 2825.3000 ;
        RECT 2.0000 2846.5800 5.0000 2847.0600 ;
        RECT 2.0000 2841.1400 5.0000 2841.6200 ;
        RECT 2.0000 2835.7000 5.0000 2836.1800 ;
        RECT 2.0000 2857.4600 5.0000 2857.9400 ;
        RECT 2.0000 2852.0200 5.0000 2852.5000 ;
        RECT 2.0000 2873.7800 5.0000 2874.2600 ;
        RECT 2.0000 2868.3400 5.0000 2868.8200 ;
        RECT 2.0000 2862.9000 5.0000 2863.3800 ;
        RECT 2.0000 2879.2200 5.0000 2879.7000 ;
        RECT 3385.2000 1497.4600 3388.2000 1497.9400 ;
        RECT 3385.2000 1453.9400 3388.2000 1454.4200 ;
        RECT 3385.2000 1448.5000 3388.2000 1448.9800 ;
        RECT 3385.2000 1470.2600 3388.2000 1470.7400 ;
        RECT 3385.2000 1464.8200 3388.2000 1465.3000 ;
        RECT 3385.2000 1459.3800 3388.2000 1459.8600 ;
        RECT 3385.2000 1481.1400 3388.2000 1481.6200 ;
        RECT 3385.2000 1475.7000 3388.2000 1476.1800 ;
        RECT 3385.2000 1492.0200 3388.2000 1492.5000 ;
        RECT 3385.2000 1486.5800 3388.2000 1487.0600 ;
        RECT 3385.2000 1508.3400 3388.2000 1508.8200 ;
        RECT 3385.2000 1502.9000 3388.2000 1503.3800 ;
        RECT 3385.2000 1519.2200 3388.2000 1519.7000 ;
        RECT 3385.2000 1513.7800 3388.2000 1514.2600 ;
        RECT 3385.2000 1535.5400 3388.2000 1536.0200 ;
        RECT 3385.2000 1530.1000 3388.2000 1530.5800 ;
        RECT 3385.2000 1524.6600 3388.2000 1525.1400 ;
        RECT 3385.2000 1546.4200 3388.2000 1546.9000 ;
        RECT 3385.2000 1540.9800 3388.2000 1541.4600 ;
        RECT 3385.2000 1562.7400 3388.2000 1563.2200 ;
        RECT 3385.2000 1557.3000 3388.2000 1557.7800 ;
        RECT 3385.2000 1551.8600 3388.2000 1552.3400 ;
        RECT 3385.2000 1573.6200 3388.2000 1574.1000 ;
        RECT 3385.2000 1568.1800 3388.2000 1568.6600 ;
        RECT 3385.2000 1589.9400 3388.2000 1590.4200 ;
        RECT 3385.2000 1584.5000 3388.2000 1584.9800 ;
        RECT 3385.2000 1579.0600 3388.2000 1579.5400 ;
        RECT 3385.2000 1600.8200 3388.2000 1601.3000 ;
        RECT 3385.2000 1595.3800 3388.2000 1595.8600 ;
        RECT 3385.2000 1611.7000 3388.2000 1612.1800 ;
        RECT 3385.2000 1606.2600 3388.2000 1606.7400 ;
        RECT 3385.2000 1628.0200 3388.2000 1628.5000 ;
        RECT 3385.2000 1622.5800 3388.2000 1623.0600 ;
        RECT 3385.2000 1617.1400 3388.2000 1617.6200 ;
        RECT 3385.2000 1638.9000 3388.2000 1639.3800 ;
        RECT 3385.2000 1633.4600 3388.2000 1633.9400 ;
        RECT 3385.2000 1655.2200 3388.2000 1655.7000 ;
        RECT 3385.2000 1649.7800 3388.2000 1650.2600 ;
        RECT 3385.2000 1644.3400 3388.2000 1644.8200 ;
        RECT 3385.2000 1709.6200 3388.2000 1710.1000 ;
        RECT 3385.2000 1666.1000 3388.2000 1666.5800 ;
        RECT 3385.2000 1660.6600 3388.2000 1661.1400 ;
        RECT 3385.2000 1682.4200 3388.2000 1682.9000 ;
        RECT 3385.2000 1676.9800 3388.2000 1677.4600 ;
        RECT 3385.2000 1671.5400 3388.2000 1672.0200 ;
        RECT 3385.2000 1693.3000 3388.2000 1693.7800 ;
        RECT 3385.2000 1687.8600 3388.2000 1688.3400 ;
        RECT 3385.2000 1704.1800 3388.2000 1704.6600 ;
        RECT 3385.2000 1698.7400 3388.2000 1699.2200 ;
        RECT 3385.2000 1720.5000 3388.2000 1720.9800 ;
        RECT 3385.2000 1715.0600 3388.2000 1715.5400 ;
        RECT 3385.2000 1731.3800 3388.2000 1731.8600 ;
        RECT 3385.2000 1725.9400 3388.2000 1726.4200 ;
        RECT 3385.2000 1747.7000 3388.2000 1748.1800 ;
        RECT 3385.2000 1742.2600 3388.2000 1742.7400 ;
        RECT 3385.2000 1736.8200 3388.2000 1737.3000 ;
        RECT 3385.2000 1758.5800 3388.2000 1759.0600 ;
        RECT 3385.2000 1753.1400 3388.2000 1753.6200 ;
        RECT 3385.2000 1774.9000 3388.2000 1775.3800 ;
        RECT 3385.2000 1769.4600 3388.2000 1769.9400 ;
        RECT 3385.2000 1764.0200 3388.2000 1764.5000 ;
        RECT 3385.2000 1785.7800 3388.2000 1786.2600 ;
        RECT 3385.2000 1780.3400 3388.2000 1780.8200 ;
        RECT 3385.2000 1802.1000 3388.2000 1802.5800 ;
        RECT 3385.2000 1796.6600 3388.2000 1797.1400 ;
        RECT 3385.2000 1791.2200 3388.2000 1791.7000 ;
        RECT 3385.2000 1812.9800 3388.2000 1813.4600 ;
        RECT 3385.2000 1807.5400 3388.2000 1808.0200 ;
        RECT 3385.2000 1823.8600 3388.2000 1824.3400 ;
        RECT 3385.2000 1818.4200 3388.2000 1818.9000 ;
        RECT 3385.2000 1840.1800 3388.2000 1840.6600 ;
        RECT 3385.2000 1834.7400 3388.2000 1835.2200 ;
        RECT 3385.2000 1829.3000 3388.2000 1829.7800 ;
        RECT 3385.2000 1851.0600 3388.2000 1851.5400 ;
        RECT 3385.2000 1845.6200 3388.2000 1846.1000 ;
        RECT 3385.2000 1867.3800 3388.2000 1867.8600 ;
        RECT 3385.2000 1861.9400 3388.2000 1862.4200 ;
        RECT 3385.2000 1856.5000 3388.2000 1856.9800 ;
        RECT 3385.2000 1878.2600 3388.2000 1878.7400 ;
        RECT 3385.2000 1872.8200 3388.2000 1873.3000 ;
        RECT 3385.2000 1894.5800 3388.2000 1895.0600 ;
        RECT 3385.2000 1889.1400 3388.2000 1889.6200 ;
        RECT 3385.2000 1883.7000 3388.2000 1884.1800 ;
        RECT 3385.2000 1905.4600 3388.2000 1905.9400 ;
        RECT 3385.2000 1900.0200 3388.2000 1900.5000 ;
        RECT 3385.2000 1916.3400 3388.2000 1916.8200 ;
        RECT 3385.2000 1910.9000 3388.2000 1911.3800 ;
        RECT 3385.2000 1932.6600 3388.2000 1933.1400 ;
        RECT 3385.2000 1927.2200 3388.2000 1927.7000 ;
        RECT 3385.2000 1921.7800 3388.2000 1922.2600 ;
        RECT 3385.2000 1943.5400 3388.2000 1944.0200 ;
        RECT 3385.2000 1938.1000 3388.2000 1938.5800 ;
        RECT 3385.2000 1959.8600 3388.2000 1960.3400 ;
        RECT 3385.2000 1954.4200 3388.2000 1954.9000 ;
        RECT 3385.2000 1948.9800 3388.2000 1949.4600 ;
        RECT 3385.2000 1970.7400 3388.2000 1971.2200 ;
        RECT 3385.2000 1965.3000 3388.2000 1965.7800 ;
        RECT 3385.2000 1987.0600 3388.2000 1987.5400 ;
        RECT 3385.2000 1981.6200 3388.2000 1982.1000 ;
        RECT 3385.2000 1976.1800 3388.2000 1976.6600 ;
        RECT 3385.2000 1997.9400 3388.2000 1998.4200 ;
        RECT 3385.2000 1992.5000 3388.2000 1992.9800 ;
        RECT 3385.2000 2014.2600 3388.2000 2014.7400 ;
        RECT 3385.2000 2008.8200 3388.2000 2009.3000 ;
        RECT 3385.2000 2003.3800 3388.2000 2003.8600 ;
        RECT 3385.2000 2025.1400 3388.2000 2025.6200 ;
        RECT 3385.2000 2019.7000 3388.2000 2020.1800 ;
        RECT 3385.2000 2036.0200 3388.2000 2036.5000 ;
        RECT 3385.2000 2030.5800 3388.2000 2031.0600 ;
        RECT 3385.2000 2052.3400 3388.2000 2052.8200 ;
        RECT 3385.2000 2046.9000 3388.2000 2047.3800 ;
        RECT 3385.2000 2041.4600 3388.2000 2041.9400 ;
        RECT 3385.2000 2063.2200 3388.2000 2063.7000 ;
        RECT 3385.2000 2057.7800 3388.2000 2058.2600 ;
        RECT 3385.2000 2079.5400 3388.2000 2080.0200 ;
        RECT 3385.2000 2074.1000 3388.2000 2074.5800 ;
        RECT 3385.2000 2068.6600 3388.2000 2069.1400 ;
        RECT 3385.2000 2106.7400 3388.2000 2107.2200 ;
        RECT 3385.2000 2090.4200 3388.2000 2090.9000 ;
        RECT 3385.2000 2084.9800 3388.2000 2085.4600 ;
        RECT 3385.2000 2101.3000 3388.2000 2101.7800 ;
        RECT 3385.2000 2095.8600 3388.2000 2096.3400 ;
        RECT 3385.2000 2117.6200 3388.2000 2118.1000 ;
        RECT 3385.2000 2112.1800 3388.2000 2112.6600 ;
        RECT 3385.2000 2128.5000 3388.2000 2128.9800 ;
        RECT 3385.2000 2123.0600 3388.2000 2123.5400 ;
        RECT 3385.2000 2144.8200 3388.2000 2145.3000 ;
        RECT 3385.2000 2139.3800 3388.2000 2139.8600 ;
        RECT 3385.2000 2133.9400 3388.2000 2134.4200 ;
        RECT 3385.2000 2155.7000 3388.2000 2156.1800 ;
        RECT 3385.2000 2150.2600 3388.2000 2150.7400 ;
        RECT 3385.2000 2172.0200 3388.2000 2172.5000 ;
        RECT 3385.2000 2166.5800 3388.2000 2167.0600 ;
        RECT 3385.2000 2161.1400 3388.2000 2161.6200 ;
        RECT 3385.2000 2182.9000 3388.2000 2183.3800 ;
        RECT 3385.2000 2177.4600 3388.2000 2177.9400 ;
        RECT 3385.2000 2199.2200 3388.2000 2199.7000 ;
        RECT 3385.2000 2193.7800 3388.2000 2194.2600 ;
        RECT 3385.2000 2188.3400 3388.2000 2188.8200 ;
        RECT 3385.2000 2210.1000 3388.2000 2210.5800 ;
        RECT 3385.2000 2204.6600 3388.2000 2205.1400 ;
        RECT 3385.2000 2220.9800 3388.2000 2221.4600 ;
        RECT 3385.2000 2215.5400 3388.2000 2216.0200 ;
        RECT 3385.2000 2237.3000 3388.2000 2237.7800 ;
        RECT 3385.2000 2231.8600 3388.2000 2232.3400 ;
        RECT 3385.2000 2226.4200 3388.2000 2226.9000 ;
        RECT 3385.2000 2248.1800 3388.2000 2248.6600 ;
        RECT 3385.2000 2242.7400 3388.2000 2243.2200 ;
        RECT 3385.2000 2264.5000 3388.2000 2264.9800 ;
        RECT 3385.2000 2259.0600 3388.2000 2259.5400 ;
        RECT 3385.2000 2253.6200 3388.2000 2254.1000 ;
        RECT 3385.2000 2275.3800 3388.2000 2275.8600 ;
        RECT 3385.2000 2269.9400 3388.2000 2270.4200 ;
        RECT 3385.2000 2291.7000 3388.2000 2292.1800 ;
        RECT 3385.2000 2286.2600 3388.2000 2286.7400 ;
        RECT 3385.2000 2280.8200 3388.2000 2281.3000 ;
        RECT 3385.2000 2716.0200 3388.2000 2716.5000 ;
        RECT 3385.2000 2503.8600 3388.2000 2504.3400 ;
        RECT 3385.2000 2302.5800 3388.2000 2303.0600 ;
        RECT 3385.2000 2297.1400 3388.2000 2297.6200 ;
        RECT 3385.2000 2313.4600 3388.2000 2313.9400 ;
        RECT 3385.2000 2308.0200 3388.2000 2308.5000 ;
        RECT 3385.2000 2329.7800 3388.2000 2330.2600 ;
        RECT 3385.2000 2324.3400 3388.2000 2324.8200 ;
        RECT 3385.2000 2318.9000 3388.2000 2319.3800 ;
        RECT 3385.2000 2340.6600 3388.2000 2341.1400 ;
        RECT 3385.2000 2335.2200 3388.2000 2335.7000 ;
        RECT 3385.2000 2356.9800 3388.2000 2357.4600 ;
        RECT 3385.2000 2351.5400 3388.2000 2352.0200 ;
        RECT 3385.2000 2346.1000 3388.2000 2346.5800 ;
        RECT 3385.2000 2367.8600 3388.2000 2368.3400 ;
        RECT 3385.2000 2362.4200 3388.2000 2362.9000 ;
        RECT 3385.2000 2384.1800 3388.2000 2384.6600 ;
        RECT 3385.2000 2378.7400 3388.2000 2379.2200 ;
        RECT 3385.2000 2373.3000 3388.2000 2373.7800 ;
        RECT 3385.2000 2395.0600 3388.2000 2395.5400 ;
        RECT 3385.2000 2389.6200 3388.2000 2390.1000 ;
        RECT 3385.2000 2411.3800 3388.2000 2411.8600 ;
        RECT 3385.2000 2405.9400 3388.2000 2406.4200 ;
        RECT 3385.2000 2400.5000 3388.2000 2400.9800 ;
        RECT 3385.2000 2422.2600 3388.2000 2422.7400 ;
        RECT 3385.2000 2416.8200 3388.2000 2417.3000 ;
        RECT 3385.2000 2433.1400 3388.2000 2433.6200 ;
        RECT 3385.2000 2427.7000 3388.2000 2428.1800 ;
        RECT 3385.2000 2449.4600 3388.2000 2449.9400 ;
        RECT 3385.2000 2444.0200 3388.2000 2444.5000 ;
        RECT 3385.2000 2438.5800 3388.2000 2439.0600 ;
        RECT 3385.2000 2460.3400 3388.2000 2460.8200 ;
        RECT 3385.2000 2454.9000 3388.2000 2455.3800 ;
        RECT 3385.2000 2476.6600 3388.2000 2477.1400 ;
        RECT 3385.2000 2471.2200 3388.2000 2471.7000 ;
        RECT 3385.2000 2465.7800 3388.2000 2466.2600 ;
        RECT 3385.2000 2487.5400 3388.2000 2488.0200 ;
        RECT 3385.2000 2482.1000 3388.2000 2482.5800 ;
        RECT 3385.2000 2498.4200 3388.2000 2498.9000 ;
        RECT 3385.2000 2492.9800 3388.2000 2493.4600 ;
        RECT 3385.2000 2514.7400 3388.2000 2515.2200 ;
        RECT 3385.2000 2509.3000 3388.2000 2509.7800 ;
        RECT 3385.2000 2525.6200 3388.2000 2526.1000 ;
        RECT 3385.2000 2520.1800 3388.2000 2520.6600 ;
        RECT 3385.2000 2541.9400 3388.2000 2542.4200 ;
        RECT 3385.2000 2536.5000 3388.2000 2536.9800 ;
        RECT 3385.2000 2531.0600 3388.2000 2531.5400 ;
        RECT 3385.2000 2552.8200 3388.2000 2553.3000 ;
        RECT 3385.2000 2547.3800 3388.2000 2547.8600 ;
        RECT 3385.2000 2569.1400 3388.2000 2569.6200 ;
        RECT 3385.2000 2563.7000 3388.2000 2564.1800 ;
        RECT 3385.2000 2558.2600 3388.2000 2558.7400 ;
        RECT 3385.2000 2580.0200 3388.2000 2580.5000 ;
        RECT 3385.2000 2574.5800 3388.2000 2575.0600 ;
        RECT 3385.2000 2596.3400 3388.2000 2596.8200 ;
        RECT 3385.2000 2590.9000 3388.2000 2591.3800 ;
        RECT 3385.2000 2585.4600 3388.2000 2585.9400 ;
        RECT 3385.2000 2607.2200 3388.2000 2607.7000 ;
        RECT 3385.2000 2601.7800 3388.2000 2602.2600 ;
        RECT 3385.2000 2618.1000 3388.2000 2618.5800 ;
        RECT 3385.2000 2612.6600 3388.2000 2613.1400 ;
        RECT 3385.2000 2634.4200 3388.2000 2634.9000 ;
        RECT 3385.2000 2628.9800 3388.2000 2629.4600 ;
        RECT 3385.2000 2623.5400 3388.2000 2624.0200 ;
        RECT 3385.2000 2645.3000 3388.2000 2645.7800 ;
        RECT 3385.2000 2639.8600 3388.2000 2640.3400 ;
        RECT 3385.2000 2661.6200 3388.2000 2662.1000 ;
        RECT 3385.2000 2656.1800 3388.2000 2656.6600 ;
        RECT 3385.2000 2650.7400 3388.2000 2651.2200 ;
        RECT 3385.2000 2672.5000 3388.2000 2672.9800 ;
        RECT 3385.2000 2667.0600 3388.2000 2667.5400 ;
        RECT 3385.2000 2688.8200 3388.2000 2689.3000 ;
        RECT 3385.2000 2683.3800 3388.2000 2683.8600 ;
        RECT 3385.2000 2677.9400 3388.2000 2678.4200 ;
        RECT 3385.2000 2699.7000 3388.2000 2700.1800 ;
        RECT 3385.2000 2694.2600 3388.2000 2694.7400 ;
        RECT 3385.2000 2710.5800 3388.2000 2711.0600 ;
        RECT 3385.2000 2705.1400 3388.2000 2705.6200 ;
        RECT 3385.2000 2726.9000 3388.2000 2727.3800 ;
        RECT 3385.2000 2721.4600 3388.2000 2721.9400 ;
        RECT 3385.2000 2737.7800 3388.2000 2738.2600 ;
        RECT 3385.2000 2732.3400 3388.2000 2732.8200 ;
        RECT 3385.2000 2754.1000 3388.2000 2754.5800 ;
        RECT 3385.2000 2748.6600 3388.2000 2749.1400 ;
        RECT 3385.2000 2743.2200 3388.2000 2743.7000 ;
        RECT 3385.2000 2764.9800 3388.2000 2765.4600 ;
        RECT 3385.2000 2759.5400 3388.2000 2760.0200 ;
        RECT 3385.2000 2781.3000 3388.2000 2781.7800 ;
        RECT 3385.2000 2775.8600 3388.2000 2776.3400 ;
        RECT 3385.2000 2770.4200 3388.2000 2770.9000 ;
        RECT 3385.2000 2792.1800 3388.2000 2792.6600 ;
        RECT 3385.2000 2786.7400 3388.2000 2787.2200 ;
        RECT 3385.2000 2808.5000 3388.2000 2808.9800 ;
        RECT 3385.2000 2803.0600 3388.2000 2803.5400 ;
        RECT 3385.2000 2797.6200 3388.2000 2798.1000 ;
        RECT 3385.2000 2819.3800 3388.2000 2819.8600 ;
        RECT 3385.2000 2813.9400 3388.2000 2814.4200 ;
        RECT 3385.2000 2830.2600 3388.2000 2830.7400 ;
        RECT 3385.2000 2824.8200 3388.2000 2825.3000 ;
        RECT 3385.2000 2846.5800 3388.2000 2847.0600 ;
        RECT 3385.2000 2841.1400 3388.2000 2841.6200 ;
        RECT 3385.2000 2835.7000 3388.2000 2836.1800 ;
        RECT 3385.2000 2857.4600 3388.2000 2857.9400 ;
        RECT 3385.2000 2852.0200 3388.2000 2852.5000 ;
        RECT 3385.2000 2873.7800 3388.2000 2874.2600 ;
        RECT 3385.2000 2868.3400 3388.2000 2868.8200 ;
        RECT 3385.2000 2862.9000 3388.2000 2863.3800 ;
        RECT 3385.2000 2879.2200 3388.2000 2879.7000 ;
      LAYER met4 ;
        RECT 3385.2000 2.0000 3388.2000 2887.6600 ;
        RECT 2.0000 2.0000 5.0000 2887.6600 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2805.7800 76.7900 2807.2800 520.5800 ;
        RECT 3308.3000 76.7900 3309.8000 520.5800 ;
      LAYER met3 ;
        RECT 3308.3000 102.5200 3309.8000 103.0000 ;
        RECT 3308.3000 97.0800 3309.8000 97.5600 ;
        RECT 3308.3000 91.6400 3309.8000 92.1200 ;
        RECT 3308.3000 86.2000 3309.8000 86.6800 ;
        RECT 2805.7800 102.5200 2807.2800 103.0000 ;
        RECT 2805.7800 97.0800 2807.2800 97.5600 ;
        RECT 2805.7800 91.6400 2807.2800 92.1200 ;
        RECT 2805.7800 86.2000 2807.2800 86.6800 ;
        RECT 2805.7800 519.0800 3309.8000 520.5800 ;
        RECT 2805.7800 76.7900 3309.8000 78.2900 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2805.7800 536.0700 2807.2800 979.8600 ;
        RECT 3308.3000 536.0700 3309.8000 979.8600 ;
      LAYER met3 ;
        RECT 3308.3000 561.8000 3309.8000 562.2800 ;
        RECT 3308.3000 556.3600 3309.8000 556.8400 ;
        RECT 3308.3000 550.9200 3309.8000 551.4000 ;
        RECT 3308.3000 545.4800 3309.8000 545.9600 ;
        RECT 2805.7800 561.8000 2807.2800 562.2800 ;
        RECT 2805.7800 556.3600 2807.2800 556.8400 ;
        RECT 2805.7800 550.9200 2807.2800 551.4000 ;
        RECT 2805.7800 545.4800 2807.2800 545.9600 ;
        RECT 2805.7800 978.3600 3309.8000 979.8600 ;
        RECT 2805.7800 536.0700 3309.8000 537.5700 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2805.7800 995.3500 2807.2800 1439.1400 ;
        RECT 3308.3000 995.3500 3309.8000 1439.1400 ;
      LAYER met3 ;
        RECT 3308.3000 1021.0800 3309.8000 1021.5600 ;
        RECT 3308.3000 1015.6400 3309.8000 1016.1200 ;
        RECT 3308.3000 1010.2000 3309.8000 1010.6800 ;
        RECT 3308.3000 1004.7600 3309.8000 1005.2400 ;
        RECT 2805.7800 1021.0800 2807.2800 1021.5600 ;
        RECT 2805.7800 1015.6400 2807.2800 1016.1200 ;
        RECT 2805.7800 1010.2000 2807.2800 1010.6800 ;
        RECT 2805.7800 1004.7600 2807.2800 1005.2400 ;
        RECT 2805.7800 1437.6400 3309.8000 1439.1400 ;
        RECT 2805.7800 995.3500 3309.8000 996.8500 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2805.7800 1454.6300 2807.2800 1898.4200 ;
        RECT 3308.3000 1454.6300 3309.8000 1898.4200 ;
      LAYER met3 ;
        RECT 3308.3000 1480.3600 3309.8000 1480.8400 ;
        RECT 3308.3000 1474.9200 3309.8000 1475.4000 ;
        RECT 3308.3000 1469.4800 3309.8000 1469.9600 ;
        RECT 3308.3000 1464.0400 3309.8000 1464.5200 ;
        RECT 2805.7800 1480.3600 2807.2800 1480.8400 ;
        RECT 2805.7800 1474.9200 2807.2800 1475.4000 ;
        RECT 2805.7800 1469.4800 2807.2800 1469.9600 ;
        RECT 2805.7800 1464.0400 2807.2800 1464.5200 ;
        RECT 2805.7800 1896.9200 3309.8000 1898.4200 ;
        RECT 2805.7800 1454.6300 3309.8000 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2805.7800 1913.9100 2807.2800 2357.7000 ;
        RECT 3308.3000 1913.9100 3309.8000 2357.7000 ;
      LAYER met3 ;
        RECT 3308.3000 1939.6400 3309.8000 1940.1200 ;
        RECT 3308.3000 1934.2000 3309.8000 1934.6800 ;
        RECT 3308.3000 1928.7600 3309.8000 1929.2400 ;
        RECT 3308.3000 1923.3200 3309.8000 1923.8000 ;
        RECT 2805.7800 1939.6400 2807.2800 1940.1200 ;
        RECT 2805.7800 1934.2000 2807.2800 1934.6800 ;
        RECT 2805.7800 1928.7600 2807.2800 1929.2400 ;
        RECT 2805.7800 1923.3200 2807.2800 1923.8000 ;
        RECT 2805.7800 2356.2000 3309.8000 2357.7000 ;
        RECT 2805.7800 1913.9100 3309.8000 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2805.7800 2373.1900 2807.2800 2816.9800 ;
        RECT 3308.3000 2373.1900 3309.8000 2816.9800 ;
      LAYER met3 ;
        RECT 3308.3000 2398.9200 3309.8000 2399.4000 ;
        RECT 3308.3000 2393.4800 3309.8000 2393.9600 ;
        RECT 3308.3000 2388.0400 3309.8000 2388.5200 ;
        RECT 3308.3000 2382.6000 3309.8000 2383.0800 ;
        RECT 2805.7800 2398.9200 2807.2800 2399.4000 ;
        RECT 2805.7800 2393.4800 2807.2800 2393.9600 ;
        RECT 2805.7800 2388.0400 2807.2800 2388.5200 ;
        RECT 2805.7800 2382.6000 2807.2800 2383.0800 ;
        RECT 2805.7800 2815.4800 3309.8000 2816.9800 ;
        RECT 2805.7800 2373.1900 3309.8000 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 538.7300 226.6500 747.0300 ;
        RECT 163.5100 538.7300 164.5100 747.0300 ;
      LAYER met3 ;
        RECT 225.6500 741.5800 226.6500 742.0600 ;
        RECT 225.6500 730.7000 226.6500 731.1800 ;
        RECT 225.6500 736.1400 226.6500 736.6200 ;
        RECT 225.6500 714.3800 226.6500 714.8600 ;
        RECT 225.6500 719.8200 226.6500 720.3000 ;
        RECT 225.6500 703.5000 226.6500 703.9800 ;
        RECT 225.6500 708.9400 226.6500 709.4200 ;
        RECT 225.6500 725.2600 226.6500 725.7400 ;
        RECT 225.6500 687.1800 226.6500 687.6600 ;
        RECT 225.6500 692.6200 226.6500 693.1000 ;
        RECT 225.6500 670.8600 226.6500 671.3400 ;
        RECT 225.6500 676.3000 226.6500 676.7800 ;
        RECT 225.6500 681.7400 226.6500 682.2200 ;
        RECT 225.6500 659.9800 226.6500 660.4600 ;
        RECT 225.6500 665.4200 226.6500 665.9000 ;
        RECT 225.6500 643.6600 226.6500 644.1400 ;
        RECT 225.6500 649.1000 226.6500 649.5800 ;
        RECT 225.6500 654.5400 226.6500 655.0200 ;
        RECT 225.6500 698.0600 226.6500 698.5400 ;
        RECT 163.5100 741.5800 164.5100 742.0600 ;
        RECT 163.5100 730.7000 164.5100 731.1800 ;
        RECT 163.5100 736.1400 164.5100 736.6200 ;
        RECT 163.5100 714.3800 164.5100 714.8600 ;
        RECT 163.5100 719.8200 164.5100 720.3000 ;
        RECT 163.5100 703.5000 164.5100 703.9800 ;
        RECT 163.5100 708.9400 164.5100 709.4200 ;
        RECT 163.5100 725.2600 164.5100 725.7400 ;
        RECT 163.5100 687.1800 164.5100 687.6600 ;
        RECT 163.5100 692.6200 164.5100 693.1000 ;
        RECT 163.5100 670.8600 164.5100 671.3400 ;
        RECT 163.5100 676.3000 164.5100 676.7800 ;
        RECT 163.5100 681.7400 164.5100 682.2200 ;
        RECT 163.5100 659.9800 164.5100 660.4600 ;
        RECT 163.5100 665.4200 164.5100 665.9000 ;
        RECT 163.5100 643.6600 164.5100 644.1400 ;
        RECT 163.5100 649.1000 164.5100 649.5800 ;
        RECT 163.5100 654.5400 164.5100 655.0200 ;
        RECT 163.5100 698.0600 164.5100 698.5400 ;
        RECT 225.6500 632.7800 226.6500 633.2600 ;
        RECT 225.6500 638.2200 226.6500 638.7000 ;
        RECT 225.6500 616.4600 226.6500 616.9400 ;
        RECT 225.6500 621.9000 226.6500 622.3800 ;
        RECT 225.6500 627.3400 226.6500 627.8200 ;
        RECT 225.6500 605.5800 226.6500 606.0600 ;
        RECT 225.6500 611.0200 226.6500 611.5000 ;
        RECT 225.6500 589.2600 226.6500 589.7400 ;
        RECT 225.6500 594.7000 226.6500 595.1800 ;
        RECT 225.6500 600.1400 226.6500 600.6200 ;
        RECT 225.6500 578.3800 226.6500 578.8600 ;
        RECT 225.6500 583.8200 226.6500 584.3000 ;
        RECT 225.6500 562.0600 226.6500 562.5400 ;
        RECT 225.6500 567.5000 226.6500 567.9800 ;
        RECT 225.6500 572.9400 226.6500 573.4200 ;
        RECT 225.6500 551.1800 226.6500 551.6600 ;
        RECT 225.6500 556.6200 226.6500 557.1000 ;
        RECT 225.6500 545.7400 226.6500 546.2200 ;
        RECT 163.5100 632.7800 164.5100 633.2600 ;
        RECT 163.5100 638.2200 164.5100 638.7000 ;
        RECT 163.5100 616.4600 164.5100 616.9400 ;
        RECT 163.5100 621.9000 164.5100 622.3800 ;
        RECT 163.5100 627.3400 164.5100 627.8200 ;
        RECT 163.5100 605.5800 164.5100 606.0600 ;
        RECT 163.5100 611.0200 164.5100 611.5000 ;
        RECT 163.5100 589.2600 164.5100 589.7400 ;
        RECT 163.5100 594.7000 164.5100 595.1800 ;
        RECT 163.5100 600.1400 164.5100 600.6200 ;
        RECT 163.5100 578.3800 164.5100 578.8600 ;
        RECT 163.5100 583.8200 164.5100 584.3000 ;
        RECT 163.5100 562.0600 164.5100 562.5400 ;
        RECT 163.5100 567.5000 164.5100 567.9800 ;
        RECT 163.5100 572.9400 164.5100 573.4200 ;
        RECT 163.5100 551.1800 164.5100 551.6600 ;
        RECT 163.5100 556.6200 164.5100 557.1000 ;
        RECT 163.5100 545.7400 164.5100 546.2200 ;
        RECT 163.5100 746.0300 226.6500 747.0300 ;
        RECT 163.5100 538.7300 226.6500 539.7300 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 309.0900 226.6500 517.3900 ;
        RECT 163.5100 309.0900 164.5100 517.3900 ;
      LAYER met3 ;
        RECT 225.6500 511.9400 226.6500 512.4200 ;
        RECT 225.6500 501.0600 226.6500 501.5400 ;
        RECT 225.6500 506.5000 226.6500 506.9800 ;
        RECT 225.6500 484.7400 226.6500 485.2200 ;
        RECT 225.6500 490.1800 226.6500 490.6600 ;
        RECT 225.6500 473.8600 226.6500 474.3400 ;
        RECT 225.6500 479.3000 226.6500 479.7800 ;
        RECT 225.6500 495.6200 226.6500 496.1000 ;
        RECT 225.6500 457.5400 226.6500 458.0200 ;
        RECT 225.6500 462.9800 226.6500 463.4600 ;
        RECT 225.6500 441.2200 226.6500 441.7000 ;
        RECT 225.6500 446.6600 226.6500 447.1400 ;
        RECT 225.6500 452.1000 226.6500 452.5800 ;
        RECT 225.6500 430.3400 226.6500 430.8200 ;
        RECT 225.6500 435.7800 226.6500 436.2600 ;
        RECT 225.6500 414.0200 226.6500 414.5000 ;
        RECT 225.6500 419.4600 226.6500 419.9400 ;
        RECT 225.6500 424.9000 226.6500 425.3800 ;
        RECT 225.6500 468.4200 226.6500 468.9000 ;
        RECT 163.5100 511.9400 164.5100 512.4200 ;
        RECT 163.5100 501.0600 164.5100 501.5400 ;
        RECT 163.5100 506.5000 164.5100 506.9800 ;
        RECT 163.5100 484.7400 164.5100 485.2200 ;
        RECT 163.5100 490.1800 164.5100 490.6600 ;
        RECT 163.5100 473.8600 164.5100 474.3400 ;
        RECT 163.5100 479.3000 164.5100 479.7800 ;
        RECT 163.5100 495.6200 164.5100 496.1000 ;
        RECT 163.5100 457.5400 164.5100 458.0200 ;
        RECT 163.5100 462.9800 164.5100 463.4600 ;
        RECT 163.5100 441.2200 164.5100 441.7000 ;
        RECT 163.5100 446.6600 164.5100 447.1400 ;
        RECT 163.5100 452.1000 164.5100 452.5800 ;
        RECT 163.5100 430.3400 164.5100 430.8200 ;
        RECT 163.5100 435.7800 164.5100 436.2600 ;
        RECT 163.5100 414.0200 164.5100 414.5000 ;
        RECT 163.5100 419.4600 164.5100 419.9400 ;
        RECT 163.5100 424.9000 164.5100 425.3800 ;
        RECT 163.5100 468.4200 164.5100 468.9000 ;
        RECT 225.6500 403.1400 226.6500 403.6200 ;
        RECT 225.6500 408.5800 226.6500 409.0600 ;
        RECT 225.6500 386.8200 226.6500 387.3000 ;
        RECT 225.6500 392.2600 226.6500 392.7400 ;
        RECT 225.6500 397.7000 226.6500 398.1800 ;
        RECT 225.6500 375.9400 226.6500 376.4200 ;
        RECT 225.6500 381.3800 226.6500 381.8600 ;
        RECT 225.6500 359.6200 226.6500 360.1000 ;
        RECT 225.6500 365.0600 226.6500 365.5400 ;
        RECT 225.6500 370.5000 226.6500 370.9800 ;
        RECT 225.6500 348.7400 226.6500 349.2200 ;
        RECT 225.6500 354.1800 226.6500 354.6600 ;
        RECT 225.6500 332.4200 226.6500 332.9000 ;
        RECT 225.6500 337.8600 226.6500 338.3400 ;
        RECT 225.6500 343.3000 226.6500 343.7800 ;
        RECT 225.6500 321.5400 226.6500 322.0200 ;
        RECT 225.6500 326.9800 226.6500 327.4600 ;
        RECT 225.6500 316.1000 226.6500 316.5800 ;
        RECT 163.5100 403.1400 164.5100 403.6200 ;
        RECT 163.5100 408.5800 164.5100 409.0600 ;
        RECT 163.5100 386.8200 164.5100 387.3000 ;
        RECT 163.5100 392.2600 164.5100 392.7400 ;
        RECT 163.5100 397.7000 164.5100 398.1800 ;
        RECT 163.5100 375.9400 164.5100 376.4200 ;
        RECT 163.5100 381.3800 164.5100 381.8600 ;
        RECT 163.5100 359.6200 164.5100 360.1000 ;
        RECT 163.5100 365.0600 164.5100 365.5400 ;
        RECT 163.5100 370.5000 164.5100 370.9800 ;
        RECT 163.5100 348.7400 164.5100 349.2200 ;
        RECT 163.5100 354.1800 164.5100 354.6600 ;
        RECT 163.5100 332.4200 164.5100 332.9000 ;
        RECT 163.5100 337.8600 164.5100 338.3400 ;
        RECT 163.5100 343.3000 164.5100 343.7800 ;
        RECT 163.5100 321.5400 164.5100 322.0200 ;
        RECT 163.5100 326.9800 164.5100 327.4600 ;
        RECT 163.5100 316.1000 164.5100 316.5800 ;
        RECT 163.5100 516.3900 226.6500 517.3900 ;
        RECT 163.5100 309.0900 226.6500 310.0900 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 79.4500 226.6500 287.7500 ;
        RECT 163.5100 79.4500 164.5100 287.7500 ;
      LAYER met3 ;
        RECT 225.6500 282.3000 226.6500 282.7800 ;
        RECT 225.6500 271.4200 226.6500 271.9000 ;
        RECT 225.6500 276.8600 226.6500 277.3400 ;
        RECT 225.6500 255.1000 226.6500 255.5800 ;
        RECT 225.6500 260.5400 226.6500 261.0200 ;
        RECT 225.6500 244.2200 226.6500 244.7000 ;
        RECT 225.6500 249.6600 226.6500 250.1400 ;
        RECT 225.6500 265.9800 226.6500 266.4600 ;
        RECT 225.6500 227.9000 226.6500 228.3800 ;
        RECT 225.6500 233.3400 226.6500 233.8200 ;
        RECT 225.6500 211.5800 226.6500 212.0600 ;
        RECT 225.6500 217.0200 226.6500 217.5000 ;
        RECT 225.6500 222.4600 226.6500 222.9400 ;
        RECT 225.6500 200.7000 226.6500 201.1800 ;
        RECT 225.6500 206.1400 226.6500 206.6200 ;
        RECT 225.6500 184.3800 226.6500 184.8600 ;
        RECT 225.6500 189.8200 226.6500 190.3000 ;
        RECT 225.6500 195.2600 226.6500 195.7400 ;
        RECT 225.6500 238.7800 226.6500 239.2600 ;
        RECT 163.5100 282.3000 164.5100 282.7800 ;
        RECT 163.5100 271.4200 164.5100 271.9000 ;
        RECT 163.5100 276.8600 164.5100 277.3400 ;
        RECT 163.5100 255.1000 164.5100 255.5800 ;
        RECT 163.5100 260.5400 164.5100 261.0200 ;
        RECT 163.5100 244.2200 164.5100 244.7000 ;
        RECT 163.5100 249.6600 164.5100 250.1400 ;
        RECT 163.5100 265.9800 164.5100 266.4600 ;
        RECT 163.5100 227.9000 164.5100 228.3800 ;
        RECT 163.5100 233.3400 164.5100 233.8200 ;
        RECT 163.5100 211.5800 164.5100 212.0600 ;
        RECT 163.5100 217.0200 164.5100 217.5000 ;
        RECT 163.5100 222.4600 164.5100 222.9400 ;
        RECT 163.5100 200.7000 164.5100 201.1800 ;
        RECT 163.5100 206.1400 164.5100 206.6200 ;
        RECT 163.5100 184.3800 164.5100 184.8600 ;
        RECT 163.5100 189.8200 164.5100 190.3000 ;
        RECT 163.5100 195.2600 164.5100 195.7400 ;
        RECT 163.5100 238.7800 164.5100 239.2600 ;
        RECT 225.6500 173.5000 226.6500 173.9800 ;
        RECT 225.6500 178.9400 226.6500 179.4200 ;
        RECT 225.6500 157.1800 226.6500 157.6600 ;
        RECT 225.6500 162.6200 226.6500 163.1000 ;
        RECT 225.6500 168.0600 226.6500 168.5400 ;
        RECT 225.6500 146.3000 226.6500 146.7800 ;
        RECT 225.6500 151.7400 226.6500 152.2200 ;
        RECT 225.6500 129.9800 226.6500 130.4600 ;
        RECT 225.6500 135.4200 226.6500 135.9000 ;
        RECT 225.6500 140.8600 226.6500 141.3400 ;
        RECT 225.6500 119.1000 226.6500 119.5800 ;
        RECT 225.6500 124.5400 226.6500 125.0200 ;
        RECT 225.6500 102.7800 226.6500 103.2600 ;
        RECT 225.6500 108.2200 226.6500 108.7000 ;
        RECT 225.6500 113.6600 226.6500 114.1400 ;
        RECT 225.6500 91.9000 226.6500 92.3800 ;
        RECT 225.6500 97.3400 226.6500 97.8200 ;
        RECT 225.6500 86.4600 226.6500 86.9400 ;
        RECT 163.5100 173.5000 164.5100 173.9800 ;
        RECT 163.5100 178.9400 164.5100 179.4200 ;
        RECT 163.5100 157.1800 164.5100 157.6600 ;
        RECT 163.5100 162.6200 164.5100 163.1000 ;
        RECT 163.5100 168.0600 164.5100 168.5400 ;
        RECT 163.5100 146.3000 164.5100 146.7800 ;
        RECT 163.5100 151.7400 164.5100 152.2200 ;
        RECT 163.5100 129.9800 164.5100 130.4600 ;
        RECT 163.5100 135.4200 164.5100 135.9000 ;
        RECT 163.5100 140.8600 164.5100 141.3400 ;
        RECT 163.5100 119.1000 164.5100 119.5800 ;
        RECT 163.5100 124.5400 164.5100 125.0200 ;
        RECT 163.5100 102.7800 164.5100 103.2600 ;
        RECT 163.5100 108.2200 164.5100 108.7000 ;
        RECT 163.5100 113.6600 164.5100 114.1400 ;
        RECT 163.5100 91.9000 164.5100 92.3800 ;
        RECT 163.5100 97.3400 164.5100 97.8200 ;
        RECT 163.5100 86.4600 164.5100 86.9400 ;
        RECT 163.5100 286.7500 226.6500 287.7500 ;
        RECT 163.5100 79.4500 226.6500 80.4500 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 2605.4900 226.6500 2813.7900 ;
        RECT 163.5100 2605.4900 164.5100 2813.7900 ;
      LAYER met3 ;
        RECT 225.6500 2808.3400 226.6500 2808.8200 ;
        RECT 225.6500 2797.4600 226.6500 2797.9400 ;
        RECT 225.6500 2802.9000 226.6500 2803.3800 ;
        RECT 225.6500 2781.1400 226.6500 2781.6200 ;
        RECT 225.6500 2786.5800 226.6500 2787.0600 ;
        RECT 225.6500 2770.2600 226.6500 2770.7400 ;
        RECT 225.6500 2775.7000 226.6500 2776.1800 ;
        RECT 225.6500 2792.0200 226.6500 2792.5000 ;
        RECT 225.6500 2753.9400 226.6500 2754.4200 ;
        RECT 225.6500 2759.3800 226.6500 2759.8600 ;
        RECT 225.6500 2737.6200 226.6500 2738.1000 ;
        RECT 225.6500 2743.0600 226.6500 2743.5400 ;
        RECT 225.6500 2748.5000 226.6500 2748.9800 ;
        RECT 225.6500 2726.7400 226.6500 2727.2200 ;
        RECT 225.6500 2732.1800 226.6500 2732.6600 ;
        RECT 225.6500 2710.4200 226.6500 2710.9000 ;
        RECT 225.6500 2715.8600 226.6500 2716.3400 ;
        RECT 225.6500 2721.3000 226.6500 2721.7800 ;
        RECT 225.6500 2764.8200 226.6500 2765.3000 ;
        RECT 163.5100 2808.3400 164.5100 2808.8200 ;
        RECT 163.5100 2797.4600 164.5100 2797.9400 ;
        RECT 163.5100 2802.9000 164.5100 2803.3800 ;
        RECT 163.5100 2781.1400 164.5100 2781.6200 ;
        RECT 163.5100 2786.5800 164.5100 2787.0600 ;
        RECT 163.5100 2770.2600 164.5100 2770.7400 ;
        RECT 163.5100 2775.7000 164.5100 2776.1800 ;
        RECT 163.5100 2792.0200 164.5100 2792.5000 ;
        RECT 163.5100 2753.9400 164.5100 2754.4200 ;
        RECT 163.5100 2759.3800 164.5100 2759.8600 ;
        RECT 163.5100 2737.6200 164.5100 2738.1000 ;
        RECT 163.5100 2743.0600 164.5100 2743.5400 ;
        RECT 163.5100 2748.5000 164.5100 2748.9800 ;
        RECT 163.5100 2726.7400 164.5100 2727.2200 ;
        RECT 163.5100 2732.1800 164.5100 2732.6600 ;
        RECT 163.5100 2710.4200 164.5100 2710.9000 ;
        RECT 163.5100 2715.8600 164.5100 2716.3400 ;
        RECT 163.5100 2721.3000 164.5100 2721.7800 ;
        RECT 163.5100 2764.8200 164.5100 2765.3000 ;
        RECT 225.6500 2699.5400 226.6500 2700.0200 ;
        RECT 225.6500 2704.9800 226.6500 2705.4600 ;
        RECT 225.6500 2683.2200 226.6500 2683.7000 ;
        RECT 225.6500 2688.6600 226.6500 2689.1400 ;
        RECT 225.6500 2694.1000 226.6500 2694.5800 ;
        RECT 225.6500 2672.3400 226.6500 2672.8200 ;
        RECT 225.6500 2677.7800 226.6500 2678.2600 ;
        RECT 225.6500 2656.0200 226.6500 2656.5000 ;
        RECT 225.6500 2661.4600 226.6500 2661.9400 ;
        RECT 225.6500 2666.9000 226.6500 2667.3800 ;
        RECT 225.6500 2645.1400 226.6500 2645.6200 ;
        RECT 225.6500 2650.5800 226.6500 2651.0600 ;
        RECT 225.6500 2628.8200 226.6500 2629.3000 ;
        RECT 225.6500 2634.2600 226.6500 2634.7400 ;
        RECT 225.6500 2639.7000 226.6500 2640.1800 ;
        RECT 225.6500 2617.9400 226.6500 2618.4200 ;
        RECT 225.6500 2623.3800 226.6500 2623.8600 ;
        RECT 225.6500 2612.5000 226.6500 2612.9800 ;
        RECT 163.5100 2699.5400 164.5100 2700.0200 ;
        RECT 163.5100 2704.9800 164.5100 2705.4600 ;
        RECT 163.5100 2683.2200 164.5100 2683.7000 ;
        RECT 163.5100 2688.6600 164.5100 2689.1400 ;
        RECT 163.5100 2694.1000 164.5100 2694.5800 ;
        RECT 163.5100 2672.3400 164.5100 2672.8200 ;
        RECT 163.5100 2677.7800 164.5100 2678.2600 ;
        RECT 163.5100 2656.0200 164.5100 2656.5000 ;
        RECT 163.5100 2661.4600 164.5100 2661.9400 ;
        RECT 163.5100 2666.9000 164.5100 2667.3800 ;
        RECT 163.5100 2645.1400 164.5100 2645.6200 ;
        RECT 163.5100 2650.5800 164.5100 2651.0600 ;
        RECT 163.5100 2628.8200 164.5100 2629.3000 ;
        RECT 163.5100 2634.2600 164.5100 2634.7400 ;
        RECT 163.5100 2639.7000 164.5100 2640.1800 ;
        RECT 163.5100 2617.9400 164.5100 2618.4200 ;
        RECT 163.5100 2623.3800 164.5100 2623.8600 ;
        RECT 163.5100 2612.5000 164.5100 2612.9800 ;
        RECT 163.5100 2812.7900 226.6500 2813.7900 ;
        RECT 163.5100 2605.4900 226.6500 2606.4900 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 2375.8500 226.6500 2584.1500 ;
        RECT 163.5100 2375.8500 164.5100 2584.1500 ;
      LAYER met3 ;
        RECT 225.6500 2578.7000 226.6500 2579.1800 ;
        RECT 225.6500 2567.8200 226.6500 2568.3000 ;
        RECT 225.6500 2573.2600 226.6500 2573.7400 ;
        RECT 225.6500 2551.5000 226.6500 2551.9800 ;
        RECT 225.6500 2556.9400 226.6500 2557.4200 ;
        RECT 225.6500 2540.6200 226.6500 2541.1000 ;
        RECT 225.6500 2546.0600 226.6500 2546.5400 ;
        RECT 225.6500 2562.3800 226.6500 2562.8600 ;
        RECT 225.6500 2524.3000 226.6500 2524.7800 ;
        RECT 225.6500 2529.7400 226.6500 2530.2200 ;
        RECT 225.6500 2507.9800 226.6500 2508.4600 ;
        RECT 225.6500 2513.4200 226.6500 2513.9000 ;
        RECT 225.6500 2518.8600 226.6500 2519.3400 ;
        RECT 225.6500 2497.1000 226.6500 2497.5800 ;
        RECT 225.6500 2502.5400 226.6500 2503.0200 ;
        RECT 225.6500 2480.7800 226.6500 2481.2600 ;
        RECT 225.6500 2486.2200 226.6500 2486.7000 ;
        RECT 225.6500 2491.6600 226.6500 2492.1400 ;
        RECT 225.6500 2535.1800 226.6500 2535.6600 ;
        RECT 163.5100 2578.7000 164.5100 2579.1800 ;
        RECT 163.5100 2567.8200 164.5100 2568.3000 ;
        RECT 163.5100 2573.2600 164.5100 2573.7400 ;
        RECT 163.5100 2551.5000 164.5100 2551.9800 ;
        RECT 163.5100 2556.9400 164.5100 2557.4200 ;
        RECT 163.5100 2540.6200 164.5100 2541.1000 ;
        RECT 163.5100 2546.0600 164.5100 2546.5400 ;
        RECT 163.5100 2562.3800 164.5100 2562.8600 ;
        RECT 163.5100 2524.3000 164.5100 2524.7800 ;
        RECT 163.5100 2529.7400 164.5100 2530.2200 ;
        RECT 163.5100 2507.9800 164.5100 2508.4600 ;
        RECT 163.5100 2513.4200 164.5100 2513.9000 ;
        RECT 163.5100 2518.8600 164.5100 2519.3400 ;
        RECT 163.5100 2497.1000 164.5100 2497.5800 ;
        RECT 163.5100 2502.5400 164.5100 2503.0200 ;
        RECT 163.5100 2480.7800 164.5100 2481.2600 ;
        RECT 163.5100 2486.2200 164.5100 2486.7000 ;
        RECT 163.5100 2491.6600 164.5100 2492.1400 ;
        RECT 163.5100 2535.1800 164.5100 2535.6600 ;
        RECT 225.6500 2469.9000 226.6500 2470.3800 ;
        RECT 225.6500 2475.3400 226.6500 2475.8200 ;
        RECT 225.6500 2453.5800 226.6500 2454.0600 ;
        RECT 225.6500 2459.0200 226.6500 2459.5000 ;
        RECT 225.6500 2464.4600 226.6500 2464.9400 ;
        RECT 225.6500 2442.7000 226.6500 2443.1800 ;
        RECT 225.6500 2448.1400 226.6500 2448.6200 ;
        RECT 225.6500 2426.3800 226.6500 2426.8600 ;
        RECT 225.6500 2431.8200 226.6500 2432.3000 ;
        RECT 225.6500 2437.2600 226.6500 2437.7400 ;
        RECT 225.6500 2415.5000 226.6500 2415.9800 ;
        RECT 225.6500 2420.9400 226.6500 2421.4200 ;
        RECT 225.6500 2399.1800 226.6500 2399.6600 ;
        RECT 225.6500 2404.6200 226.6500 2405.1000 ;
        RECT 225.6500 2410.0600 226.6500 2410.5400 ;
        RECT 225.6500 2388.3000 226.6500 2388.7800 ;
        RECT 225.6500 2393.7400 226.6500 2394.2200 ;
        RECT 225.6500 2382.8600 226.6500 2383.3400 ;
        RECT 163.5100 2469.9000 164.5100 2470.3800 ;
        RECT 163.5100 2475.3400 164.5100 2475.8200 ;
        RECT 163.5100 2453.5800 164.5100 2454.0600 ;
        RECT 163.5100 2459.0200 164.5100 2459.5000 ;
        RECT 163.5100 2464.4600 164.5100 2464.9400 ;
        RECT 163.5100 2442.7000 164.5100 2443.1800 ;
        RECT 163.5100 2448.1400 164.5100 2448.6200 ;
        RECT 163.5100 2426.3800 164.5100 2426.8600 ;
        RECT 163.5100 2431.8200 164.5100 2432.3000 ;
        RECT 163.5100 2437.2600 164.5100 2437.7400 ;
        RECT 163.5100 2415.5000 164.5100 2415.9800 ;
        RECT 163.5100 2420.9400 164.5100 2421.4200 ;
        RECT 163.5100 2399.1800 164.5100 2399.6600 ;
        RECT 163.5100 2404.6200 164.5100 2405.1000 ;
        RECT 163.5100 2410.0600 164.5100 2410.5400 ;
        RECT 163.5100 2388.3000 164.5100 2388.7800 ;
        RECT 163.5100 2393.7400 164.5100 2394.2200 ;
        RECT 163.5100 2382.8600 164.5100 2383.3400 ;
        RECT 163.5100 2583.1500 226.6500 2584.1500 ;
        RECT 163.5100 2375.8500 226.6500 2376.8500 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 2146.2100 226.6500 2354.5100 ;
        RECT 163.5100 2146.2100 164.5100 2354.5100 ;
      LAYER met3 ;
        RECT 225.6500 2349.0600 226.6500 2349.5400 ;
        RECT 225.6500 2338.1800 226.6500 2338.6600 ;
        RECT 225.6500 2343.6200 226.6500 2344.1000 ;
        RECT 225.6500 2321.8600 226.6500 2322.3400 ;
        RECT 225.6500 2327.3000 226.6500 2327.7800 ;
        RECT 225.6500 2310.9800 226.6500 2311.4600 ;
        RECT 225.6500 2316.4200 226.6500 2316.9000 ;
        RECT 225.6500 2332.7400 226.6500 2333.2200 ;
        RECT 225.6500 2294.6600 226.6500 2295.1400 ;
        RECT 225.6500 2300.1000 226.6500 2300.5800 ;
        RECT 225.6500 2278.3400 226.6500 2278.8200 ;
        RECT 225.6500 2283.7800 226.6500 2284.2600 ;
        RECT 225.6500 2289.2200 226.6500 2289.7000 ;
        RECT 225.6500 2267.4600 226.6500 2267.9400 ;
        RECT 225.6500 2272.9000 226.6500 2273.3800 ;
        RECT 225.6500 2251.1400 226.6500 2251.6200 ;
        RECT 225.6500 2256.5800 226.6500 2257.0600 ;
        RECT 225.6500 2262.0200 226.6500 2262.5000 ;
        RECT 225.6500 2305.5400 226.6500 2306.0200 ;
        RECT 163.5100 2349.0600 164.5100 2349.5400 ;
        RECT 163.5100 2338.1800 164.5100 2338.6600 ;
        RECT 163.5100 2343.6200 164.5100 2344.1000 ;
        RECT 163.5100 2321.8600 164.5100 2322.3400 ;
        RECT 163.5100 2327.3000 164.5100 2327.7800 ;
        RECT 163.5100 2310.9800 164.5100 2311.4600 ;
        RECT 163.5100 2316.4200 164.5100 2316.9000 ;
        RECT 163.5100 2332.7400 164.5100 2333.2200 ;
        RECT 163.5100 2294.6600 164.5100 2295.1400 ;
        RECT 163.5100 2300.1000 164.5100 2300.5800 ;
        RECT 163.5100 2278.3400 164.5100 2278.8200 ;
        RECT 163.5100 2283.7800 164.5100 2284.2600 ;
        RECT 163.5100 2289.2200 164.5100 2289.7000 ;
        RECT 163.5100 2267.4600 164.5100 2267.9400 ;
        RECT 163.5100 2272.9000 164.5100 2273.3800 ;
        RECT 163.5100 2251.1400 164.5100 2251.6200 ;
        RECT 163.5100 2256.5800 164.5100 2257.0600 ;
        RECT 163.5100 2262.0200 164.5100 2262.5000 ;
        RECT 163.5100 2305.5400 164.5100 2306.0200 ;
        RECT 225.6500 2240.2600 226.6500 2240.7400 ;
        RECT 225.6500 2245.7000 226.6500 2246.1800 ;
        RECT 225.6500 2223.9400 226.6500 2224.4200 ;
        RECT 225.6500 2229.3800 226.6500 2229.8600 ;
        RECT 225.6500 2234.8200 226.6500 2235.3000 ;
        RECT 225.6500 2213.0600 226.6500 2213.5400 ;
        RECT 225.6500 2218.5000 226.6500 2218.9800 ;
        RECT 225.6500 2196.7400 226.6500 2197.2200 ;
        RECT 225.6500 2202.1800 226.6500 2202.6600 ;
        RECT 225.6500 2207.6200 226.6500 2208.1000 ;
        RECT 225.6500 2185.8600 226.6500 2186.3400 ;
        RECT 225.6500 2191.3000 226.6500 2191.7800 ;
        RECT 225.6500 2169.5400 226.6500 2170.0200 ;
        RECT 225.6500 2174.9800 226.6500 2175.4600 ;
        RECT 225.6500 2180.4200 226.6500 2180.9000 ;
        RECT 225.6500 2158.6600 226.6500 2159.1400 ;
        RECT 225.6500 2164.1000 226.6500 2164.5800 ;
        RECT 225.6500 2153.2200 226.6500 2153.7000 ;
        RECT 163.5100 2240.2600 164.5100 2240.7400 ;
        RECT 163.5100 2245.7000 164.5100 2246.1800 ;
        RECT 163.5100 2223.9400 164.5100 2224.4200 ;
        RECT 163.5100 2229.3800 164.5100 2229.8600 ;
        RECT 163.5100 2234.8200 164.5100 2235.3000 ;
        RECT 163.5100 2213.0600 164.5100 2213.5400 ;
        RECT 163.5100 2218.5000 164.5100 2218.9800 ;
        RECT 163.5100 2196.7400 164.5100 2197.2200 ;
        RECT 163.5100 2202.1800 164.5100 2202.6600 ;
        RECT 163.5100 2207.6200 164.5100 2208.1000 ;
        RECT 163.5100 2185.8600 164.5100 2186.3400 ;
        RECT 163.5100 2191.3000 164.5100 2191.7800 ;
        RECT 163.5100 2169.5400 164.5100 2170.0200 ;
        RECT 163.5100 2174.9800 164.5100 2175.4600 ;
        RECT 163.5100 2180.4200 164.5100 2180.9000 ;
        RECT 163.5100 2158.6600 164.5100 2159.1400 ;
        RECT 163.5100 2164.1000 164.5100 2164.5800 ;
        RECT 163.5100 2153.2200 164.5100 2153.7000 ;
        RECT 163.5100 2353.5100 226.6500 2354.5100 ;
        RECT 163.5100 2146.2100 226.6500 2147.2100 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 1916.5700 226.6500 2124.8700 ;
        RECT 163.5100 1916.5700 164.5100 2124.8700 ;
      LAYER met3 ;
        RECT 225.6500 2119.4200 226.6500 2119.9000 ;
        RECT 225.6500 2108.5400 226.6500 2109.0200 ;
        RECT 225.6500 2113.9800 226.6500 2114.4600 ;
        RECT 225.6500 2092.2200 226.6500 2092.7000 ;
        RECT 225.6500 2097.6600 226.6500 2098.1400 ;
        RECT 225.6500 2081.3400 226.6500 2081.8200 ;
        RECT 225.6500 2086.7800 226.6500 2087.2600 ;
        RECT 225.6500 2103.1000 226.6500 2103.5800 ;
        RECT 225.6500 2065.0200 226.6500 2065.5000 ;
        RECT 225.6500 2070.4600 226.6500 2070.9400 ;
        RECT 225.6500 2048.7000 226.6500 2049.1800 ;
        RECT 225.6500 2054.1400 226.6500 2054.6200 ;
        RECT 225.6500 2059.5800 226.6500 2060.0600 ;
        RECT 225.6500 2037.8200 226.6500 2038.3000 ;
        RECT 225.6500 2043.2600 226.6500 2043.7400 ;
        RECT 225.6500 2021.5000 226.6500 2021.9800 ;
        RECT 225.6500 2026.9400 226.6500 2027.4200 ;
        RECT 225.6500 2032.3800 226.6500 2032.8600 ;
        RECT 225.6500 2075.9000 226.6500 2076.3800 ;
        RECT 163.5100 2119.4200 164.5100 2119.9000 ;
        RECT 163.5100 2108.5400 164.5100 2109.0200 ;
        RECT 163.5100 2113.9800 164.5100 2114.4600 ;
        RECT 163.5100 2092.2200 164.5100 2092.7000 ;
        RECT 163.5100 2097.6600 164.5100 2098.1400 ;
        RECT 163.5100 2081.3400 164.5100 2081.8200 ;
        RECT 163.5100 2086.7800 164.5100 2087.2600 ;
        RECT 163.5100 2103.1000 164.5100 2103.5800 ;
        RECT 163.5100 2065.0200 164.5100 2065.5000 ;
        RECT 163.5100 2070.4600 164.5100 2070.9400 ;
        RECT 163.5100 2048.7000 164.5100 2049.1800 ;
        RECT 163.5100 2054.1400 164.5100 2054.6200 ;
        RECT 163.5100 2059.5800 164.5100 2060.0600 ;
        RECT 163.5100 2037.8200 164.5100 2038.3000 ;
        RECT 163.5100 2043.2600 164.5100 2043.7400 ;
        RECT 163.5100 2021.5000 164.5100 2021.9800 ;
        RECT 163.5100 2026.9400 164.5100 2027.4200 ;
        RECT 163.5100 2032.3800 164.5100 2032.8600 ;
        RECT 163.5100 2075.9000 164.5100 2076.3800 ;
        RECT 225.6500 2010.6200 226.6500 2011.1000 ;
        RECT 225.6500 2016.0600 226.6500 2016.5400 ;
        RECT 225.6500 1994.3000 226.6500 1994.7800 ;
        RECT 225.6500 1999.7400 226.6500 2000.2200 ;
        RECT 225.6500 2005.1800 226.6500 2005.6600 ;
        RECT 225.6500 1983.4200 226.6500 1983.9000 ;
        RECT 225.6500 1988.8600 226.6500 1989.3400 ;
        RECT 225.6500 1967.1000 226.6500 1967.5800 ;
        RECT 225.6500 1972.5400 226.6500 1973.0200 ;
        RECT 225.6500 1977.9800 226.6500 1978.4600 ;
        RECT 225.6500 1956.2200 226.6500 1956.7000 ;
        RECT 225.6500 1961.6600 226.6500 1962.1400 ;
        RECT 225.6500 1939.9000 226.6500 1940.3800 ;
        RECT 225.6500 1945.3400 226.6500 1945.8200 ;
        RECT 225.6500 1950.7800 226.6500 1951.2600 ;
        RECT 225.6500 1929.0200 226.6500 1929.5000 ;
        RECT 225.6500 1934.4600 226.6500 1934.9400 ;
        RECT 225.6500 1923.5800 226.6500 1924.0600 ;
        RECT 163.5100 2010.6200 164.5100 2011.1000 ;
        RECT 163.5100 2016.0600 164.5100 2016.5400 ;
        RECT 163.5100 1994.3000 164.5100 1994.7800 ;
        RECT 163.5100 1999.7400 164.5100 2000.2200 ;
        RECT 163.5100 2005.1800 164.5100 2005.6600 ;
        RECT 163.5100 1983.4200 164.5100 1983.9000 ;
        RECT 163.5100 1988.8600 164.5100 1989.3400 ;
        RECT 163.5100 1967.1000 164.5100 1967.5800 ;
        RECT 163.5100 1972.5400 164.5100 1973.0200 ;
        RECT 163.5100 1977.9800 164.5100 1978.4600 ;
        RECT 163.5100 1956.2200 164.5100 1956.7000 ;
        RECT 163.5100 1961.6600 164.5100 1962.1400 ;
        RECT 163.5100 1939.9000 164.5100 1940.3800 ;
        RECT 163.5100 1945.3400 164.5100 1945.8200 ;
        RECT 163.5100 1950.7800 164.5100 1951.2600 ;
        RECT 163.5100 1929.0200 164.5100 1929.5000 ;
        RECT 163.5100 1934.4600 164.5100 1934.9400 ;
        RECT 163.5100 1923.5800 164.5100 1924.0600 ;
        RECT 163.5100 2123.8700 226.6500 2124.8700 ;
        RECT 163.5100 1916.5700 226.6500 1917.5700 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 1686.9300 226.6500 1895.2300 ;
        RECT 163.5100 1686.9300 164.5100 1895.2300 ;
      LAYER met3 ;
        RECT 225.6500 1889.7800 226.6500 1890.2600 ;
        RECT 225.6500 1878.9000 226.6500 1879.3800 ;
        RECT 225.6500 1884.3400 226.6500 1884.8200 ;
        RECT 225.6500 1862.5800 226.6500 1863.0600 ;
        RECT 225.6500 1868.0200 226.6500 1868.5000 ;
        RECT 225.6500 1851.7000 226.6500 1852.1800 ;
        RECT 225.6500 1857.1400 226.6500 1857.6200 ;
        RECT 225.6500 1873.4600 226.6500 1873.9400 ;
        RECT 225.6500 1835.3800 226.6500 1835.8600 ;
        RECT 225.6500 1840.8200 226.6500 1841.3000 ;
        RECT 225.6500 1819.0600 226.6500 1819.5400 ;
        RECT 225.6500 1824.5000 226.6500 1824.9800 ;
        RECT 225.6500 1829.9400 226.6500 1830.4200 ;
        RECT 225.6500 1808.1800 226.6500 1808.6600 ;
        RECT 225.6500 1813.6200 226.6500 1814.1000 ;
        RECT 225.6500 1791.8600 226.6500 1792.3400 ;
        RECT 225.6500 1797.3000 226.6500 1797.7800 ;
        RECT 225.6500 1802.7400 226.6500 1803.2200 ;
        RECT 225.6500 1846.2600 226.6500 1846.7400 ;
        RECT 163.5100 1889.7800 164.5100 1890.2600 ;
        RECT 163.5100 1878.9000 164.5100 1879.3800 ;
        RECT 163.5100 1884.3400 164.5100 1884.8200 ;
        RECT 163.5100 1862.5800 164.5100 1863.0600 ;
        RECT 163.5100 1868.0200 164.5100 1868.5000 ;
        RECT 163.5100 1851.7000 164.5100 1852.1800 ;
        RECT 163.5100 1857.1400 164.5100 1857.6200 ;
        RECT 163.5100 1873.4600 164.5100 1873.9400 ;
        RECT 163.5100 1835.3800 164.5100 1835.8600 ;
        RECT 163.5100 1840.8200 164.5100 1841.3000 ;
        RECT 163.5100 1819.0600 164.5100 1819.5400 ;
        RECT 163.5100 1824.5000 164.5100 1824.9800 ;
        RECT 163.5100 1829.9400 164.5100 1830.4200 ;
        RECT 163.5100 1808.1800 164.5100 1808.6600 ;
        RECT 163.5100 1813.6200 164.5100 1814.1000 ;
        RECT 163.5100 1791.8600 164.5100 1792.3400 ;
        RECT 163.5100 1797.3000 164.5100 1797.7800 ;
        RECT 163.5100 1802.7400 164.5100 1803.2200 ;
        RECT 163.5100 1846.2600 164.5100 1846.7400 ;
        RECT 225.6500 1780.9800 226.6500 1781.4600 ;
        RECT 225.6500 1786.4200 226.6500 1786.9000 ;
        RECT 225.6500 1764.6600 226.6500 1765.1400 ;
        RECT 225.6500 1770.1000 226.6500 1770.5800 ;
        RECT 225.6500 1775.5400 226.6500 1776.0200 ;
        RECT 225.6500 1753.7800 226.6500 1754.2600 ;
        RECT 225.6500 1759.2200 226.6500 1759.7000 ;
        RECT 225.6500 1737.4600 226.6500 1737.9400 ;
        RECT 225.6500 1742.9000 226.6500 1743.3800 ;
        RECT 225.6500 1748.3400 226.6500 1748.8200 ;
        RECT 225.6500 1726.5800 226.6500 1727.0600 ;
        RECT 225.6500 1732.0200 226.6500 1732.5000 ;
        RECT 225.6500 1710.2600 226.6500 1710.7400 ;
        RECT 225.6500 1715.7000 226.6500 1716.1800 ;
        RECT 225.6500 1721.1400 226.6500 1721.6200 ;
        RECT 225.6500 1699.3800 226.6500 1699.8600 ;
        RECT 225.6500 1704.8200 226.6500 1705.3000 ;
        RECT 225.6500 1693.9400 226.6500 1694.4200 ;
        RECT 163.5100 1780.9800 164.5100 1781.4600 ;
        RECT 163.5100 1786.4200 164.5100 1786.9000 ;
        RECT 163.5100 1764.6600 164.5100 1765.1400 ;
        RECT 163.5100 1770.1000 164.5100 1770.5800 ;
        RECT 163.5100 1775.5400 164.5100 1776.0200 ;
        RECT 163.5100 1753.7800 164.5100 1754.2600 ;
        RECT 163.5100 1759.2200 164.5100 1759.7000 ;
        RECT 163.5100 1737.4600 164.5100 1737.9400 ;
        RECT 163.5100 1742.9000 164.5100 1743.3800 ;
        RECT 163.5100 1748.3400 164.5100 1748.8200 ;
        RECT 163.5100 1726.5800 164.5100 1727.0600 ;
        RECT 163.5100 1732.0200 164.5100 1732.5000 ;
        RECT 163.5100 1710.2600 164.5100 1710.7400 ;
        RECT 163.5100 1715.7000 164.5100 1716.1800 ;
        RECT 163.5100 1721.1400 164.5100 1721.6200 ;
        RECT 163.5100 1699.3800 164.5100 1699.8600 ;
        RECT 163.5100 1704.8200 164.5100 1705.3000 ;
        RECT 163.5100 1693.9400 164.5100 1694.4200 ;
        RECT 163.5100 1894.2300 226.6500 1895.2300 ;
        RECT 163.5100 1686.9300 226.6500 1687.9300 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 1457.2900 226.6500 1665.5900 ;
        RECT 163.5100 1457.2900 164.5100 1665.5900 ;
      LAYER met3 ;
        RECT 225.6500 1660.1400 226.6500 1660.6200 ;
        RECT 225.6500 1649.2600 226.6500 1649.7400 ;
        RECT 225.6500 1654.7000 226.6500 1655.1800 ;
        RECT 225.6500 1632.9400 226.6500 1633.4200 ;
        RECT 225.6500 1638.3800 226.6500 1638.8600 ;
        RECT 225.6500 1622.0600 226.6500 1622.5400 ;
        RECT 225.6500 1627.5000 226.6500 1627.9800 ;
        RECT 225.6500 1643.8200 226.6500 1644.3000 ;
        RECT 225.6500 1605.7400 226.6500 1606.2200 ;
        RECT 225.6500 1611.1800 226.6500 1611.6600 ;
        RECT 225.6500 1589.4200 226.6500 1589.9000 ;
        RECT 225.6500 1594.8600 226.6500 1595.3400 ;
        RECT 225.6500 1600.3000 226.6500 1600.7800 ;
        RECT 225.6500 1578.5400 226.6500 1579.0200 ;
        RECT 225.6500 1583.9800 226.6500 1584.4600 ;
        RECT 225.6500 1562.2200 226.6500 1562.7000 ;
        RECT 225.6500 1567.6600 226.6500 1568.1400 ;
        RECT 225.6500 1573.1000 226.6500 1573.5800 ;
        RECT 225.6500 1616.6200 226.6500 1617.1000 ;
        RECT 163.5100 1660.1400 164.5100 1660.6200 ;
        RECT 163.5100 1649.2600 164.5100 1649.7400 ;
        RECT 163.5100 1654.7000 164.5100 1655.1800 ;
        RECT 163.5100 1632.9400 164.5100 1633.4200 ;
        RECT 163.5100 1638.3800 164.5100 1638.8600 ;
        RECT 163.5100 1622.0600 164.5100 1622.5400 ;
        RECT 163.5100 1627.5000 164.5100 1627.9800 ;
        RECT 163.5100 1643.8200 164.5100 1644.3000 ;
        RECT 163.5100 1605.7400 164.5100 1606.2200 ;
        RECT 163.5100 1611.1800 164.5100 1611.6600 ;
        RECT 163.5100 1589.4200 164.5100 1589.9000 ;
        RECT 163.5100 1594.8600 164.5100 1595.3400 ;
        RECT 163.5100 1600.3000 164.5100 1600.7800 ;
        RECT 163.5100 1578.5400 164.5100 1579.0200 ;
        RECT 163.5100 1583.9800 164.5100 1584.4600 ;
        RECT 163.5100 1562.2200 164.5100 1562.7000 ;
        RECT 163.5100 1567.6600 164.5100 1568.1400 ;
        RECT 163.5100 1573.1000 164.5100 1573.5800 ;
        RECT 163.5100 1616.6200 164.5100 1617.1000 ;
        RECT 225.6500 1551.3400 226.6500 1551.8200 ;
        RECT 225.6500 1556.7800 226.6500 1557.2600 ;
        RECT 225.6500 1535.0200 226.6500 1535.5000 ;
        RECT 225.6500 1540.4600 226.6500 1540.9400 ;
        RECT 225.6500 1545.9000 226.6500 1546.3800 ;
        RECT 225.6500 1524.1400 226.6500 1524.6200 ;
        RECT 225.6500 1529.5800 226.6500 1530.0600 ;
        RECT 225.6500 1507.8200 226.6500 1508.3000 ;
        RECT 225.6500 1513.2600 226.6500 1513.7400 ;
        RECT 225.6500 1518.7000 226.6500 1519.1800 ;
        RECT 225.6500 1496.9400 226.6500 1497.4200 ;
        RECT 225.6500 1502.3800 226.6500 1502.8600 ;
        RECT 225.6500 1480.6200 226.6500 1481.1000 ;
        RECT 225.6500 1486.0600 226.6500 1486.5400 ;
        RECT 225.6500 1491.5000 226.6500 1491.9800 ;
        RECT 225.6500 1469.7400 226.6500 1470.2200 ;
        RECT 225.6500 1475.1800 226.6500 1475.6600 ;
        RECT 225.6500 1464.3000 226.6500 1464.7800 ;
        RECT 163.5100 1551.3400 164.5100 1551.8200 ;
        RECT 163.5100 1556.7800 164.5100 1557.2600 ;
        RECT 163.5100 1535.0200 164.5100 1535.5000 ;
        RECT 163.5100 1540.4600 164.5100 1540.9400 ;
        RECT 163.5100 1545.9000 164.5100 1546.3800 ;
        RECT 163.5100 1524.1400 164.5100 1524.6200 ;
        RECT 163.5100 1529.5800 164.5100 1530.0600 ;
        RECT 163.5100 1507.8200 164.5100 1508.3000 ;
        RECT 163.5100 1513.2600 164.5100 1513.7400 ;
        RECT 163.5100 1518.7000 164.5100 1519.1800 ;
        RECT 163.5100 1496.9400 164.5100 1497.4200 ;
        RECT 163.5100 1502.3800 164.5100 1502.8600 ;
        RECT 163.5100 1480.6200 164.5100 1481.1000 ;
        RECT 163.5100 1486.0600 164.5100 1486.5400 ;
        RECT 163.5100 1491.5000 164.5100 1491.9800 ;
        RECT 163.5100 1469.7400 164.5100 1470.2200 ;
        RECT 163.5100 1475.1800 164.5100 1475.6600 ;
        RECT 163.5100 1464.3000 164.5100 1464.7800 ;
        RECT 163.5100 1664.5900 226.6500 1665.5900 ;
        RECT 163.5100 1457.2900 226.6500 1458.2900 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 1227.6500 226.6500 1435.9500 ;
        RECT 163.5100 1227.6500 164.5100 1435.9500 ;
      LAYER met3 ;
        RECT 225.6500 1430.5000 226.6500 1430.9800 ;
        RECT 225.6500 1419.6200 226.6500 1420.1000 ;
        RECT 225.6500 1425.0600 226.6500 1425.5400 ;
        RECT 225.6500 1403.3000 226.6500 1403.7800 ;
        RECT 225.6500 1408.7400 226.6500 1409.2200 ;
        RECT 225.6500 1392.4200 226.6500 1392.9000 ;
        RECT 225.6500 1397.8600 226.6500 1398.3400 ;
        RECT 225.6500 1414.1800 226.6500 1414.6600 ;
        RECT 225.6500 1376.1000 226.6500 1376.5800 ;
        RECT 225.6500 1381.5400 226.6500 1382.0200 ;
        RECT 225.6500 1359.7800 226.6500 1360.2600 ;
        RECT 225.6500 1365.2200 226.6500 1365.7000 ;
        RECT 225.6500 1370.6600 226.6500 1371.1400 ;
        RECT 225.6500 1348.9000 226.6500 1349.3800 ;
        RECT 225.6500 1354.3400 226.6500 1354.8200 ;
        RECT 225.6500 1332.5800 226.6500 1333.0600 ;
        RECT 225.6500 1338.0200 226.6500 1338.5000 ;
        RECT 225.6500 1343.4600 226.6500 1343.9400 ;
        RECT 225.6500 1386.9800 226.6500 1387.4600 ;
        RECT 163.5100 1430.5000 164.5100 1430.9800 ;
        RECT 163.5100 1419.6200 164.5100 1420.1000 ;
        RECT 163.5100 1425.0600 164.5100 1425.5400 ;
        RECT 163.5100 1403.3000 164.5100 1403.7800 ;
        RECT 163.5100 1408.7400 164.5100 1409.2200 ;
        RECT 163.5100 1392.4200 164.5100 1392.9000 ;
        RECT 163.5100 1397.8600 164.5100 1398.3400 ;
        RECT 163.5100 1414.1800 164.5100 1414.6600 ;
        RECT 163.5100 1376.1000 164.5100 1376.5800 ;
        RECT 163.5100 1381.5400 164.5100 1382.0200 ;
        RECT 163.5100 1359.7800 164.5100 1360.2600 ;
        RECT 163.5100 1365.2200 164.5100 1365.7000 ;
        RECT 163.5100 1370.6600 164.5100 1371.1400 ;
        RECT 163.5100 1348.9000 164.5100 1349.3800 ;
        RECT 163.5100 1354.3400 164.5100 1354.8200 ;
        RECT 163.5100 1332.5800 164.5100 1333.0600 ;
        RECT 163.5100 1338.0200 164.5100 1338.5000 ;
        RECT 163.5100 1343.4600 164.5100 1343.9400 ;
        RECT 163.5100 1386.9800 164.5100 1387.4600 ;
        RECT 225.6500 1321.7000 226.6500 1322.1800 ;
        RECT 225.6500 1327.1400 226.6500 1327.6200 ;
        RECT 225.6500 1305.3800 226.6500 1305.8600 ;
        RECT 225.6500 1310.8200 226.6500 1311.3000 ;
        RECT 225.6500 1316.2600 226.6500 1316.7400 ;
        RECT 225.6500 1294.5000 226.6500 1294.9800 ;
        RECT 225.6500 1299.9400 226.6500 1300.4200 ;
        RECT 225.6500 1278.1800 226.6500 1278.6600 ;
        RECT 225.6500 1283.6200 226.6500 1284.1000 ;
        RECT 225.6500 1289.0600 226.6500 1289.5400 ;
        RECT 225.6500 1267.3000 226.6500 1267.7800 ;
        RECT 225.6500 1272.7400 226.6500 1273.2200 ;
        RECT 225.6500 1250.9800 226.6500 1251.4600 ;
        RECT 225.6500 1256.4200 226.6500 1256.9000 ;
        RECT 225.6500 1261.8600 226.6500 1262.3400 ;
        RECT 225.6500 1240.1000 226.6500 1240.5800 ;
        RECT 225.6500 1245.5400 226.6500 1246.0200 ;
        RECT 225.6500 1234.6600 226.6500 1235.1400 ;
        RECT 163.5100 1321.7000 164.5100 1322.1800 ;
        RECT 163.5100 1327.1400 164.5100 1327.6200 ;
        RECT 163.5100 1305.3800 164.5100 1305.8600 ;
        RECT 163.5100 1310.8200 164.5100 1311.3000 ;
        RECT 163.5100 1316.2600 164.5100 1316.7400 ;
        RECT 163.5100 1294.5000 164.5100 1294.9800 ;
        RECT 163.5100 1299.9400 164.5100 1300.4200 ;
        RECT 163.5100 1278.1800 164.5100 1278.6600 ;
        RECT 163.5100 1283.6200 164.5100 1284.1000 ;
        RECT 163.5100 1289.0600 164.5100 1289.5400 ;
        RECT 163.5100 1267.3000 164.5100 1267.7800 ;
        RECT 163.5100 1272.7400 164.5100 1273.2200 ;
        RECT 163.5100 1250.9800 164.5100 1251.4600 ;
        RECT 163.5100 1256.4200 164.5100 1256.9000 ;
        RECT 163.5100 1261.8600 164.5100 1262.3400 ;
        RECT 163.5100 1240.1000 164.5100 1240.5800 ;
        RECT 163.5100 1245.5400 164.5100 1246.0200 ;
        RECT 163.5100 1234.6600 164.5100 1235.1400 ;
        RECT 163.5100 1434.9500 226.6500 1435.9500 ;
        RECT 163.5100 1227.6500 226.6500 1228.6500 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 998.0100 226.6500 1206.3100 ;
        RECT 163.5100 998.0100 164.5100 1206.3100 ;
      LAYER met3 ;
        RECT 225.6500 1200.8600 226.6500 1201.3400 ;
        RECT 225.6500 1189.9800 226.6500 1190.4600 ;
        RECT 225.6500 1195.4200 226.6500 1195.9000 ;
        RECT 225.6500 1173.6600 226.6500 1174.1400 ;
        RECT 225.6500 1179.1000 226.6500 1179.5800 ;
        RECT 225.6500 1162.7800 226.6500 1163.2600 ;
        RECT 225.6500 1168.2200 226.6500 1168.7000 ;
        RECT 225.6500 1184.5400 226.6500 1185.0200 ;
        RECT 225.6500 1146.4600 226.6500 1146.9400 ;
        RECT 225.6500 1151.9000 226.6500 1152.3800 ;
        RECT 225.6500 1130.1400 226.6500 1130.6200 ;
        RECT 225.6500 1135.5800 226.6500 1136.0600 ;
        RECT 225.6500 1141.0200 226.6500 1141.5000 ;
        RECT 225.6500 1119.2600 226.6500 1119.7400 ;
        RECT 225.6500 1124.7000 226.6500 1125.1800 ;
        RECT 225.6500 1102.9400 226.6500 1103.4200 ;
        RECT 225.6500 1108.3800 226.6500 1108.8600 ;
        RECT 225.6500 1113.8200 226.6500 1114.3000 ;
        RECT 225.6500 1157.3400 226.6500 1157.8200 ;
        RECT 163.5100 1200.8600 164.5100 1201.3400 ;
        RECT 163.5100 1189.9800 164.5100 1190.4600 ;
        RECT 163.5100 1195.4200 164.5100 1195.9000 ;
        RECT 163.5100 1173.6600 164.5100 1174.1400 ;
        RECT 163.5100 1179.1000 164.5100 1179.5800 ;
        RECT 163.5100 1162.7800 164.5100 1163.2600 ;
        RECT 163.5100 1168.2200 164.5100 1168.7000 ;
        RECT 163.5100 1184.5400 164.5100 1185.0200 ;
        RECT 163.5100 1146.4600 164.5100 1146.9400 ;
        RECT 163.5100 1151.9000 164.5100 1152.3800 ;
        RECT 163.5100 1130.1400 164.5100 1130.6200 ;
        RECT 163.5100 1135.5800 164.5100 1136.0600 ;
        RECT 163.5100 1141.0200 164.5100 1141.5000 ;
        RECT 163.5100 1119.2600 164.5100 1119.7400 ;
        RECT 163.5100 1124.7000 164.5100 1125.1800 ;
        RECT 163.5100 1102.9400 164.5100 1103.4200 ;
        RECT 163.5100 1108.3800 164.5100 1108.8600 ;
        RECT 163.5100 1113.8200 164.5100 1114.3000 ;
        RECT 163.5100 1157.3400 164.5100 1157.8200 ;
        RECT 225.6500 1092.0600 226.6500 1092.5400 ;
        RECT 225.6500 1097.5000 226.6500 1097.9800 ;
        RECT 225.6500 1075.7400 226.6500 1076.2200 ;
        RECT 225.6500 1081.1800 226.6500 1081.6600 ;
        RECT 225.6500 1086.6200 226.6500 1087.1000 ;
        RECT 225.6500 1064.8600 226.6500 1065.3400 ;
        RECT 225.6500 1070.3000 226.6500 1070.7800 ;
        RECT 225.6500 1048.5400 226.6500 1049.0200 ;
        RECT 225.6500 1053.9800 226.6500 1054.4600 ;
        RECT 225.6500 1059.4200 226.6500 1059.9000 ;
        RECT 225.6500 1037.6600 226.6500 1038.1400 ;
        RECT 225.6500 1043.1000 226.6500 1043.5800 ;
        RECT 225.6500 1021.3400 226.6500 1021.8200 ;
        RECT 225.6500 1026.7800 226.6500 1027.2600 ;
        RECT 225.6500 1032.2200 226.6500 1032.7000 ;
        RECT 225.6500 1010.4600 226.6500 1010.9400 ;
        RECT 225.6500 1015.9000 226.6500 1016.3800 ;
        RECT 225.6500 1005.0200 226.6500 1005.5000 ;
        RECT 163.5100 1092.0600 164.5100 1092.5400 ;
        RECT 163.5100 1097.5000 164.5100 1097.9800 ;
        RECT 163.5100 1075.7400 164.5100 1076.2200 ;
        RECT 163.5100 1081.1800 164.5100 1081.6600 ;
        RECT 163.5100 1086.6200 164.5100 1087.1000 ;
        RECT 163.5100 1064.8600 164.5100 1065.3400 ;
        RECT 163.5100 1070.3000 164.5100 1070.7800 ;
        RECT 163.5100 1048.5400 164.5100 1049.0200 ;
        RECT 163.5100 1053.9800 164.5100 1054.4600 ;
        RECT 163.5100 1059.4200 164.5100 1059.9000 ;
        RECT 163.5100 1037.6600 164.5100 1038.1400 ;
        RECT 163.5100 1043.1000 164.5100 1043.5800 ;
        RECT 163.5100 1021.3400 164.5100 1021.8200 ;
        RECT 163.5100 1026.7800 164.5100 1027.2600 ;
        RECT 163.5100 1032.2200 164.5100 1032.7000 ;
        RECT 163.5100 1010.4600 164.5100 1010.9400 ;
        RECT 163.5100 1015.9000 164.5100 1016.3800 ;
        RECT 163.5100 1005.0200 164.5100 1005.5000 ;
        RECT 163.5100 1205.3100 226.6500 1206.3100 ;
        RECT 163.5100 998.0100 226.6500 999.0100 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 225.6500 768.3700 226.6500 976.6700 ;
        RECT 163.5100 768.3700 164.5100 976.6700 ;
      LAYER met3 ;
        RECT 225.6500 971.2200 226.6500 971.7000 ;
        RECT 225.6500 960.3400 226.6500 960.8200 ;
        RECT 225.6500 965.7800 226.6500 966.2600 ;
        RECT 225.6500 944.0200 226.6500 944.5000 ;
        RECT 225.6500 949.4600 226.6500 949.9400 ;
        RECT 225.6500 933.1400 226.6500 933.6200 ;
        RECT 225.6500 938.5800 226.6500 939.0600 ;
        RECT 225.6500 954.9000 226.6500 955.3800 ;
        RECT 225.6500 916.8200 226.6500 917.3000 ;
        RECT 225.6500 922.2600 226.6500 922.7400 ;
        RECT 225.6500 900.5000 226.6500 900.9800 ;
        RECT 225.6500 905.9400 226.6500 906.4200 ;
        RECT 225.6500 911.3800 226.6500 911.8600 ;
        RECT 225.6500 889.6200 226.6500 890.1000 ;
        RECT 225.6500 895.0600 226.6500 895.5400 ;
        RECT 225.6500 873.3000 226.6500 873.7800 ;
        RECT 225.6500 878.7400 226.6500 879.2200 ;
        RECT 225.6500 884.1800 226.6500 884.6600 ;
        RECT 225.6500 927.7000 226.6500 928.1800 ;
        RECT 163.5100 971.2200 164.5100 971.7000 ;
        RECT 163.5100 960.3400 164.5100 960.8200 ;
        RECT 163.5100 965.7800 164.5100 966.2600 ;
        RECT 163.5100 944.0200 164.5100 944.5000 ;
        RECT 163.5100 949.4600 164.5100 949.9400 ;
        RECT 163.5100 933.1400 164.5100 933.6200 ;
        RECT 163.5100 938.5800 164.5100 939.0600 ;
        RECT 163.5100 954.9000 164.5100 955.3800 ;
        RECT 163.5100 916.8200 164.5100 917.3000 ;
        RECT 163.5100 922.2600 164.5100 922.7400 ;
        RECT 163.5100 900.5000 164.5100 900.9800 ;
        RECT 163.5100 905.9400 164.5100 906.4200 ;
        RECT 163.5100 911.3800 164.5100 911.8600 ;
        RECT 163.5100 889.6200 164.5100 890.1000 ;
        RECT 163.5100 895.0600 164.5100 895.5400 ;
        RECT 163.5100 873.3000 164.5100 873.7800 ;
        RECT 163.5100 878.7400 164.5100 879.2200 ;
        RECT 163.5100 884.1800 164.5100 884.6600 ;
        RECT 163.5100 927.7000 164.5100 928.1800 ;
        RECT 225.6500 862.4200 226.6500 862.9000 ;
        RECT 225.6500 867.8600 226.6500 868.3400 ;
        RECT 225.6500 846.1000 226.6500 846.5800 ;
        RECT 225.6500 851.5400 226.6500 852.0200 ;
        RECT 225.6500 856.9800 226.6500 857.4600 ;
        RECT 225.6500 835.2200 226.6500 835.7000 ;
        RECT 225.6500 840.6600 226.6500 841.1400 ;
        RECT 225.6500 818.9000 226.6500 819.3800 ;
        RECT 225.6500 824.3400 226.6500 824.8200 ;
        RECT 225.6500 829.7800 226.6500 830.2600 ;
        RECT 225.6500 808.0200 226.6500 808.5000 ;
        RECT 225.6500 813.4600 226.6500 813.9400 ;
        RECT 225.6500 791.7000 226.6500 792.1800 ;
        RECT 225.6500 797.1400 226.6500 797.6200 ;
        RECT 225.6500 802.5800 226.6500 803.0600 ;
        RECT 225.6500 780.8200 226.6500 781.3000 ;
        RECT 225.6500 786.2600 226.6500 786.7400 ;
        RECT 225.6500 775.3800 226.6500 775.8600 ;
        RECT 163.5100 862.4200 164.5100 862.9000 ;
        RECT 163.5100 867.8600 164.5100 868.3400 ;
        RECT 163.5100 846.1000 164.5100 846.5800 ;
        RECT 163.5100 851.5400 164.5100 852.0200 ;
        RECT 163.5100 856.9800 164.5100 857.4600 ;
        RECT 163.5100 835.2200 164.5100 835.7000 ;
        RECT 163.5100 840.6600 164.5100 841.1400 ;
        RECT 163.5100 818.9000 164.5100 819.3800 ;
        RECT 163.5100 824.3400 164.5100 824.8200 ;
        RECT 163.5100 829.7800 164.5100 830.2600 ;
        RECT 163.5100 808.0200 164.5100 808.5000 ;
        RECT 163.5100 813.4600 164.5100 813.9400 ;
        RECT 163.5100 791.7000 164.5100 792.1800 ;
        RECT 163.5100 797.1400 164.5100 797.6200 ;
        RECT 163.5100 802.5800 164.5100 803.0600 ;
        RECT 163.5100 780.8200 164.5100 781.3000 ;
        RECT 163.5100 786.2600 164.5100 786.7400 ;
        RECT 163.5100 775.3800 164.5100 775.8600 ;
        RECT 163.5100 975.6700 226.6500 976.6700 ;
        RECT 163.5100 768.3700 226.6500 769.3700 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 2257.5600 2833.6100 2259.5600 2854.5400 ;
        RECT 2454.6600 2833.6100 2456.6600 2854.5400 ;
      LAYER met3 ;
        RECT 2454.6600 2850.0400 2456.6600 2850.5200 ;
        RECT 2257.5600 2850.0400 2259.5600 2850.5200 ;
        RECT 2454.6600 2839.1600 2456.6600 2839.6400 ;
        RECT 2257.5600 2839.1600 2259.5600 2839.6400 ;
        RECT 2454.6600 2844.6000 2456.6600 2845.0800 ;
        RECT 2257.5600 2844.6000 2259.5600 2845.0800 ;
        RECT 2257.5600 2852.5400 2456.6600 2854.5400 ;
        RECT 2257.5600 2833.6100 2456.6600 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 538.5700 2443.7200 746.6700 ;
        RECT 2397.1200 538.5700 2398.7200 746.6700 ;
        RECT 2352.1200 538.5700 2353.7200 746.6700 ;
        RECT 2307.1200 538.5700 2308.7200 746.6700 ;
        RECT 2453.6600 538.5700 2456.6600 746.6700 ;
        RECT 2257.5600 538.5700 2260.5600 746.6700 ;
      LAYER met3 ;
        RECT 2453.6600 741.3200 2456.6600 741.8000 ;
        RECT 2442.1200 741.3200 2443.7200 741.8000 ;
        RECT 2453.6600 730.4400 2456.6600 730.9200 ;
        RECT 2453.6600 735.8800 2456.6600 736.3600 ;
        RECT 2442.1200 730.4400 2443.7200 730.9200 ;
        RECT 2442.1200 735.8800 2443.7200 736.3600 ;
        RECT 2453.6600 714.1200 2456.6600 714.6000 ;
        RECT 2453.6600 719.5600 2456.6600 720.0400 ;
        RECT 2442.1200 714.1200 2443.7200 714.6000 ;
        RECT 2442.1200 719.5600 2443.7200 720.0400 ;
        RECT 2453.6600 703.2400 2456.6600 703.7200 ;
        RECT 2453.6600 708.6800 2456.6600 709.1600 ;
        RECT 2442.1200 703.2400 2443.7200 703.7200 ;
        RECT 2442.1200 708.6800 2443.7200 709.1600 ;
        RECT 2453.6600 725.0000 2456.6600 725.4800 ;
        RECT 2442.1200 725.0000 2443.7200 725.4800 ;
        RECT 2397.1200 730.4400 2398.7200 730.9200 ;
        RECT 2397.1200 735.8800 2398.7200 736.3600 ;
        RECT 2397.1200 741.3200 2398.7200 741.8000 ;
        RECT 2397.1200 714.1200 2398.7200 714.6000 ;
        RECT 2397.1200 719.5600 2398.7200 720.0400 ;
        RECT 2397.1200 708.6800 2398.7200 709.1600 ;
        RECT 2397.1200 703.2400 2398.7200 703.7200 ;
        RECT 2397.1200 725.0000 2398.7200 725.4800 ;
        RECT 2453.6600 686.9200 2456.6600 687.4000 ;
        RECT 2453.6600 692.3600 2456.6600 692.8400 ;
        RECT 2442.1200 686.9200 2443.7200 687.4000 ;
        RECT 2442.1200 692.3600 2443.7200 692.8400 ;
        RECT 2453.6600 670.6000 2456.6600 671.0800 ;
        RECT 2453.6600 676.0400 2456.6600 676.5200 ;
        RECT 2453.6600 681.4800 2456.6600 681.9600 ;
        RECT 2442.1200 670.6000 2443.7200 671.0800 ;
        RECT 2442.1200 676.0400 2443.7200 676.5200 ;
        RECT 2442.1200 681.4800 2443.7200 681.9600 ;
        RECT 2453.6600 659.7200 2456.6600 660.2000 ;
        RECT 2453.6600 665.1600 2456.6600 665.6400 ;
        RECT 2442.1200 659.7200 2443.7200 660.2000 ;
        RECT 2442.1200 665.1600 2443.7200 665.6400 ;
        RECT 2453.6600 643.4000 2456.6600 643.8800 ;
        RECT 2453.6600 648.8400 2456.6600 649.3200 ;
        RECT 2453.6600 654.2800 2456.6600 654.7600 ;
        RECT 2442.1200 643.4000 2443.7200 643.8800 ;
        RECT 2442.1200 648.8400 2443.7200 649.3200 ;
        RECT 2442.1200 654.2800 2443.7200 654.7600 ;
        RECT 2397.1200 686.9200 2398.7200 687.4000 ;
        RECT 2397.1200 692.3600 2398.7200 692.8400 ;
        RECT 2397.1200 670.6000 2398.7200 671.0800 ;
        RECT 2397.1200 676.0400 2398.7200 676.5200 ;
        RECT 2397.1200 681.4800 2398.7200 681.9600 ;
        RECT 2397.1200 659.7200 2398.7200 660.2000 ;
        RECT 2397.1200 665.1600 2398.7200 665.6400 ;
        RECT 2397.1200 643.4000 2398.7200 643.8800 ;
        RECT 2397.1200 648.8400 2398.7200 649.3200 ;
        RECT 2397.1200 654.2800 2398.7200 654.7600 ;
        RECT 2453.6600 697.8000 2456.6600 698.2800 ;
        RECT 2397.1200 697.8000 2398.7200 698.2800 ;
        RECT 2442.1200 697.8000 2443.7200 698.2800 ;
        RECT 2352.1200 730.4400 2353.7200 730.9200 ;
        RECT 2352.1200 735.8800 2353.7200 736.3600 ;
        RECT 2352.1200 741.3200 2353.7200 741.8000 ;
        RECT 2307.1200 730.4400 2308.7200 730.9200 ;
        RECT 2307.1200 735.8800 2308.7200 736.3600 ;
        RECT 2307.1200 741.3200 2308.7200 741.8000 ;
        RECT 2352.1200 714.1200 2353.7200 714.6000 ;
        RECT 2352.1200 719.5600 2353.7200 720.0400 ;
        RECT 2352.1200 703.2400 2353.7200 703.7200 ;
        RECT 2352.1200 708.6800 2353.7200 709.1600 ;
        RECT 2307.1200 714.1200 2308.7200 714.6000 ;
        RECT 2307.1200 719.5600 2308.7200 720.0400 ;
        RECT 2307.1200 703.2400 2308.7200 703.7200 ;
        RECT 2307.1200 708.6800 2308.7200 709.1600 ;
        RECT 2307.1200 725.0000 2308.7200 725.4800 ;
        RECT 2352.1200 725.0000 2353.7200 725.4800 ;
        RECT 2257.5600 741.3200 2260.5600 741.8000 ;
        RECT 2257.5600 735.8800 2260.5600 736.3600 ;
        RECT 2257.5600 730.4400 2260.5600 730.9200 ;
        RECT 2257.5600 719.5600 2260.5600 720.0400 ;
        RECT 2257.5600 714.1200 2260.5600 714.6000 ;
        RECT 2257.5600 708.6800 2260.5600 709.1600 ;
        RECT 2257.5600 703.2400 2260.5600 703.7200 ;
        RECT 2257.5600 725.0000 2260.5600 725.4800 ;
        RECT 2352.1200 686.9200 2353.7200 687.4000 ;
        RECT 2352.1200 692.3600 2353.7200 692.8400 ;
        RECT 2352.1200 670.6000 2353.7200 671.0800 ;
        RECT 2352.1200 676.0400 2353.7200 676.5200 ;
        RECT 2352.1200 681.4800 2353.7200 681.9600 ;
        RECT 2307.1200 686.9200 2308.7200 687.4000 ;
        RECT 2307.1200 692.3600 2308.7200 692.8400 ;
        RECT 2307.1200 670.6000 2308.7200 671.0800 ;
        RECT 2307.1200 676.0400 2308.7200 676.5200 ;
        RECT 2307.1200 681.4800 2308.7200 681.9600 ;
        RECT 2352.1200 659.7200 2353.7200 660.2000 ;
        RECT 2352.1200 665.1600 2353.7200 665.6400 ;
        RECT 2352.1200 643.4000 2353.7200 643.8800 ;
        RECT 2352.1200 648.8400 2353.7200 649.3200 ;
        RECT 2352.1200 654.2800 2353.7200 654.7600 ;
        RECT 2307.1200 659.7200 2308.7200 660.2000 ;
        RECT 2307.1200 665.1600 2308.7200 665.6400 ;
        RECT 2307.1200 643.4000 2308.7200 643.8800 ;
        RECT 2307.1200 648.8400 2308.7200 649.3200 ;
        RECT 2307.1200 654.2800 2308.7200 654.7600 ;
        RECT 2257.5600 686.9200 2260.5600 687.4000 ;
        RECT 2257.5600 692.3600 2260.5600 692.8400 ;
        RECT 2257.5600 676.0400 2260.5600 676.5200 ;
        RECT 2257.5600 670.6000 2260.5600 671.0800 ;
        RECT 2257.5600 681.4800 2260.5600 681.9600 ;
        RECT 2257.5600 659.7200 2260.5600 660.2000 ;
        RECT 2257.5600 665.1600 2260.5600 665.6400 ;
        RECT 2257.5600 648.8400 2260.5600 649.3200 ;
        RECT 2257.5600 643.4000 2260.5600 643.8800 ;
        RECT 2257.5600 654.2800 2260.5600 654.7600 ;
        RECT 2257.5600 697.8000 2260.5600 698.2800 ;
        RECT 2307.1200 697.8000 2308.7200 698.2800 ;
        RECT 2352.1200 697.8000 2353.7200 698.2800 ;
        RECT 2453.6600 632.5200 2456.6600 633.0000 ;
        RECT 2453.6600 637.9600 2456.6600 638.4400 ;
        RECT 2442.1200 632.5200 2443.7200 633.0000 ;
        RECT 2442.1200 637.9600 2443.7200 638.4400 ;
        RECT 2453.6600 616.2000 2456.6600 616.6800 ;
        RECT 2453.6600 621.6400 2456.6600 622.1200 ;
        RECT 2453.6600 627.0800 2456.6600 627.5600 ;
        RECT 2442.1200 616.2000 2443.7200 616.6800 ;
        RECT 2442.1200 621.6400 2443.7200 622.1200 ;
        RECT 2442.1200 627.0800 2443.7200 627.5600 ;
        RECT 2453.6600 605.3200 2456.6600 605.8000 ;
        RECT 2453.6600 610.7600 2456.6600 611.2400 ;
        RECT 2442.1200 605.3200 2443.7200 605.8000 ;
        RECT 2442.1200 610.7600 2443.7200 611.2400 ;
        RECT 2453.6600 589.0000 2456.6600 589.4800 ;
        RECT 2453.6600 594.4400 2456.6600 594.9200 ;
        RECT 2453.6600 599.8800 2456.6600 600.3600 ;
        RECT 2442.1200 589.0000 2443.7200 589.4800 ;
        RECT 2442.1200 594.4400 2443.7200 594.9200 ;
        RECT 2442.1200 599.8800 2443.7200 600.3600 ;
        RECT 2397.1200 632.5200 2398.7200 633.0000 ;
        RECT 2397.1200 637.9600 2398.7200 638.4400 ;
        RECT 2397.1200 616.2000 2398.7200 616.6800 ;
        RECT 2397.1200 621.6400 2398.7200 622.1200 ;
        RECT 2397.1200 627.0800 2398.7200 627.5600 ;
        RECT 2397.1200 605.3200 2398.7200 605.8000 ;
        RECT 2397.1200 610.7600 2398.7200 611.2400 ;
        RECT 2397.1200 589.0000 2398.7200 589.4800 ;
        RECT 2397.1200 594.4400 2398.7200 594.9200 ;
        RECT 2397.1200 599.8800 2398.7200 600.3600 ;
        RECT 2453.6600 578.1200 2456.6600 578.6000 ;
        RECT 2453.6600 583.5600 2456.6600 584.0400 ;
        RECT 2442.1200 578.1200 2443.7200 578.6000 ;
        RECT 2442.1200 583.5600 2443.7200 584.0400 ;
        RECT 2453.6600 561.8000 2456.6600 562.2800 ;
        RECT 2453.6600 567.2400 2456.6600 567.7200 ;
        RECT 2453.6600 572.6800 2456.6600 573.1600 ;
        RECT 2442.1200 561.8000 2443.7200 562.2800 ;
        RECT 2442.1200 567.2400 2443.7200 567.7200 ;
        RECT 2442.1200 572.6800 2443.7200 573.1600 ;
        RECT 2453.6600 550.9200 2456.6600 551.4000 ;
        RECT 2453.6600 556.3600 2456.6600 556.8400 ;
        RECT 2442.1200 550.9200 2443.7200 551.4000 ;
        RECT 2442.1200 556.3600 2443.7200 556.8400 ;
        RECT 2453.6600 545.4800 2456.6600 545.9600 ;
        RECT 2442.1200 545.4800 2443.7200 545.9600 ;
        RECT 2397.1200 578.1200 2398.7200 578.6000 ;
        RECT 2397.1200 583.5600 2398.7200 584.0400 ;
        RECT 2397.1200 561.8000 2398.7200 562.2800 ;
        RECT 2397.1200 567.2400 2398.7200 567.7200 ;
        RECT 2397.1200 572.6800 2398.7200 573.1600 ;
        RECT 2397.1200 550.9200 2398.7200 551.4000 ;
        RECT 2397.1200 556.3600 2398.7200 556.8400 ;
        RECT 2397.1200 545.4800 2398.7200 545.9600 ;
        RECT 2352.1200 632.5200 2353.7200 633.0000 ;
        RECT 2352.1200 637.9600 2353.7200 638.4400 ;
        RECT 2352.1200 616.2000 2353.7200 616.6800 ;
        RECT 2352.1200 621.6400 2353.7200 622.1200 ;
        RECT 2352.1200 627.0800 2353.7200 627.5600 ;
        RECT 2307.1200 632.5200 2308.7200 633.0000 ;
        RECT 2307.1200 637.9600 2308.7200 638.4400 ;
        RECT 2307.1200 616.2000 2308.7200 616.6800 ;
        RECT 2307.1200 621.6400 2308.7200 622.1200 ;
        RECT 2307.1200 627.0800 2308.7200 627.5600 ;
        RECT 2352.1200 605.3200 2353.7200 605.8000 ;
        RECT 2352.1200 610.7600 2353.7200 611.2400 ;
        RECT 2352.1200 589.0000 2353.7200 589.4800 ;
        RECT 2352.1200 594.4400 2353.7200 594.9200 ;
        RECT 2352.1200 599.8800 2353.7200 600.3600 ;
        RECT 2307.1200 605.3200 2308.7200 605.8000 ;
        RECT 2307.1200 610.7600 2308.7200 611.2400 ;
        RECT 2307.1200 589.0000 2308.7200 589.4800 ;
        RECT 2307.1200 594.4400 2308.7200 594.9200 ;
        RECT 2307.1200 599.8800 2308.7200 600.3600 ;
        RECT 2257.5600 632.5200 2260.5600 633.0000 ;
        RECT 2257.5600 637.9600 2260.5600 638.4400 ;
        RECT 2257.5600 621.6400 2260.5600 622.1200 ;
        RECT 2257.5600 616.2000 2260.5600 616.6800 ;
        RECT 2257.5600 627.0800 2260.5600 627.5600 ;
        RECT 2257.5600 605.3200 2260.5600 605.8000 ;
        RECT 2257.5600 610.7600 2260.5600 611.2400 ;
        RECT 2257.5600 594.4400 2260.5600 594.9200 ;
        RECT 2257.5600 589.0000 2260.5600 589.4800 ;
        RECT 2257.5600 599.8800 2260.5600 600.3600 ;
        RECT 2352.1200 578.1200 2353.7200 578.6000 ;
        RECT 2352.1200 583.5600 2353.7200 584.0400 ;
        RECT 2352.1200 561.8000 2353.7200 562.2800 ;
        RECT 2352.1200 567.2400 2353.7200 567.7200 ;
        RECT 2352.1200 572.6800 2353.7200 573.1600 ;
        RECT 2307.1200 578.1200 2308.7200 578.6000 ;
        RECT 2307.1200 583.5600 2308.7200 584.0400 ;
        RECT 2307.1200 561.8000 2308.7200 562.2800 ;
        RECT 2307.1200 567.2400 2308.7200 567.7200 ;
        RECT 2307.1200 572.6800 2308.7200 573.1600 ;
        RECT 2352.1200 556.3600 2353.7200 556.8400 ;
        RECT 2352.1200 550.9200 2353.7200 551.4000 ;
        RECT 2352.1200 545.4800 2353.7200 545.9600 ;
        RECT 2307.1200 556.3600 2308.7200 556.8400 ;
        RECT 2307.1200 550.9200 2308.7200 551.4000 ;
        RECT 2307.1200 545.4800 2308.7200 545.9600 ;
        RECT 2257.5600 578.1200 2260.5600 578.6000 ;
        RECT 2257.5600 583.5600 2260.5600 584.0400 ;
        RECT 2257.5600 567.2400 2260.5600 567.7200 ;
        RECT 2257.5600 561.8000 2260.5600 562.2800 ;
        RECT 2257.5600 572.6800 2260.5600 573.1600 ;
        RECT 2257.5600 550.9200 2260.5600 551.4000 ;
        RECT 2257.5600 556.3600 2260.5600 556.8400 ;
        RECT 2257.5600 545.4800 2260.5600 545.9600 ;
        RECT 2257.5600 743.6700 2456.6600 746.6700 ;
        RECT 2257.5600 538.5700 2456.6600 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 308.9300 2443.7200 517.0300 ;
        RECT 2397.1200 308.9300 2398.7200 517.0300 ;
        RECT 2352.1200 308.9300 2353.7200 517.0300 ;
        RECT 2307.1200 308.9300 2308.7200 517.0300 ;
        RECT 2453.6600 308.9300 2456.6600 517.0300 ;
        RECT 2257.5600 308.9300 2260.5600 517.0300 ;
      LAYER met3 ;
        RECT 2453.6600 511.6800 2456.6600 512.1600 ;
        RECT 2442.1200 511.6800 2443.7200 512.1600 ;
        RECT 2453.6600 500.8000 2456.6600 501.2800 ;
        RECT 2453.6600 506.2400 2456.6600 506.7200 ;
        RECT 2442.1200 500.8000 2443.7200 501.2800 ;
        RECT 2442.1200 506.2400 2443.7200 506.7200 ;
        RECT 2453.6600 484.4800 2456.6600 484.9600 ;
        RECT 2453.6600 489.9200 2456.6600 490.4000 ;
        RECT 2442.1200 484.4800 2443.7200 484.9600 ;
        RECT 2442.1200 489.9200 2443.7200 490.4000 ;
        RECT 2453.6600 473.6000 2456.6600 474.0800 ;
        RECT 2453.6600 479.0400 2456.6600 479.5200 ;
        RECT 2442.1200 473.6000 2443.7200 474.0800 ;
        RECT 2442.1200 479.0400 2443.7200 479.5200 ;
        RECT 2453.6600 495.3600 2456.6600 495.8400 ;
        RECT 2442.1200 495.3600 2443.7200 495.8400 ;
        RECT 2397.1200 500.8000 2398.7200 501.2800 ;
        RECT 2397.1200 506.2400 2398.7200 506.7200 ;
        RECT 2397.1200 511.6800 2398.7200 512.1600 ;
        RECT 2397.1200 484.4800 2398.7200 484.9600 ;
        RECT 2397.1200 489.9200 2398.7200 490.4000 ;
        RECT 2397.1200 479.0400 2398.7200 479.5200 ;
        RECT 2397.1200 473.6000 2398.7200 474.0800 ;
        RECT 2397.1200 495.3600 2398.7200 495.8400 ;
        RECT 2453.6600 457.2800 2456.6600 457.7600 ;
        RECT 2453.6600 462.7200 2456.6600 463.2000 ;
        RECT 2442.1200 457.2800 2443.7200 457.7600 ;
        RECT 2442.1200 462.7200 2443.7200 463.2000 ;
        RECT 2453.6600 440.9600 2456.6600 441.4400 ;
        RECT 2453.6600 446.4000 2456.6600 446.8800 ;
        RECT 2453.6600 451.8400 2456.6600 452.3200 ;
        RECT 2442.1200 440.9600 2443.7200 441.4400 ;
        RECT 2442.1200 446.4000 2443.7200 446.8800 ;
        RECT 2442.1200 451.8400 2443.7200 452.3200 ;
        RECT 2453.6600 430.0800 2456.6600 430.5600 ;
        RECT 2453.6600 435.5200 2456.6600 436.0000 ;
        RECT 2442.1200 430.0800 2443.7200 430.5600 ;
        RECT 2442.1200 435.5200 2443.7200 436.0000 ;
        RECT 2453.6600 413.7600 2456.6600 414.2400 ;
        RECT 2453.6600 419.2000 2456.6600 419.6800 ;
        RECT 2453.6600 424.6400 2456.6600 425.1200 ;
        RECT 2442.1200 413.7600 2443.7200 414.2400 ;
        RECT 2442.1200 419.2000 2443.7200 419.6800 ;
        RECT 2442.1200 424.6400 2443.7200 425.1200 ;
        RECT 2397.1200 457.2800 2398.7200 457.7600 ;
        RECT 2397.1200 462.7200 2398.7200 463.2000 ;
        RECT 2397.1200 440.9600 2398.7200 441.4400 ;
        RECT 2397.1200 446.4000 2398.7200 446.8800 ;
        RECT 2397.1200 451.8400 2398.7200 452.3200 ;
        RECT 2397.1200 430.0800 2398.7200 430.5600 ;
        RECT 2397.1200 435.5200 2398.7200 436.0000 ;
        RECT 2397.1200 413.7600 2398.7200 414.2400 ;
        RECT 2397.1200 419.2000 2398.7200 419.6800 ;
        RECT 2397.1200 424.6400 2398.7200 425.1200 ;
        RECT 2453.6600 468.1600 2456.6600 468.6400 ;
        RECT 2397.1200 468.1600 2398.7200 468.6400 ;
        RECT 2442.1200 468.1600 2443.7200 468.6400 ;
        RECT 2352.1200 500.8000 2353.7200 501.2800 ;
        RECT 2352.1200 506.2400 2353.7200 506.7200 ;
        RECT 2352.1200 511.6800 2353.7200 512.1600 ;
        RECT 2307.1200 500.8000 2308.7200 501.2800 ;
        RECT 2307.1200 506.2400 2308.7200 506.7200 ;
        RECT 2307.1200 511.6800 2308.7200 512.1600 ;
        RECT 2352.1200 484.4800 2353.7200 484.9600 ;
        RECT 2352.1200 489.9200 2353.7200 490.4000 ;
        RECT 2352.1200 473.6000 2353.7200 474.0800 ;
        RECT 2352.1200 479.0400 2353.7200 479.5200 ;
        RECT 2307.1200 484.4800 2308.7200 484.9600 ;
        RECT 2307.1200 489.9200 2308.7200 490.4000 ;
        RECT 2307.1200 473.6000 2308.7200 474.0800 ;
        RECT 2307.1200 479.0400 2308.7200 479.5200 ;
        RECT 2307.1200 495.3600 2308.7200 495.8400 ;
        RECT 2352.1200 495.3600 2353.7200 495.8400 ;
        RECT 2257.5600 511.6800 2260.5600 512.1600 ;
        RECT 2257.5600 506.2400 2260.5600 506.7200 ;
        RECT 2257.5600 500.8000 2260.5600 501.2800 ;
        RECT 2257.5600 489.9200 2260.5600 490.4000 ;
        RECT 2257.5600 484.4800 2260.5600 484.9600 ;
        RECT 2257.5600 479.0400 2260.5600 479.5200 ;
        RECT 2257.5600 473.6000 2260.5600 474.0800 ;
        RECT 2257.5600 495.3600 2260.5600 495.8400 ;
        RECT 2352.1200 457.2800 2353.7200 457.7600 ;
        RECT 2352.1200 462.7200 2353.7200 463.2000 ;
        RECT 2352.1200 440.9600 2353.7200 441.4400 ;
        RECT 2352.1200 446.4000 2353.7200 446.8800 ;
        RECT 2352.1200 451.8400 2353.7200 452.3200 ;
        RECT 2307.1200 457.2800 2308.7200 457.7600 ;
        RECT 2307.1200 462.7200 2308.7200 463.2000 ;
        RECT 2307.1200 440.9600 2308.7200 441.4400 ;
        RECT 2307.1200 446.4000 2308.7200 446.8800 ;
        RECT 2307.1200 451.8400 2308.7200 452.3200 ;
        RECT 2352.1200 430.0800 2353.7200 430.5600 ;
        RECT 2352.1200 435.5200 2353.7200 436.0000 ;
        RECT 2352.1200 413.7600 2353.7200 414.2400 ;
        RECT 2352.1200 419.2000 2353.7200 419.6800 ;
        RECT 2352.1200 424.6400 2353.7200 425.1200 ;
        RECT 2307.1200 430.0800 2308.7200 430.5600 ;
        RECT 2307.1200 435.5200 2308.7200 436.0000 ;
        RECT 2307.1200 413.7600 2308.7200 414.2400 ;
        RECT 2307.1200 419.2000 2308.7200 419.6800 ;
        RECT 2307.1200 424.6400 2308.7200 425.1200 ;
        RECT 2257.5600 457.2800 2260.5600 457.7600 ;
        RECT 2257.5600 462.7200 2260.5600 463.2000 ;
        RECT 2257.5600 446.4000 2260.5600 446.8800 ;
        RECT 2257.5600 440.9600 2260.5600 441.4400 ;
        RECT 2257.5600 451.8400 2260.5600 452.3200 ;
        RECT 2257.5600 430.0800 2260.5600 430.5600 ;
        RECT 2257.5600 435.5200 2260.5600 436.0000 ;
        RECT 2257.5600 419.2000 2260.5600 419.6800 ;
        RECT 2257.5600 413.7600 2260.5600 414.2400 ;
        RECT 2257.5600 424.6400 2260.5600 425.1200 ;
        RECT 2257.5600 468.1600 2260.5600 468.6400 ;
        RECT 2307.1200 468.1600 2308.7200 468.6400 ;
        RECT 2352.1200 468.1600 2353.7200 468.6400 ;
        RECT 2453.6600 402.8800 2456.6600 403.3600 ;
        RECT 2453.6600 408.3200 2456.6600 408.8000 ;
        RECT 2442.1200 402.8800 2443.7200 403.3600 ;
        RECT 2442.1200 408.3200 2443.7200 408.8000 ;
        RECT 2453.6600 386.5600 2456.6600 387.0400 ;
        RECT 2453.6600 392.0000 2456.6600 392.4800 ;
        RECT 2453.6600 397.4400 2456.6600 397.9200 ;
        RECT 2442.1200 386.5600 2443.7200 387.0400 ;
        RECT 2442.1200 392.0000 2443.7200 392.4800 ;
        RECT 2442.1200 397.4400 2443.7200 397.9200 ;
        RECT 2453.6600 375.6800 2456.6600 376.1600 ;
        RECT 2453.6600 381.1200 2456.6600 381.6000 ;
        RECT 2442.1200 375.6800 2443.7200 376.1600 ;
        RECT 2442.1200 381.1200 2443.7200 381.6000 ;
        RECT 2453.6600 359.3600 2456.6600 359.8400 ;
        RECT 2453.6600 364.8000 2456.6600 365.2800 ;
        RECT 2453.6600 370.2400 2456.6600 370.7200 ;
        RECT 2442.1200 359.3600 2443.7200 359.8400 ;
        RECT 2442.1200 364.8000 2443.7200 365.2800 ;
        RECT 2442.1200 370.2400 2443.7200 370.7200 ;
        RECT 2397.1200 402.8800 2398.7200 403.3600 ;
        RECT 2397.1200 408.3200 2398.7200 408.8000 ;
        RECT 2397.1200 386.5600 2398.7200 387.0400 ;
        RECT 2397.1200 392.0000 2398.7200 392.4800 ;
        RECT 2397.1200 397.4400 2398.7200 397.9200 ;
        RECT 2397.1200 375.6800 2398.7200 376.1600 ;
        RECT 2397.1200 381.1200 2398.7200 381.6000 ;
        RECT 2397.1200 359.3600 2398.7200 359.8400 ;
        RECT 2397.1200 364.8000 2398.7200 365.2800 ;
        RECT 2397.1200 370.2400 2398.7200 370.7200 ;
        RECT 2453.6600 348.4800 2456.6600 348.9600 ;
        RECT 2453.6600 353.9200 2456.6600 354.4000 ;
        RECT 2442.1200 348.4800 2443.7200 348.9600 ;
        RECT 2442.1200 353.9200 2443.7200 354.4000 ;
        RECT 2453.6600 332.1600 2456.6600 332.6400 ;
        RECT 2453.6600 337.6000 2456.6600 338.0800 ;
        RECT 2453.6600 343.0400 2456.6600 343.5200 ;
        RECT 2442.1200 332.1600 2443.7200 332.6400 ;
        RECT 2442.1200 337.6000 2443.7200 338.0800 ;
        RECT 2442.1200 343.0400 2443.7200 343.5200 ;
        RECT 2453.6600 321.2800 2456.6600 321.7600 ;
        RECT 2453.6600 326.7200 2456.6600 327.2000 ;
        RECT 2442.1200 321.2800 2443.7200 321.7600 ;
        RECT 2442.1200 326.7200 2443.7200 327.2000 ;
        RECT 2453.6600 315.8400 2456.6600 316.3200 ;
        RECT 2442.1200 315.8400 2443.7200 316.3200 ;
        RECT 2397.1200 348.4800 2398.7200 348.9600 ;
        RECT 2397.1200 353.9200 2398.7200 354.4000 ;
        RECT 2397.1200 332.1600 2398.7200 332.6400 ;
        RECT 2397.1200 337.6000 2398.7200 338.0800 ;
        RECT 2397.1200 343.0400 2398.7200 343.5200 ;
        RECT 2397.1200 321.2800 2398.7200 321.7600 ;
        RECT 2397.1200 326.7200 2398.7200 327.2000 ;
        RECT 2397.1200 315.8400 2398.7200 316.3200 ;
        RECT 2352.1200 402.8800 2353.7200 403.3600 ;
        RECT 2352.1200 408.3200 2353.7200 408.8000 ;
        RECT 2352.1200 386.5600 2353.7200 387.0400 ;
        RECT 2352.1200 392.0000 2353.7200 392.4800 ;
        RECT 2352.1200 397.4400 2353.7200 397.9200 ;
        RECT 2307.1200 402.8800 2308.7200 403.3600 ;
        RECT 2307.1200 408.3200 2308.7200 408.8000 ;
        RECT 2307.1200 386.5600 2308.7200 387.0400 ;
        RECT 2307.1200 392.0000 2308.7200 392.4800 ;
        RECT 2307.1200 397.4400 2308.7200 397.9200 ;
        RECT 2352.1200 375.6800 2353.7200 376.1600 ;
        RECT 2352.1200 381.1200 2353.7200 381.6000 ;
        RECT 2352.1200 359.3600 2353.7200 359.8400 ;
        RECT 2352.1200 364.8000 2353.7200 365.2800 ;
        RECT 2352.1200 370.2400 2353.7200 370.7200 ;
        RECT 2307.1200 375.6800 2308.7200 376.1600 ;
        RECT 2307.1200 381.1200 2308.7200 381.6000 ;
        RECT 2307.1200 359.3600 2308.7200 359.8400 ;
        RECT 2307.1200 364.8000 2308.7200 365.2800 ;
        RECT 2307.1200 370.2400 2308.7200 370.7200 ;
        RECT 2257.5600 402.8800 2260.5600 403.3600 ;
        RECT 2257.5600 408.3200 2260.5600 408.8000 ;
        RECT 2257.5600 392.0000 2260.5600 392.4800 ;
        RECT 2257.5600 386.5600 2260.5600 387.0400 ;
        RECT 2257.5600 397.4400 2260.5600 397.9200 ;
        RECT 2257.5600 375.6800 2260.5600 376.1600 ;
        RECT 2257.5600 381.1200 2260.5600 381.6000 ;
        RECT 2257.5600 364.8000 2260.5600 365.2800 ;
        RECT 2257.5600 359.3600 2260.5600 359.8400 ;
        RECT 2257.5600 370.2400 2260.5600 370.7200 ;
        RECT 2352.1200 348.4800 2353.7200 348.9600 ;
        RECT 2352.1200 353.9200 2353.7200 354.4000 ;
        RECT 2352.1200 332.1600 2353.7200 332.6400 ;
        RECT 2352.1200 337.6000 2353.7200 338.0800 ;
        RECT 2352.1200 343.0400 2353.7200 343.5200 ;
        RECT 2307.1200 348.4800 2308.7200 348.9600 ;
        RECT 2307.1200 353.9200 2308.7200 354.4000 ;
        RECT 2307.1200 332.1600 2308.7200 332.6400 ;
        RECT 2307.1200 337.6000 2308.7200 338.0800 ;
        RECT 2307.1200 343.0400 2308.7200 343.5200 ;
        RECT 2352.1200 326.7200 2353.7200 327.2000 ;
        RECT 2352.1200 321.2800 2353.7200 321.7600 ;
        RECT 2352.1200 315.8400 2353.7200 316.3200 ;
        RECT 2307.1200 326.7200 2308.7200 327.2000 ;
        RECT 2307.1200 321.2800 2308.7200 321.7600 ;
        RECT 2307.1200 315.8400 2308.7200 316.3200 ;
        RECT 2257.5600 348.4800 2260.5600 348.9600 ;
        RECT 2257.5600 353.9200 2260.5600 354.4000 ;
        RECT 2257.5600 337.6000 2260.5600 338.0800 ;
        RECT 2257.5600 332.1600 2260.5600 332.6400 ;
        RECT 2257.5600 343.0400 2260.5600 343.5200 ;
        RECT 2257.5600 321.2800 2260.5600 321.7600 ;
        RECT 2257.5600 326.7200 2260.5600 327.2000 ;
        RECT 2257.5600 315.8400 2260.5600 316.3200 ;
        RECT 2257.5600 514.0300 2456.6600 517.0300 ;
        RECT 2257.5600 308.9300 2456.6600 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 79.2900 2443.7200 287.3900 ;
        RECT 2397.1200 79.2900 2398.7200 287.3900 ;
        RECT 2352.1200 79.2900 2353.7200 287.3900 ;
        RECT 2307.1200 79.2900 2308.7200 287.3900 ;
        RECT 2453.6600 79.2900 2456.6600 287.3900 ;
        RECT 2257.5600 79.2900 2260.5600 287.3900 ;
      LAYER met3 ;
        RECT 2453.6600 282.0400 2456.6600 282.5200 ;
        RECT 2442.1200 282.0400 2443.7200 282.5200 ;
        RECT 2453.6600 271.1600 2456.6600 271.6400 ;
        RECT 2453.6600 276.6000 2456.6600 277.0800 ;
        RECT 2442.1200 271.1600 2443.7200 271.6400 ;
        RECT 2442.1200 276.6000 2443.7200 277.0800 ;
        RECT 2453.6600 254.8400 2456.6600 255.3200 ;
        RECT 2453.6600 260.2800 2456.6600 260.7600 ;
        RECT 2442.1200 254.8400 2443.7200 255.3200 ;
        RECT 2442.1200 260.2800 2443.7200 260.7600 ;
        RECT 2453.6600 243.9600 2456.6600 244.4400 ;
        RECT 2453.6600 249.4000 2456.6600 249.8800 ;
        RECT 2442.1200 243.9600 2443.7200 244.4400 ;
        RECT 2442.1200 249.4000 2443.7200 249.8800 ;
        RECT 2453.6600 265.7200 2456.6600 266.2000 ;
        RECT 2442.1200 265.7200 2443.7200 266.2000 ;
        RECT 2397.1200 271.1600 2398.7200 271.6400 ;
        RECT 2397.1200 276.6000 2398.7200 277.0800 ;
        RECT 2397.1200 282.0400 2398.7200 282.5200 ;
        RECT 2397.1200 254.8400 2398.7200 255.3200 ;
        RECT 2397.1200 260.2800 2398.7200 260.7600 ;
        RECT 2397.1200 249.4000 2398.7200 249.8800 ;
        RECT 2397.1200 243.9600 2398.7200 244.4400 ;
        RECT 2397.1200 265.7200 2398.7200 266.2000 ;
        RECT 2453.6600 227.6400 2456.6600 228.1200 ;
        RECT 2453.6600 233.0800 2456.6600 233.5600 ;
        RECT 2442.1200 227.6400 2443.7200 228.1200 ;
        RECT 2442.1200 233.0800 2443.7200 233.5600 ;
        RECT 2453.6600 211.3200 2456.6600 211.8000 ;
        RECT 2453.6600 216.7600 2456.6600 217.2400 ;
        RECT 2453.6600 222.2000 2456.6600 222.6800 ;
        RECT 2442.1200 211.3200 2443.7200 211.8000 ;
        RECT 2442.1200 216.7600 2443.7200 217.2400 ;
        RECT 2442.1200 222.2000 2443.7200 222.6800 ;
        RECT 2453.6600 200.4400 2456.6600 200.9200 ;
        RECT 2453.6600 205.8800 2456.6600 206.3600 ;
        RECT 2442.1200 200.4400 2443.7200 200.9200 ;
        RECT 2442.1200 205.8800 2443.7200 206.3600 ;
        RECT 2453.6600 184.1200 2456.6600 184.6000 ;
        RECT 2453.6600 189.5600 2456.6600 190.0400 ;
        RECT 2453.6600 195.0000 2456.6600 195.4800 ;
        RECT 2442.1200 184.1200 2443.7200 184.6000 ;
        RECT 2442.1200 189.5600 2443.7200 190.0400 ;
        RECT 2442.1200 195.0000 2443.7200 195.4800 ;
        RECT 2397.1200 227.6400 2398.7200 228.1200 ;
        RECT 2397.1200 233.0800 2398.7200 233.5600 ;
        RECT 2397.1200 211.3200 2398.7200 211.8000 ;
        RECT 2397.1200 216.7600 2398.7200 217.2400 ;
        RECT 2397.1200 222.2000 2398.7200 222.6800 ;
        RECT 2397.1200 200.4400 2398.7200 200.9200 ;
        RECT 2397.1200 205.8800 2398.7200 206.3600 ;
        RECT 2397.1200 184.1200 2398.7200 184.6000 ;
        RECT 2397.1200 189.5600 2398.7200 190.0400 ;
        RECT 2397.1200 195.0000 2398.7200 195.4800 ;
        RECT 2453.6600 238.5200 2456.6600 239.0000 ;
        RECT 2397.1200 238.5200 2398.7200 239.0000 ;
        RECT 2442.1200 238.5200 2443.7200 239.0000 ;
        RECT 2352.1200 271.1600 2353.7200 271.6400 ;
        RECT 2352.1200 276.6000 2353.7200 277.0800 ;
        RECT 2352.1200 282.0400 2353.7200 282.5200 ;
        RECT 2307.1200 271.1600 2308.7200 271.6400 ;
        RECT 2307.1200 276.6000 2308.7200 277.0800 ;
        RECT 2307.1200 282.0400 2308.7200 282.5200 ;
        RECT 2352.1200 254.8400 2353.7200 255.3200 ;
        RECT 2352.1200 260.2800 2353.7200 260.7600 ;
        RECT 2352.1200 243.9600 2353.7200 244.4400 ;
        RECT 2352.1200 249.4000 2353.7200 249.8800 ;
        RECT 2307.1200 254.8400 2308.7200 255.3200 ;
        RECT 2307.1200 260.2800 2308.7200 260.7600 ;
        RECT 2307.1200 243.9600 2308.7200 244.4400 ;
        RECT 2307.1200 249.4000 2308.7200 249.8800 ;
        RECT 2307.1200 265.7200 2308.7200 266.2000 ;
        RECT 2352.1200 265.7200 2353.7200 266.2000 ;
        RECT 2257.5600 282.0400 2260.5600 282.5200 ;
        RECT 2257.5600 276.6000 2260.5600 277.0800 ;
        RECT 2257.5600 271.1600 2260.5600 271.6400 ;
        RECT 2257.5600 260.2800 2260.5600 260.7600 ;
        RECT 2257.5600 254.8400 2260.5600 255.3200 ;
        RECT 2257.5600 249.4000 2260.5600 249.8800 ;
        RECT 2257.5600 243.9600 2260.5600 244.4400 ;
        RECT 2257.5600 265.7200 2260.5600 266.2000 ;
        RECT 2352.1200 227.6400 2353.7200 228.1200 ;
        RECT 2352.1200 233.0800 2353.7200 233.5600 ;
        RECT 2352.1200 211.3200 2353.7200 211.8000 ;
        RECT 2352.1200 216.7600 2353.7200 217.2400 ;
        RECT 2352.1200 222.2000 2353.7200 222.6800 ;
        RECT 2307.1200 227.6400 2308.7200 228.1200 ;
        RECT 2307.1200 233.0800 2308.7200 233.5600 ;
        RECT 2307.1200 211.3200 2308.7200 211.8000 ;
        RECT 2307.1200 216.7600 2308.7200 217.2400 ;
        RECT 2307.1200 222.2000 2308.7200 222.6800 ;
        RECT 2352.1200 200.4400 2353.7200 200.9200 ;
        RECT 2352.1200 205.8800 2353.7200 206.3600 ;
        RECT 2352.1200 184.1200 2353.7200 184.6000 ;
        RECT 2352.1200 189.5600 2353.7200 190.0400 ;
        RECT 2352.1200 195.0000 2353.7200 195.4800 ;
        RECT 2307.1200 200.4400 2308.7200 200.9200 ;
        RECT 2307.1200 205.8800 2308.7200 206.3600 ;
        RECT 2307.1200 184.1200 2308.7200 184.6000 ;
        RECT 2307.1200 189.5600 2308.7200 190.0400 ;
        RECT 2307.1200 195.0000 2308.7200 195.4800 ;
        RECT 2257.5600 227.6400 2260.5600 228.1200 ;
        RECT 2257.5600 233.0800 2260.5600 233.5600 ;
        RECT 2257.5600 216.7600 2260.5600 217.2400 ;
        RECT 2257.5600 211.3200 2260.5600 211.8000 ;
        RECT 2257.5600 222.2000 2260.5600 222.6800 ;
        RECT 2257.5600 200.4400 2260.5600 200.9200 ;
        RECT 2257.5600 205.8800 2260.5600 206.3600 ;
        RECT 2257.5600 189.5600 2260.5600 190.0400 ;
        RECT 2257.5600 184.1200 2260.5600 184.6000 ;
        RECT 2257.5600 195.0000 2260.5600 195.4800 ;
        RECT 2257.5600 238.5200 2260.5600 239.0000 ;
        RECT 2307.1200 238.5200 2308.7200 239.0000 ;
        RECT 2352.1200 238.5200 2353.7200 239.0000 ;
        RECT 2453.6600 173.2400 2456.6600 173.7200 ;
        RECT 2453.6600 178.6800 2456.6600 179.1600 ;
        RECT 2442.1200 173.2400 2443.7200 173.7200 ;
        RECT 2442.1200 178.6800 2443.7200 179.1600 ;
        RECT 2453.6600 156.9200 2456.6600 157.4000 ;
        RECT 2453.6600 162.3600 2456.6600 162.8400 ;
        RECT 2453.6600 167.8000 2456.6600 168.2800 ;
        RECT 2442.1200 156.9200 2443.7200 157.4000 ;
        RECT 2442.1200 162.3600 2443.7200 162.8400 ;
        RECT 2442.1200 167.8000 2443.7200 168.2800 ;
        RECT 2453.6600 146.0400 2456.6600 146.5200 ;
        RECT 2453.6600 151.4800 2456.6600 151.9600 ;
        RECT 2442.1200 146.0400 2443.7200 146.5200 ;
        RECT 2442.1200 151.4800 2443.7200 151.9600 ;
        RECT 2453.6600 129.7200 2456.6600 130.2000 ;
        RECT 2453.6600 135.1600 2456.6600 135.6400 ;
        RECT 2453.6600 140.6000 2456.6600 141.0800 ;
        RECT 2442.1200 129.7200 2443.7200 130.2000 ;
        RECT 2442.1200 135.1600 2443.7200 135.6400 ;
        RECT 2442.1200 140.6000 2443.7200 141.0800 ;
        RECT 2397.1200 173.2400 2398.7200 173.7200 ;
        RECT 2397.1200 178.6800 2398.7200 179.1600 ;
        RECT 2397.1200 156.9200 2398.7200 157.4000 ;
        RECT 2397.1200 162.3600 2398.7200 162.8400 ;
        RECT 2397.1200 167.8000 2398.7200 168.2800 ;
        RECT 2397.1200 146.0400 2398.7200 146.5200 ;
        RECT 2397.1200 151.4800 2398.7200 151.9600 ;
        RECT 2397.1200 129.7200 2398.7200 130.2000 ;
        RECT 2397.1200 135.1600 2398.7200 135.6400 ;
        RECT 2397.1200 140.6000 2398.7200 141.0800 ;
        RECT 2453.6600 118.8400 2456.6600 119.3200 ;
        RECT 2453.6600 124.2800 2456.6600 124.7600 ;
        RECT 2442.1200 118.8400 2443.7200 119.3200 ;
        RECT 2442.1200 124.2800 2443.7200 124.7600 ;
        RECT 2453.6600 102.5200 2456.6600 103.0000 ;
        RECT 2453.6600 107.9600 2456.6600 108.4400 ;
        RECT 2453.6600 113.4000 2456.6600 113.8800 ;
        RECT 2442.1200 102.5200 2443.7200 103.0000 ;
        RECT 2442.1200 107.9600 2443.7200 108.4400 ;
        RECT 2442.1200 113.4000 2443.7200 113.8800 ;
        RECT 2453.6600 91.6400 2456.6600 92.1200 ;
        RECT 2453.6600 97.0800 2456.6600 97.5600 ;
        RECT 2442.1200 91.6400 2443.7200 92.1200 ;
        RECT 2442.1200 97.0800 2443.7200 97.5600 ;
        RECT 2453.6600 86.2000 2456.6600 86.6800 ;
        RECT 2442.1200 86.2000 2443.7200 86.6800 ;
        RECT 2397.1200 118.8400 2398.7200 119.3200 ;
        RECT 2397.1200 124.2800 2398.7200 124.7600 ;
        RECT 2397.1200 102.5200 2398.7200 103.0000 ;
        RECT 2397.1200 107.9600 2398.7200 108.4400 ;
        RECT 2397.1200 113.4000 2398.7200 113.8800 ;
        RECT 2397.1200 91.6400 2398.7200 92.1200 ;
        RECT 2397.1200 97.0800 2398.7200 97.5600 ;
        RECT 2397.1200 86.2000 2398.7200 86.6800 ;
        RECT 2352.1200 173.2400 2353.7200 173.7200 ;
        RECT 2352.1200 178.6800 2353.7200 179.1600 ;
        RECT 2352.1200 156.9200 2353.7200 157.4000 ;
        RECT 2352.1200 162.3600 2353.7200 162.8400 ;
        RECT 2352.1200 167.8000 2353.7200 168.2800 ;
        RECT 2307.1200 173.2400 2308.7200 173.7200 ;
        RECT 2307.1200 178.6800 2308.7200 179.1600 ;
        RECT 2307.1200 156.9200 2308.7200 157.4000 ;
        RECT 2307.1200 162.3600 2308.7200 162.8400 ;
        RECT 2307.1200 167.8000 2308.7200 168.2800 ;
        RECT 2352.1200 146.0400 2353.7200 146.5200 ;
        RECT 2352.1200 151.4800 2353.7200 151.9600 ;
        RECT 2352.1200 129.7200 2353.7200 130.2000 ;
        RECT 2352.1200 135.1600 2353.7200 135.6400 ;
        RECT 2352.1200 140.6000 2353.7200 141.0800 ;
        RECT 2307.1200 146.0400 2308.7200 146.5200 ;
        RECT 2307.1200 151.4800 2308.7200 151.9600 ;
        RECT 2307.1200 129.7200 2308.7200 130.2000 ;
        RECT 2307.1200 135.1600 2308.7200 135.6400 ;
        RECT 2307.1200 140.6000 2308.7200 141.0800 ;
        RECT 2257.5600 173.2400 2260.5600 173.7200 ;
        RECT 2257.5600 178.6800 2260.5600 179.1600 ;
        RECT 2257.5600 162.3600 2260.5600 162.8400 ;
        RECT 2257.5600 156.9200 2260.5600 157.4000 ;
        RECT 2257.5600 167.8000 2260.5600 168.2800 ;
        RECT 2257.5600 146.0400 2260.5600 146.5200 ;
        RECT 2257.5600 151.4800 2260.5600 151.9600 ;
        RECT 2257.5600 135.1600 2260.5600 135.6400 ;
        RECT 2257.5600 129.7200 2260.5600 130.2000 ;
        RECT 2257.5600 140.6000 2260.5600 141.0800 ;
        RECT 2352.1200 118.8400 2353.7200 119.3200 ;
        RECT 2352.1200 124.2800 2353.7200 124.7600 ;
        RECT 2352.1200 102.5200 2353.7200 103.0000 ;
        RECT 2352.1200 107.9600 2353.7200 108.4400 ;
        RECT 2352.1200 113.4000 2353.7200 113.8800 ;
        RECT 2307.1200 118.8400 2308.7200 119.3200 ;
        RECT 2307.1200 124.2800 2308.7200 124.7600 ;
        RECT 2307.1200 102.5200 2308.7200 103.0000 ;
        RECT 2307.1200 107.9600 2308.7200 108.4400 ;
        RECT 2307.1200 113.4000 2308.7200 113.8800 ;
        RECT 2352.1200 97.0800 2353.7200 97.5600 ;
        RECT 2352.1200 91.6400 2353.7200 92.1200 ;
        RECT 2352.1200 86.2000 2353.7200 86.6800 ;
        RECT 2307.1200 97.0800 2308.7200 97.5600 ;
        RECT 2307.1200 91.6400 2308.7200 92.1200 ;
        RECT 2307.1200 86.2000 2308.7200 86.6800 ;
        RECT 2257.5600 118.8400 2260.5600 119.3200 ;
        RECT 2257.5600 124.2800 2260.5600 124.7600 ;
        RECT 2257.5600 107.9600 2260.5600 108.4400 ;
        RECT 2257.5600 102.5200 2260.5600 103.0000 ;
        RECT 2257.5600 113.4000 2260.5600 113.8800 ;
        RECT 2257.5600 91.6400 2260.5600 92.1200 ;
        RECT 2257.5600 97.0800 2260.5600 97.5600 ;
        RECT 2257.5600 86.2000 2260.5600 86.6800 ;
        RECT 2257.5600 284.3900 2456.6600 287.3900 ;
        RECT 2257.5600 79.2900 2456.6600 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 2257.5600 37.6700 2259.5600 58.6000 ;
        RECT 2454.6600 37.6700 2456.6600 58.6000 ;
      LAYER met3 ;
        RECT 2454.6600 54.1000 2456.6600 54.5800 ;
        RECT 2257.5600 54.1000 2259.5600 54.5800 ;
        RECT 2454.6600 43.2200 2456.6600 43.7000 ;
        RECT 2257.5600 43.2200 2259.5600 43.7000 ;
        RECT 2454.6600 48.6600 2456.6600 49.1400 ;
        RECT 2257.5600 48.6600 2259.5600 49.1400 ;
        RECT 2257.5600 56.6000 2456.6600 58.6000 ;
        RECT 2257.5600 37.6700 2456.6600 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 2605.3300 2443.7200 2813.4300 ;
        RECT 2397.1200 2605.3300 2398.7200 2813.4300 ;
        RECT 2352.1200 2605.3300 2353.7200 2813.4300 ;
        RECT 2307.1200 2605.3300 2308.7200 2813.4300 ;
        RECT 2453.6600 2605.3300 2456.6600 2813.4300 ;
        RECT 2257.5600 2605.3300 2260.5600 2813.4300 ;
      LAYER met3 ;
        RECT 2453.6600 2808.0800 2456.6600 2808.5600 ;
        RECT 2442.1200 2808.0800 2443.7200 2808.5600 ;
        RECT 2453.6600 2797.2000 2456.6600 2797.6800 ;
        RECT 2453.6600 2802.6400 2456.6600 2803.1200 ;
        RECT 2442.1200 2797.2000 2443.7200 2797.6800 ;
        RECT 2442.1200 2802.6400 2443.7200 2803.1200 ;
        RECT 2453.6600 2780.8800 2456.6600 2781.3600 ;
        RECT 2453.6600 2786.3200 2456.6600 2786.8000 ;
        RECT 2442.1200 2780.8800 2443.7200 2781.3600 ;
        RECT 2442.1200 2786.3200 2443.7200 2786.8000 ;
        RECT 2453.6600 2770.0000 2456.6600 2770.4800 ;
        RECT 2453.6600 2775.4400 2456.6600 2775.9200 ;
        RECT 2442.1200 2770.0000 2443.7200 2770.4800 ;
        RECT 2442.1200 2775.4400 2443.7200 2775.9200 ;
        RECT 2453.6600 2791.7600 2456.6600 2792.2400 ;
        RECT 2442.1200 2791.7600 2443.7200 2792.2400 ;
        RECT 2397.1200 2797.2000 2398.7200 2797.6800 ;
        RECT 2397.1200 2802.6400 2398.7200 2803.1200 ;
        RECT 2397.1200 2808.0800 2398.7200 2808.5600 ;
        RECT 2397.1200 2780.8800 2398.7200 2781.3600 ;
        RECT 2397.1200 2786.3200 2398.7200 2786.8000 ;
        RECT 2397.1200 2775.4400 2398.7200 2775.9200 ;
        RECT 2397.1200 2770.0000 2398.7200 2770.4800 ;
        RECT 2397.1200 2791.7600 2398.7200 2792.2400 ;
        RECT 2453.6600 2753.6800 2456.6600 2754.1600 ;
        RECT 2453.6600 2759.1200 2456.6600 2759.6000 ;
        RECT 2442.1200 2753.6800 2443.7200 2754.1600 ;
        RECT 2442.1200 2759.1200 2443.7200 2759.6000 ;
        RECT 2453.6600 2737.3600 2456.6600 2737.8400 ;
        RECT 2453.6600 2742.8000 2456.6600 2743.2800 ;
        RECT 2453.6600 2748.2400 2456.6600 2748.7200 ;
        RECT 2442.1200 2737.3600 2443.7200 2737.8400 ;
        RECT 2442.1200 2742.8000 2443.7200 2743.2800 ;
        RECT 2442.1200 2748.2400 2443.7200 2748.7200 ;
        RECT 2453.6600 2726.4800 2456.6600 2726.9600 ;
        RECT 2453.6600 2731.9200 2456.6600 2732.4000 ;
        RECT 2442.1200 2726.4800 2443.7200 2726.9600 ;
        RECT 2442.1200 2731.9200 2443.7200 2732.4000 ;
        RECT 2453.6600 2710.1600 2456.6600 2710.6400 ;
        RECT 2453.6600 2715.6000 2456.6600 2716.0800 ;
        RECT 2453.6600 2721.0400 2456.6600 2721.5200 ;
        RECT 2442.1200 2710.1600 2443.7200 2710.6400 ;
        RECT 2442.1200 2715.6000 2443.7200 2716.0800 ;
        RECT 2442.1200 2721.0400 2443.7200 2721.5200 ;
        RECT 2397.1200 2753.6800 2398.7200 2754.1600 ;
        RECT 2397.1200 2759.1200 2398.7200 2759.6000 ;
        RECT 2397.1200 2737.3600 2398.7200 2737.8400 ;
        RECT 2397.1200 2742.8000 2398.7200 2743.2800 ;
        RECT 2397.1200 2748.2400 2398.7200 2748.7200 ;
        RECT 2397.1200 2726.4800 2398.7200 2726.9600 ;
        RECT 2397.1200 2731.9200 2398.7200 2732.4000 ;
        RECT 2397.1200 2710.1600 2398.7200 2710.6400 ;
        RECT 2397.1200 2715.6000 2398.7200 2716.0800 ;
        RECT 2397.1200 2721.0400 2398.7200 2721.5200 ;
        RECT 2453.6600 2764.5600 2456.6600 2765.0400 ;
        RECT 2397.1200 2764.5600 2398.7200 2765.0400 ;
        RECT 2442.1200 2764.5600 2443.7200 2765.0400 ;
        RECT 2352.1200 2797.2000 2353.7200 2797.6800 ;
        RECT 2352.1200 2802.6400 2353.7200 2803.1200 ;
        RECT 2352.1200 2808.0800 2353.7200 2808.5600 ;
        RECT 2307.1200 2797.2000 2308.7200 2797.6800 ;
        RECT 2307.1200 2802.6400 2308.7200 2803.1200 ;
        RECT 2307.1200 2808.0800 2308.7200 2808.5600 ;
        RECT 2352.1200 2780.8800 2353.7200 2781.3600 ;
        RECT 2352.1200 2786.3200 2353.7200 2786.8000 ;
        RECT 2352.1200 2770.0000 2353.7200 2770.4800 ;
        RECT 2352.1200 2775.4400 2353.7200 2775.9200 ;
        RECT 2307.1200 2780.8800 2308.7200 2781.3600 ;
        RECT 2307.1200 2786.3200 2308.7200 2786.8000 ;
        RECT 2307.1200 2770.0000 2308.7200 2770.4800 ;
        RECT 2307.1200 2775.4400 2308.7200 2775.9200 ;
        RECT 2307.1200 2791.7600 2308.7200 2792.2400 ;
        RECT 2352.1200 2791.7600 2353.7200 2792.2400 ;
        RECT 2257.5600 2808.0800 2260.5600 2808.5600 ;
        RECT 2257.5600 2802.6400 2260.5600 2803.1200 ;
        RECT 2257.5600 2797.2000 2260.5600 2797.6800 ;
        RECT 2257.5600 2786.3200 2260.5600 2786.8000 ;
        RECT 2257.5600 2780.8800 2260.5600 2781.3600 ;
        RECT 2257.5600 2775.4400 2260.5600 2775.9200 ;
        RECT 2257.5600 2770.0000 2260.5600 2770.4800 ;
        RECT 2257.5600 2791.7600 2260.5600 2792.2400 ;
        RECT 2352.1200 2753.6800 2353.7200 2754.1600 ;
        RECT 2352.1200 2759.1200 2353.7200 2759.6000 ;
        RECT 2352.1200 2737.3600 2353.7200 2737.8400 ;
        RECT 2352.1200 2742.8000 2353.7200 2743.2800 ;
        RECT 2352.1200 2748.2400 2353.7200 2748.7200 ;
        RECT 2307.1200 2753.6800 2308.7200 2754.1600 ;
        RECT 2307.1200 2759.1200 2308.7200 2759.6000 ;
        RECT 2307.1200 2737.3600 2308.7200 2737.8400 ;
        RECT 2307.1200 2742.8000 2308.7200 2743.2800 ;
        RECT 2307.1200 2748.2400 2308.7200 2748.7200 ;
        RECT 2352.1200 2726.4800 2353.7200 2726.9600 ;
        RECT 2352.1200 2731.9200 2353.7200 2732.4000 ;
        RECT 2352.1200 2710.1600 2353.7200 2710.6400 ;
        RECT 2352.1200 2715.6000 2353.7200 2716.0800 ;
        RECT 2352.1200 2721.0400 2353.7200 2721.5200 ;
        RECT 2307.1200 2726.4800 2308.7200 2726.9600 ;
        RECT 2307.1200 2731.9200 2308.7200 2732.4000 ;
        RECT 2307.1200 2710.1600 2308.7200 2710.6400 ;
        RECT 2307.1200 2715.6000 2308.7200 2716.0800 ;
        RECT 2307.1200 2721.0400 2308.7200 2721.5200 ;
        RECT 2257.5600 2753.6800 2260.5600 2754.1600 ;
        RECT 2257.5600 2759.1200 2260.5600 2759.6000 ;
        RECT 2257.5600 2742.8000 2260.5600 2743.2800 ;
        RECT 2257.5600 2737.3600 2260.5600 2737.8400 ;
        RECT 2257.5600 2748.2400 2260.5600 2748.7200 ;
        RECT 2257.5600 2726.4800 2260.5600 2726.9600 ;
        RECT 2257.5600 2731.9200 2260.5600 2732.4000 ;
        RECT 2257.5600 2715.6000 2260.5600 2716.0800 ;
        RECT 2257.5600 2710.1600 2260.5600 2710.6400 ;
        RECT 2257.5600 2721.0400 2260.5600 2721.5200 ;
        RECT 2257.5600 2764.5600 2260.5600 2765.0400 ;
        RECT 2307.1200 2764.5600 2308.7200 2765.0400 ;
        RECT 2352.1200 2764.5600 2353.7200 2765.0400 ;
        RECT 2453.6600 2699.2800 2456.6600 2699.7600 ;
        RECT 2453.6600 2704.7200 2456.6600 2705.2000 ;
        RECT 2442.1200 2699.2800 2443.7200 2699.7600 ;
        RECT 2442.1200 2704.7200 2443.7200 2705.2000 ;
        RECT 2453.6600 2682.9600 2456.6600 2683.4400 ;
        RECT 2453.6600 2688.4000 2456.6600 2688.8800 ;
        RECT 2453.6600 2693.8400 2456.6600 2694.3200 ;
        RECT 2442.1200 2682.9600 2443.7200 2683.4400 ;
        RECT 2442.1200 2688.4000 2443.7200 2688.8800 ;
        RECT 2442.1200 2693.8400 2443.7200 2694.3200 ;
        RECT 2453.6600 2672.0800 2456.6600 2672.5600 ;
        RECT 2453.6600 2677.5200 2456.6600 2678.0000 ;
        RECT 2442.1200 2672.0800 2443.7200 2672.5600 ;
        RECT 2442.1200 2677.5200 2443.7200 2678.0000 ;
        RECT 2453.6600 2655.7600 2456.6600 2656.2400 ;
        RECT 2453.6600 2661.2000 2456.6600 2661.6800 ;
        RECT 2453.6600 2666.6400 2456.6600 2667.1200 ;
        RECT 2442.1200 2655.7600 2443.7200 2656.2400 ;
        RECT 2442.1200 2661.2000 2443.7200 2661.6800 ;
        RECT 2442.1200 2666.6400 2443.7200 2667.1200 ;
        RECT 2397.1200 2699.2800 2398.7200 2699.7600 ;
        RECT 2397.1200 2704.7200 2398.7200 2705.2000 ;
        RECT 2397.1200 2682.9600 2398.7200 2683.4400 ;
        RECT 2397.1200 2688.4000 2398.7200 2688.8800 ;
        RECT 2397.1200 2693.8400 2398.7200 2694.3200 ;
        RECT 2397.1200 2672.0800 2398.7200 2672.5600 ;
        RECT 2397.1200 2677.5200 2398.7200 2678.0000 ;
        RECT 2397.1200 2655.7600 2398.7200 2656.2400 ;
        RECT 2397.1200 2661.2000 2398.7200 2661.6800 ;
        RECT 2397.1200 2666.6400 2398.7200 2667.1200 ;
        RECT 2453.6600 2644.8800 2456.6600 2645.3600 ;
        RECT 2453.6600 2650.3200 2456.6600 2650.8000 ;
        RECT 2442.1200 2644.8800 2443.7200 2645.3600 ;
        RECT 2442.1200 2650.3200 2443.7200 2650.8000 ;
        RECT 2453.6600 2628.5600 2456.6600 2629.0400 ;
        RECT 2453.6600 2634.0000 2456.6600 2634.4800 ;
        RECT 2453.6600 2639.4400 2456.6600 2639.9200 ;
        RECT 2442.1200 2628.5600 2443.7200 2629.0400 ;
        RECT 2442.1200 2634.0000 2443.7200 2634.4800 ;
        RECT 2442.1200 2639.4400 2443.7200 2639.9200 ;
        RECT 2453.6600 2617.6800 2456.6600 2618.1600 ;
        RECT 2453.6600 2623.1200 2456.6600 2623.6000 ;
        RECT 2442.1200 2617.6800 2443.7200 2618.1600 ;
        RECT 2442.1200 2623.1200 2443.7200 2623.6000 ;
        RECT 2453.6600 2612.2400 2456.6600 2612.7200 ;
        RECT 2442.1200 2612.2400 2443.7200 2612.7200 ;
        RECT 2397.1200 2644.8800 2398.7200 2645.3600 ;
        RECT 2397.1200 2650.3200 2398.7200 2650.8000 ;
        RECT 2397.1200 2628.5600 2398.7200 2629.0400 ;
        RECT 2397.1200 2634.0000 2398.7200 2634.4800 ;
        RECT 2397.1200 2639.4400 2398.7200 2639.9200 ;
        RECT 2397.1200 2617.6800 2398.7200 2618.1600 ;
        RECT 2397.1200 2623.1200 2398.7200 2623.6000 ;
        RECT 2397.1200 2612.2400 2398.7200 2612.7200 ;
        RECT 2352.1200 2699.2800 2353.7200 2699.7600 ;
        RECT 2352.1200 2704.7200 2353.7200 2705.2000 ;
        RECT 2352.1200 2682.9600 2353.7200 2683.4400 ;
        RECT 2352.1200 2688.4000 2353.7200 2688.8800 ;
        RECT 2352.1200 2693.8400 2353.7200 2694.3200 ;
        RECT 2307.1200 2699.2800 2308.7200 2699.7600 ;
        RECT 2307.1200 2704.7200 2308.7200 2705.2000 ;
        RECT 2307.1200 2682.9600 2308.7200 2683.4400 ;
        RECT 2307.1200 2688.4000 2308.7200 2688.8800 ;
        RECT 2307.1200 2693.8400 2308.7200 2694.3200 ;
        RECT 2352.1200 2672.0800 2353.7200 2672.5600 ;
        RECT 2352.1200 2677.5200 2353.7200 2678.0000 ;
        RECT 2352.1200 2655.7600 2353.7200 2656.2400 ;
        RECT 2352.1200 2661.2000 2353.7200 2661.6800 ;
        RECT 2352.1200 2666.6400 2353.7200 2667.1200 ;
        RECT 2307.1200 2672.0800 2308.7200 2672.5600 ;
        RECT 2307.1200 2677.5200 2308.7200 2678.0000 ;
        RECT 2307.1200 2655.7600 2308.7200 2656.2400 ;
        RECT 2307.1200 2661.2000 2308.7200 2661.6800 ;
        RECT 2307.1200 2666.6400 2308.7200 2667.1200 ;
        RECT 2257.5600 2699.2800 2260.5600 2699.7600 ;
        RECT 2257.5600 2704.7200 2260.5600 2705.2000 ;
        RECT 2257.5600 2688.4000 2260.5600 2688.8800 ;
        RECT 2257.5600 2682.9600 2260.5600 2683.4400 ;
        RECT 2257.5600 2693.8400 2260.5600 2694.3200 ;
        RECT 2257.5600 2672.0800 2260.5600 2672.5600 ;
        RECT 2257.5600 2677.5200 2260.5600 2678.0000 ;
        RECT 2257.5600 2661.2000 2260.5600 2661.6800 ;
        RECT 2257.5600 2655.7600 2260.5600 2656.2400 ;
        RECT 2257.5600 2666.6400 2260.5600 2667.1200 ;
        RECT 2352.1200 2644.8800 2353.7200 2645.3600 ;
        RECT 2352.1200 2650.3200 2353.7200 2650.8000 ;
        RECT 2352.1200 2628.5600 2353.7200 2629.0400 ;
        RECT 2352.1200 2634.0000 2353.7200 2634.4800 ;
        RECT 2352.1200 2639.4400 2353.7200 2639.9200 ;
        RECT 2307.1200 2644.8800 2308.7200 2645.3600 ;
        RECT 2307.1200 2650.3200 2308.7200 2650.8000 ;
        RECT 2307.1200 2628.5600 2308.7200 2629.0400 ;
        RECT 2307.1200 2634.0000 2308.7200 2634.4800 ;
        RECT 2307.1200 2639.4400 2308.7200 2639.9200 ;
        RECT 2352.1200 2623.1200 2353.7200 2623.6000 ;
        RECT 2352.1200 2617.6800 2353.7200 2618.1600 ;
        RECT 2352.1200 2612.2400 2353.7200 2612.7200 ;
        RECT 2307.1200 2623.1200 2308.7200 2623.6000 ;
        RECT 2307.1200 2617.6800 2308.7200 2618.1600 ;
        RECT 2307.1200 2612.2400 2308.7200 2612.7200 ;
        RECT 2257.5600 2644.8800 2260.5600 2645.3600 ;
        RECT 2257.5600 2650.3200 2260.5600 2650.8000 ;
        RECT 2257.5600 2634.0000 2260.5600 2634.4800 ;
        RECT 2257.5600 2628.5600 2260.5600 2629.0400 ;
        RECT 2257.5600 2639.4400 2260.5600 2639.9200 ;
        RECT 2257.5600 2617.6800 2260.5600 2618.1600 ;
        RECT 2257.5600 2623.1200 2260.5600 2623.6000 ;
        RECT 2257.5600 2612.2400 2260.5600 2612.7200 ;
        RECT 2257.5600 2810.4300 2456.6600 2813.4300 ;
        RECT 2257.5600 2605.3300 2456.6600 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 2375.6900 2443.7200 2583.7900 ;
        RECT 2397.1200 2375.6900 2398.7200 2583.7900 ;
        RECT 2352.1200 2375.6900 2353.7200 2583.7900 ;
        RECT 2307.1200 2375.6900 2308.7200 2583.7900 ;
        RECT 2453.6600 2375.6900 2456.6600 2583.7900 ;
        RECT 2257.5600 2375.6900 2260.5600 2583.7900 ;
      LAYER met3 ;
        RECT 2453.6600 2578.4400 2456.6600 2578.9200 ;
        RECT 2442.1200 2578.4400 2443.7200 2578.9200 ;
        RECT 2453.6600 2567.5600 2456.6600 2568.0400 ;
        RECT 2453.6600 2573.0000 2456.6600 2573.4800 ;
        RECT 2442.1200 2567.5600 2443.7200 2568.0400 ;
        RECT 2442.1200 2573.0000 2443.7200 2573.4800 ;
        RECT 2453.6600 2551.2400 2456.6600 2551.7200 ;
        RECT 2453.6600 2556.6800 2456.6600 2557.1600 ;
        RECT 2442.1200 2551.2400 2443.7200 2551.7200 ;
        RECT 2442.1200 2556.6800 2443.7200 2557.1600 ;
        RECT 2453.6600 2540.3600 2456.6600 2540.8400 ;
        RECT 2453.6600 2545.8000 2456.6600 2546.2800 ;
        RECT 2442.1200 2540.3600 2443.7200 2540.8400 ;
        RECT 2442.1200 2545.8000 2443.7200 2546.2800 ;
        RECT 2453.6600 2562.1200 2456.6600 2562.6000 ;
        RECT 2442.1200 2562.1200 2443.7200 2562.6000 ;
        RECT 2397.1200 2567.5600 2398.7200 2568.0400 ;
        RECT 2397.1200 2573.0000 2398.7200 2573.4800 ;
        RECT 2397.1200 2578.4400 2398.7200 2578.9200 ;
        RECT 2397.1200 2551.2400 2398.7200 2551.7200 ;
        RECT 2397.1200 2556.6800 2398.7200 2557.1600 ;
        RECT 2397.1200 2545.8000 2398.7200 2546.2800 ;
        RECT 2397.1200 2540.3600 2398.7200 2540.8400 ;
        RECT 2397.1200 2562.1200 2398.7200 2562.6000 ;
        RECT 2453.6600 2524.0400 2456.6600 2524.5200 ;
        RECT 2453.6600 2529.4800 2456.6600 2529.9600 ;
        RECT 2442.1200 2524.0400 2443.7200 2524.5200 ;
        RECT 2442.1200 2529.4800 2443.7200 2529.9600 ;
        RECT 2453.6600 2507.7200 2456.6600 2508.2000 ;
        RECT 2453.6600 2513.1600 2456.6600 2513.6400 ;
        RECT 2453.6600 2518.6000 2456.6600 2519.0800 ;
        RECT 2442.1200 2507.7200 2443.7200 2508.2000 ;
        RECT 2442.1200 2513.1600 2443.7200 2513.6400 ;
        RECT 2442.1200 2518.6000 2443.7200 2519.0800 ;
        RECT 2453.6600 2496.8400 2456.6600 2497.3200 ;
        RECT 2453.6600 2502.2800 2456.6600 2502.7600 ;
        RECT 2442.1200 2496.8400 2443.7200 2497.3200 ;
        RECT 2442.1200 2502.2800 2443.7200 2502.7600 ;
        RECT 2453.6600 2480.5200 2456.6600 2481.0000 ;
        RECT 2453.6600 2485.9600 2456.6600 2486.4400 ;
        RECT 2453.6600 2491.4000 2456.6600 2491.8800 ;
        RECT 2442.1200 2480.5200 2443.7200 2481.0000 ;
        RECT 2442.1200 2485.9600 2443.7200 2486.4400 ;
        RECT 2442.1200 2491.4000 2443.7200 2491.8800 ;
        RECT 2397.1200 2524.0400 2398.7200 2524.5200 ;
        RECT 2397.1200 2529.4800 2398.7200 2529.9600 ;
        RECT 2397.1200 2507.7200 2398.7200 2508.2000 ;
        RECT 2397.1200 2513.1600 2398.7200 2513.6400 ;
        RECT 2397.1200 2518.6000 2398.7200 2519.0800 ;
        RECT 2397.1200 2496.8400 2398.7200 2497.3200 ;
        RECT 2397.1200 2502.2800 2398.7200 2502.7600 ;
        RECT 2397.1200 2480.5200 2398.7200 2481.0000 ;
        RECT 2397.1200 2485.9600 2398.7200 2486.4400 ;
        RECT 2397.1200 2491.4000 2398.7200 2491.8800 ;
        RECT 2453.6600 2534.9200 2456.6600 2535.4000 ;
        RECT 2397.1200 2534.9200 2398.7200 2535.4000 ;
        RECT 2442.1200 2534.9200 2443.7200 2535.4000 ;
        RECT 2352.1200 2567.5600 2353.7200 2568.0400 ;
        RECT 2352.1200 2573.0000 2353.7200 2573.4800 ;
        RECT 2352.1200 2578.4400 2353.7200 2578.9200 ;
        RECT 2307.1200 2567.5600 2308.7200 2568.0400 ;
        RECT 2307.1200 2573.0000 2308.7200 2573.4800 ;
        RECT 2307.1200 2578.4400 2308.7200 2578.9200 ;
        RECT 2352.1200 2551.2400 2353.7200 2551.7200 ;
        RECT 2352.1200 2556.6800 2353.7200 2557.1600 ;
        RECT 2352.1200 2540.3600 2353.7200 2540.8400 ;
        RECT 2352.1200 2545.8000 2353.7200 2546.2800 ;
        RECT 2307.1200 2551.2400 2308.7200 2551.7200 ;
        RECT 2307.1200 2556.6800 2308.7200 2557.1600 ;
        RECT 2307.1200 2540.3600 2308.7200 2540.8400 ;
        RECT 2307.1200 2545.8000 2308.7200 2546.2800 ;
        RECT 2307.1200 2562.1200 2308.7200 2562.6000 ;
        RECT 2352.1200 2562.1200 2353.7200 2562.6000 ;
        RECT 2257.5600 2578.4400 2260.5600 2578.9200 ;
        RECT 2257.5600 2573.0000 2260.5600 2573.4800 ;
        RECT 2257.5600 2567.5600 2260.5600 2568.0400 ;
        RECT 2257.5600 2556.6800 2260.5600 2557.1600 ;
        RECT 2257.5600 2551.2400 2260.5600 2551.7200 ;
        RECT 2257.5600 2545.8000 2260.5600 2546.2800 ;
        RECT 2257.5600 2540.3600 2260.5600 2540.8400 ;
        RECT 2257.5600 2562.1200 2260.5600 2562.6000 ;
        RECT 2352.1200 2524.0400 2353.7200 2524.5200 ;
        RECT 2352.1200 2529.4800 2353.7200 2529.9600 ;
        RECT 2352.1200 2507.7200 2353.7200 2508.2000 ;
        RECT 2352.1200 2513.1600 2353.7200 2513.6400 ;
        RECT 2352.1200 2518.6000 2353.7200 2519.0800 ;
        RECT 2307.1200 2524.0400 2308.7200 2524.5200 ;
        RECT 2307.1200 2529.4800 2308.7200 2529.9600 ;
        RECT 2307.1200 2507.7200 2308.7200 2508.2000 ;
        RECT 2307.1200 2513.1600 2308.7200 2513.6400 ;
        RECT 2307.1200 2518.6000 2308.7200 2519.0800 ;
        RECT 2352.1200 2496.8400 2353.7200 2497.3200 ;
        RECT 2352.1200 2502.2800 2353.7200 2502.7600 ;
        RECT 2352.1200 2480.5200 2353.7200 2481.0000 ;
        RECT 2352.1200 2485.9600 2353.7200 2486.4400 ;
        RECT 2352.1200 2491.4000 2353.7200 2491.8800 ;
        RECT 2307.1200 2496.8400 2308.7200 2497.3200 ;
        RECT 2307.1200 2502.2800 2308.7200 2502.7600 ;
        RECT 2307.1200 2480.5200 2308.7200 2481.0000 ;
        RECT 2307.1200 2485.9600 2308.7200 2486.4400 ;
        RECT 2307.1200 2491.4000 2308.7200 2491.8800 ;
        RECT 2257.5600 2524.0400 2260.5600 2524.5200 ;
        RECT 2257.5600 2529.4800 2260.5600 2529.9600 ;
        RECT 2257.5600 2513.1600 2260.5600 2513.6400 ;
        RECT 2257.5600 2507.7200 2260.5600 2508.2000 ;
        RECT 2257.5600 2518.6000 2260.5600 2519.0800 ;
        RECT 2257.5600 2496.8400 2260.5600 2497.3200 ;
        RECT 2257.5600 2502.2800 2260.5600 2502.7600 ;
        RECT 2257.5600 2485.9600 2260.5600 2486.4400 ;
        RECT 2257.5600 2480.5200 2260.5600 2481.0000 ;
        RECT 2257.5600 2491.4000 2260.5600 2491.8800 ;
        RECT 2257.5600 2534.9200 2260.5600 2535.4000 ;
        RECT 2307.1200 2534.9200 2308.7200 2535.4000 ;
        RECT 2352.1200 2534.9200 2353.7200 2535.4000 ;
        RECT 2453.6600 2469.6400 2456.6600 2470.1200 ;
        RECT 2453.6600 2475.0800 2456.6600 2475.5600 ;
        RECT 2442.1200 2469.6400 2443.7200 2470.1200 ;
        RECT 2442.1200 2475.0800 2443.7200 2475.5600 ;
        RECT 2453.6600 2453.3200 2456.6600 2453.8000 ;
        RECT 2453.6600 2458.7600 2456.6600 2459.2400 ;
        RECT 2453.6600 2464.2000 2456.6600 2464.6800 ;
        RECT 2442.1200 2453.3200 2443.7200 2453.8000 ;
        RECT 2442.1200 2458.7600 2443.7200 2459.2400 ;
        RECT 2442.1200 2464.2000 2443.7200 2464.6800 ;
        RECT 2453.6600 2442.4400 2456.6600 2442.9200 ;
        RECT 2453.6600 2447.8800 2456.6600 2448.3600 ;
        RECT 2442.1200 2442.4400 2443.7200 2442.9200 ;
        RECT 2442.1200 2447.8800 2443.7200 2448.3600 ;
        RECT 2453.6600 2426.1200 2456.6600 2426.6000 ;
        RECT 2453.6600 2431.5600 2456.6600 2432.0400 ;
        RECT 2453.6600 2437.0000 2456.6600 2437.4800 ;
        RECT 2442.1200 2426.1200 2443.7200 2426.6000 ;
        RECT 2442.1200 2431.5600 2443.7200 2432.0400 ;
        RECT 2442.1200 2437.0000 2443.7200 2437.4800 ;
        RECT 2397.1200 2469.6400 2398.7200 2470.1200 ;
        RECT 2397.1200 2475.0800 2398.7200 2475.5600 ;
        RECT 2397.1200 2453.3200 2398.7200 2453.8000 ;
        RECT 2397.1200 2458.7600 2398.7200 2459.2400 ;
        RECT 2397.1200 2464.2000 2398.7200 2464.6800 ;
        RECT 2397.1200 2442.4400 2398.7200 2442.9200 ;
        RECT 2397.1200 2447.8800 2398.7200 2448.3600 ;
        RECT 2397.1200 2426.1200 2398.7200 2426.6000 ;
        RECT 2397.1200 2431.5600 2398.7200 2432.0400 ;
        RECT 2397.1200 2437.0000 2398.7200 2437.4800 ;
        RECT 2453.6600 2415.2400 2456.6600 2415.7200 ;
        RECT 2453.6600 2420.6800 2456.6600 2421.1600 ;
        RECT 2442.1200 2415.2400 2443.7200 2415.7200 ;
        RECT 2442.1200 2420.6800 2443.7200 2421.1600 ;
        RECT 2453.6600 2398.9200 2456.6600 2399.4000 ;
        RECT 2453.6600 2404.3600 2456.6600 2404.8400 ;
        RECT 2453.6600 2409.8000 2456.6600 2410.2800 ;
        RECT 2442.1200 2398.9200 2443.7200 2399.4000 ;
        RECT 2442.1200 2404.3600 2443.7200 2404.8400 ;
        RECT 2442.1200 2409.8000 2443.7200 2410.2800 ;
        RECT 2453.6600 2388.0400 2456.6600 2388.5200 ;
        RECT 2453.6600 2393.4800 2456.6600 2393.9600 ;
        RECT 2442.1200 2388.0400 2443.7200 2388.5200 ;
        RECT 2442.1200 2393.4800 2443.7200 2393.9600 ;
        RECT 2453.6600 2382.6000 2456.6600 2383.0800 ;
        RECT 2442.1200 2382.6000 2443.7200 2383.0800 ;
        RECT 2397.1200 2415.2400 2398.7200 2415.7200 ;
        RECT 2397.1200 2420.6800 2398.7200 2421.1600 ;
        RECT 2397.1200 2398.9200 2398.7200 2399.4000 ;
        RECT 2397.1200 2404.3600 2398.7200 2404.8400 ;
        RECT 2397.1200 2409.8000 2398.7200 2410.2800 ;
        RECT 2397.1200 2388.0400 2398.7200 2388.5200 ;
        RECT 2397.1200 2393.4800 2398.7200 2393.9600 ;
        RECT 2397.1200 2382.6000 2398.7200 2383.0800 ;
        RECT 2352.1200 2469.6400 2353.7200 2470.1200 ;
        RECT 2352.1200 2475.0800 2353.7200 2475.5600 ;
        RECT 2352.1200 2453.3200 2353.7200 2453.8000 ;
        RECT 2352.1200 2458.7600 2353.7200 2459.2400 ;
        RECT 2352.1200 2464.2000 2353.7200 2464.6800 ;
        RECT 2307.1200 2469.6400 2308.7200 2470.1200 ;
        RECT 2307.1200 2475.0800 2308.7200 2475.5600 ;
        RECT 2307.1200 2453.3200 2308.7200 2453.8000 ;
        RECT 2307.1200 2458.7600 2308.7200 2459.2400 ;
        RECT 2307.1200 2464.2000 2308.7200 2464.6800 ;
        RECT 2352.1200 2442.4400 2353.7200 2442.9200 ;
        RECT 2352.1200 2447.8800 2353.7200 2448.3600 ;
        RECT 2352.1200 2426.1200 2353.7200 2426.6000 ;
        RECT 2352.1200 2431.5600 2353.7200 2432.0400 ;
        RECT 2352.1200 2437.0000 2353.7200 2437.4800 ;
        RECT 2307.1200 2442.4400 2308.7200 2442.9200 ;
        RECT 2307.1200 2447.8800 2308.7200 2448.3600 ;
        RECT 2307.1200 2426.1200 2308.7200 2426.6000 ;
        RECT 2307.1200 2431.5600 2308.7200 2432.0400 ;
        RECT 2307.1200 2437.0000 2308.7200 2437.4800 ;
        RECT 2257.5600 2469.6400 2260.5600 2470.1200 ;
        RECT 2257.5600 2475.0800 2260.5600 2475.5600 ;
        RECT 2257.5600 2458.7600 2260.5600 2459.2400 ;
        RECT 2257.5600 2453.3200 2260.5600 2453.8000 ;
        RECT 2257.5600 2464.2000 2260.5600 2464.6800 ;
        RECT 2257.5600 2442.4400 2260.5600 2442.9200 ;
        RECT 2257.5600 2447.8800 2260.5600 2448.3600 ;
        RECT 2257.5600 2431.5600 2260.5600 2432.0400 ;
        RECT 2257.5600 2426.1200 2260.5600 2426.6000 ;
        RECT 2257.5600 2437.0000 2260.5600 2437.4800 ;
        RECT 2352.1200 2415.2400 2353.7200 2415.7200 ;
        RECT 2352.1200 2420.6800 2353.7200 2421.1600 ;
        RECT 2352.1200 2398.9200 2353.7200 2399.4000 ;
        RECT 2352.1200 2404.3600 2353.7200 2404.8400 ;
        RECT 2352.1200 2409.8000 2353.7200 2410.2800 ;
        RECT 2307.1200 2415.2400 2308.7200 2415.7200 ;
        RECT 2307.1200 2420.6800 2308.7200 2421.1600 ;
        RECT 2307.1200 2398.9200 2308.7200 2399.4000 ;
        RECT 2307.1200 2404.3600 2308.7200 2404.8400 ;
        RECT 2307.1200 2409.8000 2308.7200 2410.2800 ;
        RECT 2352.1200 2393.4800 2353.7200 2393.9600 ;
        RECT 2352.1200 2388.0400 2353.7200 2388.5200 ;
        RECT 2352.1200 2382.6000 2353.7200 2383.0800 ;
        RECT 2307.1200 2393.4800 2308.7200 2393.9600 ;
        RECT 2307.1200 2388.0400 2308.7200 2388.5200 ;
        RECT 2307.1200 2382.6000 2308.7200 2383.0800 ;
        RECT 2257.5600 2415.2400 2260.5600 2415.7200 ;
        RECT 2257.5600 2420.6800 2260.5600 2421.1600 ;
        RECT 2257.5600 2404.3600 2260.5600 2404.8400 ;
        RECT 2257.5600 2398.9200 2260.5600 2399.4000 ;
        RECT 2257.5600 2409.8000 2260.5600 2410.2800 ;
        RECT 2257.5600 2388.0400 2260.5600 2388.5200 ;
        RECT 2257.5600 2393.4800 2260.5600 2393.9600 ;
        RECT 2257.5600 2382.6000 2260.5600 2383.0800 ;
        RECT 2257.5600 2580.7900 2456.6600 2583.7900 ;
        RECT 2257.5600 2375.6900 2456.6600 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 2146.0500 2443.7200 2354.1500 ;
        RECT 2397.1200 2146.0500 2398.7200 2354.1500 ;
        RECT 2352.1200 2146.0500 2353.7200 2354.1500 ;
        RECT 2307.1200 2146.0500 2308.7200 2354.1500 ;
        RECT 2453.6600 2146.0500 2456.6600 2354.1500 ;
        RECT 2257.5600 2146.0500 2260.5600 2354.1500 ;
      LAYER met3 ;
        RECT 2453.6600 2348.8000 2456.6600 2349.2800 ;
        RECT 2442.1200 2348.8000 2443.7200 2349.2800 ;
        RECT 2453.6600 2337.9200 2456.6600 2338.4000 ;
        RECT 2453.6600 2343.3600 2456.6600 2343.8400 ;
        RECT 2442.1200 2337.9200 2443.7200 2338.4000 ;
        RECT 2442.1200 2343.3600 2443.7200 2343.8400 ;
        RECT 2453.6600 2321.6000 2456.6600 2322.0800 ;
        RECT 2453.6600 2327.0400 2456.6600 2327.5200 ;
        RECT 2442.1200 2321.6000 2443.7200 2322.0800 ;
        RECT 2442.1200 2327.0400 2443.7200 2327.5200 ;
        RECT 2453.6600 2310.7200 2456.6600 2311.2000 ;
        RECT 2453.6600 2316.1600 2456.6600 2316.6400 ;
        RECT 2442.1200 2310.7200 2443.7200 2311.2000 ;
        RECT 2442.1200 2316.1600 2443.7200 2316.6400 ;
        RECT 2453.6600 2332.4800 2456.6600 2332.9600 ;
        RECT 2442.1200 2332.4800 2443.7200 2332.9600 ;
        RECT 2397.1200 2337.9200 2398.7200 2338.4000 ;
        RECT 2397.1200 2343.3600 2398.7200 2343.8400 ;
        RECT 2397.1200 2348.8000 2398.7200 2349.2800 ;
        RECT 2397.1200 2321.6000 2398.7200 2322.0800 ;
        RECT 2397.1200 2327.0400 2398.7200 2327.5200 ;
        RECT 2397.1200 2316.1600 2398.7200 2316.6400 ;
        RECT 2397.1200 2310.7200 2398.7200 2311.2000 ;
        RECT 2397.1200 2332.4800 2398.7200 2332.9600 ;
        RECT 2453.6600 2294.4000 2456.6600 2294.8800 ;
        RECT 2453.6600 2299.8400 2456.6600 2300.3200 ;
        RECT 2442.1200 2294.4000 2443.7200 2294.8800 ;
        RECT 2442.1200 2299.8400 2443.7200 2300.3200 ;
        RECT 2453.6600 2278.0800 2456.6600 2278.5600 ;
        RECT 2453.6600 2283.5200 2456.6600 2284.0000 ;
        RECT 2453.6600 2288.9600 2456.6600 2289.4400 ;
        RECT 2442.1200 2278.0800 2443.7200 2278.5600 ;
        RECT 2442.1200 2283.5200 2443.7200 2284.0000 ;
        RECT 2442.1200 2288.9600 2443.7200 2289.4400 ;
        RECT 2453.6600 2267.2000 2456.6600 2267.6800 ;
        RECT 2453.6600 2272.6400 2456.6600 2273.1200 ;
        RECT 2442.1200 2267.2000 2443.7200 2267.6800 ;
        RECT 2442.1200 2272.6400 2443.7200 2273.1200 ;
        RECT 2453.6600 2250.8800 2456.6600 2251.3600 ;
        RECT 2453.6600 2256.3200 2456.6600 2256.8000 ;
        RECT 2453.6600 2261.7600 2456.6600 2262.2400 ;
        RECT 2442.1200 2250.8800 2443.7200 2251.3600 ;
        RECT 2442.1200 2256.3200 2443.7200 2256.8000 ;
        RECT 2442.1200 2261.7600 2443.7200 2262.2400 ;
        RECT 2397.1200 2294.4000 2398.7200 2294.8800 ;
        RECT 2397.1200 2299.8400 2398.7200 2300.3200 ;
        RECT 2397.1200 2278.0800 2398.7200 2278.5600 ;
        RECT 2397.1200 2283.5200 2398.7200 2284.0000 ;
        RECT 2397.1200 2288.9600 2398.7200 2289.4400 ;
        RECT 2397.1200 2267.2000 2398.7200 2267.6800 ;
        RECT 2397.1200 2272.6400 2398.7200 2273.1200 ;
        RECT 2397.1200 2250.8800 2398.7200 2251.3600 ;
        RECT 2397.1200 2256.3200 2398.7200 2256.8000 ;
        RECT 2397.1200 2261.7600 2398.7200 2262.2400 ;
        RECT 2453.6600 2305.2800 2456.6600 2305.7600 ;
        RECT 2397.1200 2305.2800 2398.7200 2305.7600 ;
        RECT 2442.1200 2305.2800 2443.7200 2305.7600 ;
        RECT 2352.1200 2337.9200 2353.7200 2338.4000 ;
        RECT 2352.1200 2343.3600 2353.7200 2343.8400 ;
        RECT 2352.1200 2348.8000 2353.7200 2349.2800 ;
        RECT 2307.1200 2337.9200 2308.7200 2338.4000 ;
        RECT 2307.1200 2343.3600 2308.7200 2343.8400 ;
        RECT 2307.1200 2348.8000 2308.7200 2349.2800 ;
        RECT 2352.1200 2321.6000 2353.7200 2322.0800 ;
        RECT 2352.1200 2327.0400 2353.7200 2327.5200 ;
        RECT 2352.1200 2310.7200 2353.7200 2311.2000 ;
        RECT 2352.1200 2316.1600 2353.7200 2316.6400 ;
        RECT 2307.1200 2321.6000 2308.7200 2322.0800 ;
        RECT 2307.1200 2327.0400 2308.7200 2327.5200 ;
        RECT 2307.1200 2310.7200 2308.7200 2311.2000 ;
        RECT 2307.1200 2316.1600 2308.7200 2316.6400 ;
        RECT 2307.1200 2332.4800 2308.7200 2332.9600 ;
        RECT 2352.1200 2332.4800 2353.7200 2332.9600 ;
        RECT 2257.5600 2348.8000 2260.5600 2349.2800 ;
        RECT 2257.5600 2343.3600 2260.5600 2343.8400 ;
        RECT 2257.5600 2337.9200 2260.5600 2338.4000 ;
        RECT 2257.5600 2327.0400 2260.5600 2327.5200 ;
        RECT 2257.5600 2321.6000 2260.5600 2322.0800 ;
        RECT 2257.5600 2316.1600 2260.5600 2316.6400 ;
        RECT 2257.5600 2310.7200 2260.5600 2311.2000 ;
        RECT 2257.5600 2332.4800 2260.5600 2332.9600 ;
        RECT 2352.1200 2294.4000 2353.7200 2294.8800 ;
        RECT 2352.1200 2299.8400 2353.7200 2300.3200 ;
        RECT 2352.1200 2278.0800 2353.7200 2278.5600 ;
        RECT 2352.1200 2283.5200 2353.7200 2284.0000 ;
        RECT 2352.1200 2288.9600 2353.7200 2289.4400 ;
        RECT 2307.1200 2294.4000 2308.7200 2294.8800 ;
        RECT 2307.1200 2299.8400 2308.7200 2300.3200 ;
        RECT 2307.1200 2278.0800 2308.7200 2278.5600 ;
        RECT 2307.1200 2283.5200 2308.7200 2284.0000 ;
        RECT 2307.1200 2288.9600 2308.7200 2289.4400 ;
        RECT 2352.1200 2267.2000 2353.7200 2267.6800 ;
        RECT 2352.1200 2272.6400 2353.7200 2273.1200 ;
        RECT 2352.1200 2250.8800 2353.7200 2251.3600 ;
        RECT 2352.1200 2256.3200 2353.7200 2256.8000 ;
        RECT 2352.1200 2261.7600 2353.7200 2262.2400 ;
        RECT 2307.1200 2267.2000 2308.7200 2267.6800 ;
        RECT 2307.1200 2272.6400 2308.7200 2273.1200 ;
        RECT 2307.1200 2250.8800 2308.7200 2251.3600 ;
        RECT 2307.1200 2256.3200 2308.7200 2256.8000 ;
        RECT 2307.1200 2261.7600 2308.7200 2262.2400 ;
        RECT 2257.5600 2294.4000 2260.5600 2294.8800 ;
        RECT 2257.5600 2299.8400 2260.5600 2300.3200 ;
        RECT 2257.5600 2283.5200 2260.5600 2284.0000 ;
        RECT 2257.5600 2278.0800 2260.5600 2278.5600 ;
        RECT 2257.5600 2288.9600 2260.5600 2289.4400 ;
        RECT 2257.5600 2267.2000 2260.5600 2267.6800 ;
        RECT 2257.5600 2272.6400 2260.5600 2273.1200 ;
        RECT 2257.5600 2256.3200 2260.5600 2256.8000 ;
        RECT 2257.5600 2250.8800 2260.5600 2251.3600 ;
        RECT 2257.5600 2261.7600 2260.5600 2262.2400 ;
        RECT 2257.5600 2305.2800 2260.5600 2305.7600 ;
        RECT 2307.1200 2305.2800 2308.7200 2305.7600 ;
        RECT 2352.1200 2305.2800 2353.7200 2305.7600 ;
        RECT 2453.6600 2240.0000 2456.6600 2240.4800 ;
        RECT 2453.6600 2245.4400 2456.6600 2245.9200 ;
        RECT 2442.1200 2240.0000 2443.7200 2240.4800 ;
        RECT 2442.1200 2245.4400 2443.7200 2245.9200 ;
        RECT 2453.6600 2223.6800 2456.6600 2224.1600 ;
        RECT 2453.6600 2229.1200 2456.6600 2229.6000 ;
        RECT 2453.6600 2234.5600 2456.6600 2235.0400 ;
        RECT 2442.1200 2223.6800 2443.7200 2224.1600 ;
        RECT 2442.1200 2229.1200 2443.7200 2229.6000 ;
        RECT 2442.1200 2234.5600 2443.7200 2235.0400 ;
        RECT 2453.6600 2212.8000 2456.6600 2213.2800 ;
        RECT 2453.6600 2218.2400 2456.6600 2218.7200 ;
        RECT 2442.1200 2212.8000 2443.7200 2213.2800 ;
        RECT 2442.1200 2218.2400 2443.7200 2218.7200 ;
        RECT 2453.6600 2196.4800 2456.6600 2196.9600 ;
        RECT 2453.6600 2201.9200 2456.6600 2202.4000 ;
        RECT 2453.6600 2207.3600 2456.6600 2207.8400 ;
        RECT 2442.1200 2196.4800 2443.7200 2196.9600 ;
        RECT 2442.1200 2201.9200 2443.7200 2202.4000 ;
        RECT 2442.1200 2207.3600 2443.7200 2207.8400 ;
        RECT 2397.1200 2240.0000 2398.7200 2240.4800 ;
        RECT 2397.1200 2245.4400 2398.7200 2245.9200 ;
        RECT 2397.1200 2223.6800 2398.7200 2224.1600 ;
        RECT 2397.1200 2229.1200 2398.7200 2229.6000 ;
        RECT 2397.1200 2234.5600 2398.7200 2235.0400 ;
        RECT 2397.1200 2212.8000 2398.7200 2213.2800 ;
        RECT 2397.1200 2218.2400 2398.7200 2218.7200 ;
        RECT 2397.1200 2196.4800 2398.7200 2196.9600 ;
        RECT 2397.1200 2201.9200 2398.7200 2202.4000 ;
        RECT 2397.1200 2207.3600 2398.7200 2207.8400 ;
        RECT 2453.6600 2185.6000 2456.6600 2186.0800 ;
        RECT 2453.6600 2191.0400 2456.6600 2191.5200 ;
        RECT 2442.1200 2185.6000 2443.7200 2186.0800 ;
        RECT 2442.1200 2191.0400 2443.7200 2191.5200 ;
        RECT 2453.6600 2169.2800 2456.6600 2169.7600 ;
        RECT 2453.6600 2174.7200 2456.6600 2175.2000 ;
        RECT 2453.6600 2180.1600 2456.6600 2180.6400 ;
        RECT 2442.1200 2169.2800 2443.7200 2169.7600 ;
        RECT 2442.1200 2174.7200 2443.7200 2175.2000 ;
        RECT 2442.1200 2180.1600 2443.7200 2180.6400 ;
        RECT 2453.6600 2158.4000 2456.6600 2158.8800 ;
        RECT 2453.6600 2163.8400 2456.6600 2164.3200 ;
        RECT 2442.1200 2158.4000 2443.7200 2158.8800 ;
        RECT 2442.1200 2163.8400 2443.7200 2164.3200 ;
        RECT 2453.6600 2152.9600 2456.6600 2153.4400 ;
        RECT 2442.1200 2152.9600 2443.7200 2153.4400 ;
        RECT 2397.1200 2185.6000 2398.7200 2186.0800 ;
        RECT 2397.1200 2191.0400 2398.7200 2191.5200 ;
        RECT 2397.1200 2169.2800 2398.7200 2169.7600 ;
        RECT 2397.1200 2174.7200 2398.7200 2175.2000 ;
        RECT 2397.1200 2180.1600 2398.7200 2180.6400 ;
        RECT 2397.1200 2158.4000 2398.7200 2158.8800 ;
        RECT 2397.1200 2163.8400 2398.7200 2164.3200 ;
        RECT 2397.1200 2152.9600 2398.7200 2153.4400 ;
        RECT 2352.1200 2240.0000 2353.7200 2240.4800 ;
        RECT 2352.1200 2245.4400 2353.7200 2245.9200 ;
        RECT 2352.1200 2223.6800 2353.7200 2224.1600 ;
        RECT 2352.1200 2229.1200 2353.7200 2229.6000 ;
        RECT 2352.1200 2234.5600 2353.7200 2235.0400 ;
        RECT 2307.1200 2240.0000 2308.7200 2240.4800 ;
        RECT 2307.1200 2245.4400 2308.7200 2245.9200 ;
        RECT 2307.1200 2223.6800 2308.7200 2224.1600 ;
        RECT 2307.1200 2229.1200 2308.7200 2229.6000 ;
        RECT 2307.1200 2234.5600 2308.7200 2235.0400 ;
        RECT 2352.1200 2212.8000 2353.7200 2213.2800 ;
        RECT 2352.1200 2218.2400 2353.7200 2218.7200 ;
        RECT 2352.1200 2196.4800 2353.7200 2196.9600 ;
        RECT 2352.1200 2201.9200 2353.7200 2202.4000 ;
        RECT 2352.1200 2207.3600 2353.7200 2207.8400 ;
        RECT 2307.1200 2212.8000 2308.7200 2213.2800 ;
        RECT 2307.1200 2218.2400 2308.7200 2218.7200 ;
        RECT 2307.1200 2196.4800 2308.7200 2196.9600 ;
        RECT 2307.1200 2201.9200 2308.7200 2202.4000 ;
        RECT 2307.1200 2207.3600 2308.7200 2207.8400 ;
        RECT 2257.5600 2240.0000 2260.5600 2240.4800 ;
        RECT 2257.5600 2245.4400 2260.5600 2245.9200 ;
        RECT 2257.5600 2229.1200 2260.5600 2229.6000 ;
        RECT 2257.5600 2223.6800 2260.5600 2224.1600 ;
        RECT 2257.5600 2234.5600 2260.5600 2235.0400 ;
        RECT 2257.5600 2212.8000 2260.5600 2213.2800 ;
        RECT 2257.5600 2218.2400 2260.5600 2218.7200 ;
        RECT 2257.5600 2201.9200 2260.5600 2202.4000 ;
        RECT 2257.5600 2196.4800 2260.5600 2196.9600 ;
        RECT 2257.5600 2207.3600 2260.5600 2207.8400 ;
        RECT 2352.1200 2185.6000 2353.7200 2186.0800 ;
        RECT 2352.1200 2191.0400 2353.7200 2191.5200 ;
        RECT 2352.1200 2169.2800 2353.7200 2169.7600 ;
        RECT 2352.1200 2174.7200 2353.7200 2175.2000 ;
        RECT 2352.1200 2180.1600 2353.7200 2180.6400 ;
        RECT 2307.1200 2185.6000 2308.7200 2186.0800 ;
        RECT 2307.1200 2191.0400 2308.7200 2191.5200 ;
        RECT 2307.1200 2169.2800 2308.7200 2169.7600 ;
        RECT 2307.1200 2174.7200 2308.7200 2175.2000 ;
        RECT 2307.1200 2180.1600 2308.7200 2180.6400 ;
        RECT 2352.1200 2163.8400 2353.7200 2164.3200 ;
        RECT 2352.1200 2158.4000 2353.7200 2158.8800 ;
        RECT 2352.1200 2152.9600 2353.7200 2153.4400 ;
        RECT 2307.1200 2163.8400 2308.7200 2164.3200 ;
        RECT 2307.1200 2158.4000 2308.7200 2158.8800 ;
        RECT 2307.1200 2152.9600 2308.7200 2153.4400 ;
        RECT 2257.5600 2185.6000 2260.5600 2186.0800 ;
        RECT 2257.5600 2191.0400 2260.5600 2191.5200 ;
        RECT 2257.5600 2174.7200 2260.5600 2175.2000 ;
        RECT 2257.5600 2169.2800 2260.5600 2169.7600 ;
        RECT 2257.5600 2180.1600 2260.5600 2180.6400 ;
        RECT 2257.5600 2158.4000 2260.5600 2158.8800 ;
        RECT 2257.5600 2163.8400 2260.5600 2164.3200 ;
        RECT 2257.5600 2152.9600 2260.5600 2153.4400 ;
        RECT 2257.5600 2351.1500 2456.6600 2354.1500 ;
        RECT 2257.5600 2146.0500 2456.6600 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 1916.4100 2443.7200 2124.5100 ;
        RECT 2397.1200 1916.4100 2398.7200 2124.5100 ;
        RECT 2352.1200 1916.4100 2353.7200 2124.5100 ;
        RECT 2307.1200 1916.4100 2308.7200 2124.5100 ;
        RECT 2453.6600 1916.4100 2456.6600 2124.5100 ;
        RECT 2257.5600 1916.4100 2260.5600 2124.5100 ;
      LAYER met3 ;
        RECT 2453.6600 2119.1600 2456.6600 2119.6400 ;
        RECT 2442.1200 2119.1600 2443.7200 2119.6400 ;
        RECT 2453.6600 2108.2800 2456.6600 2108.7600 ;
        RECT 2453.6600 2113.7200 2456.6600 2114.2000 ;
        RECT 2442.1200 2108.2800 2443.7200 2108.7600 ;
        RECT 2442.1200 2113.7200 2443.7200 2114.2000 ;
        RECT 2453.6600 2091.9600 2456.6600 2092.4400 ;
        RECT 2453.6600 2097.4000 2456.6600 2097.8800 ;
        RECT 2442.1200 2091.9600 2443.7200 2092.4400 ;
        RECT 2442.1200 2097.4000 2443.7200 2097.8800 ;
        RECT 2453.6600 2081.0800 2456.6600 2081.5600 ;
        RECT 2453.6600 2086.5200 2456.6600 2087.0000 ;
        RECT 2442.1200 2081.0800 2443.7200 2081.5600 ;
        RECT 2442.1200 2086.5200 2443.7200 2087.0000 ;
        RECT 2453.6600 2102.8400 2456.6600 2103.3200 ;
        RECT 2442.1200 2102.8400 2443.7200 2103.3200 ;
        RECT 2397.1200 2108.2800 2398.7200 2108.7600 ;
        RECT 2397.1200 2113.7200 2398.7200 2114.2000 ;
        RECT 2397.1200 2119.1600 2398.7200 2119.6400 ;
        RECT 2397.1200 2091.9600 2398.7200 2092.4400 ;
        RECT 2397.1200 2097.4000 2398.7200 2097.8800 ;
        RECT 2397.1200 2086.5200 2398.7200 2087.0000 ;
        RECT 2397.1200 2081.0800 2398.7200 2081.5600 ;
        RECT 2397.1200 2102.8400 2398.7200 2103.3200 ;
        RECT 2453.6600 2064.7600 2456.6600 2065.2400 ;
        RECT 2453.6600 2070.2000 2456.6600 2070.6800 ;
        RECT 2442.1200 2064.7600 2443.7200 2065.2400 ;
        RECT 2442.1200 2070.2000 2443.7200 2070.6800 ;
        RECT 2453.6600 2048.4400 2456.6600 2048.9200 ;
        RECT 2453.6600 2053.8800 2456.6600 2054.3600 ;
        RECT 2453.6600 2059.3200 2456.6600 2059.8000 ;
        RECT 2442.1200 2048.4400 2443.7200 2048.9200 ;
        RECT 2442.1200 2053.8800 2443.7200 2054.3600 ;
        RECT 2442.1200 2059.3200 2443.7200 2059.8000 ;
        RECT 2453.6600 2037.5600 2456.6600 2038.0400 ;
        RECT 2453.6600 2043.0000 2456.6600 2043.4800 ;
        RECT 2442.1200 2037.5600 2443.7200 2038.0400 ;
        RECT 2442.1200 2043.0000 2443.7200 2043.4800 ;
        RECT 2453.6600 2021.2400 2456.6600 2021.7200 ;
        RECT 2453.6600 2026.6800 2456.6600 2027.1600 ;
        RECT 2453.6600 2032.1200 2456.6600 2032.6000 ;
        RECT 2442.1200 2021.2400 2443.7200 2021.7200 ;
        RECT 2442.1200 2026.6800 2443.7200 2027.1600 ;
        RECT 2442.1200 2032.1200 2443.7200 2032.6000 ;
        RECT 2397.1200 2064.7600 2398.7200 2065.2400 ;
        RECT 2397.1200 2070.2000 2398.7200 2070.6800 ;
        RECT 2397.1200 2048.4400 2398.7200 2048.9200 ;
        RECT 2397.1200 2053.8800 2398.7200 2054.3600 ;
        RECT 2397.1200 2059.3200 2398.7200 2059.8000 ;
        RECT 2397.1200 2037.5600 2398.7200 2038.0400 ;
        RECT 2397.1200 2043.0000 2398.7200 2043.4800 ;
        RECT 2397.1200 2021.2400 2398.7200 2021.7200 ;
        RECT 2397.1200 2026.6800 2398.7200 2027.1600 ;
        RECT 2397.1200 2032.1200 2398.7200 2032.6000 ;
        RECT 2453.6600 2075.6400 2456.6600 2076.1200 ;
        RECT 2397.1200 2075.6400 2398.7200 2076.1200 ;
        RECT 2442.1200 2075.6400 2443.7200 2076.1200 ;
        RECT 2352.1200 2108.2800 2353.7200 2108.7600 ;
        RECT 2352.1200 2113.7200 2353.7200 2114.2000 ;
        RECT 2352.1200 2119.1600 2353.7200 2119.6400 ;
        RECT 2307.1200 2108.2800 2308.7200 2108.7600 ;
        RECT 2307.1200 2113.7200 2308.7200 2114.2000 ;
        RECT 2307.1200 2119.1600 2308.7200 2119.6400 ;
        RECT 2352.1200 2091.9600 2353.7200 2092.4400 ;
        RECT 2352.1200 2097.4000 2353.7200 2097.8800 ;
        RECT 2352.1200 2081.0800 2353.7200 2081.5600 ;
        RECT 2352.1200 2086.5200 2353.7200 2087.0000 ;
        RECT 2307.1200 2091.9600 2308.7200 2092.4400 ;
        RECT 2307.1200 2097.4000 2308.7200 2097.8800 ;
        RECT 2307.1200 2081.0800 2308.7200 2081.5600 ;
        RECT 2307.1200 2086.5200 2308.7200 2087.0000 ;
        RECT 2307.1200 2102.8400 2308.7200 2103.3200 ;
        RECT 2352.1200 2102.8400 2353.7200 2103.3200 ;
        RECT 2257.5600 2119.1600 2260.5600 2119.6400 ;
        RECT 2257.5600 2113.7200 2260.5600 2114.2000 ;
        RECT 2257.5600 2108.2800 2260.5600 2108.7600 ;
        RECT 2257.5600 2097.4000 2260.5600 2097.8800 ;
        RECT 2257.5600 2091.9600 2260.5600 2092.4400 ;
        RECT 2257.5600 2086.5200 2260.5600 2087.0000 ;
        RECT 2257.5600 2081.0800 2260.5600 2081.5600 ;
        RECT 2257.5600 2102.8400 2260.5600 2103.3200 ;
        RECT 2352.1200 2064.7600 2353.7200 2065.2400 ;
        RECT 2352.1200 2070.2000 2353.7200 2070.6800 ;
        RECT 2352.1200 2048.4400 2353.7200 2048.9200 ;
        RECT 2352.1200 2053.8800 2353.7200 2054.3600 ;
        RECT 2352.1200 2059.3200 2353.7200 2059.8000 ;
        RECT 2307.1200 2064.7600 2308.7200 2065.2400 ;
        RECT 2307.1200 2070.2000 2308.7200 2070.6800 ;
        RECT 2307.1200 2048.4400 2308.7200 2048.9200 ;
        RECT 2307.1200 2053.8800 2308.7200 2054.3600 ;
        RECT 2307.1200 2059.3200 2308.7200 2059.8000 ;
        RECT 2352.1200 2037.5600 2353.7200 2038.0400 ;
        RECT 2352.1200 2043.0000 2353.7200 2043.4800 ;
        RECT 2352.1200 2021.2400 2353.7200 2021.7200 ;
        RECT 2352.1200 2026.6800 2353.7200 2027.1600 ;
        RECT 2352.1200 2032.1200 2353.7200 2032.6000 ;
        RECT 2307.1200 2037.5600 2308.7200 2038.0400 ;
        RECT 2307.1200 2043.0000 2308.7200 2043.4800 ;
        RECT 2307.1200 2021.2400 2308.7200 2021.7200 ;
        RECT 2307.1200 2026.6800 2308.7200 2027.1600 ;
        RECT 2307.1200 2032.1200 2308.7200 2032.6000 ;
        RECT 2257.5600 2064.7600 2260.5600 2065.2400 ;
        RECT 2257.5600 2070.2000 2260.5600 2070.6800 ;
        RECT 2257.5600 2053.8800 2260.5600 2054.3600 ;
        RECT 2257.5600 2048.4400 2260.5600 2048.9200 ;
        RECT 2257.5600 2059.3200 2260.5600 2059.8000 ;
        RECT 2257.5600 2037.5600 2260.5600 2038.0400 ;
        RECT 2257.5600 2043.0000 2260.5600 2043.4800 ;
        RECT 2257.5600 2026.6800 2260.5600 2027.1600 ;
        RECT 2257.5600 2021.2400 2260.5600 2021.7200 ;
        RECT 2257.5600 2032.1200 2260.5600 2032.6000 ;
        RECT 2257.5600 2075.6400 2260.5600 2076.1200 ;
        RECT 2307.1200 2075.6400 2308.7200 2076.1200 ;
        RECT 2352.1200 2075.6400 2353.7200 2076.1200 ;
        RECT 2453.6600 2010.3600 2456.6600 2010.8400 ;
        RECT 2453.6600 2015.8000 2456.6600 2016.2800 ;
        RECT 2442.1200 2010.3600 2443.7200 2010.8400 ;
        RECT 2442.1200 2015.8000 2443.7200 2016.2800 ;
        RECT 2453.6600 1994.0400 2456.6600 1994.5200 ;
        RECT 2453.6600 1999.4800 2456.6600 1999.9600 ;
        RECT 2453.6600 2004.9200 2456.6600 2005.4000 ;
        RECT 2442.1200 1994.0400 2443.7200 1994.5200 ;
        RECT 2442.1200 1999.4800 2443.7200 1999.9600 ;
        RECT 2442.1200 2004.9200 2443.7200 2005.4000 ;
        RECT 2453.6600 1983.1600 2456.6600 1983.6400 ;
        RECT 2453.6600 1988.6000 2456.6600 1989.0800 ;
        RECT 2442.1200 1983.1600 2443.7200 1983.6400 ;
        RECT 2442.1200 1988.6000 2443.7200 1989.0800 ;
        RECT 2453.6600 1966.8400 2456.6600 1967.3200 ;
        RECT 2453.6600 1972.2800 2456.6600 1972.7600 ;
        RECT 2453.6600 1977.7200 2456.6600 1978.2000 ;
        RECT 2442.1200 1966.8400 2443.7200 1967.3200 ;
        RECT 2442.1200 1972.2800 2443.7200 1972.7600 ;
        RECT 2442.1200 1977.7200 2443.7200 1978.2000 ;
        RECT 2397.1200 2010.3600 2398.7200 2010.8400 ;
        RECT 2397.1200 2015.8000 2398.7200 2016.2800 ;
        RECT 2397.1200 1994.0400 2398.7200 1994.5200 ;
        RECT 2397.1200 1999.4800 2398.7200 1999.9600 ;
        RECT 2397.1200 2004.9200 2398.7200 2005.4000 ;
        RECT 2397.1200 1983.1600 2398.7200 1983.6400 ;
        RECT 2397.1200 1988.6000 2398.7200 1989.0800 ;
        RECT 2397.1200 1966.8400 2398.7200 1967.3200 ;
        RECT 2397.1200 1972.2800 2398.7200 1972.7600 ;
        RECT 2397.1200 1977.7200 2398.7200 1978.2000 ;
        RECT 2453.6600 1955.9600 2456.6600 1956.4400 ;
        RECT 2453.6600 1961.4000 2456.6600 1961.8800 ;
        RECT 2442.1200 1955.9600 2443.7200 1956.4400 ;
        RECT 2442.1200 1961.4000 2443.7200 1961.8800 ;
        RECT 2453.6600 1939.6400 2456.6600 1940.1200 ;
        RECT 2453.6600 1945.0800 2456.6600 1945.5600 ;
        RECT 2453.6600 1950.5200 2456.6600 1951.0000 ;
        RECT 2442.1200 1939.6400 2443.7200 1940.1200 ;
        RECT 2442.1200 1945.0800 2443.7200 1945.5600 ;
        RECT 2442.1200 1950.5200 2443.7200 1951.0000 ;
        RECT 2453.6600 1928.7600 2456.6600 1929.2400 ;
        RECT 2453.6600 1934.2000 2456.6600 1934.6800 ;
        RECT 2442.1200 1928.7600 2443.7200 1929.2400 ;
        RECT 2442.1200 1934.2000 2443.7200 1934.6800 ;
        RECT 2453.6600 1923.3200 2456.6600 1923.8000 ;
        RECT 2442.1200 1923.3200 2443.7200 1923.8000 ;
        RECT 2397.1200 1955.9600 2398.7200 1956.4400 ;
        RECT 2397.1200 1961.4000 2398.7200 1961.8800 ;
        RECT 2397.1200 1939.6400 2398.7200 1940.1200 ;
        RECT 2397.1200 1945.0800 2398.7200 1945.5600 ;
        RECT 2397.1200 1950.5200 2398.7200 1951.0000 ;
        RECT 2397.1200 1928.7600 2398.7200 1929.2400 ;
        RECT 2397.1200 1934.2000 2398.7200 1934.6800 ;
        RECT 2397.1200 1923.3200 2398.7200 1923.8000 ;
        RECT 2352.1200 2010.3600 2353.7200 2010.8400 ;
        RECT 2352.1200 2015.8000 2353.7200 2016.2800 ;
        RECT 2352.1200 1994.0400 2353.7200 1994.5200 ;
        RECT 2352.1200 1999.4800 2353.7200 1999.9600 ;
        RECT 2352.1200 2004.9200 2353.7200 2005.4000 ;
        RECT 2307.1200 2010.3600 2308.7200 2010.8400 ;
        RECT 2307.1200 2015.8000 2308.7200 2016.2800 ;
        RECT 2307.1200 1994.0400 2308.7200 1994.5200 ;
        RECT 2307.1200 1999.4800 2308.7200 1999.9600 ;
        RECT 2307.1200 2004.9200 2308.7200 2005.4000 ;
        RECT 2352.1200 1983.1600 2353.7200 1983.6400 ;
        RECT 2352.1200 1988.6000 2353.7200 1989.0800 ;
        RECT 2352.1200 1966.8400 2353.7200 1967.3200 ;
        RECT 2352.1200 1972.2800 2353.7200 1972.7600 ;
        RECT 2352.1200 1977.7200 2353.7200 1978.2000 ;
        RECT 2307.1200 1983.1600 2308.7200 1983.6400 ;
        RECT 2307.1200 1988.6000 2308.7200 1989.0800 ;
        RECT 2307.1200 1966.8400 2308.7200 1967.3200 ;
        RECT 2307.1200 1972.2800 2308.7200 1972.7600 ;
        RECT 2307.1200 1977.7200 2308.7200 1978.2000 ;
        RECT 2257.5600 2010.3600 2260.5600 2010.8400 ;
        RECT 2257.5600 2015.8000 2260.5600 2016.2800 ;
        RECT 2257.5600 1999.4800 2260.5600 1999.9600 ;
        RECT 2257.5600 1994.0400 2260.5600 1994.5200 ;
        RECT 2257.5600 2004.9200 2260.5600 2005.4000 ;
        RECT 2257.5600 1983.1600 2260.5600 1983.6400 ;
        RECT 2257.5600 1988.6000 2260.5600 1989.0800 ;
        RECT 2257.5600 1972.2800 2260.5600 1972.7600 ;
        RECT 2257.5600 1966.8400 2260.5600 1967.3200 ;
        RECT 2257.5600 1977.7200 2260.5600 1978.2000 ;
        RECT 2352.1200 1955.9600 2353.7200 1956.4400 ;
        RECT 2352.1200 1961.4000 2353.7200 1961.8800 ;
        RECT 2352.1200 1939.6400 2353.7200 1940.1200 ;
        RECT 2352.1200 1945.0800 2353.7200 1945.5600 ;
        RECT 2352.1200 1950.5200 2353.7200 1951.0000 ;
        RECT 2307.1200 1955.9600 2308.7200 1956.4400 ;
        RECT 2307.1200 1961.4000 2308.7200 1961.8800 ;
        RECT 2307.1200 1939.6400 2308.7200 1940.1200 ;
        RECT 2307.1200 1945.0800 2308.7200 1945.5600 ;
        RECT 2307.1200 1950.5200 2308.7200 1951.0000 ;
        RECT 2352.1200 1934.2000 2353.7200 1934.6800 ;
        RECT 2352.1200 1928.7600 2353.7200 1929.2400 ;
        RECT 2352.1200 1923.3200 2353.7200 1923.8000 ;
        RECT 2307.1200 1934.2000 2308.7200 1934.6800 ;
        RECT 2307.1200 1928.7600 2308.7200 1929.2400 ;
        RECT 2307.1200 1923.3200 2308.7200 1923.8000 ;
        RECT 2257.5600 1955.9600 2260.5600 1956.4400 ;
        RECT 2257.5600 1961.4000 2260.5600 1961.8800 ;
        RECT 2257.5600 1945.0800 2260.5600 1945.5600 ;
        RECT 2257.5600 1939.6400 2260.5600 1940.1200 ;
        RECT 2257.5600 1950.5200 2260.5600 1951.0000 ;
        RECT 2257.5600 1928.7600 2260.5600 1929.2400 ;
        RECT 2257.5600 1934.2000 2260.5600 1934.6800 ;
        RECT 2257.5600 1923.3200 2260.5600 1923.8000 ;
        RECT 2257.5600 2121.5100 2456.6600 2124.5100 ;
        RECT 2257.5600 1916.4100 2456.6600 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 1686.7700 2443.7200 1894.8700 ;
        RECT 2397.1200 1686.7700 2398.7200 1894.8700 ;
        RECT 2352.1200 1686.7700 2353.7200 1894.8700 ;
        RECT 2307.1200 1686.7700 2308.7200 1894.8700 ;
        RECT 2453.6600 1686.7700 2456.6600 1894.8700 ;
        RECT 2257.5600 1686.7700 2260.5600 1894.8700 ;
      LAYER met3 ;
        RECT 2453.6600 1889.5200 2456.6600 1890.0000 ;
        RECT 2442.1200 1889.5200 2443.7200 1890.0000 ;
        RECT 2453.6600 1878.6400 2456.6600 1879.1200 ;
        RECT 2453.6600 1884.0800 2456.6600 1884.5600 ;
        RECT 2442.1200 1878.6400 2443.7200 1879.1200 ;
        RECT 2442.1200 1884.0800 2443.7200 1884.5600 ;
        RECT 2453.6600 1862.3200 2456.6600 1862.8000 ;
        RECT 2453.6600 1867.7600 2456.6600 1868.2400 ;
        RECT 2442.1200 1862.3200 2443.7200 1862.8000 ;
        RECT 2442.1200 1867.7600 2443.7200 1868.2400 ;
        RECT 2453.6600 1851.4400 2456.6600 1851.9200 ;
        RECT 2453.6600 1856.8800 2456.6600 1857.3600 ;
        RECT 2442.1200 1851.4400 2443.7200 1851.9200 ;
        RECT 2442.1200 1856.8800 2443.7200 1857.3600 ;
        RECT 2453.6600 1873.2000 2456.6600 1873.6800 ;
        RECT 2442.1200 1873.2000 2443.7200 1873.6800 ;
        RECT 2397.1200 1878.6400 2398.7200 1879.1200 ;
        RECT 2397.1200 1884.0800 2398.7200 1884.5600 ;
        RECT 2397.1200 1889.5200 2398.7200 1890.0000 ;
        RECT 2397.1200 1862.3200 2398.7200 1862.8000 ;
        RECT 2397.1200 1867.7600 2398.7200 1868.2400 ;
        RECT 2397.1200 1856.8800 2398.7200 1857.3600 ;
        RECT 2397.1200 1851.4400 2398.7200 1851.9200 ;
        RECT 2397.1200 1873.2000 2398.7200 1873.6800 ;
        RECT 2453.6600 1835.1200 2456.6600 1835.6000 ;
        RECT 2453.6600 1840.5600 2456.6600 1841.0400 ;
        RECT 2442.1200 1835.1200 2443.7200 1835.6000 ;
        RECT 2442.1200 1840.5600 2443.7200 1841.0400 ;
        RECT 2453.6600 1818.8000 2456.6600 1819.2800 ;
        RECT 2453.6600 1824.2400 2456.6600 1824.7200 ;
        RECT 2453.6600 1829.6800 2456.6600 1830.1600 ;
        RECT 2442.1200 1818.8000 2443.7200 1819.2800 ;
        RECT 2442.1200 1824.2400 2443.7200 1824.7200 ;
        RECT 2442.1200 1829.6800 2443.7200 1830.1600 ;
        RECT 2453.6600 1807.9200 2456.6600 1808.4000 ;
        RECT 2453.6600 1813.3600 2456.6600 1813.8400 ;
        RECT 2442.1200 1807.9200 2443.7200 1808.4000 ;
        RECT 2442.1200 1813.3600 2443.7200 1813.8400 ;
        RECT 2453.6600 1791.6000 2456.6600 1792.0800 ;
        RECT 2453.6600 1797.0400 2456.6600 1797.5200 ;
        RECT 2453.6600 1802.4800 2456.6600 1802.9600 ;
        RECT 2442.1200 1791.6000 2443.7200 1792.0800 ;
        RECT 2442.1200 1797.0400 2443.7200 1797.5200 ;
        RECT 2442.1200 1802.4800 2443.7200 1802.9600 ;
        RECT 2397.1200 1835.1200 2398.7200 1835.6000 ;
        RECT 2397.1200 1840.5600 2398.7200 1841.0400 ;
        RECT 2397.1200 1818.8000 2398.7200 1819.2800 ;
        RECT 2397.1200 1824.2400 2398.7200 1824.7200 ;
        RECT 2397.1200 1829.6800 2398.7200 1830.1600 ;
        RECT 2397.1200 1807.9200 2398.7200 1808.4000 ;
        RECT 2397.1200 1813.3600 2398.7200 1813.8400 ;
        RECT 2397.1200 1791.6000 2398.7200 1792.0800 ;
        RECT 2397.1200 1797.0400 2398.7200 1797.5200 ;
        RECT 2397.1200 1802.4800 2398.7200 1802.9600 ;
        RECT 2453.6600 1846.0000 2456.6600 1846.4800 ;
        RECT 2397.1200 1846.0000 2398.7200 1846.4800 ;
        RECT 2442.1200 1846.0000 2443.7200 1846.4800 ;
        RECT 2352.1200 1878.6400 2353.7200 1879.1200 ;
        RECT 2352.1200 1884.0800 2353.7200 1884.5600 ;
        RECT 2352.1200 1889.5200 2353.7200 1890.0000 ;
        RECT 2307.1200 1878.6400 2308.7200 1879.1200 ;
        RECT 2307.1200 1884.0800 2308.7200 1884.5600 ;
        RECT 2307.1200 1889.5200 2308.7200 1890.0000 ;
        RECT 2352.1200 1862.3200 2353.7200 1862.8000 ;
        RECT 2352.1200 1867.7600 2353.7200 1868.2400 ;
        RECT 2352.1200 1851.4400 2353.7200 1851.9200 ;
        RECT 2352.1200 1856.8800 2353.7200 1857.3600 ;
        RECT 2307.1200 1862.3200 2308.7200 1862.8000 ;
        RECT 2307.1200 1867.7600 2308.7200 1868.2400 ;
        RECT 2307.1200 1851.4400 2308.7200 1851.9200 ;
        RECT 2307.1200 1856.8800 2308.7200 1857.3600 ;
        RECT 2307.1200 1873.2000 2308.7200 1873.6800 ;
        RECT 2352.1200 1873.2000 2353.7200 1873.6800 ;
        RECT 2257.5600 1889.5200 2260.5600 1890.0000 ;
        RECT 2257.5600 1884.0800 2260.5600 1884.5600 ;
        RECT 2257.5600 1878.6400 2260.5600 1879.1200 ;
        RECT 2257.5600 1867.7600 2260.5600 1868.2400 ;
        RECT 2257.5600 1862.3200 2260.5600 1862.8000 ;
        RECT 2257.5600 1856.8800 2260.5600 1857.3600 ;
        RECT 2257.5600 1851.4400 2260.5600 1851.9200 ;
        RECT 2257.5600 1873.2000 2260.5600 1873.6800 ;
        RECT 2352.1200 1835.1200 2353.7200 1835.6000 ;
        RECT 2352.1200 1840.5600 2353.7200 1841.0400 ;
        RECT 2352.1200 1818.8000 2353.7200 1819.2800 ;
        RECT 2352.1200 1824.2400 2353.7200 1824.7200 ;
        RECT 2352.1200 1829.6800 2353.7200 1830.1600 ;
        RECT 2307.1200 1835.1200 2308.7200 1835.6000 ;
        RECT 2307.1200 1840.5600 2308.7200 1841.0400 ;
        RECT 2307.1200 1818.8000 2308.7200 1819.2800 ;
        RECT 2307.1200 1824.2400 2308.7200 1824.7200 ;
        RECT 2307.1200 1829.6800 2308.7200 1830.1600 ;
        RECT 2352.1200 1807.9200 2353.7200 1808.4000 ;
        RECT 2352.1200 1813.3600 2353.7200 1813.8400 ;
        RECT 2352.1200 1791.6000 2353.7200 1792.0800 ;
        RECT 2352.1200 1797.0400 2353.7200 1797.5200 ;
        RECT 2352.1200 1802.4800 2353.7200 1802.9600 ;
        RECT 2307.1200 1807.9200 2308.7200 1808.4000 ;
        RECT 2307.1200 1813.3600 2308.7200 1813.8400 ;
        RECT 2307.1200 1791.6000 2308.7200 1792.0800 ;
        RECT 2307.1200 1797.0400 2308.7200 1797.5200 ;
        RECT 2307.1200 1802.4800 2308.7200 1802.9600 ;
        RECT 2257.5600 1835.1200 2260.5600 1835.6000 ;
        RECT 2257.5600 1840.5600 2260.5600 1841.0400 ;
        RECT 2257.5600 1824.2400 2260.5600 1824.7200 ;
        RECT 2257.5600 1818.8000 2260.5600 1819.2800 ;
        RECT 2257.5600 1829.6800 2260.5600 1830.1600 ;
        RECT 2257.5600 1807.9200 2260.5600 1808.4000 ;
        RECT 2257.5600 1813.3600 2260.5600 1813.8400 ;
        RECT 2257.5600 1797.0400 2260.5600 1797.5200 ;
        RECT 2257.5600 1791.6000 2260.5600 1792.0800 ;
        RECT 2257.5600 1802.4800 2260.5600 1802.9600 ;
        RECT 2257.5600 1846.0000 2260.5600 1846.4800 ;
        RECT 2307.1200 1846.0000 2308.7200 1846.4800 ;
        RECT 2352.1200 1846.0000 2353.7200 1846.4800 ;
        RECT 2453.6600 1780.7200 2456.6600 1781.2000 ;
        RECT 2453.6600 1786.1600 2456.6600 1786.6400 ;
        RECT 2442.1200 1780.7200 2443.7200 1781.2000 ;
        RECT 2442.1200 1786.1600 2443.7200 1786.6400 ;
        RECT 2453.6600 1764.4000 2456.6600 1764.8800 ;
        RECT 2453.6600 1769.8400 2456.6600 1770.3200 ;
        RECT 2453.6600 1775.2800 2456.6600 1775.7600 ;
        RECT 2442.1200 1764.4000 2443.7200 1764.8800 ;
        RECT 2442.1200 1769.8400 2443.7200 1770.3200 ;
        RECT 2442.1200 1775.2800 2443.7200 1775.7600 ;
        RECT 2453.6600 1753.5200 2456.6600 1754.0000 ;
        RECT 2453.6600 1758.9600 2456.6600 1759.4400 ;
        RECT 2442.1200 1753.5200 2443.7200 1754.0000 ;
        RECT 2442.1200 1758.9600 2443.7200 1759.4400 ;
        RECT 2453.6600 1737.2000 2456.6600 1737.6800 ;
        RECT 2453.6600 1742.6400 2456.6600 1743.1200 ;
        RECT 2453.6600 1748.0800 2456.6600 1748.5600 ;
        RECT 2442.1200 1737.2000 2443.7200 1737.6800 ;
        RECT 2442.1200 1742.6400 2443.7200 1743.1200 ;
        RECT 2442.1200 1748.0800 2443.7200 1748.5600 ;
        RECT 2397.1200 1780.7200 2398.7200 1781.2000 ;
        RECT 2397.1200 1786.1600 2398.7200 1786.6400 ;
        RECT 2397.1200 1764.4000 2398.7200 1764.8800 ;
        RECT 2397.1200 1769.8400 2398.7200 1770.3200 ;
        RECT 2397.1200 1775.2800 2398.7200 1775.7600 ;
        RECT 2397.1200 1753.5200 2398.7200 1754.0000 ;
        RECT 2397.1200 1758.9600 2398.7200 1759.4400 ;
        RECT 2397.1200 1737.2000 2398.7200 1737.6800 ;
        RECT 2397.1200 1742.6400 2398.7200 1743.1200 ;
        RECT 2397.1200 1748.0800 2398.7200 1748.5600 ;
        RECT 2453.6600 1726.3200 2456.6600 1726.8000 ;
        RECT 2453.6600 1731.7600 2456.6600 1732.2400 ;
        RECT 2442.1200 1726.3200 2443.7200 1726.8000 ;
        RECT 2442.1200 1731.7600 2443.7200 1732.2400 ;
        RECT 2453.6600 1710.0000 2456.6600 1710.4800 ;
        RECT 2453.6600 1715.4400 2456.6600 1715.9200 ;
        RECT 2453.6600 1720.8800 2456.6600 1721.3600 ;
        RECT 2442.1200 1710.0000 2443.7200 1710.4800 ;
        RECT 2442.1200 1715.4400 2443.7200 1715.9200 ;
        RECT 2442.1200 1720.8800 2443.7200 1721.3600 ;
        RECT 2453.6600 1699.1200 2456.6600 1699.6000 ;
        RECT 2453.6600 1704.5600 2456.6600 1705.0400 ;
        RECT 2442.1200 1699.1200 2443.7200 1699.6000 ;
        RECT 2442.1200 1704.5600 2443.7200 1705.0400 ;
        RECT 2453.6600 1693.6800 2456.6600 1694.1600 ;
        RECT 2442.1200 1693.6800 2443.7200 1694.1600 ;
        RECT 2397.1200 1726.3200 2398.7200 1726.8000 ;
        RECT 2397.1200 1731.7600 2398.7200 1732.2400 ;
        RECT 2397.1200 1710.0000 2398.7200 1710.4800 ;
        RECT 2397.1200 1715.4400 2398.7200 1715.9200 ;
        RECT 2397.1200 1720.8800 2398.7200 1721.3600 ;
        RECT 2397.1200 1699.1200 2398.7200 1699.6000 ;
        RECT 2397.1200 1704.5600 2398.7200 1705.0400 ;
        RECT 2397.1200 1693.6800 2398.7200 1694.1600 ;
        RECT 2352.1200 1780.7200 2353.7200 1781.2000 ;
        RECT 2352.1200 1786.1600 2353.7200 1786.6400 ;
        RECT 2352.1200 1764.4000 2353.7200 1764.8800 ;
        RECT 2352.1200 1769.8400 2353.7200 1770.3200 ;
        RECT 2352.1200 1775.2800 2353.7200 1775.7600 ;
        RECT 2307.1200 1780.7200 2308.7200 1781.2000 ;
        RECT 2307.1200 1786.1600 2308.7200 1786.6400 ;
        RECT 2307.1200 1764.4000 2308.7200 1764.8800 ;
        RECT 2307.1200 1769.8400 2308.7200 1770.3200 ;
        RECT 2307.1200 1775.2800 2308.7200 1775.7600 ;
        RECT 2352.1200 1753.5200 2353.7200 1754.0000 ;
        RECT 2352.1200 1758.9600 2353.7200 1759.4400 ;
        RECT 2352.1200 1737.2000 2353.7200 1737.6800 ;
        RECT 2352.1200 1742.6400 2353.7200 1743.1200 ;
        RECT 2352.1200 1748.0800 2353.7200 1748.5600 ;
        RECT 2307.1200 1753.5200 2308.7200 1754.0000 ;
        RECT 2307.1200 1758.9600 2308.7200 1759.4400 ;
        RECT 2307.1200 1737.2000 2308.7200 1737.6800 ;
        RECT 2307.1200 1742.6400 2308.7200 1743.1200 ;
        RECT 2307.1200 1748.0800 2308.7200 1748.5600 ;
        RECT 2257.5600 1780.7200 2260.5600 1781.2000 ;
        RECT 2257.5600 1786.1600 2260.5600 1786.6400 ;
        RECT 2257.5600 1769.8400 2260.5600 1770.3200 ;
        RECT 2257.5600 1764.4000 2260.5600 1764.8800 ;
        RECT 2257.5600 1775.2800 2260.5600 1775.7600 ;
        RECT 2257.5600 1753.5200 2260.5600 1754.0000 ;
        RECT 2257.5600 1758.9600 2260.5600 1759.4400 ;
        RECT 2257.5600 1742.6400 2260.5600 1743.1200 ;
        RECT 2257.5600 1737.2000 2260.5600 1737.6800 ;
        RECT 2257.5600 1748.0800 2260.5600 1748.5600 ;
        RECT 2352.1200 1726.3200 2353.7200 1726.8000 ;
        RECT 2352.1200 1731.7600 2353.7200 1732.2400 ;
        RECT 2352.1200 1710.0000 2353.7200 1710.4800 ;
        RECT 2352.1200 1715.4400 2353.7200 1715.9200 ;
        RECT 2352.1200 1720.8800 2353.7200 1721.3600 ;
        RECT 2307.1200 1726.3200 2308.7200 1726.8000 ;
        RECT 2307.1200 1731.7600 2308.7200 1732.2400 ;
        RECT 2307.1200 1710.0000 2308.7200 1710.4800 ;
        RECT 2307.1200 1715.4400 2308.7200 1715.9200 ;
        RECT 2307.1200 1720.8800 2308.7200 1721.3600 ;
        RECT 2352.1200 1704.5600 2353.7200 1705.0400 ;
        RECT 2352.1200 1699.1200 2353.7200 1699.6000 ;
        RECT 2352.1200 1693.6800 2353.7200 1694.1600 ;
        RECT 2307.1200 1704.5600 2308.7200 1705.0400 ;
        RECT 2307.1200 1699.1200 2308.7200 1699.6000 ;
        RECT 2307.1200 1693.6800 2308.7200 1694.1600 ;
        RECT 2257.5600 1726.3200 2260.5600 1726.8000 ;
        RECT 2257.5600 1731.7600 2260.5600 1732.2400 ;
        RECT 2257.5600 1715.4400 2260.5600 1715.9200 ;
        RECT 2257.5600 1710.0000 2260.5600 1710.4800 ;
        RECT 2257.5600 1720.8800 2260.5600 1721.3600 ;
        RECT 2257.5600 1699.1200 2260.5600 1699.6000 ;
        RECT 2257.5600 1704.5600 2260.5600 1705.0400 ;
        RECT 2257.5600 1693.6800 2260.5600 1694.1600 ;
        RECT 2257.5600 1891.8700 2456.6600 1894.8700 ;
        RECT 2257.5600 1686.7700 2456.6600 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 1457.1300 2443.7200 1665.2300 ;
        RECT 2397.1200 1457.1300 2398.7200 1665.2300 ;
        RECT 2352.1200 1457.1300 2353.7200 1665.2300 ;
        RECT 2307.1200 1457.1300 2308.7200 1665.2300 ;
        RECT 2453.6600 1457.1300 2456.6600 1665.2300 ;
        RECT 2257.5600 1457.1300 2260.5600 1665.2300 ;
      LAYER met3 ;
        RECT 2453.6600 1659.8800 2456.6600 1660.3600 ;
        RECT 2442.1200 1659.8800 2443.7200 1660.3600 ;
        RECT 2453.6600 1649.0000 2456.6600 1649.4800 ;
        RECT 2453.6600 1654.4400 2456.6600 1654.9200 ;
        RECT 2442.1200 1649.0000 2443.7200 1649.4800 ;
        RECT 2442.1200 1654.4400 2443.7200 1654.9200 ;
        RECT 2453.6600 1632.6800 2456.6600 1633.1600 ;
        RECT 2453.6600 1638.1200 2456.6600 1638.6000 ;
        RECT 2442.1200 1632.6800 2443.7200 1633.1600 ;
        RECT 2442.1200 1638.1200 2443.7200 1638.6000 ;
        RECT 2453.6600 1621.8000 2456.6600 1622.2800 ;
        RECT 2453.6600 1627.2400 2456.6600 1627.7200 ;
        RECT 2442.1200 1621.8000 2443.7200 1622.2800 ;
        RECT 2442.1200 1627.2400 2443.7200 1627.7200 ;
        RECT 2453.6600 1643.5600 2456.6600 1644.0400 ;
        RECT 2442.1200 1643.5600 2443.7200 1644.0400 ;
        RECT 2397.1200 1649.0000 2398.7200 1649.4800 ;
        RECT 2397.1200 1654.4400 2398.7200 1654.9200 ;
        RECT 2397.1200 1659.8800 2398.7200 1660.3600 ;
        RECT 2397.1200 1632.6800 2398.7200 1633.1600 ;
        RECT 2397.1200 1638.1200 2398.7200 1638.6000 ;
        RECT 2397.1200 1627.2400 2398.7200 1627.7200 ;
        RECT 2397.1200 1621.8000 2398.7200 1622.2800 ;
        RECT 2397.1200 1643.5600 2398.7200 1644.0400 ;
        RECT 2453.6600 1605.4800 2456.6600 1605.9600 ;
        RECT 2453.6600 1610.9200 2456.6600 1611.4000 ;
        RECT 2442.1200 1605.4800 2443.7200 1605.9600 ;
        RECT 2442.1200 1610.9200 2443.7200 1611.4000 ;
        RECT 2453.6600 1589.1600 2456.6600 1589.6400 ;
        RECT 2453.6600 1594.6000 2456.6600 1595.0800 ;
        RECT 2453.6600 1600.0400 2456.6600 1600.5200 ;
        RECT 2442.1200 1589.1600 2443.7200 1589.6400 ;
        RECT 2442.1200 1594.6000 2443.7200 1595.0800 ;
        RECT 2442.1200 1600.0400 2443.7200 1600.5200 ;
        RECT 2453.6600 1578.2800 2456.6600 1578.7600 ;
        RECT 2453.6600 1583.7200 2456.6600 1584.2000 ;
        RECT 2442.1200 1578.2800 2443.7200 1578.7600 ;
        RECT 2442.1200 1583.7200 2443.7200 1584.2000 ;
        RECT 2453.6600 1561.9600 2456.6600 1562.4400 ;
        RECT 2453.6600 1567.4000 2456.6600 1567.8800 ;
        RECT 2453.6600 1572.8400 2456.6600 1573.3200 ;
        RECT 2442.1200 1561.9600 2443.7200 1562.4400 ;
        RECT 2442.1200 1567.4000 2443.7200 1567.8800 ;
        RECT 2442.1200 1572.8400 2443.7200 1573.3200 ;
        RECT 2397.1200 1605.4800 2398.7200 1605.9600 ;
        RECT 2397.1200 1610.9200 2398.7200 1611.4000 ;
        RECT 2397.1200 1589.1600 2398.7200 1589.6400 ;
        RECT 2397.1200 1594.6000 2398.7200 1595.0800 ;
        RECT 2397.1200 1600.0400 2398.7200 1600.5200 ;
        RECT 2397.1200 1578.2800 2398.7200 1578.7600 ;
        RECT 2397.1200 1583.7200 2398.7200 1584.2000 ;
        RECT 2397.1200 1561.9600 2398.7200 1562.4400 ;
        RECT 2397.1200 1567.4000 2398.7200 1567.8800 ;
        RECT 2397.1200 1572.8400 2398.7200 1573.3200 ;
        RECT 2453.6600 1616.3600 2456.6600 1616.8400 ;
        RECT 2397.1200 1616.3600 2398.7200 1616.8400 ;
        RECT 2442.1200 1616.3600 2443.7200 1616.8400 ;
        RECT 2352.1200 1649.0000 2353.7200 1649.4800 ;
        RECT 2352.1200 1654.4400 2353.7200 1654.9200 ;
        RECT 2352.1200 1659.8800 2353.7200 1660.3600 ;
        RECT 2307.1200 1649.0000 2308.7200 1649.4800 ;
        RECT 2307.1200 1654.4400 2308.7200 1654.9200 ;
        RECT 2307.1200 1659.8800 2308.7200 1660.3600 ;
        RECT 2352.1200 1632.6800 2353.7200 1633.1600 ;
        RECT 2352.1200 1638.1200 2353.7200 1638.6000 ;
        RECT 2352.1200 1621.8000 2353.7200 1622.2800 ;
        RECT 2352.1200 1627.2400 2353.7200 1627.7200 ;
        RECT 2307.1200 1632.6800 2308.7200 1633.1600 ;
        RECT 2307.1200 1638.1200 2308.7200 1638.6000 ;
        RECT 2307.1200 1621.8000 2308.7200 1622.2800 ;
        RECT 2307.1200 1627.2400 2308.7200 1627.7200 ;
        RECT 2307.1200 1643.5600 2308.7200 1644.0400 ;
        RECT 2352.1200 1643.5600 2353.7200 1644.0400 ;
        RECT 2257.5600 1659.8800 2260.5600 1660.3600 ;
        RECT 2257.5600 1654.4400 2260.5600 1654.9200 ;
        RECT 2257.5600 1649.0000 2260.5600 1649.4800 ;
        RECT 2257.5600 1638.1200 2260.5600 1638.6000 ;
        RECT 2257.5600 1632.6800 2260.5600 1633.1600 ;
        RECT 2257.5600 1627.2400 2260.5600 1627.7200 ;
        RECT 2257.5600 1621.8000 2260.5600 1622.2800 ;
        RECT 2257.5600 1643.5600 2260.5600 1644.0400 ;
        RECT 2352.1200 1605.4800 2353.7200 1605.9600 ;
        RECT 2352.1200 1610.9200 2353.7200 1611.4000 ;
        RECT 2352.1200 1589.1600 2353.7200 1589.6400 ;
        RECT 2352.1200 1594.6000 2353.7200 1595.0800 ;
        RECT 2352.1200 1600.0400 2353.7200 1600.5200 ;
        RECT 2307.1200 1605.4800 2308.7200 1605.9600 ;
        RECT 2307.1200 1610.9200 2308.7200 1611.4000 ;
        RECT 2307.1200 1589.1600 2308.7200 1589.6400 ;
        RECT 2307.1200 1594.6000 2308.7200 1595.0800 ;
        RECT 2307.1200 1600.0400 2308.7200 1600.5200 ;
        RECT 2352.1200 1578.2800 2353.7200 1578.7600 ;
        RECT 2352.1200 1583.7200 2353.7200 1584.2000 ;
        RECT 2352.1200 1561.9600 2353.7200 1562.4400 ;
        RECT 2352.1200 1567.4000 2353.7200 1567.8800 ;
        RECT 2352.1200 1572.8400 2353.7200 1573.3200 ;
        RECT 2307.1200 1578.2800 2308.7200 1578.7600 ;
        RECT 2307.1200 1583.7200 2308.7200 1584.2000 ;
        RECT 2307.1200 1561.9600 2308.7200 1562.4400 ;
        RECT 2307.1200 1567.4000 2308.7200 1567.8800 ;
        RECT 2307.1200 1572.8400 2308.7200 1573.3200 ;
        RECT 2257.5600 1605.4800 2260.5600 1605.9600 ;
        RECT 2257.5600 1610.9200 2260.5600 1611.4000 ;
        RECT 2257.5600 1594.6000 2260.5600 1595.0800 ;
        RECT 2257.5600 1589.1600 2260.5600 1589.6400 ;
        RECT 2257.5600 1600.0400 2260.5600 1600.5200 ;
        RECT 2257.5600 1578.2800 2260.5600 1578.7600 ;
        RECT 2257.5600 1583.7200 2260.5600 1584.2000 ;
        RECT 2257.5600 1567.4000 2260.5600 1567.8800 ;
        RECT 2257.5600 1561.9600 2260.5600 1562.4400 ;
        RECT 2257.5600 1572.8400 2260.5600 1573.3200 ;
        RECT 2257.5600 1616.3600 2260.5600 1616.8400 ;
        RECT 2307.1200 1616.3600 2308.7200 1616.8400 ;
        RECT 2352.1200 1616.3600 2353.7200 1616.8400 ;
        RECT 2453.6600 1551.0800 2456.6600 1551.5600 ;
        RECT 2453.6600 1556.5200 2456.6600 1557.0000 ;
        RECT 2442.1200 1551.0800 2443.7200 1551.5600 ;
        RECT 2442.1200 1556.5200 2443.7200 1557.0000 ;
        RECT 2453.6600 1534.7600 2456.6600 1535.2400 ;
        RECT 2453.6600 1540.2000 2456.6600 1540.6800 ;
        RECT 2453.6600 1545.6400 2456.6600 1546.1200 ;
        RECT 2442.1200 1534.7600 2443.7200 1535.2400 ;
        RECT 2442.1200 1540.2000 2443.7200 1540.6800 ;
        RECT 2442.1200 1545.6400 2443.7200 1546.1200 ;
        RECT 2453.6600 1523.8800 2456.6600 1524.3600 ;
        RECT 2453.6600 1529.3200 2456.6600 1529.8000 ;
        RECT 2442.1200 1523.8800 2443.7200 1524.3600 ;
        RECT 2442.1200 1529.3200 2443.7200 1529.8000 ;
        RECT 2453.6600 1507.5600 2456.6600 1508.0400 ;
        RECT 2453.6600 1513.0000 2456.6600 1513.4800 ;
        RECT 2453.6600 1518.4400 2456.6600 1518.9200 ;
        RECT 2442.1200 1507.5600 2443.7200 1508.0400 ;
        RECT 2442.1200 1513.0000 2443.7200 1513.4800 ;
        RECT 2442.1200 1518.4400 2443.7200 1518.9200 ;
        RECT 2397.1200 1551.0800 2398.7200 1551.5600 ;
        RECT 2397.1200 1556.5200 2398.7200 1557.0000 ;
        RECT 2397.1200 1534.7600 2398.7200 1535.2400 ;
        RECT 2397.1200 1540.2000 2398.7200 1540.6800 ;
        RECT 2397.1200 1545.6400 2398.7200 1546.1200 ;
        RECT 2397.1200 1523.8800 2398.7200 1524.3600 ;
        RECT 2397.1200 1529.3200 2398.7200 1529.8000 ;
        RECT 2397.1200 1507.5600 2398.7200 1508.0400 ;
        RECT 2397.1200 1513.0000 2398.7200 1513.4800 ;
        RECT 2397.1200 1518.4400 2398.7200 1518.9200 ;
        RECT 2453.6600 1496.6800 2456.6600 1497.1600 ;
        RECT 2453.6600 1502.1200 2456.6600 1502.6000 ;
        RECT 2442.1200 1496.6800 2443.7200 1497.1600 ;
        RECT 2442.1200 1502.1200 2443.7200 1502.6000 ;
        RECT 2453.6600 1480.3600 2456.6600 1480.8400 ;
        RECT 2453.6600 1485.8000 2456.6600 1486.2800 ;
        RECT 2453.6600 1491.2400 2456.6600 1491.7200 ;
        RECT 2442.1200 1480.3600 2443.7200 1480.8400 ;
        RECT 2442.1200 1485.8000 2443.7200 1486.2800 ;
        RECT 2442.1200 1491.2400 2443.7200 1491.7200 ;
        RECT 2453.6600 1469.4800 2456.6600 1469.9600 ;
        RECT 2453.6600 1474.9200 2456.6600 1475.4000 ;
        RECT 2442.1200 1469.4800 2443.7200 1469.9600 ;
        RECT 2442.1200 1474.9200 2443.7200 1475.4000 ;
        RECT 2453.6600 1464.0400 2456.6600 1464.5200 ;
        RECT 2442.1200 1464.0400 2443.7200 1464.5200 ;
        RECT 2397.1200 1496.6800 2398.7200 1497.1600 ;
        RECT 2397.1200 1502.1200 2398.7200 1502.6000 ;
        RECT 2397.1200 1480.3600 2398.7200 1480.8400 ;
        RECT 2397.1200 1485.8000 2398.7200 1486.2800 ;
        RECT 2397.1200 1491.2400 2398.7200 1491.7200 ;
        RECT 2397.1200 1469.4800 2398.7200 1469.9600 ;
        RECT 2397.1200 1474.9200 2398.7200 1475.4000 ;
        RECT 2397.1200 1464.0400 2398.7200 1464.5200 ;
        RECT 2352.1200 1551.0800 2353.7200 1551.5600 ;
        RECT 2352.1200 1556.5200 2353.7200 1557.0000 ;
        RECT 2352.1200 1534.7600 2353.7200 1535.2400 ;
        RECT 2352.1200 1540.2000 2353.7200 1540.6800 ;
        RECT 2352.1200 1545.6400 2353.7200 1546.1200 ;
        RECT 2307.1200 1551.0800 2308.7200 1551.5600 ;
        RECT 2307.1200 1556.5200 2308.7200 1557.0000 ;
        RECT 2307.1200 1534.7600 2308.7200 1535.2400 ;
        RECT 2307.1200 1540.2000 2308.7200 1540.6800 ;
        RECT 2307.1200 1545.6400 2308.7200 1546.1200 ;
        RECT 2352.1200 1523.8800 2353.7200 1524.3600 ;
        RECT 2352.1200 1529.3200 2353.7200 1529.8000 ;
        RECT 2352.1200 1507.5600 2353.7200 1508.0400 ;
        RECT 2352.1200 1513.0000 2353.7200 1513.4800 ;
        RECT 2352.1200 1518.4400 2353.7200 1518.9200 ;
        RECT 2307.1200 1523.8800 2308.7200 1524.3600 ;
        RECT 2307.1200 1529.3200 2308.7200 1529.8000 ;
        RECT 2307.1200 1507.5600 2308.7200 1508.0400 ;
        RECT 2307.1200 1513.0000 2308.7200 1513.4800 ;
        RECT 2307.1200 1518.4400 2308.7200 1518.9200 ;
        RECT 2257.5600 1551.0800 2260.5600 1551.5600 ;
        RECT 2257.5600 1556.5200 2260.5600 1557.0000 ;
        RECT 2257.5600 1540.2000 2260.5600 1540.6800 ;
        RECT 2257.5600 1534.7600 2260.5600 1535.2400 ;
        RECT 2257.5600 1545.6400 2260.5600 1546.1200 ;
        RECT 2257.5600 1523.8800 2260.5600 1524.3600 ;
        RECT 2257.5600 1529.3200 2260.5600 1529.8000 ;
        RECT 2257.5600 1513.0000 2260.5600 1513.4800 ;
        RECT 2257.5600 1507.5600 2260.5600 1508.0400 ;
        RECT 2257.5600 1518.4400 2260.5600 1518.9200 ;
        RECT 2352.1200 1496.6800 2353.7200 1497.1600 ;
        RECT 2352.1200 1502.1200 2353.7200 1502.6000 ;
        RECT 2352.1200 1480.3600 2353.7200 1480.8400 ;
        RECT 2352.1200 1485.8000 2353.7200 1486.2800 ;
        RECT 2352.1200 1491.2400 2353.7200 1491.7200 ;
        RECT 2307.1200 1496.6800 2308.7200 1497.1600 ;
        RECT 2307.1200 1502.1200 2308.7200 1502.6000 ;
        RECT 2307.1200 1480.3600 2308.7200 1480.8400 ;
        RECT 2307.1200 1485.8000 2308.7200 1486.2800 ;
        RECT 2307.1200 1491.2400 2308.7200 1491.7200 ;
        RECT 2352.1200 1474.9200 2353.7200 1475.4000 ;
        RECT 2352.1200 1469.4800 2353.7200 1469.9600 ;
        RECT 2352.1200 1464.0400 2353.7200 1464.5200 ;
        RECT 2307.1200 1474.9200 2308.7200 1475.4000 ;
        RECT 2307.1200 1469.4800 2308.7200 1469.9600 ;
        RECT 2307.1200 1464.0400 2308.7200 1464.5200 ;
        RECT 2257.5600 1496.6800 2260.5600 1497.1600 ;
        RECT 2257.5600 1502.1200 2260.5600 1502.6000 ;
        RECT 2257.5600 1485.8000 2260.5600 1486.2800 ;
        RECT 2257.5600 1480.3600 2260.5600 1480.8400 ;
        RECT 2257.5600 1491.2400 2260.5600 1491.7200 ;
        RECT 2257.5600 1469.4800 2260.5600 1469.9600 ;
        RECT 2257.5600 1474.9200 2260.5600 1475.4000 ;
        RECT 2257.5600 1464.0400 2260.5600 1464.5200 ;
        RECT 2257.5600 1662.2300 2456.6600 1665.2300 ;
        RECT 2257.5600 1457.1300 2456.6600 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 1227.4900 2443.7200 1435.5900 ;
        RECT 2397.1200 1227.4900 2398.7200 1435.5900 ;
        RECT 2352.1200 1227.4900 2353.7200 1435.5900 ;
        RECT 2307.1200 1227.4900 2308.7200 1435.5900 ;
        RECT 2453.6600 1227.4900 2456.6600 1435.5900 ;
        RECT 2257.5600 1227.4900 2260.5600 1435.5900 ;
      LAYER met3 ;
        RECT 2453.6600 1430.2400 2456.6600 1430.7200 ;
        RECT 2442.1200 1430.2400 2443.7200 1430.7200 ;
        RECT 2453.6600 1419.3600 2456.6600 1419.8400 ;
        RECT 2453.6600 1424.8000 2456.6600 1425.2800 ;
        RECT 2442.1200 1419.3600 2443.7200 1419.8400 ;
        RECT 2442.1200 1424.8000 2443.7200 1425.2800 ;
        RECT 2453.6600 1403.0400 2456.6600 1403.5200 ;
        RECT 2453.6600 1408.4800 2456.6600 1408.9600 ;
        RECT 2442.1200 1403.0400 2443.7200 1403.5200 ;
        RECT 2442.1200 1408.4800 2443.7200 1408.9600 ;
        RECT 2453.6600 1392.1600 2456.6600 1392.6400 ;
        RECT 2453.6600 1397.6000 2456.6600 1398.0800 ;
        RECT 2442.1200 1392.1600 2443.7200 1392.6400 ;
        RECT 2442.1200 1397.6000 2443.7200 1398.0800 ;
        RECT 2453.6600 1413.9200 2456.6600 1414.4000 ;
        RECT 2442.1200 1413.9200 2443.7200 1414.4000 ;
        RECT 2397.1200 1419.3600 2398.7200 1419.8400 ;
        RECT 2397.1200 1424.8000 2398.7200 1425.2800 ;
        RECT 2397.1200 1430.2400 2398.7200 1430.7200 ;
        RECT 2397.1200 1403.0400 2398.7200 1403.5200 ;
        RECT 2397.1200 1408.4800 2398.7200 1408.9600 ;
        RECT 2397.1200 1397.6000 2398.7200 1398.0800 ;
        RECT 2397.1200 1392.1600 2398.7200 1392.6400 ;
        RECT 2397.1200 1413.9200 2398.7200 1414.4000 ;
        RECT 2453.6600 1375.8400 2456.6600 1376.3200 ;
        RECT 2453.6600 1381.2800 2456.6600 1381.7600 ;
        RECT 2442.1200 1375.8400 2443.7200 1376.3200 ;
        RECT 2442.1200 1381.2800 2443.7200 1381.7600 ;
        RECT 2453.6600 1359.5200 2456.6600 1360.0000 ;
        RECT 2453.6600 1364.9600 2456.6600 1365.4400 ;
        RECT 2453.6600 1370.4000 2456.6600 1370.8800 ;
        RECT 2442.1200 1359.5200 2443.7200 1360.0000 ;
        RECT 2442.1200 1364.9600 2443.7200 1365.4400 ;
        RECT 2442.1200 1370.4000 2443.7200 1370.8800 ;
        RECT 2453.6600 1348.6400 2456.6600 1349.1200 ;
        RECT 2453.6600 1354.0800 2456.6600 1354.5600 ;
        RECT 2442.1200 1348.6400 2443.7200 1349.1200 ;
        RECT 2442.1200 1354.0800 2443.7200 1354.5600 ;
        RECT 2453.6600 1332.3200 2456.6600 1332.8000 ;
        RECT 2453.6600 1337.7600 2456.6600 1338.2400 ;
        RECT 2453.6600 1343.2000 2456.6600 1343.6800 ;
        RECT 2442.1200 1332.3200 2443.7200 1332.8000 ;
        RECT 2442.1200 1337.7600 2443.7200 1338.2400 ;
        RECT 2442.1200 1343.2000 2443.7200 1343.6800 ;
        RECT 2397.1200 1375.8400 2398.7200 1376.3200 ;
        RECT 2397.1200 1381.2800 2398.7200 1381.7600 ;
        RECT 2397.1200 1359.5200 2398.7200 1360.0000 ;
        RECT 2397.1200 1364.9600 2398.7200 1365.4400 ;
        RECT 2397.1200 1370.4000 2398.7200 1370.8800 ;
        RECT 2397.1200 1348.6400 2398.7200 1349.1200 ;
        RECT 2397.1200 1354.0800 2398.7200 1354.5600 ;
        RECT 2397.1200 1332.3200 2398.7200 1332.8000 ;
        RECT 2397.1200 1337.7600 2398.7200 1338.2400 ;
        RECT 2397.1200 1343.2000 2398.7200 1343.6800 ;
        RECT 2453.6600 1386.7200 2456.6600 1387.2000 ;
        RECT 2397.1200 1386.7200 2398.7200 1387.2000 ;
        RECT 2442.1200 1386.7200 2443.7200 1387.2000 ;
        RECT 2352.1200 1419.3600 2353.7200 1419.8400 ;
        RECT 2352.1200 1424.8000 2353.7200 1425.2800 ;
        RECT 2352.1200 1430.2400 2353.7200 1430.7200 ;
        RECT 2307.1200 1419.3600 2308.7200 1419.8400 ;
        RECT 2307.1200 1424.8000 2308.7200 1425.2800 ;
        RECT 2307.1200 1430.2400 2308.7200 1430.7200 ;
        RECT 2352.1200 1403.0400 2353.7200 1403.5200 ;
        RECT 2352.1200 1408.4800 2353.7200 1408.9600 ;
        RECT 2352.1200 1392.1600 2353.7200 1392.6400 ;
        RECT 2352.1200 1397.6000 2353.7200 1398.0800 ;
        RECT 2307.1200 1403.0400 2308.7200 1403.5200 ;
        RECT 2307.1200 1408.4800 2308.7200 1408.9600 ;
        RECT 2307.1200 1392.1600 2308.7200 1392.6400 ;
        RECT 2307.1200 1397.6000 2308.7200 1398.0800 ;
        RECT 2307.1200 1413.9200 2308.7200 1414.4000 ;
        RECT 2352.1200 1413.9200 2353.7200 1414.4000 ;
        RECT 2257.5600 1430.2400 2260.5600 1430.7200 ;
        RECT 2257.5600 1424.8000 2260.5600 1425.2800 ;
        RECT 2257.5600 1419.3600 2260.5600 1419.8400 ;
        RECT 2257.5600 1408.4800 2260.5600 1408.9600 ;
        RECT 2257.5600 1403.0400 2260.5600 1403.5200 ;
        RECT 2257.5600 1397.6000 2260.5600 1398.0800 ;
        RECT 2257.5600 1392.1600 2260.5600 1392.6400 ;
        RECT 2257.5600 1413.9200 2260.5600 1414.4000 ;
        RECT 2352.1200 1375.8400 2353.7200 1376.3200 ;
        RECT 2352.1200 1381.2800 2353.7200 1381.7600 ;
        RECT 2352.1200 1359.5200 2353.7200 1360.0000 ;
        RECT 2352.1200 1364.9600 2353.7200 1365.4400 ;
        RECT 2352.1200 1370.4000 2353.7200 1370.8800 ;
        RECT 2307.1200 1375.8400 2308.7200 1376.3200 ;
        RECT 2307.1200 1381.2800 2308.7200 1381.7600 ;
        RECT 2307.1200 1359.5200 2308.7200 1360.0000 ;
        RECT 2307.1200 1364.9600 2308.7200 1365.4400 ;
        RECT 2307.1200 1370.4000 2308.7200 1370.8800 ;
        RECT 2352.1200 1348.6400 2353.7200 1349.1200 ;
        RECT 2352.1200 1354.0800 2353.7200 1354.5600 ;
        RECT 2352.1200 1332.3200 2353.7200 1332.8000 ;
        RECT 2352.1200 1337.7600 2353.7200 1338.2400 ;
        RECT 2352.1200 1343.2000 2353.7200 1343.6800 ;
        RECT 2307.1200 1348.6400 2308.7200 1349.1200 ;
        RECT 2307.1200 1354.0800 2308.7200 1354.5600 ;
        RECT 2307.1200 1332.3200 2308.7200 1332.8000 ;
        RECT 2307.1200 1337.7600 2308.7200 1338.2400 ;
        RECT 2307.1200 1343.2000 2308.7200 1343.6800 ;
        RECT 2257.5600 1375.8400 2260.5600 1376.3200 ;
        RECT 2257.5600 1381.2800 2260.5600 1381.7600 ;
        RECT 2257.5600 1364.9600 2260.5600 1365.4400 ;
        RECT 2257.5600 1359.5200 2260.5600 1360.0000 ;
        RECT 2257.5600 1370.4000 2260.5600 1370.8800 ;
        RECT 2257.5600 1348.6400 2260.5600 1349.1200 ;
        RECT 2257.5600 1354.0800 2260.5600 1354.5600 ;
        RECT 2257.5600 1337.7600 2260.5600 1338.2400 ;
        RECT 2257.5600 1332.3200 2260.5600 1332.8000 ;
        RECT 2257.5600 1343.2000 2260.5600 1343.6800 ;
        RECT 2257.5600 1386.7200 2260.5600 1387.2000 ;
        RECT 2307.1200 1386.7200 2308.7200 1387.2000 ;
        RECT 2352.1200 1386.7200 2353.7200 1387.2000 ;
        RECT 2453.6600 1321.4400 2456.6600 1321.9200 ;
        RECT 2453.6600 1326.8800 2456.6600 1327.3600 ;
        RECT 2442.1200 1321.4400 2443.7200 1321.9200 ;
        RECT 2442.1200 1326.8800 2443.7200 1327.3600 ;
        RECT 2453.6600 1305.1200 2456.6600 1305.6000 ;
        RECT 2453.6600 1310.5600 2456.6600 1311.0400 ;
        RECT 2453.6600 1316.0000 2456.6600 1316.4800 ;
        RECT 2442.1200 1305.1200 2443.7200 1305.6000 ;
        RECT 2442.1200 1310.5600 2443.7200 1311.0400 ;
        RECT 2442.1200 1316.0000 2443.7200 1316.4800 ;
        RECT 2453.6600 1294.2400 2456.6600 1294.7200 ;
        RECT 2453.6600 1299.6800 2456.6600 1300.1600 ;
        RECT 2442.1200 1294.2400 2443.7200 1294.7200 ;
        RECT 2442.1200 1299.6800 2443.7200 1300.1600 ;
        RECT 2453.6600 1277.9200 2456.6600 1278.4000 ;
        RECT 2453.6600 1283.3600 2456.6600 1283.8400 ;
        RECT 2453.6600 1288.8000 2456.6600 1289.2800 ;
        RECT 2442.1200 1277.9200 2443.7200 1278.4000 ;
        RECT 2442.1200 1283.3600 2443.7200 1283.8400 ;
        RECT 2442.1200 1288.8000 2443.7200 1289.2800 ;
        RECT 2397.1200 1321.4400 2398.7200 1321.9200 ;
        RECT 2397.1200 1326.8800 2398.7200 1327.3600 ;
        RECT 2397.1200 1305.1200 2398.7200 1305.6000 ;
        RECT 2397.1200 1310.5600 2398.7200 1311.0400 ;
        RECT 2397.1200 1316.0000 2398.7200 1316.4800 ;
        RECT 2397.1200 1294.2400 2398.7200 1294.7200 ;
        RECT 2397.1200 1299.6800 2398.7200 1300.1600 ;
        RECT 2397.1200 1277.9200 2398.7200 1278.4000 ;
        RECT 2397.1200 1283.3600 2398.7200 1283.8400 ;
        RECT 2397.1200 1288.8000 2398.7200 1289.2800 ;
        RECT 2453.6600 1267.0400 2456.6600 1267.5200 ;
        RECT 2453.6600 1272.4800 2456.6600 1272.9600 ;
        RECT 2442.1200 1267.0400 2443.7200 1267.5200 ;
        RECT 2442.1200 1272.4800 2443.7200 1272.9600 ;
        RECT 2453.6600 1250.7200 2456.6600 1251.2000 ;
        RECT 2453.6600 1256.1600 2456.6600 1256.6400 ;
        RECT 2453.6600 1261.6000 2456.6600 1262.0800 ;
        RECT 2442.1200 1250.7200 2443.7200 1251.2000 ;
        RECT 2442.1200 1256.1600 2443.7200 1256.6400 ;
        RECT 2442.1200 1261.6000 2443.7200 1262.0800 ;
        RECT 2453.6600 1239.8400 2456.6600 1240.3200 ;
        RECT 2453.6600 1245.2800 2456.6600 1245.7600 ;
        RECT 2442.1200 1239.8400 2443.7200 1240.3200 ;
        RECT 2442.1200 1245.2800 2443.7200 1245.7600 ;
        RECT 2453.6600 1234.4000 2456.6600 1234.8800 ;
        RECT 2442.1200 1234.4000 2443.7200 1234.8800 ;
        RECT 2397.1200 1267.0400 2398.7200 1267.5200 ;
        RECT 2397.1200 1272.4800 2398.7200 1272.9600 ;
        RECT 2397.1200 1250.7200 2398.7200 1251.2000 ;
        RECT 2397.1200 1256.1600 2398.7200 1256.6400 ;
        RECT 2397.1200 1261.6000 2398.7200 1262.0800 ;
        RECT 2397.1200 1239.8400 2398.7200 1240.3200 ;
        RECT 2397.1200 1245.2800 2398.7200 1245.7600 ;
        RECT 2397.1200 1234.4000 2398.7200 1234.8800 ;
        RECT 2352.1200 1321.4400 2353.7200 1321.9200 ;
        RECT 2352.1200 1326.8800 2353.7200 1327.3600 ;
        RECT 2352.1200 1305.1200 2353.7200 1305.6000 ;
        RECT 2352.1200 1310.5600 2353.7200 1311.0400 ;
        RECT 2352.1200 1316.0000 2353.7200 1316.4800 ;
        RECT 2307.1200 1321.4400 2308.7200 1321.9200 ;
        RECT 2307.1200 1326.8800 2308.7200 1327.3600 ;
        RECT 2307.1200 1305.1200 2308.7200 1305.6000 ;
        RECT 2307.1200 1310.5600 2308.7200 1311.0400 ;
        RECT 2307.1200 1316.0000 2308.7200 1316.4800 ;
        RECT 2352.1200 1294.2400 2353.7200 1294.7200 ;
        RECT 2352.1200 1299.6800 2353.7200 1300.1600 ;
        RECT 2352.1200 1277.9200 2353.7200 1278.4000 ;
        RECT 2352.1200 1283.3600 2353.7200 1283.8400 ;
        RECT 2352.1200 1288.8000 2353.7200 1289.2800 ;
        RECT 2307.1200 1294.2400 2308.7200 1294.7200 ;
        RECT 2307.1200 1299.6800 2308.7200 1300.1600 ;
        RECT 2307.1200 1277.9200 2308.7200 1278.4000 ;
        RECT 2307.1200 1283.3600 2308.7200 1283.8400 ;
        RECT 2307.1200 1288.8000 2308.7200 1289.2800 ;
        RECT 2257.5600 1321.4400 2260.5600 1321.9200 ;
        RECT 2257.5600 1326.8800 2260.5600 1327.3600 ;
        RECT 2257.5600 1310.5600 2260.5600 1311.0400 ;
        RECT 2257.5600 1305.1200 2260.5600 1305.6000 ;
        RECT 2257.5600 1316.0000 2260.5600 1316.4800 ;
        RECT 2257.5600 1294.2400 2260.5600 1294.7200 ;
        RECT 2257.5600 1299.6800 2260.5600 1300.1600 ;
        RECT 2257.5600 1283.3600 2260.5600 1283.8400 ;
        RECT 2257.5600 1277.9200 2260.5600 1278.4000 ;
        RECT 2257.5600 1288.8000 2260.5600 1289.2800 ;
        RECT 2352.1200 1267.0400 2353.7200 1267.5200 ;
        RECT 2352.1200 1272.4800 2353.7200 1272.9600 ;
        RECT 2352.1200 1250.7200 2353.7200 1251.2000 ;
        RECT 2352.1200 1256.1600 2353.7200 1256.6400 ;
        RECT 2352.1200 1261.6000 2353.7200 1262.0800 ;
        RECT 2307.1200 1267.0400 2308.7200 1267.5200 ;
        RECT 2307.1200 1272.4800 2308.7200 1272.9600 ;
        RECT 2307.1200 1250.7200 2308.7200 1251.2000 ;
        RECT 2307.1200 1256.1600 2308.7200 1256.6400 ;
        RECT 2307.1200 1261.6000 2308.7200 1262.0800 ;
        RECT 2352.1200 1245.2800 2353.7200 1245.7600 ;
        RECT 2352.1200 1239.8400 2353.7200 1240.3200 ;
        RECT 2352.1200 1234.4000 2353.7200 1234.8800 ;
        RECT 2307.1200 1245.2800 2308.7200 1245.7600 ;
        RECT 2307.1200 1239.8400 2308.7200 1240.3200 ;
        RECT 2307.1200 1234.4000 2308.7200 1234.8800 ;
        RECT 2257.5600 1267.0400 2260.5600 1267.5200 ;
        RECT 2257.5600 1272.4800 2260.5600 1272.9600 ;
        RECT 2257.5600 1256.1600 2260.5600 1256.6400 ;
        RECT 2257.5600 1250.7200 2260.5600 1251.2000 ;
        RECT 2257.5600 1261.6000 2260.5600 1262.0800 ;
        RECT 2257.5600 1239.8400 2260.5600 1240.3200 ;
        RECT 2257.5600 1245.2800 2260.5600 1245.7600 ;
        RECT 2257.5600 1234.4000 2260.5600 1234.8800 ;
        RECT 2257.5600 1432.5900 2456.6600 1435.5900 ;
        RECT 2257.5600 1227.4900 2456.6600 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 997.8500 2443.7200 1205.9500 ;
        RECT 2397.1200 997.8500 2398.7200 1205.9500 ;
        RECT 2352.1200 997.8500 2353.7200 1205.9500 ;
        RECT 2307.1200 997.8500 2308.7200 1205.9500 ;
        RECT 2453.6600 997.8500 2456.6600 1205.9500 ;
        RECT 2257.5600 997.8500 2260.5600 1205.9500 ;
      LAYER met3 ;
        RECT 2453.6600 1200.6000 2456.6600 1201.0800 ;
        RECT 2442.1200 1200.6000 2443.7200 1201.0800 ;
        RECT 2453.6600 1189.7200 2456.6600 1190.2000 ;
        RECT 2453.6600 1195.1600 2456.6600 1195.6400 ;
        RECT 2442.1200 1189.7200 2443.7200 1190.2000 ;
        RECT 2442.1200 1195.1600 2443.7200 1195.6400 ;
        RECT 2453.6600 1173.4000 2456.6600 1173.8800 ;
        RECT 2453.6600 1178.8400 2456.6600 1179.3200 ;
        RECT 2442.1200 1173.4000 2443.7200 1173.8800 ;
        RECT 2442.1200 1178.8400 2443.7200 1179.3200 ;
        RECT 2453.6600 1162.5200 2456.6600 1163.0000 ;
        RECT 2453.6600 1167.9600 2456.6600 1168.4400 ;
        RECT 2442.1200 1162.5200 2443.7200 1163.0000 ;
        RECT 2442.1200 1167.9600 2443.7200 1168.4400 ;
        RECT 2453.6600 1184.2800 2456.6600 1184.7600 ;
        RECT 2442.1200 1184.2800 2443.7200 1184.7600 ;
        RECT 2397.1200 1189.7200 2398.7200 1190.2000 ;
        RECT 2397.1200 1195.1600 2398.7200 1195.6400 ;
        RECT 2397.1200 1200.6000 2398.7200 1201.0800 ;
        RECT 2397.1200 1173.4000 2398.7200 1173.8800 ;
        RECT 2397.1200 1178.8400 2398.7200 1179.3200 ;
        RECT 2397.1200 1167.9600 2398.7200 1168.4400 ;
        RECT 2397.1200 1162.5200 2398.7200 1163.0000 ;
        RECT 2397.1200 1184.2800 2398.7200 1184.7600 ;
        RECT 2453.6600 1146.2000 2456.6600 1146.6800 ;
        RECT 2453.6600 1151.6400 2456.6600 1152.1200 ;
        RECT 2442.1200 1146.2000 2443.7200 1146.6800 ;
        RECT 2442.1200 1151.6400 2443.7200 1152.1200 ;
        RECT 2453.6600 1129.8800 2456.6600 1130.3600 ;
        RECT 2453.6600 1135.3200 2456.6600 1135.8000 ;
        RECT 2453.6600 1140.7600 2456.6600 1141.2400 ;
        RECT 2442.1200 1129.8800 2443.7200 1130.3600 ;
        RECT 2442.1200 1135.3200 2443.7200 1135.8000 ;
        RECT 2442.1200 1140.7600 2443.7200 1141.2400 ;
        RECT 2453.6600 1119.0000 2456.6600 1119.4800 ;
        RECT 2453.6600 1124.4400 2456.6600 1124.9200 ;
        RECT 2442.1200 1119.0000 2443.7200 1119.4800 ;
        RECT 2442.1200 1124.4400 2443.7200 1124.9200 ;
        RECT 2453.6600 1102.6800 2456.6600 1103.1600 ;
        RECT 2453.6600 1108.1200 2456.6600 1108.6000 ;
        RECT 2453.6600 1113.5600 2456.6600 1114.0400 ;
        RECT 2442.1200 1102.6800 2443.7200 1103.1600 ;
        RECT 2442.1200 1108.1200 2443.7200 1108.6000 ;
        RECT 2442.1200 1113.5600 2443.7200 1114.0400 ;
        RECT 2397.1200 1146.2000 2398.7200 1146.6800 ;
        RECT 2397.1200 1151.6400 2398.7200 1152.1200 ;
        RECT 2397.1200 1129.8800 2398.7200 1130.3600 ;
        RECT 2397.1200 1135.3200 2398.7200 1135.8000 ;
        RECT 2397.1200 1140.7600 2398.7200 1141.2400 ;
        RECT 2397.1200 1119.0000 2398.7200 1119.4800 ;
        RECT 2397.1200 1124.4400 2398.7200 1124.9200 ;
        RECT 2397.1200 1102.6800 2398.7200 1103.1600 ;
        RECT 2397.1200 1108.1200 2398.7200 1108.6000 ;
        RECT 2397.1200 1113.5600 2398.7200 1114.0400 ;
        RECT 2453.6600 1157.0800 2456.6600 1157.5600 ;
        RECT 2397.1200 1157.0800 2398.7200 1157.5600 ;
        RECT 2442.1200 1157.0800 2443.7200 1157.5600 ;
        RECT 2352.1200 1189.7200 2353.7200 1190.2000 ;
        RECT 2352.1200 1195.1600 2353.7200 1195.6400 ;
        RECT 2352.1200 1200.6000 2353.7200 1201.0800 ;
        RECT 2307.1200 1189.7200 2308.7200 1190.2000 ;
        RECT 2307.1200 1195.1600 2308.7200 1195.6400 ;
        RECT 2307.1200 1200.6000 2308.7200 1201.0800 ;
        RECT 2352.1200 1173.4000 2353.7200 1173.8800 ;
        RECT 2352.1200 1178.8400 2353.7200 1179.3200 ;
        RECT 2352.1200 1162.5200 2353.7200 1163.0000 ;
        RECT 2352.1200 1167.9600 2353.7200 1168.4400 ;
        RECT 2307.1200 1173.4000 2308.7200 1173.8800 ;
        RECT 2307.1200 1178.8400 2308.7200 1179.3200 ;
        RECT 2307.1200 1162.5200 2308.7200 1163.0000 ;
        RECT 2307.1200 1167.9600 2308.7200 1168.4400 ;
        RECT 2307.1200 1184.2800 2308.7200 1184.7600 ;
        RECT 2352.1200 1184.2800 2353.7200 1184.7600 ;
        RECT 2257.5600 1200.6000 2260.5600 1201.0800 ;
        RECT 2257.5600 1195.1600 2260.5600 1195.6400 ;
        RECT 2257.5600 1189.7200 2260.5600 1190.2000 ;
        RECT 2257.5600 1178.8400 2260.5600 1179.3200 ;
        RECT 2257.5600 1173.4000 2260.5600 1173.8800 ;
        RECT 2257.5600 1167.9600 2260.5600 1168.4400 ;
        RECT 2257.5600 1162.5200 2260.5600 1163.0000 ;
        RECT 2257.5600 1184.2800 2260.5600 1184.7600 ;
        RECT 2352.1200 1146.2000 2353.7200 1146.6800 ;
        RECT 2352.1200 1151.6400 2353.7200 1152.1200 ;
        RECT 2352.1200 1129.8800 2353.7200 1130.3600 ;
        RECT 2352.1200 1135.3200 2353.7200 1135.8000 ;
        RECT 2352.1200 1140.7600 2353.7200 1141.2400 ;
        RECT 2307.1200 1146.2000 2308.7200 1146.6800 ;
        RECT 2307.1200 1151.6400 2308.7200 1152.1200 ;
        RECT 2307.1200 1129.8800 2308.7200 1130.3600 ;
        RECT 2307.1200 1135.3200 2308.7200 1135.8000 ;
        RECT 2307.1200 1140.7600 2308.7200 1141.2400 ;
        RECT 2352.1200 1119.0000 2353.7200 1119.4800 ;
        RECT 2352.1200 1124.4400 2353.7200 1124.9200 ;
        RECT 2352.1200 1102.6800 2353.7200 1103.1600 ;
        RECT 2352.1200 1108.1200 2353.7200 1108.6000 ;
        RECT 2352.1200 1113.5600 2353.7200 1114.0400 ;
        RECT 2307.1200 1119.0000 2308.7200 1119.4800 ;
        RECT 2307.1200 1124.4400 2308.7200 1124.9200 ;
        RECT 2307.1200 1102.6800 2308.7200 1103.1600 ;
        RECT 2307.1200 1108.1200 2308.7200 1108.6000 ;
        RECT 2307.1200 1113.5600 2308.7200 1114.0400 ;
        RECT 2257.5600 1146.2000 2260.5600 1146.6800 ;
        RECT 2257.5600 1151.6400 2260.5600 1152.1200 ;
        RECT 2257.5600 1135.3200 2260.5600 1135.8000 ;
        RECT 2257.5600 1129.8800 2260.5600 1130.3600 ;
        RECT 2257.5600 1140.7600 2260.5600 1141.2400 ;
        RECT 2257.5600 1119.0000 2260.5600 1119.4800 ;
        RECT 2257.5600 1124.4400 2260.5600 1124.9200 ;
        RECT 2257.5600 1108.1200 2260.5600 1108.6000 ;
        RECT 2257.5600 1102.6800 2260.5600 1103.1600 ;
        RECT 2257.5600 1113.5600 2260.5600 1114.0400 ;
        RECT 2257.5600 1157.0800 2260.5600 1157.5600 ;
        RECT 2307.1200 1157.0800 2308.7200 1157.5600 ;
        RECT 2352.1200 1157.0800 2353.7200 1157.5600 ;
        RECT 2453.6600 1091.8000 2456.6600 1092.2800 ;
        RECT 2453.6600 1097.2400 2456.6600 1097.7200 ;
        RECT 2442.1200 1091.8000 2443.7200 1092.2800 ;
        RECT 2442.1200 1097.2400 2443.7200 1097.7200 ;
        RECT 2453.6600 1075.4800 2456.6600 1075.9600 ;
        RECT 2453.6600 1080.9200 2456.6600 1081.4000 ;
        RECT 2453.6600 1086.3600 2456.6600 1086.8400 ;
        RECT 2442.1200 1075.4800 2443.7200 1075.9600 ;
        RECT 2442.1200 1080.9200 2443.7200 1081.4000 ;
        RECT 2442.1200 1086.3600 2443.7200 1086.8400 ;
        RECT 2453.6600 1064.6000 2456.6600 1065.0800 ;
        RECT 2453.6600 1070.0400 2456.6600 1070.5200 ;
        RECT 2442.1200 1064.6000 2443.7200 1065.0800 ;
        RECT 2442.1200 1070.0400 2443.7200 1070.5200 ;
        RECT 2453.6600 1048.2800 2456.6600 1048.7600 ;
        RECT 2453.6600 1053.7200 2456.6600 1054.2000 ;
        RECT 2453.6600 1059.1600 2456.6600 1059.6400 ;
        RECT 2442.1200 1048.2800 2443.7200 1048.7600 ;
        RECT 2442.1200 1053.7200 2443.7200 1054.2000 ;
        RECT 2442.1200 1059.1600 2443.7200 1059.6400 ;
        RECT 2397.1200 1091.8000 2398.7200 1092.2800 ;
        RECT 2397.1200 1097.2400 2398.7200 1097.7200 ;
        RECT 2397.1200 1075.4800 2398.7200 1075.9600 ;
        RECT 2397.1200 1080.9200 2398.7200 1081.4000 ;
        RECT 2397.1200 1086.3600 2398.7200 1086.8400 ;
        RECT 2397.1200 1064.6000 2398.7200 1065.0800 ;
        RECT 2397.1200 1070.0400 2398.7200 1070.5200 ;
        RECT 2397.1200 1048.2800 2398.7200 1048.7600 ;
        RECT 2397.1200 1053.7200 2398.7200 1054.2000 ;
        RECT 2397.1200 1059.1600 2398.7200 1059.6400 ;
        RECT 2453.6600 1037.4000 2456.6600 1037.8800 ;
        RECT 2453.6600 1042.8400 2456.6600 1043.3200 ;
        RECT 2442.1200 1037.4000 2443.7200 1037.8800 ;
        RECT 2442.1200 1042.8400 2443.7200 1043.3200 ;
        RECT 2453.6600 1021.0800 2456.6600 1021.5600 ;
        RECT 2453.6600 1026.5200 2456.6600 1027.0000 ;
        RECT 2453.6600 1031.9600 2456.6600 1032.4400 ;
        RECT 2442.1200 1021.0800 2443.7200 1021.5600 ;
        RECT 2442.1200 1026.5200 2443.7200 1027.0000 ;
        RECT 2442.1200 1031.9600 2443.7200 1032.4400 ;
        RECT 2453.6600 1010.2000 2456.6600 1010.6800 ;
        RECT 2453.6600 1015.6400 2456.6600 1016.1200 ;
        RECT 2442.1200 1010.2000 2443.7200 1010.6800 ;
        RECT 2442.1200 1015.6400 2443.7200 1016.1200 ;
        RECT 2453.6600 1004.7600 2456.6600 1005.2400 ;
        RECT 2442.1200 1004.7600 2443.7200 1005.2400 ;
        RECT 2397.1200 1037.4000 2398.7200 1037.8800 ;
        RECT 2397.1200 1042.8400 2398.7200 1043.3200 ;
        RECT 2397.1200 1021.0800 2398.7200 1021.5600 ;
        RECT 2397.1200 1026.5200 2398.7200 1027.0000 ;
        RECT 2397.1200 1031.9600 2398.7200 1032.4400 ;
        RECT 2397.1200 1010.2000 2398.7200 1010.6800 ;
        RECT 2397.1200 1015.6400 2398.7200 1016.1200 ;
        RECT 2397.1200 1004.7600 2398.7200 1005.2400 ;
        RECT 2352.1200 1091.8000 2353.7200 1092.2800 ;
        RECT 2352.1200 1097.2400 2353.7200 1097.7200 ;
        RECT 2352.1200 1075.4800 2353.7200 1075.9600 ;
        RECT 2352.1200 1080.9200 2353.7200 1081.4000 ;
        RECT 2352.1200 1086.3600 2353.7200 1086.8400 ;
        RECT 2307.1200 1091.8000 2308.7200 1092.2800 ;
        RECT 2307.1200 1097.2400 2308.7200 1097.7200 ;
        RECT 2307.1200 1075.4800 2308.7200 1075.9600 ;
        RECT 2307.1200 1080.9200 2308.7200 1081.4000 ;
        RECT 2307.1200 1086.3600 2308.7200 1086.8400 ;
        RECT 2352.1200 1064.6000 2353.7200 1065.0800 ;
        RECT 2352.1200 1070.0400 2353.7200 1070.5200 ;
        RECT 2352.1200 1048.2800 2353.7200 1048.7600 ;
        RECT 2352.1200 1053.7200 2353.7200 1054.2000 ;
        RECT 2352.1200 1059.1600 2353.7200 1059.6400 ;
        RECT 2307.1200 1064.6000 2308.7200 1065.0800 ;
        RECT 2307.1200 1070.0400 2308.7200 1070.5200 ;
        RECT 2307.1200 1048.2800 2308.7200 1048.7600 ;
        RECT 2307.1200 1053.7200 2308.7200 1054.2000 ;
        RECT 2307.1200 1059.1600 2308.7200 1059.6400 ;
        RECT 2257.5600 1091.8000 2260.5600 1092.2800 ;
        RECT 2257.5600 1097.2400 2260.5600 1097.7200 ;
        RECT 2257.5600 1080.9200 2260.5600 1081.4000 ;
        RECT 2257.5600 1075.4800 2260.5600 1075.9600 ;
        RECT 2257.5600 1086.3600 2260.5600 1086.8400 ;
        RECT 2257.5600 1064.6000 2260.5600 1065.0800 ;
        RECT 2257.5600 1070.0400 2260.5600 1070.5200 ;
        RECT 2257.5600 1053.7200 2260.5600 1054.2000 ;
        RECT 2257.5600 1048.2800 2260.5600 1048.7600 ;
        RECT 2257.5600 1059.1600 2260.5600 1059.6400 ;
        RECT 2352.1200 1037.4000 2353.7200 1037.8800 ;
        RECT 2352.1200 1042.8400 2353.7200 1043.3200 ;
        RECT 2352.1200 1021.0800 2353.7200 1021.5600 ;
        RECT 2352.1200 1026.5200 2353.7200 1027.0000 ;
        RECT 2352.1200 1031.9600 2353.7200 1032.4400 ;
        RECT 2307.1200 1037.4000 2308.7200 1037.8800 ;
        RECT 2307.1200 1042.8400 2308.7200 1043.3200 ;
        RECT 2307.1200 1021.0800 2308.7200 1021.5600 ;
        RECT 2307.1200 1026.5200 2308.7200 1027.0000 ;
        RECT 2307.1200 1031.9600 2308.7200 1032.4400 ;
        RECT 2352.1200 1015.6400 2353.7200 1016.1200 ;
        RECT 2352.1200 1010.2000 2353.7200 1010.6800 ;
        RECT 2352.1200 1004.7600 2353.7200 1005.2400 ;
        RECT 2307.1200 1015.6400 2308.7200 1016.1200 ;
        RECT 2307.1200 1010.2000 2308.7200 1010.6800 ;
        RECT 2307.1200 1004.7600 2308.7200 1005.2400 ;
        RECT 2257.5600 1037.4000 2260.5600 1037.8800 ;
        RECT 2257.5600 1042.8400 2260.5600 1043.3200 ;
        RECT 2257.5600 1026.5200 2260.5600 1027.0000 ;
        RECT 2257.5600 1021.0800 2260.5600 1021.5600 ;
        RECT 2257.5600 1031.9600 2260.5600 1032.4400 ;
        RECT 2257.5600 1010.2000 2260.5600 1010.6800 ;
        RECT 2257.5600 1015.6400 2260.5600 1016.1200 ;
        RECT 2257.5600 1004.7600 2260.5600 1005.2400 ;
        RECT 2257.5600 1202.9500 2456.6600 1205.9500 ;
        RECT 2257.5600 997.8500 2456.6600 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2442.1200 768.2100 2443.7200 976.3100 ;
        RECT 2397.1200 768.2100 2398.7200 976.3100 ;
        RECT 2352.1200 768.2100 2353.7200 976.3100 ;
        RECT 2307.1200 768.2100 2308.7200 976.3100 ;
        RECT 2453.6600 768.2100 2456.6600 976.3100 ;
        RECT 2257.5600 768.2100 2260.5600 976.3100 ;
      LAYER met3 ;
        RECT 2453.6600 970.9600 2456.6600 971.4400 ;
        RECT 2442.1200 970.9600 2443.7200 971.4400 ;
        RECT 2453.6600 960.0800 2456.6600 960.5600 ;
        RECT 2453.6600 965.5200 2456.6600 966.0000 ;
        RECT 2442.1200 960.0800 2443.7200 960.5600 ;
        RECT 2442.1200 965.5200 2443.7200 966.0000 ;
        RECT 2453.6600 943.7600 2456.6600 944.2400 ;
        RECT 2453.6600 949.2000 2456.6600 949.6800 ;
        RECT 2442.1200 943.7600 2443.7200 944.2400 ;
        RECT 2442.1200 949.2000 2443.7200 949.6800 ;
        RECT 2453.6600 932.8800 2456.6600 933.3600 ;
        RECT 2453.6600 938.3200 2456.6600 938.8000 ;
        RECT 2442.1200 932.8800 2443.7200 933.3600 ;
        RECT 2442.1200 938.3200 2443.7200 938.8000 ;
        RECT 2453.6600 954.6400 2456.6600 955.1200 ;
        RECT 2442.1200 954.6400 2443.7200 955.1200 ;
        RECT 2397.1200 960.0800 2398.7200 960.5600 ;
        RECT 2397.1200 965.5200 2398.7200 966.0000 ;
        RECT 2397.1200 970.9600 2398.7200 971.4400 ;
        RECT 2397.1200 943.7600 2398.7200 944.2400 ;
        RECT 2397.1200 949.2000 2398.7200 949.6800 ;
        RECT 2397.1200 938.3200 2398.7200 938.8000 ;
        RECT 2397.1200 932.8800 2398.7200 933.3600 ;
        RECT 2397.1200 954.6400 2398.7200 955.1200 ;
        RECT 2453.6600 916.5600 2456.6600 917.0400 ;
        RECT 2453.6600 922.0000 2456.6600 922.4800 ;
        RECT 2442.1200 916.5600 2443.7200 917.0400 ;
        RECT 2442.1200 922.0000 2443.7200 922.4800 ;
        RECT 2453.6600 900.2400 2456.6600 900.7200 ;
        RECT 2453.6600 905.6800 2456.6600 906.1600 ;
        RECT 2453.6600 911.1200 2456.6600 911.6000 ;
        RECT 2442.1200 900.2400 2443.7200 900.7200 ;
        RECT 2442.1200 905.6800 2443.7200 906.1600 ;
        RECT 2442.1200 911.1200 2443.7200 911.6000 ;
        RECT 2453.6600 889.3600 2456.6600 889.8400 ;
        RECT 2453.6600 894.8000 2456.6600 895.2800 ;
        RECT 2442.1200 889.3600 2443.7200 889.8400 ;
        RECT 2442.1200 894.8000 2443.7200 895.2800 ;
        RECT 2453.6600 873.0400 2456.6600 873.5200 ;
        RECT 2453.6600 878.4800 2456.6600 878.9600 ;
        RECT 2453.6600 883.9200 2456.6600 884.4000 ;
        RECT 2442.1200 873.0400 2443.7200 873.5200 ;
        RECT 2442.1200 878.4800 2443.7200 878.9600 ;
        RECT 2442.1200 883.9200 2443.7200 884.4000 ;
        RECT 2397.1200 916.5600 2398.7200 917.0400 ;
        RECT 2397.1200 922.0000 2398.7200 922.4800 ;
        RECT 2397.1200 900.2400 2398.7200 900.7200 ;
        RECT 2397.1200 905.6800 2398.7200 906.1600 ;
        RECT 2397.1200 911.1200 2398.7200 911.6000 ;
        RECT 2397.1200 889.3600 2398.7200 889.8400 ;
        RECT 2397.1200 894.8000 2398.7200 895.2800 ;
        RECT 2397.1200 873.0400 2398.7200 873.5200 ;
        RECT 2397.1200 878.4800 2398.7200 878.9600 ;
        RECT 2397.1200 883.9200 2398.7200 884.4000 ;
        RECT 2453.6600 927.4400 2456.6600 927.9200 ;
        RECT 2397.1200 927.4400 2398.7200 927.9200 ;
        RECT 2442.1200 927.4400 2443.7200 927.9200 ;
        RECT 2352.1200 960.0800 2353.7200 960.5600 ;
        RECT 2352.1200 965.5200 2353.7200 966.0000 ;
        RECT 2352.1200 970.9600 2353.7200 971.4400 ;
        RECT 2307.1200 960.0800 2308.7200 960.5600 ;
        RECT 2307.1200 965.5200 2308.7200 966.0000 ;
        RECT 2307.1200 970.9600 2308.7200 971.4400 ;
        RECT 2352.1200 943.7600 2353.7200 944.2400 ;
        RECT 2352.1200 949.2000 2353.7200 949.6800 ;
        RECT 2352.1200 932.8800 2353.7200 933.3600 ;
        RECT 2352.1200 938.3200 2353.7200 938.8000 ;
        RECT 2307.1200 943.7600 2308.7200 944.2400 ;
        RECT 2307.1200 949.2000 2308.7200 949.6800 ;
        RECT 2307.1200 932.8800 2308.7200 933.3600 ;
        RECT 2307.1200 938.3200 2308.7200 938.8000 ;
        RECT 2307.1200 954.6400 2308.7200 955.1200 ;
        RECT 2352.1200 954.6400 2353.7200 955.1200 ;
        RECT 2257.5600 970.9600 2260.5600 971.4400 ;
        RECT 2257.5600 965.5200 2260.5600 966.0000 ;
        RECT 2257.5600 960.0800 2260.5600 960.5600 ;
        RECT 2257.5600 949.2000 2260.5600 949.6800 ;
        RECT 2257.5600 943.7600 2260.5600 944.2400 ;
        RECT 2257.5600 938.3200 2260.5600 938.8000 ;
        RECT 2257.5600 932.8800 2260.5600 933.3600 ;
        RECT 2257.5600 954.6400 2260.5600 955.1200 ;
        RECT 2352.1200 916.5600 2353.7200 917.0400 ;
        RECT 2352.1200 922.0000 2353.7200 922.4800 ;
        RECT 2352.1200 900.2400 2353.7200 900.7200 ;
        RECT 2352.1200 905.6800 2353.7200 906.1600 ;
        RECT 2352.1200 911.1200 2353.7200 911.6000 ;
        RECT 2307.1200 916.5600 2308.7200 917.0400 ;
        RECT 2307.1200 922.0000 2308.7200 922.4800 ;
        RECT 2307.1200 900.2400 2308.7200 900.7200 ;
        RECT 2307.1200 905.6800 2308.7200 906.1600 ;
        RECT 2307.1200 911.1200 2308.7200 911.6000 ;
        RECT 2352.1200 889.3600 2353.7200 889.8400 ;
        RECT 2352.1200 894.8000 2353.7200 895.2800 ;
        RECT 2352.1200 873.0400 2353.7200 873.5200 ;
        RECT 2352.1200 878.4800 2353.7200 878.9600 ;
        RECT 2352.1200 883.9200 2353.7200 884.4000 ;
        RECT 2307.1200 889.3600 2308.7200 889.8400 ;
        RECT 2307.1200 894.8000 2308.7200 895.2800 ;
        RECT 2307.1200 873.0400 2308.7200 873.5200 ;
        RECT 2307.1200 878.4800 2308.7200 878.9600 ;
        RECT 2307.1200 883.9200 2308.7200 884.4000 ;
        RECT 2257.5600 916.5600 2260.5600 917.0400 ;
        RECT 2257.5600 922.0000 2260.5600 922.4800 ;
        RECT 2257.5600 905.6800 2260.5600 906.1600 ;
        RECT 2257.5600 900.2400 2260.5600 900.7200 ;
        RECT 2257.5600 911.1200 2260.5600 911.6000 ;
        RECT 2257.5600 889.3600 2260.5600 889.8400 ;
        RECT 2257.5600 894.8000 2260.5600 895.2800 ;
        RECT 2257.5600 878.4800 2260.5600 878.9600 ;
        RECT 2257.5600 873.0400 2260.5600 873.5200 ;
        RECT 2257.5600 883.9200 2260.5600 884.4000 ;
        RECT 2257.5600 927.4400 2260.5600 927.9200 ;
        RECT 2307.1200 927.4400 2308.7200 927.9200 ;
        RECT 2352.1200 927.4400 2353.7200 927.9200 ;
        RECT 2453.6600 862.1600 2456.6600 862.6400 ;
        RECT 2453.6600 867.6000 2456.6600 868.0800 ;
        RECT 2442.1200 862.1600 2443.7200 862.6400 ;
        RECT 2442.1200 867.6000 2443.7200 868.0800 ;
        RECT 2453.6600 845.8400 2456.6600 846.3200 ;
        RECT 2453.6600 851.2800 2456.6600 851.7600 ;
        RECT 2453.6600 856.7200 2456.6600 857.2000 ;
        RECT 2442.1200 845.8400 2443.7200 846.3200 ;
        RECT 2442.1200 851.2800 2443.7200 851.7600 ;
        RECT 2442.1200 856.7200 2443.7200 857.2000 ;
        RECT 2453.6600 834.9600 2456.6600 835.4400 ;
        RECT 2453.6600 840.4000 2456.6600 840.8800 ;
        RECT 2442.1200 834.9600 2443.7200 835.4400 ;
        RECT 2442.1200 840.4000 2443.7200 840.8800 ;
        RECT 2453.6600 818.6400 2456.6600 819.1200 ;
        RECT 2453.6600 824.0800 2456.6600 824.5600 ;
        RECT 2453.6600 829.5200 2456.6600 830.0000 ;
        RECT 2442.1200 818.6400 2443.7200 819.1200 ;
        RECT 2442.1200 824.0800 2443.7200 824.5600 ;
        RECT 2442.1200 829.5200 2443.7200 830.0000 ;
        RECT 2397.1200 862.1600 2398.7200 862.6400 ;
        RECT 2397.1200 867.6000 2398.7200 868.0800 ;
        RECT 2397.1200 845.8400 2398.7200 846.3200 ;
        RECT 2397.1200 851.2800 2398.7200 851.7600 ;
        RECT 2397.1200 856.7200 2398.7200 857.2000 ;
        RECT 2397.1200 834.9600 2398.7200 835.4400 ;
        RECT 2397.1200 840.4000 2398.7200 840.8800 ;
        RECT 2397.1200 818.6400 2398.7200 819.1200 ;
        RECT 2397.1200 824.0800 2398.7200 824.5600 ;
        RECT 2397.1200 829.5200 2398.7200 830.0000 ;
        RECT 2453.6600 807.7600 2456.6600 808.2400 ;
        RECT 2453.6600 813.2000 2456.6600 813.6800 ;
        RECT 2442.1200 807.7600 2443.7200 808.2400 ;
        RECT 2442.1200 813.2000 2443.7200 813.6800 ;
        RECT 2453.6600 791.4400 2456.6600 791.9200 ;
        RECT 2453.6600 796.8800 2456.6600 797.3600 ;
        RECT 2453.6600 802.3200 2456.6600 802.8000 ;
        RECT 2442.1200 791.4400 2443.7200 791.9200 ;
        RECT 2442.1200 796.8800 2443.7200 797.3600 ;
        RECT 2442.1200 802.3200 2443.7200 802.8000 ;
        RECT 2453.6600 780.5600 2456.6600 781.0400 ;
        RECT 2453.6600 786.0000 2456.6600 786.4800 ;
        RECT 2442.1200 780.5600 2443.7200 781.0400 ;
        RECT 2442.1200 786.0000 2443.7200 786.4800 ;
        RECT 2453.6600 775.1200 2456.6600 775.6000 ;
        RECT 2442.1200 775.1200 2443.7200 775.6000 ;
        RECT 2397.1200 807.7600 2398.7200 808.2400 ;
        RECT 2397.1200 813.2000 2398.7200 813.6800 ;
        RECT 2397.1200 791.4400 2398.7200 791.9200 ;
        RECT 2397.1200 796.8800 2398.7200 797.3600 ;
        RECT 2397.1200 802.3200 2398.7200 802.8000 ;
        RECT 2397.1200 780.5600 2398.7200 781.0400 ;
        RECT 2397.1200 786.0000 2398.7200 786.4800 ;
        RECT 2397.1200 775.1200 2398.7200 775.6000 ;
        RECT 2352.1200 862.1600 2353.7200 862.6400 ;
        RECT 2352.1200 867.6000 2353.7200 868.0800 ;
        RECT 2352.1200 845.8400 2353.7200 846.3200 ;
        RECT 2352.1200 851.2800 2353.7200 851.7600 ;
        RECT 2352.1200 856.7200 2353.7200 857.2000 ;
        RECT 2307.1200 862.1600 2308.7200 862.6400 ;
        RECT 2307.1200 867.6000 2308.7200 868.0800 ;
        RECT 2307.1200 845.8400 2308.7200 846.3200 ;
        RECT 2307.1200 851.2800 2308.7200 851.7600 ;
        RECT 2307.1200 856.7200 2308.7200 857.2000 ;
        RECT 2352.1200 834.9600 2353.7200 835.4400 ;
        RECT 2352.1200 840.4000 2353.7200 840.8800 ;
        RECT 2352.1200 818.6400 2353.7200 819.1200 ;
        RECT 2352.1200 824.0800 2353.7200 824.5600 ;
        RECT 2352.1200 829.5200 2353.7200 830.0000 ;
        RECT 2307.1200 834.9600 2308.7200 835.4400 ;
        RECT 2307.1200 840.4000 2308.7200 840.8800 ;
        RECT 2307.1200 818.6400 2308.7200 819.1200 ;
        RECT 2307.1200 824.0800 2308.7200 824.5600 ;
        RECT 2307.1200 829.5200 2308.7200 830.0000 ;
        RECT 2257.5600 862.1600 2260.5600 862.6400 ;
        RECT 2257.5600 867.6000 2260.5600 868.0800 ;
        RECT 2257.5600 851.2800 2260.5600 851.7600 ;
        RECT 2257.5600 845.8400 2260.5600 846.3200 ;
        RECT 2257.5600 856.7200 2260.5600 857.2000 ;
        RECT 2257.5600 834.9600 2260.5600 835.4400 ;
        RECT 2257.5600 840.4000 2260.5600 840.8800 ;
        RECT 2257.5600 824.0800 2260.5600 824.5600 ;
        RECT 2257.5600 818.6400 2260.5600 819.1200 ;
        RECT 2257.5600 829.5200 2260.5600 830.0000 ;
        RECT 2352.1200 807.7600 2353.7200 808.2400 ;
        RECT 2352.1200 813.2000 2353.7200 813.6800 ;
        RECT 2352.1200 791.4400 2353.7200 791.9200 ;
        RECT 2352.1200 796.8800 2353.7200 797.3600 ;
        RECT 2352.1200 802.3200 2353.7200 802.8000 ;
        RECT 2307.1200 807.7600 2308.7200 808.2400 ;
        RECT 2307.1200 813.2000 2308.7200 813.6800 ;
        RECT 2307.1200 791.4400 2308.7200 791.9200 ;
        RECT 2307.1200 796.8800 2308.7200 797.3600 ;
        RECT 2307.1200 802.3200 2308.7200 802.8000 ;
        RECT 2352.1200 786.0000 2353.7200 786.4800 ;
        RECT 2352.1200 780.5600 2353.7200 781.0400 ;
        RECT 2352.1200 775.1200 2353.7200 775.6000 ;
        RECT 2307.1200 786.0000 2308.7200 786.4800 ;
        RECT 2307.1200 780.5600 2308.7200 781.0400 ;
        RECT 2307.1200 775.1200 2308.7200 775.6000 ;
        RECT 2257.5600 807.7600 2260.5600 808.2400 ;
        RECT 2257.5600 813.2000 2260.5600 813.6800 ;
        RECT 2257.5600 796.8800 2260.5600 797.3600 ;
        RECT 2257.5600 791.4400 2260.5600 791.9200 ;
        RECT 2257.5600 802.3200 2260.5600 802.8000 ;
        RECT 2257.5600 780.5600 2260.5600 781.0400 ;
        RECT 2257.5600 786.0000 2260.5600 786.4800 ;
        RECT 2257.5600 775.1200 2260.5600 775.6000 ;
        RECT 2257.5600 973.3100 2456.6600 976.3100 ;
        RECT 2257.5600 768.2100 2456.6600 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 2477.7800 2833.6100 2479.7800 2854.5400 ;
        RECT 2674.8800 2833.6100 2676.8800 2854.5400 ;
      LAYER met3 ;
        RECT 2674.8800 2850.0400 2676.8800 2850.5200 ;
        RECT 2477.7800 2850.0400 2479.7800 2850.5200 ;
        RECT 2674.8800 2839.1600 2676.8800 2839.6400 ;
        RECT 2477.7800 2839.1600 2479.7800 2839.6400 ;
        RECT 2674.8800 2844.6000 2676.8800 2845.0800 ;
        RECT 2477.7800 2844.6000 2479.7800 2845.0800 ;
        RECT 2477.7800 2852.5400 2676.8800 2854.5400 ;
        RECT 2477.7800 2833.6100 2676.8800 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 538.5700 2663.9400 746.6700 ;
        RECT 2617.3400 538.5700 2618.9400 746.6700 ;
        RECT 2572.3400 538.5700 2573.9400 746.6700 ;
        RECT 2527.3400 538.5700 2528.9400 746.6700 ;
        RECT 2673.8800 538.5700 2676.8800 746.6700 ;
        RECT 2477.7800 538.5700 2480.7800 746.6700 ;
      LAYER met3 ;
        RECT 2673.8800 741.3200 2676.8800 741.8000 ;
        RECT 2662.3400 741.3200 2663.9400 741.8000 ;
        RECT 2673.8800 730.4400 2676.8800 730.9200 ;
        RECT 2673.8800 735.8800 2676.8800 736.3600 ;
        RECT 2662.3400 730.4400 2663.9400 730.9200 ;
        RECT 2662.3400 735.8800 2663.9400 736.3600 ;
        RECT 2673.8800 714.1200 2676.8800 714.6000 ;
        RECT 2673.8800 719.5600 2676.8800 720.0400 ;
        RECT 2662.3400 714.1200 2663.9400 714.6000 ;
        RECT 2662.3400 719.5600 2663.9400 720.0400 ;
        RECT 2673.8800 703.2400 2676.8800 703.7200 ;
        RECT 2673.8800 708.6800 2676.8800 709.1600 ;
        RECT 2662.3400 703.2400 2663.9400 703.7200 ;
        RECT 2662.3400 708.6800 2663.9400 709.1600 ;
        RECT 2673.8800 725.0000 2676.8800 725.4800 ;
        RECT 2662.3400 725.0000 2663.9400 725.4800 ;
        RECT 2617.3400 730.4400 2618.9400 730.9200 ;
        RECT 2617.3400 735.8800 2618.9400 736.3600 ;
        RECT 2617.3400 741.3200 2618.9400 741.8000 ;
        RECT 2617.3400 714.1200 2618.9400 714.6000 ;
        RECT 2617.3400 719.5600 2618.9400 720.0400 ;
        RECT 2617.3400 708.6800 2618.9400 709.1600 ;
        RECT 2617.3400 703.2400 2618.9400 703.7200 ;
        RECT 2617.3400 725.0000 2618.9400 725.4800 ;
        RECT 2673.8800 686.9200 2676.8800 687.4000 ;
        RECT 2673.8800 692.3600 2676.8800 692.8400 ;
        RECT 2662.3400 686.9200 2663.9400 687.4000 ;
        RECT 2662.3400 692.3600 2663.9400 692.8400 ;
        RECT 2673.8800 670.6000 2676.8800 671.0800 ;
        RECT 2673.8800 676.0400 2676.8800 676.5200 ;
        RECT 2673.8800 681.4800 2676.8800 681.9600 ;
        RECT 2662.3400 670.6000 2663.9400 671.0800 ;
        RECT 2662.3400 676.0400 2663.9400 676.5200 ;
        RECT 2662.3400 681.4800 2663.9400 681.9600 ;
        RECT 2673.8800 659.7200 2676.8800 660.2000 ;
        RECT 2673.8800 665.1600 2676.8800 665.6400 ;
        RECT 2662.3400 659.7200 2663.9400 660.2000 ;
        RECT 2662.3400 665.1600 2663.9400 665.6400 ;
        RECT 2673.8800 643.4000 2676.8800 643.8800 ;
        RECT 2673.8800 648.8400 2676.8800 649.3200 ;
        RECT 2673.8800 654.2800 2676.8800 654.7600 ;
        RECT 2662.3400 643.4000 2663.9400 643.8800 ;
        RECT 2662.3400 648.8400 2663.9400 649.3200 ;
        RECT 2662.3400 654.2800 2663.9400 654.7600 ;
        RECT 2617.3400 686.9200 2618.9400 687.4000 ;
        RECT 2617.3400 692.3600 2618.9400 692.8400 ;
        RECT 2617.3400 670.6000 2618.9400 671.0800 ;
        RECT 2617.3400 676.0400 2618.9400 676.5200 ;
        RECT 2617.3400 681.4800 2618.9400 681.9600 ;
        RECT 2617.3400 659.7200 2618.9400 660.2000 ;
        RECT 2617.3400 665.1600 2618.9400 665.6400 ;
        RECT 2617.3400 643.4000 2618.9400 643.8800 ;
        RECT 2617.3400 648.8400 2618.9400 649.3200 ;
        RECT 2617.3400 654.2800 2618.9400 654.7600 ;
        RECT 2673.8800 697.8000 2676.8800 698.2800 ;
        RECT 2617.3400 697.8000 2618.9400 698.2800 ;
        RECT 2662.3400 697.8000 2663.9400 698.2800 ;
        RECT 2572.3400 730.4400 2573.9400 730.9200 ;
        RECT 2572.3400 735.8800 2573.9400 736.3600 ;
        RECT 2572.3400 741.3200 2573.9400 741.8000 ;
        RECT 2527.3400 730.4400 2528.9400 730.9200 ;
        RECT 2527.3400 735.8800 2528.9400 736.3600 ;
        RECT 2527.3400 741.3200 2528.9400 741.8000 ;
        RECT 2572.3400 714.1200 2573.9400 714.6000 ;
        RECT 2572.3400 719.5600 2573.9400 720.0400 ;
        RECT 2572.3400 703.2400 2573.9400 703.7200 ;
        RECT 2572.3400 708.6800 2573.9400 709.1600 ;
        RECT 2527.3400 714.1200 2528.9400 714.6000 ;
        RECT 2527.3400 719.5600 2528.9400 720.0400 ;
        RECT 2527.3400 703.2400 2528.9400 703.7200 ;
        RECT 2527.3400 708.6800 2528.9400 709.1600 ;
        RECT 2527.3400 725.0000 2528.9400 725.4800 ;
        RECT 2572.3400 725.0000 2573.9400 725.4800 ;
        RECT 2477.7800 741.3200 2480.7800 741.8000 ;
        RECT 2477.7800 735.8800 2480.7800 736.3600 ;
        RECT 2477.7800 730.4400 2480.7800 730.9200 ;
        RECT 2477.7800 719.5600 2480.7800 720.0400 ;
        RECT 2477.7800 714.1200 2480.7800 714.6000 ;
        RECT 2477.7800 708.6800 2480.7800 709.1600 ;
        RECT 2477.7800 703.2400 2480.7800 703.7200 ;
        RECT 2477.7800 725.0000 2480.7800 725.4800 ;
        RECT 2572.3400 686.9200 2573.9400 687.4000 ;
        RECT 2572.3400 692.3600 2573.9400 692.8400 ;
        RECT 2572.3400 670.6000 2573.9400 671.0800 ;
        RECT 2572.3400 676.0400 2573.9400 676.5200 ;
        RECT 2572.3400 681.4800 2573.9400 681.9600 ;
        RECT 2527.3400 686.9200 2528.9400 687.4000 ;
        RECT 2527.3400 692.3600 2528.9400 692.8400 ;
        RECT 2527.3400 670.6000 2528.9400 671.0800 ;
        RECT 2527.3400 676.0400 2528.9400 676.5200 ;
        RECT 2527.3400 681.4800 2528.9400 681.9600 ;
        RECT 2572.3400 659.7200 2573.9400 660.2000 ;
        RECT 2572.3400 665.1600 2573.9400 665.6400 ;
        RECT 2572.3400 643.4000 2573.9400 643.8800 ;
        RECT 2572.3400 648.8400 2573.9400 649.3200 ;
        RECT 2572.3400 654.2800 2573.9400 654.7600 ;
        RECT 2527.3400 659.7200 2528.9400 660.2000 ;
        RECT 2527.3400 665.1600 2528.9400 665.6400 ;
        RECT 2527.3400 643.4000 2528.9400 643.8800 ;
        RECT 2527.3400 648.8400 2528.9400 649.3200 ;
        RECT 2527.3400 654.2800 2528.9400 654.7600 ;
        RECT 2477.7800 686.9200 2480.7800 687.4000 ;
        RECT 2477.7800 692.3600 2480.7800 692.8400 ;
        RECT 2477.7800 676.0400 2480.7800 676.5200 ;
        RECT 2477.7800 670.6000 2480.7800 671.0800 ;
        RECT 2477.7800 681.4800 2480.7800 681.9600 ;
        RECT 2477.7800 659.7200 2480.7800 660.2000 ;
        RECT 2477.7800 665.1600 2480.7800 665.6400 ;
        RECT 2477.7800 648.8400 2480.7800 649.3200 ;
        RECT 2477.7800 643.4000 2480.7800 643.8800 ;
        RECT 2477.7800 654.2800 2480.7800 654.7600 ;
        RECT 2477.7800 697.8000 2480.7800 698.2800 ;
        RECT 2527.3400 697.8000 2528.9400 698.2800 ;
        RECT 2572.3400 697.8000 2573.9400 698.2800 ;
        RECT 2673.8800 632.5200 2676.8800 633.0000 ;
        RECT 2673.8800 637.9600 2676.8800 638.4400 ;
        RECT 2662.3400 632.5200 2663.9400 633.0000 ;
        RECT 2662.3400 637.9600 2663.9400 638.4400 ;
        RECT 2673.8800 616.2000 2676.8800 616.6800 ;
        RECT 2673.8800 621.6400 2676.8800 622.1200 ;
        RECT 2673.8800 627.0800 2676.8800 627.5600 ;
        RECT 2662.3400 616.2000 2663.9400 616.6800 ;
        RECT 2662.3400 621.6400 2663.9400 622.1200 ;
        RECT 2662.3400 627.0800 2663.9400 627.5600 ;
        RECT 2673.8800 605.3200 2676.8800 605.8000 ;
        RECT 2673.8800 610.7600 2676.8800 611.2400 ;
        RECT 2662.3400 605.3200 2663.9400 605.8000 ;
        RECT 2662.3400 610.7600 2663.9400 611.2400 ;
        RECT 2673.8800 589.0000 2676.8800 589.4800 ;
        RECT 2673.8800 594.4400 2676.8800 594.9200 ;
        RECT 2673.8800 599.8800 2676.8800 600.3600 ;
        RECT 2662.3400 589.0000 2663.9400 589.4800 ;
        RECT 2662.3400 594.4400 2663.9400 594.9200 ;
        RECT 2662.3400 599.8800 2663.9400 600.3600 ;
        RECT 2617.3400 632.5200 2618.9400 633.0000 ;
        RECT 2617.3400 637.9600 2618.9400 638.4400 ;
        RECT 2617.3400 616.2000 2618.9400 616.6800 ;
        RECT 2617.3400 621.6400 2618.9400 622.1200 ;
        RECT 2617.3400 627.0800 2618.9400 627.5600 ;
        RECT 2617.3400 605.3200 2618.9400 605.8000 ;
        RECT 2617.3400 610.7600 2618.9400 611.2400 ;
        RECT 2617.3400 589.0000 2618.9400 589.4800 ;
        RECT 2617.3400 594.4400 2618.9400 594.9200 ;
        RECT 2617.3400 599.8800 2618.9400 600.3600 ;
        RECT 2673.8800 578.1200 2676.8800 578.6000 ;
        RECT 2673.8800 583.5600 2676.8800 584.0400 ;
        RECT 2662.3400 578.1200 2663.9400 578.6000 ;
        RECT 2662.3400 583.5600 2663.9400 584.0400 ;
        RECT 2673.8800 561.8000 2676.8800 562.2800 ;
        RECT 2673.8800 567.2400 2676.8800 567.7200 ;
        RECT 2673.8800 572.6800 2676.8800 573.1600 ;
        RECT 2662.3400 561.8000 2663.9400 562.2800 ;
        RECT 2662.3400 567.2400 2663.9400 567.7200 ;
        RECT 2662.3400 572.6800 2663.9400 573.1600 ;
        RECT 2673.8800 550.9200 2676.8800 551.4000 ;
        RECT 2673.8800 556.3600 2676.8800 556.8400 ;
        RECT 2662.3400 550.9200 2663.9400 551.4000 ;
        RECT 2662.3400 556.3600 2663.9400 556.8400 ;
        RECT 2673.8800 545.4800 2676.8800 545.9600 ;
        RECT 2662.3400 545.4800 2663.9400 545.9600 ;
        RECT 2617.3400 578.1200 2618.9400 578.6000 ;
        RECT 2617.3400 583.5600 2618.9400 584.0400 ;
        RECT 2617.3400 561.8000 2618.9400 562.2800 ;
        RECT 2617.3400 567.2400 2618.9400 567.7200 ;
        RECT 2617.3400 572.6800 2618.9400 573.1600 ;
        RECT 2617.3400 550.9200 2618.9400 551.4000 ;
        RECT 2617.3400 556.3600 2618.9400 556.8400 ;
        RECT 2617.3400 545.4800 2618.9400 545.9600 ;
        RECT 2572.3400 632.5200 2573.9400 633.0000 ;
        RECT 2572.3400 637.9600 2573.9400 638.4400 ;
        RECT 2572.3400 616.2000 2573.9400 616.6800 ;
        RECT 2572.3400 621.6400 2573.9400 622.1200 ;
        RECT 2572.3400 627.0800 2573.9400 627.5600 ;
        RECT 2527.3400 632.5200 2528.9400 633.0000 ;
        RECT 2527.3400 637.9600 2528.9400 638.4400 ;
        RECT 2527.3400 616.2000 2528.9400 616.6800 ;
        RECT 2527.3400 621.6400 2528.9400 622.1200 ;
        RECT 2527.3400 627.0800 2528.9400 627.5600 ;
        RECT 2572.3400 605.3200 2573.9400 605.8000 ;
        RECT 2572.3400 610.7600 2573.9400 611.2400 ;
        RECT 2572.3400 589.0000 2573.9400 589.4800 ;
        RECT 2572.3400 594.4400 2573.9400 594.9200 ;
        RECT 2572.3400 599.8800 2573.9400 600.3600 ;
        RECT 2527.3400 605.3200 2528.9400 605.8000 ;
        RECT 2527.3400 610.7600 2528.9400 611.2400 ;
        RECT 2527.3400 589.0000 2528.9400 589.4800 ;
        RECT 2527.3400 594.4400 2528.9400 594.9200 ;
        RECT 2527.3400 599.8800 2528.9400 600.3600 ;
        RECT 2477.7800 632.5200 2480.7800 633.0000 ;
        RECT 2477.7800 637.9600 2480.7800 638.4400 ;
        RECT 2477.7800 621.6400 2480.7800 622.1200 ;
        RECT 2477.7800 616.2000 2480.7800 616.6800 ;
        RECT 2477.7800 627.0800 2480.7800 627.5600 ;
        RECT 2477.7800 605.3200 2480.7800 605.8000 ;
        RECT 2477.7800 610.7600 2480.7800 611.2400 ;
        RECT 2477.7800 594.4400 2480.7800 594.9200 ;
        RECT 2477.7800 589.0000 2480.7800 589.4800 ;
        RECT 2477.7800 599.8800 2480.7800 600.3600 ;
        RECT 2572.3400 578.1200 2573.9400 578.6000 ;
        RECT 2572.3400 583.5600 2573.9400 584.0400 ;
        RECT 2572.3400 561.8000 2573.9400 562.2800 ;
        RECT 2572.3400 567.2400 2573.9400 567.7200 ;
        RECT 2572.3400 572.6800 2573.9400 573.1600 ;
        RECT 2527.3400 578.1200 2528.9400 578.6000 ;
        RECT 2527.3400 583.5600 2528.9400 584.0400 ;
        RECT 2527.3400 561.8000 2528.9400 562.2800 ;
        RECT 2527.3400 567.2400 2528.9400 567.7200 ;
        RECT 2527.3400 572.6800 2528.9400 573.1600 ;
        RECT 2572.3400 556.3600 2573.9400 556.8400 ;
        RECT 2572.3400 550.9200 2573.9400 551.4000 ;
        RECT 2572.3400 545.4800 2573.9400 545.9600 ;
        RECT 2527.3400 556.3600 2528.9400 556.8400 ;
        RECT 2527.3400 550.9200 2528.9400 551.4000 ;
        RECT 2527.3400 545.4800 2528.9400 545.9600 ;
        RECT 2477.7800 578.1200 2480.7800 578.6000 ;
        RECT 2477.7800 583.5600 2480.7800 584.0400 ;
        RECT 2477.7800 567.2400 2480.7800 567.7200 ;
        RECT 2477.7800 561.8000 2480.7800 562.2800 ;
        RECT 2477.7800 572.6800 2480.7800 573.1600 ;
        RECT 2477.7800 550.9200 2480.7800 551.4000 ;
        RECT 2477.7800 556.3600 2480.7800 556.8400 ;
        RECT 2477.7800 545.4800 2480.7800 545.9600 ;
        RECT 2477.7800 743.6700 2676.8800 746.6700 ;
        RECT 2477.7800 538.5700 2676.8800 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 308.9300 2663.9400 517.0300 ;
        RECT 2617.3400 308.9300 2618.9400 517.0300 ;
        RECT 2572.3400 308.9300 2573.9400 517.0300 ;
        RECT 2527.3400 308.9300 2528.9400 517.0300 ;
        RECT 2673.8800 308.9300 2676.8800 517.0300 ;
        RECT 2477.7800 308.9300 2480.7800 517.0300 ;
      LAYER met3 ;
        RECT 2673.8800 511.6800 2676.8800 512.1600 ;
        RECT 2662.3400 511.6800 2663.9400 512.1600 ;
        RECT 2673.8800 500.8000 2676.8800 501.2800 ;
        RECT 2673.8800 506.2400 2676.8800 506.7200 ;
        RECT 2662.3400 500.8000 2663.9400 501.2800 ;
        RECT 2662.3400 506.2400 2663.9400 506.7200 ;
        RECT 2673.8800 484.4800 2676.8800 484.9600 ;
        RECT 2673.8800 489.9200 2676.8800 490.4000 ;
        RECT 2662.3400 484.4800 2663.9400 484.9600 ;
        RECT 2662.3400 489.9200 2663.9400 490.4000 ;
        RECT 2673.8800 473.6000 2676.8800 474.0800 ;
        RECT 2673.8800 479.0400 2676.8800 479.5200 ;
        RECT 2662.3400 473.6000 2663.9400 474.0800 ;
        RECT 2662.3400 479.0400 2663.9400 479.5200 ;
        RECT 2673.8800 495.3600 2676.8800 495.8400 ;
        RECT 2662.3400 495.3600 2663.9400 495.8400 ;
        RECT 2617.3400 500.8000 2618.9400 501.2800 ;
        RECT 2617.3400 506.2400 2618.9400 506.7200 ;
        RECT 2617.3400 511.6800 2618.9400 512.1600 ;
        RECT 2617.3400 484.4800 2618.9400 484.9600 ;
        RECT 2617.3400 489.9200 2618.9400 490.4000 ;
        RECT 2617.3400 479.0400 2618.9400 479.5200 ;
        RECT 2617.3400 473.6000 2618.9400 474.0800 ;
        RECT 2617.3400 495.3600 2618.9400 495.8400 ;
        RECT 2673.8800 457.2800 2676.8800 457.7600 ;
        RECT 2673.8800 462.7200 2676.8800 463.2000 ;
        RECT 2662.3400 457.2800 2663.9400 457.7600 ;
        RECT 2662.3400 462.7200 2663.9400 463.2000 ;
        RECT 2673.8800 440.9600 2676.8800 441.4400 ;
        RECT 2673.8800 446.4000 2676.8800 446.8800 ;
        RECT 2673.8800 451.8400 2676.8800 452.3200 ;
        RECT 2662.3400 440.9600 2663.9400 441.4400 ;
        RECT 2662.3400 446.4000 2663.9400 446.8800 ;
        RECT 2662.3400 451.8400 2663.9400 452.3200 ;
        RECT 2673.8800 430.0800 2676.8800 430.5600 ;
        RECT 2673.8800 435.5200 2676.8800 436.0000 ;
        RECT 2662.3400 430.0800 2663.9400 430.5600 ;
        RECT 2662.3400 435.5200 2663.9400 436.0000 ;
        RECT 2673.8800 413.7600 2676.8800 414.2400 ;
        RECT 2673.8800 419.2000 2676.8800 419.6800 ;
        RECT 2673.8800 424.6400 2676.8800 425.1200 ;
        RECT 2662.3400 413.7600 2663.9400 414.2400 ;
        RECT 2662.3400 419.2000 2663.9400 419.6800 ;
        RECT 2662.3400 424.6400 2663.9400 425.1200 ;
        RECT 2617.3400 457.2800 2618.9400 457.7600 ;
        RECT 2617.3400 462.7200 2618.9400 463.2000 ;
        RECT 2617.3400 440.9600 2618.9400 441.4400 ;
        RECT 2617.3400 446.4000 2618.9400 446.8800 ;
        RECT 2617.3400 451.8400 2618.9400 452.3200 ;
        RECT 2617.3400 430.0800 2618.9400 430.5600 ;
        RECT 2617.3400 435.5200 2618.9400 436.0000 ;
        RECT 2617.3400 413.7600 2618.9400 414.2400 ;
        RECT 2617.3400 419.2000 2618.9400 419.6800 ;
        RECT 2617.3400 424.6400 2618.9400 425.1200 ;
        RECT 2673.8800 468.1600 2676.8800 468.6400 ;
        RECT 2617.3400 468.1600 2618.9400 468.6400 ;
        RECT 2662.3400 468.1600 2663.9400 468.6400 ;
        RECT 2572.3400 500.8000 2573.9400 501.2800 ;
        RECT 2572.3400 506.2400 2573.9400 506.7200 ;
        RECT 2572.3400 511.6800 2573.9400 512.1600 ;
        RECT 2527.3400 500.8000 2528.9400 501.2800 ;
        RECT 2527.3400 506.2400 2528.9400 506.7200 ;
        RECT 2527.3400 511.6800 2528.9400 512.1600 ;
        RECT 2572.3400 484.4800 2573.9400 484.9600 ;
        RECT 2572.3400 489.9200 2573.9400 490.4000 ;
        RECT 2572.3400 473.6000 2573.9400 474.0800 ;
        RECT 2572.3400 479.0400 2573.9400 479.5200 ;
        RECT 2527.3400 484.4800 2528.9400 484.9600 ;
        RECT 2527.3400 489.9200 2528.9400 490.4000 ;
        RECT 2527.3400 473.6000 2528.9400 474.0800 ;
        RECT 2527.3400 479.0400 2528.9400 479.5200 ;
        RECT 2527.3400 495.3600 2528.9400 495.8400 ;
        RECT 2572.3400 495.3600 2573.9400 495.8400 ;
        RECT 2477.7800 511.6800 2480.7800 512.1600 ;
        RECT 2477.7800 506.2400 2480.7800 506.7200 ;
        RECT 2477.7800 500.8000 2480.7800 501.2800 ;
        RECT 2477.7800 489.9200 2480.7800 490.4000 ;
        RECT 2477.7800 484.4800 2480.7800 484.9600 ;
        RECT 2477.7800 479.0400 2480.7800 479.5200 ;
        RECT 2477.7800 473.6000 2480.7800 474.0800 ;
        RECT 2477.7800 495.3600 2480.7800 495.8400 ;
        RECT 2572.3400 457.2800 2573.9400 457.7600 ;
        RECT 2572.3400 462.7200 2573.9400 463.2000 ;
        RECT 2572.3400 440.9600 2573.9400 441.4400 ;
        RECT 2572.3400 446.4000 2573.9400 446.8800 ;
        RECT 2572.3400 451.8400 2573.9400 452.3200 ;
        RECT 2527.3400 457.2800 2528.9400 457.7600 ;
        RECT 2527.3400 462.7200 2528.9400 463.2000 ;
        RECT 2527.3400 440.9600 2528.9400 441.4400 ;
        RECT 2527.3400 446.4000 2528.9400 446.8800 ;
        RECT 2527.3400 451.8400 2528.9400 452.3200 ;
        RECT 2572.3400 430.0800 2573.9400 430.5600 ;
        RECT 2572.3400 435.5200 2573.9400 436.0000 ;
        RECT 2572.3400 413.7600 2573.9400 414.2400 ;
        RECT 2572.3400 419.2000 2573.9400 419.6800 ;
        RECT 2572.3400 424.6400 2573.9400 425.1200 ;
        RECT 2527.3400 430.0800 2528.9400 430.5600 ;
        RECT 2527.3400 435.5200 2528.9400 436.0000 ;
        RECT 2527.3400 413.7600 2528.9400 414.2400 ;
        RECT 2527.3400 419.2000 2528.9400 419.6800 ;
        RECT 2527.3400 424.6400 2528.9400 425.1200 ;
        RECT 2477.7800 457.2800 2480.7800 457.7600 ;
        RECT 2477.7800 462.7200 2480.7800 463.2000 ;
        RECT 2477.7800 446.4000 2480.7800 446.8800 ;
        RECT 2477.7800 440.9600 2480.7800 441.4400 ;
        RECT 2477.7800 451.8400 2480.7800 452.3200 ;
        RECT 2477.7800 430.0800 2480.7800 430.5600 ;
        RECT 2477.7800 435.5200 2480.7800 436.0000 ;
        RECT 2477.7800 419.2000 2480.7800 419.6800 ;
        RECT 2477.7800 413.7600 2480.7800 414.2400 ;
        RECT 2477.7800 424.6400 2480.7800 425.1200 ;
        RECT 2477.7800 468.1600 2480.7800 468.6400 ;
        RECT 2527.3400 468.1600 2528.9400 468.6400 ;
        RECT 2572.3400 468.1600 2573.9400 468.6400 ;
        RECT 2673.8800 402.8800 2676.8800 403.3600 ;
        RECT 2673.8800 408.3200 2676.8800 408.8000 ;
        RECT 2662.3400 402.8800 2663.9400 403.3600 ;
        RECT 2662.3400 408.3200 2663.9400 408.8000 ;
        RECT 2673.8800 386.5600 2676.8800 387.0400 ;
        RECT 2673.8800 392.0000 2676.8800 392.4800 ;
        RECT 2673.8800 397.4400 2676.8800 397.9200 ;
        RECT 2662.3400 386.5600 2663.9400 387.0400 ;
        RECT 2662.3400 392.0000 2663.9400 392.4800 ;
        RECT 2662.3400 397.4400 2663.9400 397.9200 ;
        RECT 2673.8800 375.6800 2676.8800 376.1600 ;
        RECT 2673.8800 381.1200 2676.8800 381.6000 ;
        RECT 2662.3400 375.6800 2663.9400 376.1600 ;
        RECT 2662.3400 381.1200 2663.9400 381.6000 ;
        RECT 2673.8800 359.3600 2676.8800 359.8400 ;
        RECT 2673.8800 364.8000 2676.8800 365.2800 ;
        RECT 2673.8800 370.2400 2676.8800 370.7200 ;
        RECT 2662.3400 359.3600 2663.9400 359.8400 ;
        RECT 2662.3400 364.8000 2663.9400 365.2800 ;
        RECT 2662.3400 370.2400 2663.9400 370.7200 ;
        RECT 2617.3400 402.8800 2618.9400 403.3600 ;
        RECT 2617.3400 408.3200 2618.9400 408.8000 ;
        RECT 2617.3400 386.5600 2618.9400 387.0400 ;
        RECT 2617.3400 392.0000 2618.9400 392.4800 ;
        RECT 2617.3400 397.4400 2618.9400 397.9200 ;
        RECT 2617.3400 375.6800 2618.9400 376.1600 ;
        RECT 2617.3400 381.1200 2618.9400 381.6000 ;
        RECT 2617.3400 359.3600 2618.9400 359.8400 ;
        RECT 2617.3400 364.8000 2618.9400 365.2800 ;
        RECT 2617.3400 370.2400 2618.9400 370.7200 ;
        RECT 2673.8800 348.4800 2676.8800 348.9600 ;
        RECT 2673.8800 353.9200 2676.8800 354.4000 ;
        RECT 2662.3400 348.4800 2663.9400 348.9600 ;
        RECT 2662.3400 353.9200 2663.9400 354.4000 ;
        RECT 2673.8800 332.1600 2676.8800 332.6400 ;
        RECT 2673.8800 337.6000 2676.8800 338.0800 ;
        RECT 2673.8800 343.0400 2676.8800 343.5200 ;
        RECT 2662.3400 332.1600 2663.9400 332.6400 ;
        RECT 2662.3400 337.6000 2663.9400 338.0800 ;
        RECT 2662.3400 343.0400 2663.9400 343.5200 ;
        RECT 2673.8800 321.2800 2676.8800 321.7600 ;
        RECT 2673.8800 326.7200 2676.8800 327.2000 ;
        RECT 2662.3400 321.2800 2663.9400 321.7600 ;
        RECT 2662.3400 326.7200 2663.9400 327.2000 ;
        RECT 2673.8800 315.8400 2676.8800 316.3200 ;
        RECT 2662.3400 315.8400 2663.9400 316.3200 ;
        RECT 2617.3400 348.4800 2618.9400 348.9600 ;
        RECT 2617.3400 353.9200 2618.9400 354.4000 ;
        RECT 2617.3400 332.1600 2618.9400 332.6400 ;
        RECT 2617.3400 337.6000 2618.9400 338.0800 ;
        RECT 2617.3400 343.0400 2618.9400 343.5200 ;
        RECT 2617.3400 321.2800 2618.9400 321.7600 ;
        RECT 2617.3400 326.7200 2618.9400 327.2000 ;
        RECT 2617.3400 315.8400 2618.9400 316.3200 ;
        RECT 2572.3400 402.8800 2573.9400 403.3600 ;
        RECT 2572.3400 408.3200 2573.9400 408.8000 ;
        RECT 2572.3400 386.5600 2573.9400 387.0400 ;
        RECT 2572.3400 392.0000 2573.9400 392.4800 ;
        RECT 2572.3400 397.4400 2573.9400 397.9200 ;
        RECT 2527.3400 402.8800 2528.9400 403.3600 ;
        RECT 2527.3400 408.3200 2528.9400 408.8000 ;
        RECT 2527.3400 386.5600 2528.9400 387.0400 ;
        RECT 2527.3400 392.0000 2528.9400 392.4800 ;
        RECT 2527.3400 397.4400 2528.9400 397.9200 ;
        RECT 2572.3400 375.6800 2573.9400 376.1600 ;
        RECT 2572.3400 381.1200 2573.9400 381.6000 ;
        RECT 2572.3400 359.3600 2573.9400 359.8400 ;
        RECT 2572.3400 364.8000 2573.9400 365.2800 ;
        RECT 2572.3400 370.2400 2573.9400 370.7200 ;
        RECT 2527.3400 375.6800 2528.9400 376.1600 ;
        RECT 2527.3400 381.1200 2528.9400 381.6000 ;
        RECT 2527.3400 359.3600 2528.9400 359.8400 ;
        RECT 2527.3400 364.8000 2528.9400 365.2800 ;
        RECT 2527.3400 370.2400 2528.9400 370.7200 ;
        RECT 2477.7800 402.8800 2480.7800 403.3600 ;
        RECT 2477.7800 408.3200 2480.7800 408.8000 ;
        RECT 2477.7800 392.0000 2480.7800 392.4800 ;
        RECT 2477.7800 386.5600 2480.7800 387.0400 ;
        RECT 2477.7800 397.4400 2480.7800 397.9200 ;
        RECT 2477.7800 375.6800 2480.7800 376.1600 ;
        RECT 2477.7800 381.1200 2480.7800 381.6000 ;
        RECT 2477.7800 364.8000 2480.7800 365.2800 ;
        RECT 2477.7800 359.3600 2480.7800 359.8400 ;
        RECT 2477.7800 370.2400 2480.7800 370.7200 ;
        RECT 2572.3400 348.4800 2573.9400 348.9600 ;
        RECT 2572.3400 353.9200 2573.9400 354.4000 ;
        RECT 2572.3400 332.1600 2573.9400 332.6400 ;
        RECT 2572.3400 337.6000 2573.9400 338.0800 ;
        RECT 2572.3400 343.0400 2573.9400 343.5200 ;
        RECT 2527.3400 348.4800 2528.9400 348.9600 ;
        RECT 2527.3400 353.9200 2528.9400 354.4000 ;
        RECT 2527.3400 332.1600 2528.9400 332.6400 ;
        RECT 2527.3400 337.6000 2528.9400 338.0800 ;
        RECT 2527.3400 343.0400 2528.9400 343.5200 ;
        RECT 2572.3400 326.7200 2573.9400 327.2000 ;
        RECT 2572.3400 321.2800 2573.9400 321.7600 ;
        RECT 2572.3400 315.8400 2573.9400 316.3200 ;
        RECT 2527.3400 326.7200 2528.9400 327.2000 ;
        RECT 2527.3400 321.2800 2528.9400 321.7600 ;
        RECT 2527.3400 315.8400 2528.9400 316.3200 ;
        RECT 2477.7800 348.4800 2480.7800 348.9600 ;
        RECT 2477.7800 353.9200 2480.7800 354.4000 ;
        RECT 2477.7800 337.6000 2480.7800 338.0800 ;
        RECT 2477.7800 332.1600 2480.7800 332.6400 ;
        RECT 2477.7800 343.0400 2480.7800 343.5200 ;
        RECT 2477.7800 321.2800 2480.7800 321.7600 ;
        RECT 2477.7800 326.7200 2480.7800 327.2000 ;
        RECT 2477.7800 315.8400 2480.7800 316.3200 ;
        RECT 2477.7800 514.0300 2676.8800 517.0300 ;
        RECT 2477.7800 308.9300 2676.8800 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 79.2900 2663.9400 287.3900 ;
        RECT 2617.3400 79.2900 2618.9400 287.3900 ;
        RECT 2572.3400 79.2900 2573.9400 287.3900 ;
        RECT 2527.3400 79.2900 2528.9400 287.3900 ;
        RECT 2673.8800 79.2900 2676.8800 287.3900 ;
        RECT 2477.7800 79.2900 2480.7800 287.3900 ;
      LAYER met3 ;
        RECT 2673.8800 282.0400 2676.8800 282.5200 ;
        RECT 2662.3400 282.0400 2663.9400 282.5200 ;
        RECT 2673.8800 271.1600 2676.8800 271.6400 ;
        RECT 2673.8800 276.6000 2676.8800 277.0800 ;
        RECT 2662.3400 271.1600 2663.9400 271.6400 ;
        RECT 2662.3400 276.6000 2663.9400 277.0800 ;
        RECT 2673.8800 254.8400 2676.8800 255.3200 ;
        RECT 2673.8800 260.2800 2676.8800 260.7600 ;
        RECT 2662.3400 254.8400 2663.9400 255.3200 ;
        RECT 2662.3400 260.2800 2663.9400 260.7600 ;
        RECT 2673.8800 243.9600 2676.8800 244.4400 ;
        RECT 2673.8800 249.4000 2676.8800 249.8800 ;
        RECT 2662.3400 243.9600 2663.9400 244.4400 ;
        RECT 2662.3400 249.4000 2663.9400 249.8800 ;
        RECT 2673.8800 265.7200 2676.8800 266.2000 ;
        RECT 2662.3400 265.7200 2663.9400 266.2000 ;
        RECT 2617.3400 271.1600 2618.9400 271.6400 ;
        RECT 2617.3400 276.6000 2618.9400 277.0800 ;
        RECT 2617.3400 282.0400 2618.9400 282.5200 ;
        RECT 2617.3400 254.8400 2618.9400 255.3200 ;
        RECT 2617.3400 260.2800 2618.9400 260.7600 ;
        RECT 2617.3400 249.4000 2618.9400 249.8800 ;
        RECT 2617.3400 243.9600 2618.9400 244.4400 ;
        RECT 2617.3400 265.7200 2618.9400 266.2000 ;
        RECT 2673.8800 227.6400 2676.8800 228.1200 ;
        RECT 2673.8800 233.0800 2676.8800 233.5600 ;
        RECT 2662.3400 227.6400 2663.9400 228.1200 ;
        RECT 2662.3400 233.0800 2663.9400 233.5600 ;
        RECT 2673.8800 211.3200 2676.8800 211.8000 ;
        RECT 2673.8800 216.7600 2676.8800 217.2400 ;
        RECT 2673.8800 222.2000 2676.8800 222.6800 ;
        RECT 2662.3400 211.3200 2663.9400 211.8000 ;
        RECT 2662.3400 216.7600 2663.9400 217.2400 ;
        RECT 2662.3400 222.2000 2663.9400 222.6800 ;
        RECT 2673.8800 200.4400 2676.8800 200.9200 ;
        RECT 2673.8800 205.8800 2676.8800 206.3600 ;
        RECT 2662.3400 200.4400 2663.9400 200.9200 ;
        RECT 2662.3400 205.8800 2663.9400 206.3600 ;
        RECT 2673.8800 184.1200 2676.8800 184.6000 ;
        RECT 2673.8800 189.5600 2676.8800 190.0400 ;
        RECT 2673.8800 195.0000 2676.8800 195.4800 ;
        RECT 2662.3400 184.1200 2663.9400 184.6000 ;
        RECT 2662.3400 189.5600 2663.9400 190.0400 ;
        RECT 2662.3400 195.0000 2663.9400 195.4800 ;
        RECT 2617.3400 227.6400 2618.9400 228.1200 ;
        RECT 2617.3400 233.0800 2618.9400 233.5600 ;
        RECT 2617.3400 211.3200 2618.9400 211.8000 ;
        RECT 2617.3400 216.7600 2618.9400 217.2400 ;
        RECT 2617.3400 222.2000 2618.9400 222.6800 ;
        RECT 2617.3400 200.4400 2618.9400 200.9200 ;
        RECT 2617.3400 205.8800 2618.9400 206.3600 ;
        RECT 2617.3400 184.1200 2618.9400 184.6000 ;
        RECT 2617.3400 189.5600 2618.9400 190.0400 ;
        RECT 2617.3400 195.0000 2618.9400 195.4800 ;
        RECT 2673.8800 238.5200 2676.8800 239.0000 ;
        RECT 2617.3400 238.5200 2618.9400 239.0000 ;
        RECT 2662.3400 238.5200 2663.9400 239.0000 ;
        RECT 2572.3400 271.1600 2573.9400 271.6400 ;
        RECT 2572.3400 276.6000 2573.9400 277.0800 ;
        RECT 2572.3400 282.0400 2573.9400 282.5200 ;
        RECT 2527.3400 271.1600 2528.9400 271.6400 ;
        RECT 2527.3400 276.6000 2528.9400 277.0800 ;
        RECT 2527.3400 282.0400 2528.9400 282.5200 ;
        RECT 2572.3400 254.8400 2573.9400 255.3200 ;
        RECT 2572.3400 260.2800 2573.9400 260.7600 ;
        RECT 2572.3400 243.9600 2573.9400 244.4400 ;
        RECT 2572.3400 249.4000 2573.9400 249.8800 ;
        RECT 2527.3400 254.8400 2528.9400 255.3200 ;
        RECT 2527.3400 260.2800 2528.9400 260.7600 ;
        RECT 2527.3400 243.9600 2528.9400 244.4400 ;
        RECT 2527.3400 249.4000 2528.9400 249.8800 ;
        RECT 2527.3400 265.7200 2528.9400 266.2000 ;
        RECT 2572.3400 265.7200 2573.9400 266.2000 ;
        RECT 2477.7800 282.0400 2480.7800 282.5200 ;
        RECT 2477.7800 276.6000 2480.7800 277.0800 ;
        RECT 2477.7800 271.1600 2480.7800 271.6400 ;
        RECT 2477.7800 260.2800 2480.7800 260.7600 ;
        RECT 2477.7800 254.8400 2480.7800 255.3200 ;
        RECT 2477.7800 249.4000 2480.7800 249.8800 ;
        RECT 2477.7800 243.9600 2480.7800 244.4400 ;
        RECT 2477.7800 265.7200 2480.7800 266.2000 ;
        RECT 2572.3400 227.6400 2573.9400 228.1200 ;
        RECT 2572.3400 233.0800 2573.9400 233.5600 ;
        RECT 2572.3400 211.3200 2573.9400 211.8000 ;
        RECT 2572.3400 216.7600 2573.9400 217.2400 ;
        RECT 2572.3400 222.2000 2573.9400 222.6800 ;
        RECT 2527.3400 227.6400 2528.9400 228.1200 ;
        RECT 2527.3400 233.0800 2528.9400 233.5600 ;
        RECT 2527.3400 211.3200 2528.9400 211.8000 ;
        RECT 2527.3400 216.7600 2528.9400 217.2400 ;
        RECT 2527.3400 222.2000 2528.9400 222.6800 ;
        RECT 2572.3400 200.4400 2573.9400 200.9200 ;
        RECT 2572.3400 205.8800 2573.9400 206.3600 ;
        RECT 2572.3400 184.1200 2573.9400 184.6000 ;
        RECT 2572.3400 189.5600 2573.9400 190.0400 ;
        RECT 2572.3400 195.0000 2573.9400 195.4800 ;
        RECT 2527.3400 200.4400 2528.9400 200.9200 ;
        RECT 2527.3400 205.8800 2528.9400 206.3600 ;
        RECT 2527.3400 184.1200 2528.9400 184.6000 ;
        RECT 2527.3400 189.5600 2528.9400 190.0400 ;
        RECT 2527.3400 195.0000 2528.9400 195.4800 ;
        RECT 2477.7800 227.6400 2480.7800 228.1200 ;
        RECT 2477.7800 233.0800 2480.7800 233.5600 ;
        RECT 2477.7800 216.7600 2480.7800 217.2400 ;
        RECT 2477.7800 211.3200 2480.7800 211.8000 ;
        RECT 2477.7800 222.2000 2480.7800 222.6800 ;
        RECT 2477.7800 200.4400 2480.7800 200.9200 ;
        RECT 2477.7800 205.8800 2480.7800 206.3600 ;
        RECT 2477.7800 189.5600 2480.7800 190.0400 ;
        RECT 2477.7800 184.1200 2480.7800 184.6000 ;
        RECT 2477.7800 195.0000 2480.7800 195.4800 ;
        RECT 2477.7800 238.5200 2480.7800 239.0000 ;
        RECT 2527.3400 238.5200 2528.9400 239.0000 ;
        RECT 2572.3400 238.5200 2573.9400 239.0000 ;
        RECT 2673.8800 173.2400 2676.8800 173.7200 ;
        RECT 2673.8800 178.6800 2676.8800 179.1600 ;
        RECT 2662.3400 173.2400 2663.9400 173.7200 ;
        RECT 2662.3400 178.6800 2663.9400 179.1600 ;
        RECT 2673.8800 156.9200 2676.8800 157.4000 ;
        RECT 2673.8800 162.3600 2676.8800 162.8400 ;
        RECT 2673.8800 167.8000 2676.8800 168.2800 ;
        RECT 2662.3400 156.9200 2663.9400 157.4000 ;
        RECT 2662.3400 162.3600 2663.9400 162.8400 ;
        RECT 2662.3400 167.8000 2663.9400 168.2800 ;
        RECT 2673.8800 146.0400 2676.8800 146.5200 ;
        RECT 2673.8800 151.4800 2676.8800 151.9600 ;
        RECT 2662.3400 146.0400 2663.9400 146.5200 ;
        RECT 2662.3400 151.4800 2663.9400 151.9600 ;
        RECT 2673.8800 129.7200 2676.8800 130.2000 ;
        RECT 2673.8800 135.1600 2676.8800 135.6400 ;
        RECT 2673.8800 140.6000 2676.8800 141.0800 ;
        RECT 2662.3400 129.7200 2663.9400 130.2000 ;
        RECT 2662.3400 135.1600 2663.9400 135.6400 ;
        RECT 2662.3400 140.6000 2663.9400 141.0800 ;
        RECT 2617.3400 173.2400 2618.9400 173.7200 ;
        RECT 2617.3400 178.6800 2618.9400 179.1600 ;
        RECT 2617.3400 156.9200 2618.9400 157.4000 ;
        RECT 2617.3400 162.3600 2618.9400 162.8400 ;
        RECT 2617.3400 167.8000 2618.9400 168.2800 ;
        RECT 2617.3400 146.0400 2618.9400 146.5200 ;
        RECT 2617.3400 151.4800 2618.9400 151.9600 ;
        RECT 2617.3400 129.7200 2618.9400 130.2000 ;
        RECT 2617.3400 135.1600 2618.9400 135.6400 ;
        RECT 2617.3400 140.6000 2618.9400 141.0800 ;
        RECT 2673.8800 118.8400 2676.8800 119.3200 ;
        RECT 2673.8800 124.2800 2676.8800 124.7600 ;
        RECT 2662.3400 118.8400 2663.9400 119.3200 ;
        RECT 2662.3400 124.2800 2663.9400 124.7600 ;
        RECT 2673.8800 102.5200 2676.8800 103.0000 ;
        RECT 2673.8800 107.9600 2676.8800 108.4400 ;
        RECT 2673.8800 113.4000 2676.8800 113.8800 ;
        RECT 2662.3400 102.5200 2663.9400 103.0000 ;
        RECT 2662.3400 107.9600 2663.9400 108.4400 ;
        RECT 2662.3400 113.4000 2663.9400 113.8800 ;
        RECT 2673.8800 91.6400 2676.8800 92.1200 ;
        RECT 2673.8800 97.0800 2676.8800 97.5600 ;
        RECT 2662.3400 91.6400 2663.9400 92.1200 ;
        RECT 2662.3400 97.0800 2663.9400 97.5600 ;
        RECT 2673.8800 86.2000 2676.8800 86.6800 ;
        RECT 2662.3400 86.2000 2663.9400 86.6800 ;
        RECT 2617.3400 118.8400 2618.9400 119.3200 ;
        RECT 2617.3400 124.2800 2618.9400 124.7600 ;
        RECT 2617.3400 102.5200 2618.9400 103.0000 ;
        RECT 2617.3400 107.9600 2618.9400 108.4400 ;
        RECT 2617.3400 113.4000 2618.9400 113.8800 ;
        RECT 2617.3400 91.6400 2618.9400 92.1200 ;
        RECT 2617.3400 97.0800 2618.9400 97.5600 ;
        RECT 2617.3400 86.2000 2618.9400 86.6800 ;
        RECT 2572.3400 173.2400 2573.9400 173.7200 ;
        RECT 2572.3400 178.6800 2573.9400 179.1600 ;
        RECT 2572.3400 156.9200 2573.9400 157.4000 ;
        RECT 2572.3400 162.3600 2573.9400 162.8400 ;
        RECT 2572.3400 167.8000 2573.9400 168.2800 ;
        RECT 2527.3400 173.2400 2528.9400 173.7200 ;
        RECT 2527.3400 178.6800 2528.9400 179.1600 ;
        RECT 2527.3400 156.9200 2528.9400 157.4000 ;
        RECT 2527.3400 162.3600 2528.9400 162.8400 ;
        RECT 2527.3400 167.8000 2528.9400 168.2800 ;
        RECT 2572.3400 146.0400 2573.9400 146.5200 ;
        RECT 2572.3400 151.4800 2573.9400 151.9600 ;
        RECT 2572.3400 129.7200 2573.9400 130.2000 ;
        RECT 2572.3400 135.1600 2573.9400 135.6400 ;
        RECT 2572.3400 140.6000 2573.9400 141.0800 ;
        RECT 2527.3400 146.0400 2528.9400 146.5200 ;
        RECT 2527.3400 151.4800 2528.9400 151.9600 ;
        RECT 2527.3400 129.7200 2528.9400 130.2000 ;
        RECT 2527.3400 135.1600 2528.9400 135.6400 ;
        RECT 2527.3400 140.6000 2528.9400 141.0800 ;
        RECT 2477.7800 173.2400 2480.7800 173.7200 ;
        RECT 2477.7800 178.6800 2480.7800 179.1600 ;
        RECT 2477.7800 162.3600 2480.7800 162.8400 ;
        RECT 2477.7800 156.9200 2480.7800 157.4000 ;
        RECT 2477.7800 167.8000 2480.7800 168.2800 ;
        RECT 2477.7800 146.0400 2480.7800 146.5200 ;
        RECT 2477.7800 151.4800 2480.7800 151.9600 ;
        RECT 2477.7800 135.1600 2480.7800 135.6400 ;
        RECT 2477.7800 129.7200 2480.7800 130.2000 ;
        RECT 2477.7800 140.6000 2480.7800 141.0800 ;
        RECT 2572.3400 118.8400 2573.9400 119.3200 ;
        RECT 2572.3400 124.2800 2573.9400 124.7600 ;
        RECT 2572.3400 102.5200 2573.9400 103.0000 ;
        RECT 2572.3400 107.9600 2573.9400 108.4400 ;
        RECT 2572.3400 113.4000 2573.9400 113.8800 ;
        RECT 2527.3400 118.8400 2528.9400 119.3200 ;
        RECT 2527.3400 124.2800 2528.9400 124.7600 ;
        RECT 2527.3400 102.5200 2528.9400 103.0000 ;
        RECT 2527.3400 107.9600 2528.9400 108.4400 ;
        RECT 2527.3400 113.4000 2528.9400 113.8800 ;
        RECT 2572.3400 97.0800 2573.9400 97.5600 ;
        RECT 2572.3400 91.6400 2573.9400 92.1200 ;
        RECT 2572.3400 86.2000 2573.9400 86.6800 ;
        RECT 2527.3400 97.0800 2528.9400 97.5600 ;
        RECT 2527.3400 91.6400 2528.9400 92.1200 ;
        RECT 2527.3400 86.2000 2528.9400 86.6800 ;
        RECT 2477.7800 118.8400 2480.7800 119.3200 ;
        RECT 2477.7800 124.2800 2480.7800 124.7600 ;
        RECT 2477.7800 107.9600 2480.7800 108.4400 ;
        RECT 2477.7800 102.5200 2480.7800 103.0000 ;
        RECT 2477.7800 113.4000 2480.7800 113.8800 ;
        RECT 2477.7800 91.6400 2480.7800 92.1200 ;
        RECT 2477.7800 97.0800 2480.7800 97.5600 ;
        RECT 2477.7800 86.2000 2480.7800 86.6800 ;
        RECT 2477.7800 284.3900 2676.8800 287.3900 ;
        RECT 2477.7800 79.2900 2676.8800 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 2477.7800 37.6700 2479.7800 58.6000 ;
        RECT 2674.8800 37.6700 2676.8800 58.6000 ;
      LAYER met3 ;
        RECT 2674.8800 54.1000 2676.8800 54.5800 ;
        RECT 2477.7800 54.1000 2479.7800 54.5800 ;
        RECT 2674.8800 43.2200 2676.8800 43.7000 ;
        RECT 2477.7800 43.2200 2479.7800 43.7000 ;
        RECT 2674.8800 48.6600 2676.8800 49.1400 ;
        RECT 2477.7800 48.6600 2479.7800 49.1400 ;
        RECT 2477.7800 56.6000 2676.8800 58.6000 ;
        RECT 2477.7800 37.6700 2676.8800 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 2605.3300 2663.9400 2813.4300 ;
        RECT 2617.3400 2605.3300 2618.9400 2813.4300 ;
        RECT 2572.3400 2605.3300 2573.9400 2813.4300 ;
        RECT 2527.3400 2605.3300 2528.9400 2813.4300 ;
        RECT 2673.8800 2605.3300 2676.8800 2813.4300 ;
        RECT 2477.7800 2605.3300 2480.7800 2813.4300 ;
      LAYER met3 ;
        RECT 2673.8800 2808.0800 2676.8800 2808.5600 ;
        RECT 2662.3400 2808.0800 2663.9400 2808.5600 ;
        RECT 2673.8800 2797.2000 2676.8800 2797.6800 ;
        RECT 2673.8800 2802.6400 2676.8800 2803.1200 ;
        RECT 2662.3400 2797.2000 2663.9400 2797.6800 ;
        RECT 2662.3400 2802.6400 2663.9400 2803.1200 ;
        RECT 2673.8800 2780.8800 2676.8800 2781.3600 ;
        RECT 2673.8800 2786.3200 2676.8800 2786.8000 ;
        RECT 2662.3400 2780.8800 2663.9400 2781.3600 ;
        RECT 2662.3400 2786.3200 2663.9400 2786.8000 ;
        RECT 2673.8800 2770.0000 2676.8800 2770.4800 ;
        RECT 2673.8800 2775.4400 2676.8800 2775.9200 ;
        RECT 2662.3400 2770.0000 2663.9400 2770.4800 ;
        RECT 2662.3400 2775.4400 2663.9400 2775.9200 ;
        RECT 2673.8800 2791.7600 2676.8800 2792.2400 ;
        RECT 2662.3400 2791.7600 2663.9400 2792.2400 ;
        RECT 2617.3400 2797.2000 2618.9400 2797.6800 ;
        RECT 2617.3400 2802.6400 2618.9400 2803.1200 ;
        RECT 2617.3400 2808.0800 2618.9400 2808.5600 ;
        RECT 2617.3400 2780.8800 2618.9400 2781.3600 ;
        RECT 2617.3400 2786.3200 2618.9400 2786.8000 ;
        RECT 2617.3400 2775.4400 2618.9400 2775.9200 ;
        RECT 2617.3400 2770.0000 2618.9400 2770.4800 ;
        RECT 2617.3400 2791.7600 2618.9400 2792.2400 ;
        RECT 2673.8800 2753.6800 2676.8800 2754.1600 ;
        RECT 2673.8800 2759.1200 2676.8800 2759.6000 ;
        RECT 2662.3400 2753.6800 2663.9400 2754.1600 ;
        RECT 2662.3400 2759.1200 2663.9400 2759.6000 ;
        RECT 2673.8800 2737.3600 2676.8800 2737.8400 ;
        RECT 2673.8800 2742.8000 2676.8800 2743.2800 ;
        RECT 2673.8800 2748.2400 2676.8800 2748.7200 ;
        RECT 2662.3400 2737.3600 2663.9400 2737.8400 ;
        RECT 2662.3400 2742.8000 2663.9400 2743.2800 ;
        RECT 2662.3400 2748.2400 2663.9400 2748.7200 ;
        RECT 2673.8800 2726.4800 2676.8800 2726.9600 ;
        RECT 2673.8800 2731.9200 2676.8800 2732.4000 ;
        RECT 2662.3400 2726.4800 2663.9400 2726.9600 ;
        RECT 2662.3400 2731.9200 2663.9400 2732.4000 ;
        RECT 2673.8800 2710.1600 2676.8800 2710.6400 ;
        RECT 2673.8800 2715.6000 2676.8800 2716.0800 ;
        RECT 2673.8800 2721.0400 2676.8800 2721.5200 ;
        RECT 2662.3400 2710.1600 2663.9400 2710.6400 ;
        RECT 2662.3400 2715.6000 2663.9400 2716.0800 ;
        RECT 2662.3400 2721.0400 2663.9400 2721.5200 ;
        RECT 2617.3400 2753.6800 2618.9400 2754.1600 ;
        RECT 2617.3400 2759.1200 2618.9400 2759.6000 ;
        RECT 2617.3400 2737.3600 2618.9400 2737.8400 ;
        RECT 2617.3400 2742.8000 2618.9400 2743.2800 ;
        RECT 2617.3400 2748.2400 2618.9400 2748.7200 ;
        RECT 2617.3400 2726.4800 2618.9400 2726.9600 ;
        RECT 2617.3400 2731.9200 2618.9400 2732.4000 ;
        RECT 2617.3400 2710.1600 2618.9400 2710.6400 ;
        RECT 2617.3400 2715.6000 2618.9400 2716.0800 ;
        RECT 2617.3400 2721.0400 2618.9400 2721.5200 ;
        RECT 2673.8800 2764.5600 2676.8800 2765.0400 ;
        RECT 2617.3400 2764.5600 2618.9400 2765.0400 ;
        RECT 2662.3400 2764.5600 2663.9400 2765.0400 ;
        RECT 2572.3400 2797.2000 2573.9400 2797.6800 ;
        RECT 2572.3400 2802.6400 2573.9400 2803.1200 ;
        RECT 2572.3400 2808.0800 2573.9400 2808.5600 ;
        RECT 2527.3400 2797.2000 2528.9400 2797.6800 ;
        RECT 2527.3400 2802.6400 2528.9400 2803.1200 ;
        RECT 2527.3400 2808.0800 2528.9400 2808.5600 ;
        RECT 2572.3400 2780.8800 2573.9400 2781.3600 ;
        RECT 2572.3400 2786.3200 2573.9400 2786.8000 ;
        RECT 2572.3400 2770.0000 2573.9400 2770.4800 ;
        RECT 2572.3400 2775.4400 2573.9400 2775.9200 ;
        RECT 2527.3400 2780.8800 2528.9400 2781.3600 ;
        RECT 2527.3400 2786.3200 2528.9400 2786.8000 ;
        RECT 2527.3400 2770.0000 2528.9400 2770.4800 ;
        RECT 2527.3400 2775.4400 2528.9400 2775.9200 ;
        RECT 2527.3400 2791.7600 2528.9400 2792.2400 ;
        RECT 2572.3400 2791.7600 2573.9400 2792.2400 ;
        RECT 2477.7800 2808.0800 2480.7800 2808.5600 ;
        RECT 2477.7800 2802.6400 2480.7800 2803.1200 ;
        RECT 2477.7800 2797.2000 2480.7800 2797.6800 ;
        RECT 2477.7800 2786.3200 2480.7800 2786.8000 ;
        RECT 2477.7800 2780.8800 2480.7800 2781.3600 ;
        RECT 2477.7800 2775.4400 2480.7800 2775.9200 ;
        RECT 2477.7800 2770.0000 2480.7800 2770.4800 ;
        RECT 2477.7800 2791.7600 2480.7800 2792.2400 ;
        RECT 2572.3400 2753.6800 2573.9400 2754.1600 ;
        RECT 2572.3400 2759.1200 2573.9400 2759.6000 ;
        RECT 2572.3400 2737.3600 2573.9400 2737.8400 ;
        RECT 2572.3400 2742.8000 2573.9400 2743.2800 ;
        RECT 2572.3400 2748.2400 2573.9400 2748.7200 ;
        RECT 2527.3400 2753.6800 2528.9400 2754.1600 ;
        RECT 2527.3400 2759.1200 2528.9400 2759.6000 ;
        RECT 2527.3400 2737.3600 2528.9400 2737.8400 ;
        RECT 2527.3400 2742.8000 2528.9400 2743.2800 ;
        RECT 2527.3400 2748.2400 2528.9400 2748.7200 ;
        RECT 2572.3400 2726.4800 2573.9400 2726.9600 ;
        RECT 2572.3400 2731.9200 2573.9400 2732.4000 ;
        RECT 2572.3400 2710.1600 2573.9400 2710.6400 ;
        RECT 2572.3400 2715.6000 2573.9400 2716.0800 ;
        RECT 2572.3400 2721.0400 2573.9400 2721.5200 ;
        RECT 2527.3400 2726.4800 2528.9400 2726.9600 ;
        RECT 2527.3400 2731.9200 2528.9400 2732.4000 ;
        RECT 2527.3400 2710.1600 2528.9400 2710.6400 ;
        RECT 2527.3400 2715.6000 2528.9400 2716.0800 ;
        RECT 2527.3400 2721.0400 2528.9400 2721.5200 ;
        RECT 2477.7800 2753.6800 2480.7800 2754.1600 ;
        RECT 2477.7800 2759.1200 2480.7800 2759.6000 ;
        RECT 2477.7800 2742.8000 2480.7800 2743.2800 ;
        RECT 2477.7800 2737.3600 2480.7800 2737.8400 ;
        RECT 2477.7800 2748.2400 2480.7800 2748.7200 ;
        RECT 2477.7800 2726.4800 2480.7800 2726.9600 ;
        RECT 2477.7800 2731.9200 2480.7800 2732.4000 ;
        RECT 2477.7800 2715.6000 2480.7800 2716.0800 ;
        RECT 2477.7800 2710.1600 2480.7800 2710.6400 ;
        RECT 2477.7800 2721.0400 2480.7800 2721.5200 ;
        RECT 2477.7800 2764.5600 2480.7800 2765.0400 ;
        RECT 2527.3400 2764.5600 2528.9400 2765.0400 ;
        RECT 2572.3400 2764.5600 2573.9400 2765.0400 ;
        RECT 2673.8800 2699.2800 2676.8800 2699.7600 ;
        RECT 2673.8800 2704.7200 2676.8800 2705.2000 ;
        RECT 2662.3400 2699.2800 2663.9400 2699.7600 ;
        RECT 2662.3400 2704.7200 2663.9400 2705.2000 ;
        RECT 2673.8800 2682.9600 2676.8800 2683.4400 ;
        RECT 2673.8800 2688.4000 2676.8800 2688.8800 ;
        RECT 2673.8800 2693.8400 2676.8800 2694.3200 ;
        RECT 2662.3400 2682.9600 2663.9400 2683.4400 ;
        RECT 2662.3400 2688.4000 2663.9400 2688.8800 ;
        RECT 2662.3400 2693.8400 2663.9400 2694.3200 ;
        RECT 2673.8800 2672.0800 2676.8800 2672.5600 ;
        RECT 2673.8800 2677.5200 2676.8800 2678.0000 ;
        RECT 2662.3400 2672.0800 2663.9400 2672.5600 ;
        RECT 2662.3400 2677.5200 2663.9400 2678.0000 ;
        RECT 2673.8800 2655.7600 2676.8800 2656.2400 ;
        RECT 2673.8800 2661.2000 2676.8800 2661.6800 ;
        RECT 2673.8800 2666.6400 2676.8800 2667.1200 ;
        RECT 2662.3400 2655.7600 2663.9400 2656.2400 ;
        RECT 2662.3400 2661.2000 2663.9400 2661.6800 ;
        RECT 2662.3400 2666.6400 2663.9400 2667.1200 ;
        RECT 2617.3400 2699.2800 2618.9400 2699.7600 ;
        RECT 2617.3400 2704.7200 2618.9400 2705.2000 ;
        RECT 2617.3400 2682.9600 2618.9400 2683.4400 ;
        RECT 2617.3400 2688.4000 2618.9400 2688.8800 ;
        RECT 2617.3400 2693.8400 2618.9400 2694.3200 ;
        RECT 2617.3400 2672.0800 2618.9400 2672.5600 ;
        RECT 2617.3400 2677.5200 2618.9400 2678.0000 ;
        RECT 2617.3400 2655.7600 2618.9400 2656.2400 ;
        RECT 2617.3400 2661.2000 2618.9400 2661.6800 ;
        RECT 2617.3400 2666.6400 2618.9400 2667.1200 ;
        RECT 2673.8800 2644.8800 2676.8800 2645.3600 ;
        RECT 2673.8800 2650.3200 2676.8800 2650.8000 ;
        RECT 2662.3400 2644.8800 2663.9400 2645.3600 ;
        RECT 2662.3400 2650.3200 2663.9400 2650.8000 ;
        RECT 2673.8800 2628.5600 2676.8800 2629.0400 ;
        RECT 2673.8800 2634.0000 2676.8800 2634.4800 ;
        RECT 2673.8800 2639.4400 2676.8800 2639.9200 ;
        RECT 2662.3400 2628.5600 2663.9400 2629.0400 ;
        RECT 2662.3400 2634.0000 2663.9400 2634.4800 ;
        RECT 2662.3400 2639.4400 2663.9400 2639.9200 ;
        RECT 2673.8800 2617.6800 2676.8800 2618.1600 ;
        RECT 2673.8800 2623.1200 2676.8800 2623.6000 ;
        RECT 2662.3400 2617.6800 2663.9400 2618.1600 ;
        RECT 2662.3400 2623.1200 2663.9400 2623.6000 ;
        RECT 2673.8800 2612.2400 2676.8800 2612.7200 ;
        RECT 2662.3400 2612.2400 2663.9400 2612.7200 ;
        RECT 2617.3400 2644.8800 2618.9400 2645.3600 ;
        RECT 2617.3400 2650.3200 2618.9400 2650.8000 ;
        RECT 2617.3400 2628.5600 2618.9400 2629.0400 ;
        RECT 2617.3400 2634.0000 2618.9400 2634.4800 ;
        RECT 2617.3400 2639.4400 2618.9400 2639.9200 ;
        RECT 2617.3400 2617.6800 2618.9400 2618.1600 ;
        RECT 2617.3400 2623.1200 2618.9400 2623.6000 ;
        RECT 2617.3400 2612.2400 2618.9400 2612.7200 ;
        RECT 2572.3400 2699.2800 2573.9400 2699.7600 ;
        RECT 2572.3400 2704.7200 2573.9400 2705.2000 ;
        RECT 2572.3400 2682.9600 2573.9400 2683.4400 ;
        RECT 2572.3400 2688.4000 2573.9400 2688.8800 ;
        RECT 2572.3400 2693.8400 2573.9400 2694.3200 ;
        RECT 2527.3400 2699.2800 2528.9400 2699.7600 ;
        RECT 2527.3400 2704.7200 2528.9400 2705.2000 ;
        RECT 2527.3400 2682.9600 2528.9400 2683.4400 ;
        RECT 2527.3400 2688.4000 2528.9400 2688.8800 ;
        RECT 2527.3400 2693.8400 2528.9400 2694.3200 ;
        RECT 2572.3400 2672.0800 2573.9400 2672.5600 ;
        RECT 2572.3400 2677.5200 2573.9400 2678.0000 ;
        RECT 2572.3400 2655.7600 2573.9400 2656.2400 ;
        RECT 2572.3400 2661.2000 2573.9400 2661.6800 ;
        RECT 2572.3400 2666.6400 2573.9400 2667.1200 ;
        RECT 2527.3400 2672.0800 2528.9400 2672.5600 ;
        RECT 2527.3400 2677.5200 2528.9400 2678.0000 ;
        RECT 2527.3400 2655.7600 2528.9400 2656.2400 ;
        RECT 2527.3400 2661.2000 2528.9400 2661.6800 ;
        RECT 2527.3400 2666.6400 2528.9400 2667.1200 ;
        RECT 2477.7800 2699.2800 2480.7800 2699.7600 ;
        RECT 2477.7800 2704.7200 2480.7800 2705.2000 ;
        RECT 2477.7800 2688.4000 2480.7800 2688.8800 ;
        RECT 2477.7800 2682.9600 2480.7800 2683.4400 ;
        RECT 2477.7800 2693.8400 2480.7800 2694.3200 ;
        RECT 2477.7800 2672.0800 2480.7800 2672.5600 ;
        RECT 2477.7800 2677.5200 2480.7800 2678.0000 ;
        RECT 2477.7800 2661.2000 2480.7800 2661.6800 ;
        RECT 2477.7800 2655.7600 2480.7800 2656.2400 ;
        RECT 2477.7800 2666.6400 2480.7800 2667.1200 ;
        RECT 2572.3400 2644.8800 2573.9400 2645.3600 ;
        RECT 2572.3400 2650.3200 2573.9400 2650.8000 ;
        RECT 2572.3400 2628.5600 2573.9400 2629.0400 ;
        RECT 2572.3400 2634.0000 2573.9400 2634.4800 ;
        RECT 2572.3400 2639.4400 2573.9400 2639.9200 ;
        RECT 2527.3400 2644.8800 2528.9400 2645.3600 ;
        RECT 2527.3400 2650.3200 2528.9400 2650.8000 ;
        RECT 2527.3400 2628.5600 2528.9400 2629.0400 ;
        RECT 2527.3400 2634.0000 2528.9400 2634.4800 ;
        RECT 2527.3400 2639.4400 2528.9400 2639.9200 ;
        RECT 2572.3400 2623.1200 2573.9400 2623.6000 ;
        RECT 2572.3400 2617.6800 2573.9400 2618.1600 ;
        RECT 2572.3400 2612.2400 2573.9400 2612.7200 ;
        RECT 2527.3400 2623.1200 2528.9400 2623.6000 ;
        RECT 2527.3400 2617.6800 2528.9400 2618.1600 ;
        RECT 2527.3400 2612.2400 2528.9400 2612.7200 ;
        RECT 2477.7800 2644.8800 2480.7800 2645.3600 ;
        RECT 2477.7800 2650.3200 2480.7800 2650.8000 ;
        RECT 2477.7800 2634.0000 2480.7800 2634.4800 ;
        RECT 2477.7800 2628.5600 2480.7800 2629.0400 ;
        RECT 2477.7800 2639.4400 2480.7800 2639.9200 ;
        RECT 2477.7800 2617.6800 2480.7800 2618.1600 ;
        RECT 2477.7800 2623.1200 2480.7800 2623.6000 ;
        RECT 2477.7800 2612.2400 2480.7800 2612.7200 ;
        RECT 2477.7800 2810.4300 2676.8800 2813.4300 ;
        RECT 2477.7800 2605.3300 2676.8800 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 2375.6900 2663.9400 2583.7900 ;
        RECT 2617.3400 2375.6900 2618.9400 2583.7900 ;
        RECT 2572.3400 2375.6900 2573.9400 2583.7900 ;
        RECT 2527.3400 2375.6900 2528.9400 2583.7900 ;
        RECT 2673.8800 2375.6900 2676.8800 2583.7900 ;
        RECT 2477.7800 2375.6900 2480.7800 2583.7900 ;
      LAYER met3 ;
        RECT 2673.8800 2578.4400 2676.8800 2578.9200 ;
        RECT 2662.3400 2578.4400 2663.9400 2578.9200 ;
        RECT 2673.8800 2567.5600 2676.8800 2568.0400 ;
        RECT 2673.8800 2573.0000 2676.8800 2573.4800 ;
        RECT 2662.3400 2567.5600 2663.9400 2568.0400 ;
        RECT 2662.3400 2573.0000 2663.9400 2573.4800 ;
        RECT 2673.8800 2551.2400 2676.8800 2551.7200 ;
        RECT 2673.8800 2556.6800 2676.8800 2557.1600 ;
        RECT 2662.3400 2551.2400 2663.9400 2551.7200 ;
        RECT 2662.3400 2556.6800 2663.9400 2557.1600 ;
        RECT 2673.8800 2540.3600 2676.8800 2540.8400 ;
        RECT 2673.8800 2545.8000 2676.8800 2546.2800 ;
        RECT 2662.3400 2540.3600 2663.9400 2540.8400 ;
        RECT 2662.3400 2545.8000 2663.9400 2546.2800 ;
        RECT 2673.8800 2562.1200 2676.8800 2562.6000 ;
        RECT 2662.3400 2562.1200 2663.9400 2562.6000 ;
        RECT 2617.3400 2567.5600 2618.9400 2568.0400 ;
        RECT 2617.3400 2573.0000 2618.9400 2573.4800 ;
        RECT 2617.3400 2578.4400 2618.9400 2578.9200 ;
        RECT 2617.3400 2551.2400 2618.9400 2551.7200 ;
        RECT 2617.3400 2556.6800 2618.9400 2557.1600 ;
        RECT 2617.3400 2545.8000 2618.9400 2546.2800 ;
        RECT 2617.3400 2540.3600 2618.9400 2540.8400 ;
        RECT 2617.3400 2562.1200 2618.9400 2562.6000 ;
        RECT 2673.8800 2524.0400 2676.8800 2524.5200 ;
        RECT 2673.8800 2529.4800 2676.8800 2529.9600 ;
        RECT 2662.3400 2524.0400 2663.9400 2524.5200 ;
        RECT 2662.3400 2529.4800 2663.9400 2529.9600 ;
        RECT 2673.8800 2507.7200 2676.8800 2508.2000 ;
        RECT 2673.8800 2513.1600 2676.8800 2513.6400 ;
        RECT 2673.8800 2518.6000 2676.8800 2519.0800 ;
        RECT 2662.3400 2507.7200 2663.9400 2508.2000 ;
        RECT 2662.3400 2513.1600 2663.9400 2513.6400 ;
        RECT 2662.3400 2518.6000 2663.9400 2519.0800 ;
        RECT 2673.8800 2496.8400 2676.8800 2497.3200 ;
        RECT 2673.8800 2502.2800 2676.8800 2502.7600 ;
        RECT 2662.3400 2496.8400 2663.9400 2497.3200 ;
        RECT 2662.3400 2502.2800 2663.9400 2502.7600 ;
        RECT 2673.8800 2480.5200 2676.8800 2481.0000 ;
        RECT 2673.8800 2485.9600 2676.8800 2486.4400 ;
        RECT 2673.8800 2491.4000 2676.8800 2491.8800 ;
        RECT 2662.3400 2480.5200 2663.9400 2481.0000 ;
        RECT 2662.3400 2485.9600 2663.9400 2486.4400 ;
        RECT 2662.3400 2491.4000 2663.9400 2491.8800 ;
        RECT 2617.3400 2524.0400 2618.9400 2524.5200 ;
        RECT 2617.3400 2529.4800 2618.9400 2529.9600 ;
        RECT 2617.3400 2507.7200 2618.9400 2508.2000 ;
        RECT 2617.3400 2513.1600 2618.9400 2513.6400 ;
        RECT 2617.3400 2518.6000 2618.9400 2519.0800 ;
        RECT 2617.3400 2496.8400 2618.9400 2497.3200 ;
        RECT 2617.3400 2502.2800 2618.9400 2502.7600 ;
        RECT 2617.3400 2480.5200 2618.9400 2481.0000 ;
        RECT 2617.3400 2485.9600 2618.9400 2486.4400 ;
        RECT 2617.3400 2491.4000 2618.9400 2491.8800 ;
        RECT 2673.8800 2534.9200 2676.8800 2535.4000 ;
        RECT 2617.3400 2534.9200 2618.9400 2535.4000 ;
        RECT 2662.3400 2534.9200 2663.9400 2535.4000 ;
        RECT 2572.3400 2567.5600 2573.9400 2568.0400 ;
        RECT 2572.3400 2573.0000 2573.9400 2573.4800 ;
        RECT 2572.3400 2578.4400 2573.9400 2578.9200 ;
        RECT 2527.3400 2567.5600 2528.9400 2568.0400 ;
        RECT 2527.3400 2573.0000 2528.9400 2573.4800 ;
        RECT 2527.3400 2578.4400 2528.9400 2578.9200 ;
        RECT 2572.3400 2551.2400 2573.9400 2551.7200 ;
        RECT 2572.3400 2556.6800 2573.9400 2557.1600 ;
        RECT 2572.3400 2540.3600 2573.9400 2540.8400 ;
        RECT 2572.3400 2545.8000 2573.9400 2546.2800 ;
        RECT 2527.3400 2551.2400 2528.9400 2551.7200 ;
        RECT 2527.3400 2556.6800 2528.9400 2557.1600 ;
        RECT 2527.3400 2540.3600 2528.9400 2540.8400 ;
        RECT 2527.3400 2545.8000 2528.9400 2546.2800 ;
        RECT 2527.3400 2562.1200 2528.9400 2562.6000 ;
        RECT 2572.3400 2562.1200 2573.9400 2562.6000 ;
        RECT 2477.7800 2578.4400 2480.7800 2578.9200 ;
        RECT 2477.7800 2573.0000 2480.7800 2573.4800 ;
        RECT 2477.7800 2567.5600 2480.7800 2568.0400 ;
        RECT 2477.7800 2556.6800 2480.7800 2557.1600 ;
        RECT 2477.7800 2551.2400 2480.7800 2551.7200 ;
        RECT 2477.7800 2545.8000 2480.7800 2546.2800 ;
        RECT 2477.7800 2540.3600 2480.7800 2540.8400 ;
        RECT 2477.7800 2562.1200 2480.7800 2562.6000 ;
        RECT 2572.3400 2524.0400 2573.9400 2524.5200 ;
        RECT 2572.3400 2529.4800 2573.9400 2529.9600 ;
        RECT 2572.3400 2507.7200 2573.9400 2508.2000 ;
        RECT 2572.3400 2513.1600 2573.9400 2513.6400 ;
        RECT 2572.3400 2518.6000 2573.9400 2519.0800 ;
        RECT 2527.3400 2524.0400 2528.9400 2524.5200 ;
        RECT 2527.3400 2529.4800 2528.9400 2529.9600 ;
        RECT 2527.3400 2507.7200 2528.9400 2508.2000 ;
        RECT 2527.3400 2513.1600 2528.9400 2513.6400 ;
        RECT 2527.3400 2518.6000 2528.9400 2519.0800 ;
        RECT 2572.3400 2496.8400 2573.9400 2497.3200 ;
        RECT 2572.3400 2502.2800 2573.9400 2502.7600 ;
        RECT 2572.3400 2480.5200 2573.9400 2481.0000 ;
        RECT 2572.3400 2485.9600 2573.9400 2486.4400 ;
        RECT 2572.3400 2491.4000 2573.9400 2491.8800 ;
        RECT 2527.3400 2496.8400 2528.9400 2497.3200 ;
        RECT 2527.3400 2502.2800 2528.9400 2502.7600 ;
        RECT 2527.3400 2480.5200 2528.9400 2481.0000 ;
        RECT 2527.3400 2485.9600 2528.9400 2486.4400 ;
        RECT 2527.3400 2491.4000 2528.9400 2491.8800 ;
        RECT 2477.7800 2524.0400 2480.7800 2524.5200 ;
        RECT 2477.7800 2529.4800 2480.7800 2529.9600 ;
        RECT 2477.7800 2513.1600 2480.7800 2513.6400 ;
        RECT 2477.7800 2507.7200 2480.7800 2508.2000 ;
        RECT 2477.7800 2518.6000 2480.7800 2519.0800 ;
        RECT 2477.7800 2496.8400 2480.7800 2497.3200 ;
        RECT 2477.7800 2502.2800 2480.7800 2502.7600 ;
        RECT 2477.7800 2485.9600 2480.7800 2486.4400 ;
        RECT 2477.7800 2480.5200 2480.7800 2481.0000 ;
        RECT 2477.7800 2491.4000 2480.7800 2491.8800 ;
        RECT 2477.7800 2534.9200 2480.7800 2535.4000 ;
        RECT 2527.3400 2534.9200 2528.9400 2535.4000 ;
        RECT 2572.3400 2534.9200 2573.9400 2535.4000 ;
        RECT 2673.8800 2469.6400 2676.8800 2470.1200 ;
        RECT 2673.8800 2475.0800 2676.8800 2475.5600 ;
        RECT 2662.3400 2469.6400 2663.9400 2470.1200 ;
        RECT 2662.3400 2475.0800 2663.9400 2475.5600 ;
        RECT 2673.8800 2453.3200 2676.8800 2453.8000 ;
        RECT 2673.8800 2458.7600 2676.8800 2459.2400 ;
        RECT 2673.8800 2464.2000 2676.8800 2464.6800 ;
        RECT 2662.3400 2453.3200 2663.9400 2453.8000 ;
        RECT 2662.3400 2458.7600 2663.9400 2459.2400 ;
        RECT 2662.3400 2464.2000 2663.9400 2464.6800 ;
        RECT 2673.8800 2442.4400 2676.8800 2442.9200 ;
        RECT 2673.8800 2447.8800 2676.8800 2448.3600 ;
        RECT 2662.3400 2442.4400 2663.9400 2442.9200 ;
        RECT 2662.3400 2447.8800 2663.9400 2448.3600 ;
        RECT 2673.8800 2426.1200 2676.8800 2426.6000 ;
        RECT 2673.8800 2431.5600 2676.8800 2432.0400 ;
        RECT 2673.8800 2437.0000 2676.8800 2437.4800 ;
        RECT 2662.3400 2426.1200 2663.9400 2426.6000 ;
        RECT 2662.3400 2431.5600 2663.9400 2432.0400 ;
        RECT 2662.3400 2437.0000 2663.9400 2437.4800 ;
        RECT 2617.3400 2469.6400 2618.9400 2470.1200 ;
        RECT 2617.3400 2475.0800 2618.9400 2475.5600 ;
        RECT 2617.3400 2453.3200 2618.9400 2453.8000 ;
        RECT 2617.3400 2458.7600 2618.9400 2459.2400 ;
        RECT 2617.3400 2464.2000 2618.9400 2464.6800 ;
        RECT 2617.3400 2442.4400 2618.9400 2442.9200 ;
        RECT 2617.3400 2447.8800 2618.9400 2448.3600 ;
        RECT 2617.3400 2426.1200 2618.9400 2426.6000 ;
        RECT 2617.3400 2431.5600 2618.9400 2432.0400 ;
        RECT 2617.3400 2437.0000 2618.9400 2437.4800 ;
        RECT 2673.8800 2415.2400 2676.8800 2415.7200 ;
        RECT 2673.8800 2420.6800 2676.8800 2421.1600 ;
        RECT 2662.3400 2415.2400 2663.9400 2415.7200 ;
        RECT 2662.3400 2420.6800 2663.9400 2421.1600 ;
        RECT 2673.8800 2398.9200 2676.8800 2399.4000 ;
        RECT 2673.8800 2404.3600 2676.8800 2404.8400 ;
        RECT 2673.8800 2409.8000 2676.8800 2410.2800 ;
        RECT 2662.3400 2398.9200 2663.9400 2399.4000 ;
        RECT 2662.3400 2404.3600 2663.9400 2404.8400 ;
        RECT 2662.3400 2409.8000 2663.9400 2410.2800 ;
        RECT 2673.8800 2388.0400 2676.8800 2388.5200 ;
        RECT 2673.8800 2393.4800 2676.8800 2393.9600 ;
        RECT 2662.3400 2388.0400 2663.9400 2388.5200 ;
        RECT 2662.3400 2393.4800 2663.9400 2393.9600 ;
        RECT 2673.8800 2382.6000 2676.8800 2383.0800 ;
        RECT 2662.3400 2382.6000 2663.9400 2383.0800 ;
        RECT 2617.3400 2415.2400 2618.9400 2415.7200 ;
        RECT 2617.3400 2420.6800 2618.9400 2421.1600 ;
        RECT 2617.3400 2398.9200 2618.9400 2399.4000 ;
        RECT 2617.3400 2404.3600 2618.9400 2404.8400 ;
        RECT 2617.3400 2409.8000 2618.9400 2410.2800 ;
        RECT 2617.3400 2388.0400 2618.9400 2388.5200 ;
        RECT 2617.3400 2393.4800 2618.9400 2393.9600 ;
        RECT 2617.3400 2382.6000 2618.9400 2383.0800 ;
        RECT 2572.3400 2469.6400 2573.9400 2470.1200 ;
        RECT 2572.3400 2475.0800 2573.9400 2475.5600 ;
        RECT 2572.3400 2453.3200 2573.9400 2453.8000 ;
        RECT 2572.3400 2458.7600 2573.9400 2459.2400 ;
        RECT 2572.3400 2464.2000 2573.9400 2464.6800 ;
        RECT 2527.3400 2469.6400 2528.9400 2470.1200 ;
        RECT 2527.3400 2475.0800 2528.9400 2475.5600 ;
        RECT 2527.3400 2453.3200 2528.9400 2453.8000 ;
        RECT 2527.3400 2458.7600 2528.9400 2459.2400 ;
        RECT 2527.3400 2464.2000 2528.9400 2464.6800 ;
        RECT 2572.3400 2442.4400 2573.9400 2442.9200 ;
        RECT 2572.3400 2447.8800 2573.9400 2448.3600 ;
        RECT 2572.3400 2426.1200 2573.9400 2426.6000 ;
        RECT 2572.3400 2431.5600 2573.9400 2432.0400 ;
        RECT 2572.3400 2437.0000 2573.9400 2437.4800 ;
        RECT 2527.3400 2442.4400 2528.9400 2442.9200 ;
        RECT 2527.3400 2447.8800 2528.9400 2448.3600 ;
        RECT 2527.3400 2426.1200 2528.9400 2426.6000 ;
        RECT 2527.3400 2431.5600 2528.9400 2432.0400 ;
        RECT 2527.3400 2437.0000 2528.9400 2437.4800 ;
        RECT 2477.7800 2469.6400 2480.7800 2470.1200 ;
        RECT 2477.7800 2475.0800 2480.7800 2475.5600 ;
        RECT 2477.7800 2458.7600 2480.7800 2459.2400 ;
        RECT 2477.7800 2453.3200 2480.7800 2453.8000 ;
        RECT 2477.7800 2464.2000 2480.7800 2464.6800 ;
        RECT 2477.7800 2442.4400 2480.7800 2442.9200 ;
        RECT 2477.7800 2447.8800 2480.7800 2448.3600 ;
        RECT 2477.7800 2431.5600 2480.7800 2432.0400 ;
        RECT 2477.7800 2426.1200 2480.7800 2426.6000 ;
        RECT 2477.7800 2437.0000 2480.7800 2437.4800 ;
        RECT 2572.3400 2415.2400 2573.9400 2415.7200 ;
        RECT 2572.3400 2420.6800 2573.9400 2421.1600 ;
        RECT 2572.3400 2398.9200 2573.9400 2399.4000 ;
        RECT 2572.3400 2404.3600 2573.9400 2404.8400 ;
        RECT 2572.3400 2409.8000 2573.9400 2410.2800 ;
        RECT 2527.3400 2415.2400 2528.9400 2415.7200 ;
        RECT 2527.3400 2420.6800 2528.9400 2421.1600 ;
        RECT 2527.3400 2398.9200 2528.9400 2399.4000 ;
        RECT 2527.3400 2404.3600 2528.9400 2404.8400 ;
        RECT 2527.3400 2409.8000 2528.9400 2410.2800 ;
        RECT 2572.3400 2393.4800 2573.9400 2393.9600 ;
        RECT 2572.3400 2388.0400 2573.9400 2388.5200 ;
        RECT 2572.3400 2382.6000 2573.9400 2383.0800 ;
        RECT 2527.3400 2393.4800 2528.9400 2393.9600 ;
        RECT 2527.3400 2388.0400 2528.9400 2388.5200 ;
        RECT 2527.3400 2382.6000 2528.9400 2383.0800 ;
        RECT 2477.7800 2415.2400 2480.7800 2415.7200 ;
        RECT 2477.7800 2420.6800 2480.7800 2421.1600 ;
        RECT 2477.7800 2404.3600 2480.7800 2404.8400 ;
        RECT 2477.7800 2398.9200 2480.7800 2399.4000 ;
        RECT 2477.7800 2409.8000 2480.7800 2410.2800 ;
        RECT 2477.7800 2388.0400 2480.7800 2388.5200 ;
        RECT 2477.7800 2393.4800 2480.7800 2393.9600 ;
        RECT 2477.7800 2382.6000 2480.7800 2383.0800 ;
        RECT 2477.7800 2580.7900 2676.8800 2583.7900 ;
        RECT 2477.7800 2375.6900 2676.8800 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 2146.0500 2663.9400 2354.1500 ;
        RECT 2617.3400 2146.0500 2618.9400 2354.1500 ;
        RECT 2572.3400 2146.0500 2573.9400 2354.1500 ;
        RECT 2527.3400 2146.0500 2528.9400 2354.1500 ;
        RECT 2673.8800 2146.0500 2676.8800 2354.1500 ;
        RECT 2477.7800 2146.0500 2480.7800 2354.1500 ;
      LAYER met3 ;
        RECT 2673.8800 2348.8000 2676.8800 2349.2800 ;
        RECT 2662.3400 2348.8000 2663.9400 2349.2800 ;
        RECT 2673.8800 2337.9200 2676.8800 2338.4000 ;
        RECT 2673.8800 2343.3600 2676.8800 2343.8400 ;
        RECT 2662.3400 2337.9200 2663.9400 2338.4000 ;
        RECT 2662.3400 2343.3600 2663.9400 2343.8400 ;
        RECT 2673.8800 2321.6000 2676.8800 2322.0800 ;
        RECT 2673.8800 2327.0400 2676.8800 2327.5200 ;
        RECT 2662.3400 2321.6000 2663.9400 2322.0800 ;
        RECT 2662.3400 2327.0400 2663.9400 2327.5200 ;
        RECT 2673.8800 2310.7200 2676.8800 2311.2000 ;
        RECT 2673.8800 2316.1600 2676.8800 2316.6400 ;
        RECT 2662.3400 2310.7200 2663.9400 2311.2000 ;
        RECT 2662.3400 2316.1600 2663.9400 2316.6400 ;
        RECT 2673.8800 2332.4800 2676.8800 2332.9600 ;
        RECT 2662.3400 2332.4800 2663.9400 2332.9600 ;
        RECT 2617.3400 2337.9200 2618.9400 2338.4000 ;
        RECT 2617.3400 2343.3600 2618.9400 2343.8400 ;
        RECT 2617.3400 2348.8000 2618.9400 2349.2800 ;
        RECT 2617.3400 2321.6000 2618.9400 2322.0800 ;
        RECT 2617.3400 2327.0400 2618.9400 2327.5200 ;
        RECT 2617.3400 2316.1600 2618.9400 2316.6400 ;
        RECT 2617.3400 2310.7200 2618.9400 2311.2000 ;
        RECT 2617.3400 2332.4800 2618.9400 2332.9600 ;
        RECT 2673.8800 2294.4000 2676.8800 2294.8800 ;
        RECT 2673.8800 2299.8400 2676.8800 2300.3200 ;
        RECT 2662.3400 2294.4000 2663.9400 2294.8800 ;
        RECT 2662.3400 2299.8400 2663.9400 2300.3200 ;
        RECT 2673.8800 2278.0800 2676.8800 2278.5600 ;
        RECT 2673.8800 2283.5200 2676.8800 2284.0000 ;
        RECT 2673.8800 2288.9600 2676.8800 2289.4400 ;
        RECT 2662.3400 2278.0800 2663.9400 2278.5600 ;
        RECT 2662.3400 2283.5200 2663.9400 2284.0000 ;
        RECT 2662.3400 2288.9600 2663.9400 2289.4400 ;
        RECT 2673.8800 2267.2000 2676.8800 2267.6800 ;
        RECT 2673.8800 2272.6400 2676.8800 2273.1200 ;
        RECT 2662.3400 2267.2000 2663.9400 2267.6800 ;
        RECT 2662.3400 2272.6400 2663.9400 2273.1200 ;
        RECT 2673.8800 2250.8800 2676.8800 2251.3600 ;
        RECT 2673.8800 2256.3200 2676.8800 2256.8000 ;
        RECT 2673.8800 2261.7600 2676.8800 2262.2400 ;
        RECT 2662.3400 2250.8800 2663.9400 2251.3600 ;
        RECT 2662.3400 2256.3200 2663.9400 2256.8000 ;
        RECT 2662.3400 2261.7600 2663.9400 2262.2400 ;
        RECT 2617.3400 2294.4000 2618.9400 2294.8800 ;
        RECT 2617.3400 2299.8400 2618.9400 2300.3200 ;
        RECT 2617.3400 2278.0800 2618.9400 2278.5600 ;
        RECT 2617.3400 2283.5200 2618.9400 2284.0000 ;
        RECT 2617.3400 2288.9600 2618.9400 2289.4400 ;
        RECT 2617.3400 2267.2000 2618.9400 2267.6800 ;
        RECT 2617.3400 2272.6400 2618.9400 2273.1200 ;
        RECT 2617.3400 2250.8800 2618.9400 2251.3600 ;
        RECT 2617.3400 2256.3200 2618.9400 2256.8000 ;
        RECT 2617.3400 2261.7600 2618.9400 2262.2400 ;
        RECT 2673.8800 2305.2800 2676.8800 2305.7600 ;
        RECT 2617.3400 2305.2800 2618.9400 2305.7600 ;
        RECT 2662.3400 2305.2800 2663.9400 2305.7600 ;
        RECT 2572.3400 2337.9200 2573.9400 2338.4000 ;
        RECT 2572.3400 2343.3600 2573.9400 2343.8400 ;
        RECT 2572.3400 2348.8000 2573.9400 2349.2800 ;
        RECT 2527.3400 2337.9200 2528.9400 2338.4000 ;
        RECT 2527.3400 2343.3600 2528.9400 2343.8400 ;
        RECT 2527.3400 2348.8000 2528.9400 2349.2800 ;
        RECT 2572.3400 2321.6000 2573.9400 2322.0800 ;
        RECT 2572.3400 2327.0400 2573.9400 2327.5200 ;
        RECT 2572.3400 2310.7200 2573.9400 2311.2000 ;
        RECT 2572.3400 2316.1600 2573.9400 2316.6400 ;
        RECT 2527.3400 2321.6000 2528.9400 2322.0800 ;
        RECT 2527.3400 2327.0400 2528.9400 2327.5200 ;
        RECT 2527.3400 2310.7200 2528.9400 2311.2000 ;
        RECT 2527.3400 2316.1600 2528.9400 2316.6400 ;
        RECT 2527.3400 2332.4800 2528.9400 2332.9600 ;
        RECT 2572.3400 2332.4800 2573.9400 2332.9600 ;
        RECT 2477.7800 2348.8000 2480.7800 2349.2800 ;
        RECT 2477.7800 2343.3600 2480.7800 2343.8400 ;
        RECT 2477.7800 2337.9200 2480.7800 2338.4000 ;
        RECT 2477.7800 2327.0400 2480.7800 2327.5200 ;
        RECT 2477.7800 2321.6000 2480.7800 2322.0800 ;
        RECT 2477.7800 2316.1600 2480.7800 2316.6400 ;
        RECT 2477.7800 2310.7200 2480.7800 2311.2000 ;
        RECT 2477.7800 2332.4800 2480.7800 2332.9600 ;
        RECT 2572.3400 2294.4000 2573.9400 2294.8800 ;
        RECT 2572.3400 2299.8400 2573.9400 2300.3200 ;
        RECT 2572.3400 2278.0800 2573.9400 2278.5600 ;
        RECT 2572.3400 2283.5200 2573.9400 2284.0000 ;
        RECT 2572.3400 2288.9600 2573.9400 2289.4400 ;
        RECT 2527.3400 2294.4000 2528.9400 2294.8800 ;
        RECT 2527.3400 2299.8400 2528.9400 2300.3200 ;
        RECT 2527.3400 2278.0800 2528.9400 2278.5600 ;
        RECT 2527.3400 2283.5200 2528.9400 2284.0000 ;
        RECT 2527.3400 2288.9600 2528.9400 2289.4400 ;
        RECT 2572.3400 2267.2000 2573.9400 2267.6800 ;
        RECT 2572.3400 2272.6400 2573.9400 2273.1200 ;
        RECT 2572.3400 2250.8800 2573.9400 2251.3600 ;
        RECT 2572.3400 2256.3200 2573.9400 2256.8000 ;
        RECT 2572.3400 2261.7600 2573.9400 2262.2400 ;
        RECT 2527.3400 2267.2000 2528.9400 2267.6800 ;
        RECT 2527.3400 2272.6400 2528.9400 2273.1200 ;
        RECT 2527.3400 2250.8800 2528.9400 2251.3600 ;
        RECT 2527.3400 2256.3200 2528.9400 2256.8000 ;
        RECT 2527.3400 2261.7600 2528.9400 2262.2400 ;
        RECT 2477.7800 2294.4000 2480.7800 2294.8800 ;
        RECT 2477.7800 2299.8400 2480.7800 2300.3200 ;
        RECT 2477.7800 2283.5200 2480.7800 2284.0000 ;
        RECT 2477.7800 2278.0800 2480.7800 2278.5600 ;
        RECT 2477.7800 2288.9600 2480.7800 2289.4400 ;
        RECT 2477.7800 2267.2000 2480.7800 2267.6800 ;
        RECT 2477.7800 2272.6400 2480.7800 2273.1200 ;
        RECT 2477.7800 2256.3200 2480.7800 2256.8000 ;
        RECT 2477.7800 2250.8800 2480.7800 2251.3600 ;
        RECT 2477.7800 2261.7600 2480.7800 2262.2400 ;
        RECT 2477.7800 2305.2800 2480.7800 2305.7600 ;
        RECT 2527.3400 2305.2800 2528.9400 2305.7600 ;
        RECT 2572.3400 2305.2800 2573.9400 2305.7600 ;
        RECT 2673.8800 2240.0000 2676.8800 2240.4800 ;
        RECT 2673.8800 2245.4400 2676.8800 2245.9200 ;
        RECT 2662.3400 2240.0000 2663.9400 2240.4800 ;
        RECT 2662.3400 2245.4400 2663.9400 2245.9200 ;
        RECT 2673.8800 2223.6800 2676.8800 2224.1600 ;
        RECT 2673.8800 2229.1200 2676.8800 2229.6000 ;
        RECT 2673.8800 2234.5600 2676.8800 2235.0400 ;
        RECT 2662.3400 2223.6800 2663.9400 2224.1600 ;
        RECT 2662.3400 2229.1200 2663.9400 2229.6000 ;
        RECT 2662.3400 2234.5600 2663.9400 2235.0400 ;
        RECT 2673.8800 2212.8000 2676.8800 2213.2800 ;
        RECT 2673.8800 2218.2400 2676.8800 2218.7200 ;
        RECT 2662.3400 2212.8000 2663.9400 2213.2800 ;
        RECT 2662.3400 2218.2400 2663.9400 2218.7200 ;
        RECT 2673.8800 2196.4800 2676.8800 2196.9600 ;
        RECT 2673.8800 2201.9200 2676.8800 2202.4000 ;
        RECT 2673.8800 2207.3600 2676.8800 2207.8400 ;
        RECT 2662.3400 2196.4800 2663.9400 2196.9600 ;
        RECT 2662.3400 2201.9200 2663.9400 2202.4000 ;
        RECT 2662.3400 2207.3600 2663.9400 2207.8400 ;
        RECT 2617.3400 2240.0000 2618.9400 2240.4800 ;
        RECT 2617.3400 2245.4400 2618.9400 2245.9200 ;
        RECT 2617.3400 2223.6800 2618.9400 2224.1600 ;
        RECT 2617.3400 2229.1200 2618.9400 2229.6000 ;
        RECT 2617.3400 2234.5600 2618.9400 2235.0400 ;
        RECT 2617.3400 2212.8000 2618.9400 2213.2800 ;
        RECT 2617.3400 2218.2400 2618.9400 2218.7200 ;
        RECT 2617.3400 2196.4800 2618.9400 2196.9600 ;
        RECT 2617.3400 2201.9200 2618.9400 2202.4000 ;
        RECT 2617.3400 2207.3600 2618.9400 2207.8400 ;
        RECT 2673.8800 2185.6000 2676.8800 2186.0800 ;
        RECT 2673.8800 2191.0400 2676.8800 2191.5200 ;
        RECT 2662.3400 2185.6000 2663.9400 2186.0800 ;
        RECT 2662.3400 2191.0400 2663.9400 2191.5200 ;
        RECT 2673.8800 2169.2800 2676.8800 2169.7600 ;
        RECT 2673.8800 2174.7200 2676.8800 2175.2000 ;
        RECT 2673.8800 2180.1600 2676.8800 2180.6400 ;
        RECT 2662.3400 2169.2800 2663.9400 2169.7600 ;
        RECT 2662.3400 2174.7200 2663.9400 2175.2000 ;
        RECT 2662.3400 2180.1600 2663.9400 2180.6400 ;
        RECT 2673.8800 2158.4000 2676.8800 2158.8800 ;
        RECT 2673.8800 2163.8400 2676.8800 2164.3200 ;
        RECT 2662.3400 2158.4000 2663.9400 2158.8800 ;
        RECT 2662.3400 2163.8400 2663.9400 2164.3200 ;
        RECT 2673.8800 2152.9600 2676.8800 2153.4400 ;
        RECT 2662.3400 2152.9600 2663.9400 2153.4400 ;
        RECT 2617.3400 2185.6000 2618.9400 2186.0800 ;
        RECT 2617.3400 2191.0400 2618.9400 2191.5200 ;
        RECT 2617.3400 2169.2800 2618.9400 2169.7600 ;
        RECT 2617.3400 2174.7200 2618.9400 2175.2000 ;
        RECT 2617.3400 2180.1600 2618.9400 2180.6400 ;
        RECT 2617.3400 2158.4000 2618.9400 2158.8800 ;
        RECT 2617.3400 2163.8400 2618.9400 2164.3200 ;
        RECT 2617.3400 2152.9600 2618.9400 2153.4400 ;
        RECT 2572.3400 2240.0000 2573.9400 2240.4800 ;
        RECT 2572.3400 2245.4400 2573.9400 2245.9200 ;
        RECT 2572.3400 2223.6800 2573.9400 2224.1600 ;
        RECT 2572.3400 2229.1200 2573.9400 2229.6000 ;
        RECT 2572.3400 2234.5600 2573.9400 2235.0400 ;
        RECT 2527.3400 2240.0000 2528.9400 2240.4800 ;
        RECT 2527.3400 2245.4400 2528.9400 2245.9200 ;
        RECT 2527.3400 2223.6800 2528.9400 2224.1600 ;
        RECT 2527.3400 2229.1200 2528.9400 2229.6000 ;
        RECT 2527.3400 2234.5600 2528.9400 2235.0400 ;
        RECT 2572.3400 2212.8000 2573.9400 2213.2800 ;
        RECT 2572.3400 2218.2400 2573.9400 2218.7200 ;
        RECT 2572.3400 2196.4800 2573.9400 2196.9600 ;
        RECT 2572.3400 2201.9200 2573.9400 2202.4000 ;
        RECT 2572.3400 2207.3600 2573.9400 2207.8400 ;
        RECT 2527.3400 2212.8000 2528.9400 2213.2800 ;
        RECT 2527.3400 2218.2400 2528.9400 2218.7200 ;
        RECT 2527.3400 2196.4800 2528.9400 2196.9600 ;
        RECT 2527.3400 2201.9200 2528.9400 2202.4000 ;
        RECT 2527.3400 2207.3600 2528.9400 2207.8400 ;
        RECT 2477.7800 2240.0000 2480.7800 2240.4800 ;
        RECT 2477.7800 2245.4400 2480.7800 2245.9200 ;
        RECT 2477.7800 2229.1200 2480.7800 2229.6000 ;
        RECT 2477.7800 2223.6800 2480.7800 2224.1600 ;
        RECT 2477.7800 2234.5600 2480.7800 2235.0400 ;
        RECT 2477.7800 2212.8000 2480.7800 2213.2800 ;
        RECT 2477.7800 2218.2400 2480.7800 2218.7200 ;
        RECT 2477.7800 2201.9200 2480.7800 2202.4000 ;
        RECT 2477.7800 2196.4800 2480.7800 2196.9600 ;
        RECT 2477.7800 2207.3600 2480.7800 2207.8400 ;
        RECT 2572.3400 2185.6000 2573.9400 2186.0800 ;
        RECT 2572.3400 2191.0400 2573.9400 2191.5200 ;
        RECT 2572.3400 2169.2800 2573.9400 2169.7600 ;
        RECT 2572.3400 2174.7200 2573.9400 2175.2000 ;
        RECT 2572.3400 2180.1600 2573.9400 2180.6400 ;
        RECT 2527.3400 2185.6000 2528.9400 2186.0800 ;
        RECT 2527.3400 2191.0400 2528.9400 2191.5200 ;
        RECT 2527.3400 2169.2800 2528.9400 2169.7600 ;
        RECT 2527.3400 2174.7200 2528.9400 2175.2000 ;
        RECT 2527.3400 2180.1600 2528.9400 2180.6400 ;
        RECT 2572.3400 2163.8400 2573.9400 2164.3200 ;
        RECT 2572.3400 2158.4000 2573.9400 2158.8800 ;
        RECT 2572.3400 2152.9600 2573.9400 2153.4400 ;
        RECT 2527.3400 2163.8400 2528.9400 2164.3200 ;
        RECT 2527.3400 2158.4000 2528.9400 2158.8800 ;
        RECT 2527.3400 2152.9600 2528.9400 2153.4400 ;
        RECT 2477.7800 2185.6000 2480.7800 2186.0800 ;
        RECT 2477.7800 2191.0400 2480.7800 2191.5200 ;
        RECT 2477.7800 2174.7200 2480.7800 2175.2000 ;
        RECT 2477.7800 2169.2800 2480.7800 2169.7600 ;
        RECT 2477.7800 2180.1600 2480.7800 2180.6400 ;
        RECT 2477.7800 2158.4000 2480.7800 2158.8800 ;
        RECT 2477.7800 2163.8400 2480.7800 2164.3200 ;
        RECT 2477.7800 2152.9600 2480.7800 2153.4400 ;
        RECT 2477.7800 2351.1500 2676.8800 2354.1500 ;
        RECT 2477.7800 2146.0500 2676.8800 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 1916.4100 2663.9400 2124.5100 ;
        RECT 2617.3400 1916.4100 2618.9400 2124.5100 ;
        RECT 2572.3400 1916.4100 2573.9400 2124.5100 ;
        RECT 2527.3400 1916.4100 2528.9400 2124.5100 ;
        RECT 2673.8800 1916.4100 2676.8800 2124.5100 ;
        RECT 2477.7800 1916.4100 2480.7800 2124.5100 ;
      LAYER met3 ;
        RECT 2673.8800 2119.1600 2676.8800 2119.6400 ;
        RECT 2662.3400 2119.1600 2663.9400 2119.6400 ;
        RECT 2673.8800 2108.2800 2676.8800 2108.7600 ;
        RECT 2673.8800 2113.7200 2676.8800 2114.2000 ;
        RECT 2662.3400 2108.2800 2663.9400 2108.7600 ;
        RECT 2662.3400 2113.7200 2663.9400 2114.2000 ;
        RECT 2673.8800 2091.9600 2676.8800 2092.4400 ;
        RECT 2673.8800 2097.4000 2676.8800 2097.8800 ;
        RECT 2662.3400 2091.9600 2663.9400 2092.4400 ;
        RECT 2662.3400 2097.4000 2663.9400 2097.8800 ;
        RECT 2673.8800 2081.0800 2676.8800 2081.5600 ;
        RECT 2673.8800 2086.5200 2676.8800 2087.0000 ;
        RECT 2662.3400 2081.0800 2663.9400 2081.5600 ;
        RECT 2662.3400 2086.5200 2663.9400 2087.0000 ;
        RECT 2673.8800 2102.8400 2676.8800 2103.3200 ;
        RECT 2662.3400 2102.8400 2663.9400 2103.3200 ;
        RECT 2617.3400 2108.2800 2618.9400 2108.7600 ;
        RECT 2617.3400 2113.7200 2618.9400 2114.2000 ;
        RECT 2617.3400 2119.1600 2618.9400 2119.6400 ;
        RECT 2617.3400 2091.9600 2618.9400 2092.4400 ;
        RECT 2617.3400 2097.4000 2618.9400 2097.8800 ;
        RECT 2617.3400 2086.5200 2618.9400 2087.0000 ;
        RECT 2617.3400 2081.0800 2618.9400 2081.5600 ;
        RECT 2617.3400 2102.8400 2618.9400 2103.3200 ;
        RECT 2673.8800 2064.7600 2676.8800 2065.2400 ;
        RECT 2673.8800 2070.2000 2676.8800 2070.6800 ;
        RECT 2662.3400 2064.7600 2663.9400 2065.2400 ;
        RECT 2662.3400 2070.2000 2663.9400 2070.6800 ;
        RECT 2673.8800 2048.4400 2676.8800 2048.9200 ;
        RECT 2673.8800 2053.8800 2676.8800 2054.3600 ;
        RECT 2673.8800 2059.3200 2676.8800 2059.8000 ;
        RECT 2662.3400 2048.4400 2663.9400 2048.9200 ;
        RECT 2662.3400 2053.8800 2663.9400 2054.3600 ;
        RECT 2662.3400 2059.3200 2663.9400 2059.8000 ;
        RECT 2673.8800 2037.5600 2676.8800 2038.0400 ;
        RECT 2673.8800 2043.0000 2676.8800 2043.4800 ;
        RECT 2662.3400 2037.5600 2663.9400 2038.0400 ;
        RECT 2662.3400 2043.0000 2663.9400 2043.4800 ;
        RECT 2673.8800 2021.2400 2676.8800 2021.7200 ;
        RECT 2673.8800 2026.6800 2676.8800 2027.1600 ;
        RECT 2673.8800 2032.1200 2676.8800 2032.6000 ;
        RECT 2662.3400 2021.2400 2663.9400 2021.7200 ;
        RECT 2662.3400 2026.6800 2663.9400 2027.1600 ;
        RECT 2662.3400 2032.1200 2663.9400 2032.6000 ;
        RECT 2617.3400 2064.7600 2618.9400 2065.2400 ;
        RECT 2617.3400 2070.2000 2618.9400 2070.6800 ;
        RECT 2617.3400 2048.4400 2618.9400 2048.9200 ;
        RECT 2617.3400 2053.8800 2618.9400 2054.3600 ;
        RECT 2617.3400 2059.3200 2618.9400 2059.8000 ;
        RECT 2617.3400 2037.5600 2618.9400 2038.0400 ;
        RECT 2617.3400 2043.0000 2618.9400 2043.4800 ;
        RECT 2617.3400 2021.2400 2618.9400 2021.7200 ;
        RECT 2617.3400 2026.6800 2618.9400 2027.1600 ;
        RECT 2617.3400 2032.1200 2618.9400 2032.6000 ;
        RECT 2673.8800 2075.6400 2676.8800 2076.1200 ;
        RECT 2617.3400 2075.6400 2618.9400 2076.1200 ;
        RECT 2662.3400 2075.6400 2663.9400 2076.1200 ;
        RECT 2572.3400 2108.2800 2573.9400 2108.7600 ;
        RECT 2572.3400 2113.7200 2573.9400 2114.2000 ;
        RECT 2572.3400 2119.1600 2573.9400 2119.6400 ;
        RECT 2527.3400 2108.2800 2528.9400 2108.7600 ;
        RECT 2527.3400 2113.7200 2528.9400 2114.2000 ;
        RECT 2527.3400 2119.1600 2528.9400 2119.6400 ;
        RECT 2572.3400 2091.9600 2573.9400 2092.4400 ;
        RECT 2572.3400 2097.4000 2573.9400 2097.8800 ;
        RECT 2572.3400 2081.0800 2573.9400 2081.5600 ;
        RECT 2572.3400 2086.5200 2573.9400 2087.0000 ;
        RECT 2527.3400 2091.9600 2528.9400 2092.4400 ;
        RECT 2527.3400 2097.4000 2528.9400 2097.8800 ;
        RECT 2527.3400 2081.0800 2528.9400 2081.5600 ;
        RECT 2527.3400 2086.5200 2528.9400 2087.0000 ;
        RECT 2527.3400 2102.8400 2528.9400 2103.3200 ;
        RECT 2572.3400 2102.8400 2573.9400 2103.3200 ;
        RECT 2477.7800 2119.1600 2480.7800 2119.6400 ;
        RECT 2477.7800 2113.7200 2480.7800 2114.2000 ;
        RECT 2477.7800 2108.2800 2480.7800 2108.7600 ;
        RECT 2477.7800 2097.4000 2480.7800 2097.8800 ;
        RECT 2477.7800 2091.9600 2480.7800 2092.4400 ;
        RECT 2477.7800 2086.5200 2480.7800 2087.0000 ;
        RECT 2477.7800 2081.0800 2480.7800 2081.5600 ;
        RECT 2477.7800 2102.8400 2480.7800 2103.3200 ;
        RECT 2572.3400 2064.7600 2573.9400 2065.2400 ;
        RECT 2572.3400 2070.2000 2573.9400 2070.6800 ;
        RECT 2572.3400 2048.4400 2573.9400 2048.9200 ;
        RECT 2572.3400 2053.8800 2573.9400 2054.3600 ;
        RECT 2572.3400 2059.3200 2573.9400 2059.8000 ;
        RECT 2527.3400 2064.7600 2528.9400 2065.2400 ;
        RECT 2527.3400 2070.2000 2528.9400 2070.6800 ;
        RECT 2527.3400 2048.4400 2528.9400 2048.9200 ;
        RECT 2527.3400 2053.8800 2528.9400 2054.3600 ;
        RECT 2527.3400 2059.3200 2528.9400 2059.8000 ;
        RECT 2572.3400 2037.5600 2573.9400 2038.0400 ;
        RECT 2572.3400 2043.0000 2573.9400 2043.4800 ;
        RECT 2572.3400 2021.2400 2573.9400 2021.7200 ;
        RECT 2572.3400 2026.6800 2573.9400 2027.1600 ;
        RECT 2572.3400 2032.1200 2573.9400 2032.6000 ;
        RECT 2527.3400 2037.5600 2528.9400 2038.0400 ;
        RECT 2527.3400 2043.0000 2528.9400 2043.4800 ;
        RECT 2527.3400 2021.2400 2528.9400 2021.7200 ;
        RECT 2527.3400 2026.6800 2528.9400 2027.1600 ;
        RECT 2527.3400 2032.1200 2528.9400 2032.6000 ;
        RECT 2477.7800 2064.7600 2480.7800 2065.2400 ;
        RECT 2477.7800 2070.2000 2480.7800 2070.6800 ;
        RECT 2477.7800 2053.8800 2480.7800 2054.3600 ;
        RECT 2477.7800 2048.4400 2480.7800 2048.9200 ;
        RECT 2477.7800 2059.3200 2480.7800 2059.8000 ;
        RECT 2477.7800 2037.5600 2480.7800 2038.0400 ;
        RECT 2477.7800 2043.0000 2480.7800 2043.4800 ;
        RECT 2477.7800 2026.6800 2480.7800 2027.1600 ;
        RECT 2477.7800 2021.2400 2480.7800 2021.7200 ;
        RECT 2477.7800 2032.1200 2480.7800 2032.6000 ;
        RECT 2477.7800 2075.6400 2480.7800 2076.1200 ;
        RECT 2527.3400 2075.6400 2528.9400 2076.1200 ;
        RECT 2572.3400 2075.6400 2573.9400 2076.1200 ;
        RECT 2673.8800 2010.3600 2676.8800 2010.8400 ;
        RECT 2673.8800 2015.8000 2676.8800 2016.2800 ;
        RECT 2662.3400 2010.3600 2663.9400 2010.8400 ;
        RECT 2662.3400 2015.8000 2663.9400 2016.2800 ;
        RECT 2673.8800 1994.0400 2676.8800 1994.5200 ;
        RECT 2673.8800 1999.4800 2676.8800 1999.9600 ;
        RECT 2673.8800 2004.9200 2676.8800 2005.4000 ;
        RECT 2662.3400 1994.0400 2663.9400 1994.5200 ;
        RECT 2662.3400 1999.4800 2663.9400 1999.9600 ;
        RECT 2662.3400 2004.9200 2663.9400 2005.4000 ;
        RECT 2673.8800 1983.1600 2676.8800 1983.6400 ;
        RECT 2673.8800 1988.6000 2676.8800 1989.0800 ;
        RECT 2662.3400 1983.1600 2663.9400 1983.6400 ;
        RECT 2662.3400 1988.6000 2663.9400 1989.0800 ;
        RECT 2673.8800 1966.8400 2676.8800 1967.3200 ;
        RECT 2673.8800 1972.2800 2676.8800 1972.7600 ;
        RECT 2673.8800 1977.7200 2676.8800 1978.2000 ;
        RECT 2662.3400 1966.8400 2663.9400 1967.3200 ;
        RECT 2662.3400 1972.2800 2663.9400 1972.7600 ;
        RECT 2662.3400 1977.7200 2663.9400 1978.2000 ;
        RECT 2617.3400 2010.3600 2618.9400 2010.8400 ;
        RECT 2617.3400 2015.8000 2618.9400 2016.2800 ;
        RECT 2617.3400 1994.0400 2618.9400 1994.5200 ;
        RECT 2617.3400 1999.4800 2618.9400 1999.9600 ;
        RECT 2617.3400 2004.9200 2618.9400 2005.4000 ;
        RECT 2617.3400 1983.1600 2618.9400 1983.6400 ;
        RECT 2617.3400 1988.6000 2618.9400 1989.0800 ;
        RECT 2617.3400 1966.8400 2618.9400 1967.3200 ;
        RECT 2617.3400 1972.2800 2618.9400 1972.7600 ;
        RECT 2617.3400 1977.7200 2618.9400 1978.2000 ;
        RECT 2673.8800 1955.9600 2676.8800 1956.4400 ;
        RECT 2673.8800 1961.4000 2676.8800 1961.8800 ;
        RECT 2662.3400 1955.9600 2663.9400 1956.4400 ;
        RECT 2662.3400 1961.4000 2663.9400 1961.8800 ;
        RECT 2673.8800 1939.6400 2676.8800 1940.1200 ;
        RECT 2673.8800 1945.0800 2676.8800 1945.5600 ;
        RECT 2673.8800 1950.5200 2676.8800 1951.0000 ;
        RECT 2662.3400 1939.6400 2663.9400 1940.1200 ;
        RECT 2662.3400 1945.0800 2663.9400 1945.5600 ;
        RECT 2662.3400 1950.5200 2663.9400 1951.0000 ;
        RECT 2673.8800 1928.7600 2676.8800 1929.2400 ;
        RECT 2673.8800 1934.2000 2676.8800 1934.6800 ;
        RECT 2662.3400 1928.7600 2663.9400 1929.2400 ;
        RECT 2662.3400 1934.2000 2663.9400 1934.6800 ;
        RECT 2673.8800 1923.3200 2676.8800 1923.8000 ;
        RECT 2662.3400 1923.3200 2663.9400 1923.8000 ;
        RECT 2617.3400 1955.9600 2618.9400 1956.4400 ;
        RECT 2617.3400 1961.4000 2618.9400 1961.8800 ;
        RECT 2617.3400 1939.6400 2618.9400 1940.1200 ;
        RECT 2617.3400 1945.0800 2618.9400 1945.5600 ;
        RECT 2617.3400 1950.5200 2618.9400 1951.0000 ;
        RECT 2617.3400 1928.7600 2618.9400 1929.2400 ;
        RECT 2617.3400 1934.2000 2618.9400 1934.6800 ;
        RECT 2617.3400 1923.3200 2618.9400 1923.8000 ;
        RECT 2572.3400 2010.3600 2573.9400 2010.8400 ;
        RECT 2572.3400 2015.8000 2573.9400 2016.2800 ;
        RECT 2572.3400 1994.0400 2573.9400 1994.5200 ;
        RECT 2572.3400 1999.4800 2573.9400 1999.9600 ;
        RECT 2572.3400 2004.9200 2573.9400 2005.4000 ;
        RECT 2527.3400 2010.3600 2528.9400 2010.8400 ;
        RECT 2527.3400 2015.8000 2528.9400 2016.2800 ;
        RECT 2527.3400 1994.0400 2528.9400 1994.5200 ;
        RECT 2527.3400 1999.4800 2528.9400 1999.9600 ;
        RECT 2527.3400 2004.9200 2528.9400 2005.4000 ;
        RECT 2572.3400 1983.1600 2573.9400 1983.6400 ;
        RECT 2572.3400 1988.6000 2573.9400 1989.0800 ;
        RECT 2572.3400 1966.8400 2573.9400 1967.3200 ;
        RECT 2572.3400 1972.2800 2573.9400 1972.7600 ;
        RECT 2572.3400 1977.7200 2573.9400 1978.2000 ;
        RECT 2527.3400 1983.1600 2528.9400 1983.6400 ;
        RECT 2527.3400 1988.6000 2528.9400 1989.0800 ;
        RECT 2527.3400 1966.8400 2528.9400 1967.3200 ;
        RECT 2527.3400 1972.2800 2528.9400 1972.7600 ;
        RECT 2527.3400 1977.7200 2528.9400 1978.2000 ;
        RECT 2477.7800 2010.3600 2480.7800 2010.8400 ;
        RECT 2477.7800 2015.8000 2480.7800 2016.2800 ;
        RECT 2477.7800 1999.4800 2480.7800 1999.9600 ;
        RECT 2477.7800 1994.0400 2480.7800 1994.5200 ;
        RECT 2477.7800 2004.9200 2480.7800 2005.4000 ;
        RECT 2477.7800 1983.1600 2480.7800 1983.6400 ;
        RECT 2477.7800 1988.6000 2480.7800 1989.0800 ;
        RECT 2477.7800 1972.2800 2480.7800 1972.7600 ;
        RECT 2477.7800 1966.8400 2480.7800 1967.3200 ;
        RECT 2477.7800 1977.7200 2480.7800 1978.2000 ;
        RECT 2572.3400 1955.9600 2573.9400 1956.4400 ;
        RECT 2572.3400 1961.4000 2573.9400 1961.8800 ;
        RECT 2572.3400 1939.6400 2573.9400 1940.1200 ;
        RECT 2572.3400 1945.0800 2573.9400 1945.5600 ;
        RECT 2572.3400 1950.5200 2573.9400 1951.0000 ;
        RECT 2527.3400 1955.9600 2528.9400 1956.4400 ;
        RECT 2527.3400 1961.4000 2528.9400 1961.8800 ;
        RECT 2527.3400 1939.6400 2528.9400 1940.1200 ;
        RECT 2527.3400 1945.0800 2528.9400 1945.5600 ;
        RECT 2527.3400 1950.5200 2528.9400 1951.0000 ;
        RECT 2572.3400 1934.2000 2573.9400 1934.6800 ;
        RECT 2572.3400 1928.7600 2573.9400 1929.2400 ;
        RECT 2572.3400 1923.3200 2573.9400 1923.8000 ;
        RECT 2527.3400 1934.2000 2528.9400 1934.6800 ;
        RECT 2527.3400 1928.7600 2528.9400 1929.2400 ;
        RECT 2527.3400 1923.3200 2528.9400 1923.8000 ;
        RECT 2477.7800 1955.9600 2480.7800 1956.4400 ;
        RECT 2477.7800 1961.4000 2480.7800 1961.8800 ;
        RECT 2477.7800 1945.0800 2480.7800 1945.5600 ;
        RECT 2477.7800 1939.6400 2480.7800 1940.1200 ;
        RECT 2477.7800 1950.5200 2480.7800 1951.0000 ;
        RECT 2477.7800 1928.7600 2480.7800 1929.2400 ;
        RECT 2477.7800 1934.2000 2480.7800 1934.6800 ;
        RECT 2477.7800 1923.3200 2480.7800 1923.8000 ;
        RECT 2477.7800 2121.5100 2676.8800 2124.5100 ;
        RECT 2477.7800 1916.4100 2676.8800 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 1686.7700 2663.9400 1894.8700 ;
        RECT 2617.3400 1686.7700 2618.9400 1894.8700 ;
        RECT 2572.3400 1686.7700 2573.9400 1894.8700 ;
        RECT 2527.3400 1686.7700 2528.9400 1894.8700 ;
        RECT 2673.8800 1686.7700 2676.8800 1894.8700 ;
        RECT 2477.7800 1686.7700 2480.7800 1894.8700 ;
      LAYER met3 ;
        RECT 2673.8800 1889.5200 2676.8800 1890.0000 ;
        RECT 2662.3400 1889.5200 2663.9400 1890.0000 ;
        RECT 2673.8800 1878.6400 2676.8800 1879.1200 ;
        RECT 2673.8800 1884.0800 2676.8800 1884.5600 ;
        RECT 2662.3400 1878.6400 2663.9400 1879.1200 ;
        RECT 2662.3400 1884.0800 2663.9400 1884.5600 ;
        RECT 2673.8800 1862.3200 2676.8800 1862.8000 ;
        RECT 2673.8800 1867.7600 2676.8800 1868.2400 ;
        RECT 2662.3400 1862.3200 2663.9400 1862.8000 ;
        RECT 2662.3400 1867.7600 2663.9400 1868.2400 ;
        RECT 2673.8800 1851.4400 2676.8800 1851.9200 ;
        RECT 2673.8800 1856.8800 2676.8800 1857.3600 ;
        RECT 2662.3400 1851.4400 2663.9400 1851.9200 ;
        RECT 2662.3400 1856.8800 2663.9400 1857.3600 ;
        RECT 2673.8800 1873.2000 2676.8800 1873.6800 ;
        RECT 2662.3400 1873.2000 2663.9400 1873.6800 ;
        RECT 2617.3400 1878.6400 2618.9400 1879.1200 ;
        RECT 2617.3400 1884.0800 2618.9400 1884.5600 ;
        RECT 2617.3400 1889.5200 2618.9400 1890.0000 ;
        RECT 2617.3400 1862.3200 2618.9400 1862.8000 ;
        RECT 2617.3400 1867.7600 2618.9400 1868.2400 ;
        RECT 2617.3400 1856.8800 2618.9400 1857.3600 ;
        RECT 2617.3400 1851.4400 2618.9400 1851.9200 ;
        RECT 2617.3400 1873.2000 2618.9400 1873.6800 ;
        RECT 2673.8800 1835.1200 2676.8800 1835.6000 ;
        RECT 2673.8800 1840.5600 2676.8800 1841.0400 ;
        RECT 2662.3400 1835.1200 2663.9400 1835.6000 ;
        RECT 2662.3400 1840.5600 2663.9400 1841.0400 ;
        RECT 2673.8800 1818.8000 2676.8800 1819.2800 ;
        RECT 2673.8800 1824.2400 2676.8800 1824.7200 ;
        RECT 2673.8800 1829.6800 2676.8800 1830.1600 ;
        RECT 2662.3400 1818.8000 2663.9400 1819.2800 ;
        RECT 2662.3400 1824.2400 2663.9400 1824.7200 ;
        RECT 2662.3400 1829.6800 2663.9400 1830.1600 ;
        RECT 2673.8800 1807.9200 2676.8800 1808.4000 ;
        RECT 2673.8800 1813.3600 2676.8800 1813.8400 ;
        RECT 2662.3400 1807.9200 2663.9400 1808.4000 ;
        RECT 2662.3400 1813.3600 2663.9400 1813.8400 ;
        RECT 2673.8800 1791.6000 2676.8800 1792.0800 ;
        RECT 2673.8800 1797.0400 2676.8800 1797.5200 ;
        RECT 2673.8800 1802.4800 2676.8800 1802.9600 ;
        RECT 2662.3400 1791.6000 2663.9400 1792.0800 ;
        RECT 2662.3400 1797.0400 2663.9400 1797.5200 ;
        RECT 2662.3400 1802.4800 2663.9400 1802.9600 ;
        RECT 2617.3400 1835.1200 2618.9400 1835.6000 ;
        RECT 2617.3400 1840.5600 2618.9400 1841.0400 ;
        RECT 2617.3400 1818.8000 2618.9400 1819.2800 ;
        RECT 2617.3400 1824.2400 2618.9400 1824.7200 ;
        RECT 2617.3400 1829.6800 2618.9400 1830.1600 ;
        RECT 2617.3400 1807.9200 2618.9400 1808.4000 ;
        RECT 2617.3400 1813.3600 2618.9400 1813.8400 ;
        RECT 2617.3400 1791.6000 2618.9400 1792.0800 ;
        RECT 2617.3400 1797.0400 2618.9400 1797.5200 ;
        RECT 2617.3400 1802.4800 2618.9400 1802.9600 ;
        RECT 2673.8800 1846.0000 2676.8800 1846.4800 ;
        RECT 2617.3400 1846.0000 2618.9400 1846.4800 ;
        RECT 2662.3400 1846.0000 2663.9400 1846.4800 ;
        RECT 2572.3400 1878.6400 2573.9400 1879.1200 ;
        RECT 2572.3400 1884.0800 2573.9400 1884.5600 ;
        RECT 2572.3400 1889.5200 2573.9400 1890.0000 ;
        RECT 2527.3400 1878.6400 2528.9400 1879.1200 ;
        RECT 2527.3400 1884.0800 2528.9400 1884.5600 ;
        RECT 2527.3400 1889.5200 2528.9400 1890.0000 ;
        RECT 2572.3400 1862.3200 2573.9400 1862.8000 ;
        RECT 2572.3400 1867.7600 2573.9400 1868.2400 ;
        RECT 2572.3400 1851.4400 2573.9400 1851.9200 ;
        RECT 2572.3400 1856.8800 2573.9400 1857.3600 ;
        RECT 2527.3400 1862.3200 2528.9400 1862.8000 ;
        RECT 2527.3400 1867.7600 2528.9400 1868.2400 ;
        RECT 2527.3400 1851.4400 2528.9400 1851.9200 ;
        RECT 2527.3400 1856.8800 2528.9400 1857.3600 ;
        RECT 2527.3400 1873.2000 2528.9400 1873.6800 ;
        RECT 2572.3400 1873.2000 2573.9400 1873.6800 ;
        RECT 2477.7800 1889.5200 2480.7800 1890.0000 ;
        RECT 2477.7800 1884.0800 2480.7800 1884.5600 ;
        RECT 2477.7800 1878.6400 2480.7800 1879.1200 ;
        RECT 2477.7800 1867.7600 2480.7800 1868.2400 ;
        RECT 2477.7800 1862.3200 2480.7800 1862.8000 ;
        RECT 2477.7800 1856.8800 2480.7800 1857.3600 ;
        RECT 2477.7800 1851.4400 2480.7800 1851.9200 ;
        RECT 2477.7800 1873.2000 2480.7800 1873.6800 ;
        RECT 2572.3400 1835.1200 2573.9400 1835.6000 ;
        RECT 2572.3400 1840.5600 2573.9400 1841.0400 ;
        RECT 2572.3400 1818.8000 2573.9400 1819.2800 ;
        RECT 2572.3400 1824.2400 2573.9400 1824.7200 ;
        RECT 2572.3400 1829.6800 2573.9400 1830.1600 ;
        RECT 2527.3400 1835.1200 2528.9400 1835.6000 ;
        RECT 2527.3400 1840.5600 2528.9400 1841.0400 ;
        RECT 2527.3400 1818.8000 2528.9400 1819.2800 ;
        RECT 2527.3400 1824.2400 2528.9400 1824.7200 ;
        RECT 2527.3400 1829.6800 2528.9400 1830.1600 ;
        RECT 2572.3400 1807.9200 2573.9400 1808.4000 ;
        RECT 2572.3400 1813.3600 2573.9400 1813.8400 ;
        RECT 2572.3400 1791.6000 2573.9400 1792.0800 ;
        RECT 2572.3400 1797.0400 2573.9400 1797.5200 ;
        RECT 2572.3400 1802.4800 2573.9400 1802.9600 ;
        RECT 2527.3400 1807.9200 2528.9400 1808.4000 ;
        RECT 2527.3400 1813.3600 2528.9400 1813.8400 ;
        RECT 2527.3400 1791.6000 2528.9400 1792.0800 ;
        RECT 2527.3400 1797.0400 2528.9400 1797.5200 ;
        RECT 2527.3400 1802.4800 2528.9400 1802.9600 ;
        RECT 2477.7800 1835.1200 2480.7800 1835.6000 ;
        RECT 2477.7800 1840.5600 2480.7800 1841.0400 ;
        RECT 2477.7800 1824.2400 2480.7800 1824.7200 ;
        RECT 2477.7800 1818.8000 2480.7800 1819.2800 ;
        RECT 2477.7800 1829.6800 2480.7800 1830.1600 ;
        RECT 2477.7800 1807.9200 2480.7800 1808.4000 ;
        RECT 2477.7800 1813.3600 2480.7800 1813.8400 ;
        RECT 2477.7800 1797.0400 2480.7800 1797.5200 ;
        RECT 2477.7800 1791.6000 2480.7800 1792.0800 ;
        RECT 2477.7800 1802.4800 2480.7800 1802.9600 ;
        RECT 2477.7800 1846.0000 2480.7800 1846.4800 ;
        RECT 2527.3400 1846.0000 2528.9400 1846.4800 ;
        RECT 2572.3400 1846.0000 2573.9400 1846.4800 ;
        RECT 2673.8800 1780.7200 2676.8800 1781.2000 ;
        RECT 2673.8800 1786.1600 2676.8800 1786.6400 ;
        RECT 2662.3400 1780.7200 2663.9400 1781.2000 ;
        RECT 2662.3400 1786.1600 2663.9400 1786.6400 ;
        RECT 2673.8800 1764.4000 2676.8800 1764.8800 ;
        RECT 2673.8800 1769.8400 2676.8800 1770.3200 ;
        RECT 2673.8800 1775.2800 2676.8800 1775.7600 ;
        RECT 2662.3400 1764.4000 2663.9400 1764.8800 ;
        RECT 2662.3400 1769.8400 2663.9400 1770.3200 ;
        RECT 2662.3400 1775.2800 2663.9400 1775.7600 ;
        RECT 2673.8800 1753.5200 2676.8800 1754.0000 ;
        RECT 2673.8800 1758.9600 2676.8800 1759.4400 ;
        RECT 2662.3400 1753.5200 2663.9400 1754.0000 ;
        RECT 2662.3400 1758.9600 2663.9400 1759.4400 ;
        RECT 2673.8800 1737.2000 2676.8800 1737.6800 ;
        RECT 2673.8800 1742.6400 2676.8800 1743.1200 ;
        RECT 2673.8800 1748.0800 2676.8800 1748.5600 ;
        RECT 2662.3400 1737.2000 2663.9400 1737.6800 ;
        RECT 2662.3400 1742.6400 2663.9400 1743.1200 ;
        RECT 2662.3400 1748.0800 2663.9400 1748.5600 ;
        RECT 2617.3400 1780.7200 2618.9400 1781.2000 ;
        RECT 2617.3400 1786.1600 2618.9400 1786.6400 ;
        RECT 2617.3400 1764.4000 2618.9400 1764.8800 ;
        RECT 2617.3400 1769.8400 2618.9400 1770.3200 ;
        RECT 2617.3400 1775.2800 2618.9400 1775.7600 ;
        RECT 2617.3400 1753.5200 2618.9400 1754.0000 ;
        RECT 2617.3400 1758.9600 2618.9400 1759.4400 ;
        RECT 2617.3400 1737.2000 2618.9400 1737.6800 ;
        RECT 2617.3400 1742.6400 2618.9400 1743.1200 ;
        RECT 2617.3400 1748.0800 2618.9400 1748.5600 ;
        RECT 2673.8800 1726.3200 2676.8800 1726.8000 ;
        RECT 2673.8800 1731.7600 2676.8800 1732.2400 ;
        RECT 2662.3400 1726.3200 2663.9400 1726.8000 ;
        RECT 2662.3400 1731.7600 2663.9400 1732.2400 ;
        RECT 2673.8800 1710.0000 2676.8800 1710.4800 ;
        RECT 2673.8800 1715.4400 2676.8800 1715.9200 ;
        RECT 2673.8800 1720.8800 2676.8800 1721.3600 ;
        RECT 2662.3400 1710.0000 2663.9400 1710.4800 ;
        RECT 2662.3400 1715.4400 2663.9400 1715.9200 ;
        RECT 2662.3400 1720.8800 2663.9400 1721.3600 ;
        RECT 2673.8800 1699.1200 2676.8800 1699.6000 ;
        RECT 2673.8800 1704.5600 2676.8800 1705.0400 ;
        RECT 2662.3400 1699.1200 2663.9400 1699.6000 ;
        RECT 2662.3400 1704.5600 2663.9400 1705.0400 ;
        RECT 2673.8800 1693.6800 2676.8800 1694.1600 ;
        RECT 2662.3400 1693.6800 2663.9400 1694.1600 ;
        RECT 2617.3400 1726.3200 2618.9400 1726.8000 ;
        RECT 2617.3400 1731.7600 2618.9400 1732.2400 ;
        RECT 2617.3400 1710.0000 2618.9400 1710.4800 ;
        RECT 2617.3400 1715.4400 2618.9400 1715.9200 ;
        RECT 2617.3400 1720.8800 2618.9400 1721.3600 ;
        RECT 2617.3400 1699.1200 2618.9400 1699.6000 ;
        RECT 2617.3400 1704.5600 2618.9400 1705.0400 ;
        RECT 2617.3400 1693.6800 2618.9400 1694.1600 ;
        RECT 2572.3400 1780.7200 2573.9400 1781.2000 ;
        RECT 2572.3400 1786.1600 2573.9400 1786.6400 ;
        RECT 2572.3400 1764.4000 2573.9400 1764.8800 ;
        RECT 2572.3400 1769.8400 2573.9400 1770.3200 ;
        RECT 2572.3400 1775.2800 2573.9400 1775.7600 ;
        RECT 2527.3400 1780.7200 2528.9400 1781.2000 ;
        RECT 2527.3400 1786.1600 2528.9400 1786.6400 ;
        RECT 2527.3400 1764.4000 2528.9400 1764.8800 ;
        RECT 2527.3400 1769.8400 2528.9400 1770.3200 ;
        RECT 2527.3400 1775.2800 2528.9400 1775.7600 ;
        RECT 2572.3400 1753.5200 2573.9400 1754.0000 ;
        RECT 2572.3400 1758.9600 2573.9400 1759.4400 ;
        RECT 2572.3400 1737.2000 2573.9400 1737.6800 ;
        RECT 2572.3400 1742.6400 2573.9400 1743.1200 ;
        RECT 2572.3400 1748.0800 2573.9400 1748.5600 ;
        RECT 2527.3400 1753.5200 2528.9400 1754.0000 ;
        RECT 2527.3400 1758.9600 2528.9400 1759.4400 ;
        RECT 2527.3400 1737.2000 2528.9400 1737.6800 ;
        RECT 2527.3400 1742.6400 2528.9400 1743.1200 ;
        RECT 2527.3400 1748.0800 2528.9400 1748.5600 ;
        RECT 2477.7800 1780.7200 2480.7800 1781.2000 ;
        RECT 2477.7800 1786.1600 2480.7800 1786.6400 ;
        RECT 2477.7800 1769.8400 2480.7800 1770.3200 ;
        RECT 2477.7800 1764.4000 2480.7800 1764.8800 ;
        RECT 2477.7800 1775.2800 2480.7800 1775.7600 ;
        RECT 2477.7800 1753.5200 2480.7800 1754.0000 ;
        RECT 2477.7800 1758.9600 2480.7800 1759.4400 ;
        RECT 2477.7800 1742.6400 2480.7800 1743.1200 ;
        RECT 2477.7800 1737.2000 2480.7800 1737.6800 ;
        RECT 2477.7800 1748.0800 2480.7800 1748.5600 ;
        RECT 2572.3400 1726.3200 2573.9400 1726.8000 ;
        RECT 2572.3400 1731.7600 2573.9400 1732.2400 ;
        RECT 2572.3400 1710.0000 2573.9400 1710.4800 ;
        RECT 2572.3400 1715.4400 2573.9400 1715.9200 ;
        RECT 2572.3400 1720.8800 2573.9400 1721.3600 ;
        RECT 2527.3400 1726.3200 2528.9400 1726.8000 ;
        RECT 2527.3400 1731.7600 2528.9400 1732.2400 ;
        RECT 2527.3400 1710.0000 2528.9400 1710.4800 ;
        RECT 2527.3400 1715.4400 2528.9400 1715.9200 ;
        RECT 2527.3400 1720.8800 2528.9400 1721.3600 ;
        RECT 2572.3400 1704.5600 2573.9400 1705.0400 ;
        RECT 2572.3400 1699.1200 2573.9400 1699.6000 ;
        RECT 2572.3400 1693.6800 2573.9400 1694.1600 ;
        RECT 2527.3400 1704.5600 2528.9400 1705.0400 ;
        RECT 2527.3400 1699.1200 2528.9400 1699.6000 ;
        RECT 2527.3400 1693.6800 2528.9400 1694.1600 ;
        RECT 2477.7800 1726.3200 2480.7800 1726.8000 ;
        RECT 2477.7800 1731.7600 2480.7800 1732.2400 ;
        RECT 2477.7800 1715.4400 2480.7800 1715.9200 ;
        RECT 2477.7800 1710.0000 2480.7800 1710.4800 ;
        RECT 2477.7800 1720.8800 2480.7800 1721.3600 ;
        RECT 2477.7800 1699.1200 2480.7800 1699.6000 ;
        RECT 2477.7800 1704.5600 2480.7800 1705.0400 ;
        RECT 2477.7800 1693.6800 2480.7800 1694.1600 ;
        RECT 2477.7800 1891.8700 2676.8800 1894.8700 ;
        RECT 2477.7800 1686.7700 2676.8800 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 1457.1300 2663.9400 1665.2300 ;
        RECT 2617.3400 1457.1300 2618.9400 1665.2300 ;
        RECT 2572.3400 1457.1300 2573.9400 1665.2300 ;
        RECT 2527.3400 1457.1300 2528.9400 1665.2300 ;
        RECT 2673.8800 1457.1300 2676.8800 1665.2300 ;
        RECT 2477.7800 1457.1300 2480.7800 1665.2300 ;
      LAYER met3 ;
        RECT 2673.8800 1659.8800 2676.8800 1660.3600 ;
        RECT 2662.3400 1659.8800 2663.9400 1660.3600 ;
        RECT 2673.8800 1649.0000 2676.8800 1649.4800 ;
        RECT 2673.8800 1654.4400 2676.8800 1654.9200 ;
        RECT 2662.3400 1649.0000 2663.9400 1649.4800 ;
        RECT 2662.3400 1654.4400 2663.9400 1654.9200 ;
        RECT 2673.8800 1632.6800 2676.8800 1633.1600 ;
        RECT 2673.8800 1638.1200 2676.8800 1638.6000 ;
        RECT 2662.3400 1632.6800 2663.9400 1633.1600 ;
        RECT 2662.3400 1638.1200 2663.9400 1638.6000 ;
        RECT 2673.8800 1621.8000 2676.8800 1622.2800 ;
        RECT 2673.8800 1627.2400 2676.8800 1627.7200 ;
        RECT 2662.3400 1621.8000 2663.9400 1622.2800 ;
        RECT 2662.3400 1627.2400 2663.9400 1627.7200 ;
        RECT 2673.8800 1643.5600 2676.8800 1644.0400 ;
        RECT 2662.3400 1643.5600 2663.9400 1644.0400 ;
        RECT 2617.3400 1649.0000 2618.9400 1649.4800 ;
        RECT 2617.3400 1654.4400 2618.9400 1654.9200 ;
        RECT 2617.3400 1659.8800 2618.9400 1660.3600 ;
        RECT 2617.3400 1632.6800 2618.9400 1633.1600 ;
        RECT 2617.3400 1638.1200 2618.9400 1638.6000 ;
        RECT 2617.3400 1627.2400 2618.9400 1627.7200 ;
        RECT 2617.3400 1621.8000 2618.9400 1622.2800 ;
        RECT 2617.3400 1643.5600 2618.9400 1644.0400 ;
        RECT 2673.8800 1605.4800 2676.8800 1605.9600 ;
        RECT 2673.8800 1610.9200 2676.8800 1611.4000 ;
        RECT 2662.3400 1605.4800 2663.9400 1605.9600 ;
        RECT 2662.3400 1610.9200 2663.9400 1611.4000 ;
        RECT 2673.8800 1589.1600 2676.8800 1589.6400 ;
        RECT 2673.8800 1594.6000 2676.8800 1595.0800 ;
        RECT 2673.8800 1600.0400 2676.8800 1600.5200 ;
        RECT 2662.3400 1589.1600 2663.9400 1589.6400 ;
        RECT 2662.3400 1594.6000 2663.9400 1595.0800 ;
        RECT 2662.3400 1600.0400 2663.9400 1600.5200 ;
        RECT 2673.8800 1578.2800 2676.8800 1578.7600 ;
        RECT 2673.8800 1583.7200 2676.8800 1584.2000 ;
        RECT 2662.3400 1578.2800 2663.9400 1578.7600 ;
        RECT 2662.3400 1583.7200 2663.9400 1584.2000 ;
        RECT 2673.8800 1561.9600 2676.8800 1562.4400 ;
        RECT 2673.8800 1567.4000 2676.8800 1567.8800 ;
        RECT 2673.8800 1572.8400 2676.8800 1573.3200 ;
        RECT 2662.3400 1561.9600 2663.9400 1562.4400 ;
        RECT 2662.3400 1567.4000 2663.9400 1567.8800 ;
        RECT 2662.3400 1572.8400 2663.9400 1573.3200 ;
        RECT 2617.3400 1605.4800 2618.9400 1605.9600 ;
        RECT 2617.3400 1610.9200 2618.9400 1611.4000 ;
        RECT 2617.3400 1589.1600 2618.9400 1589.6400 ;
        RECT 2617.3400 1594.6000 2618.9400 1595.0800 ;
        RECT 2617.3400 1600.0400 2618.9400 1600.5200 ;
        RECT 2617.3400 1578.2800 2618.9400 1578.7600 ;
        RECT 2617.3400 1583.7200 2618.9400 1584.2000 ;
        RECT 2617.3400 1561.9600 2618.9400 1562.4400 ;
        RECT 2617.3400 1567.4000 2618.9400 1567.8800 ;
        RECT 2617.3400 1572.8400 2618.9400 1573.3200 ;
        RECT 2673.8800 1616.3600 2676.8800 1616.8400 ;
        RECT 2617.3400 1616.3600 2618.9400 1616.8400 ;
        RECT 2662.3400 1616.3600 2663.9400 1616.8400 ;
        RECT 2572.3400 1649.0000 2573.9400 1649.4800 ;
        RECT 2572.3400 1654.4400 2573.9400 1654.9200 ;
        RECT 2572.3400 1659.8800 2573.9400 1660.3600 ;
        RECT 2527.3400 1649.0000 2528.9400 1649.4800 ;
        RECT 2527.3400 1654.4400 2528.9400 1654.9200 ;
        RECT 2527.3400 1659.8800 2528.9400 1660.3600 ;
        RECT 2572.3400 1632.6800 2573.9400 1633.1600 ;
        RECT 2572.3400 1638.1200 2573.9400 1638.6000 ;
        RECT 2572.3400 1621.8000 2573.9400 1622.2800 ;
        RECT 2572.3400 1627.2400 2573.9400 1627.7200 ;
        RECT 2527.3400 1632.6800 2528.9400 1633.1600 ;
        RECT 2527.3400 1638.1200 2528.9400 1638.6000 ;
        RECT 2527.3400 1621.8000 2528.9400 1622.2800 ;
        RECT 2527.3400 1627.2400 2528.9400 1627.7200 ;
        RECT 2527.3400 1643.5600 2528.9400 1644.0400 ;
        RECT 2572.3400 1643.5600 2573.9400 1644.0400 ;
        RECT 2477.7800 1659.8800 2480.7800 1660.3600 ;
        RECT 2477.7800 1654.4400 2480.7800 1654.9200 ;
        RECT 2477.7800 1649.0000 2480.7800 1649.4800 ;
        RECT 2477.7800 1638.1200 2480.7800 1638.6000 ;
        RECT 2477.7800 1632.6800 2480.7800 1633.1600 ;
        RECT 2477.7800 1627.2400 2480.7800 1627.7200 ;
        RECT 2477.7800 1621.8000 2480.7800 1622.2800 ;
        RECT 2477.7800 1643.5600 2480.7800 1644.0400 ;
        RECT 2572.3400 1605.4800 2573.9400 1605.9600 ;
        RECT 2572.3400 1610.9200 2573.9400 1611.4000 ;
        RECT 2572.3400 1589.1600 2573.9400 1589.6400 ;
        RECT 2572.3400 1594.6000 2573.9400 1595.0800 ;
        RECT 2572.3400 1600.0400 2573.9400 1600.5200 ;
        RECT 2527.3400 1605.4800 2528.9400 1605.9600 ;
        RECT 2527.3400 1610.9200 2528.9400 1611.4000 ;
        RECT 2527.3400 1589.1600 2528.9400 1589.6400 ;
        RECT 2527.3400 1594.6000 2528.9400 1595.0800 ;
        RECT 2527.3400 1600.0400 2528.9400 1600.5200 ;
        RECT 2572.3400 1578.2800 2573.9400 1578.7600 ;
        RECT 2572.3400 1583.7200 2573.9400 1584.2000 ;
        RECT 2572.3400 1561.9600 2573.9400 1562.4400 ;
        RECT 2572.3400 1567.4000 2573.9400 1567.8800 ;
        RECT 2572.3400 1572.8400 2573.9400 1573.3200 ;
        RECT 2527.3400 1578.2800 2528.9400 1578.7600 ;
        RECT 2527.3400 1583.7200 2528.9400 1584.2000 ;
        RECT 2527.3400 1561.9600 2528.9400 1562.4400 ;
        RECT 2527.3400 1567.4000 2528.9400 1567.8800 ;
        RECT 2527.3400 1572.8400 2528.9400 1573.3200 ;
        RECT 2477.7800 1605.4800 2480.7800 1605.9600 ;
        RECT 2477.7800 1610.9200 2480.7800 1611.4000 ;
        RECT 2477.7800 1594.6000 2480.7800 1595.0800 ;
        RECT 2477.7800 1589.1600 2480.7800 1589.6400 ;
        RECT 2477.7800 1600.0400 2480.7800 1600.5200 ;
        RECT 2477.7800 1578.2800 2480.7800 1578.7600 ;
        RECT 2477.7800 1583.7200 2480.7800 1584.2000 ;
        RECT 2477.7800 1567.4000 2480.7800 1567.8800 ;
        RECT 2477.7800 1561.9600 2480.7800 1562.4400 ;
        RECT 2477.7800 1572.8400 2480.7800 1573.3200 ;
        RECT 2477.7800 1616.3600 2480.7800 1616.8400 ;
        RECT 2527.3400 1616.3600 2528.9400 1616.8400 ;
        RECT 2572.3400 1616.3600 2573.9400 1616.8400 ;
        RECT 2673.8800 1551.0800 2676.8800 1551.5600 ;
        RECT 2673.8800 1556.5200 2676.8800 1557.0000 ;
        RECT 2662.3400 1551.0800 2663.9400 1551.5600 ;
        RECT 2662.3400 1556.5200 2663.9400 1557.0000 ;
        RECT 2673.8800 1534.7600 2676.8800 1535.2400 ;
        RECT 2673.8800 1540.2000 2676.8800 1540.6800 ;
        RECT 2673.8800 1545.6400 2676.8800 1546.1200 ;
        RECT 2662.3400 1534.7600 2663.9400 1535.2400 ;
        RECT 2662.3400 1540.2000 2663.9400 1540.6800 ;
        RECT 2662.3400 1545.6400 2663.9400 1546.1200 ;
        RECT 2673.8800 1523.8800 2676.8800 1524.3600 ;
        RECT 2673.8800 1529.3200 2676.8800 1529.8000 ;
        RECT 2662.3400 1523.8800 2663.9400 1524.3600 ;
        RECT 2662.3400 1529.3200 2663.9400 1529.8000 ;
        RECT 2673.8800 1507.5600 2676.8800 1508.0400 ;
        RECT 2673.8800 1513.0000 2676.8800 1513.4800 ;
        RECT 2673.8800 1518.4400 2676.8800 1518.9200 ;
        RECT 2662.3400 1507.5600 2663.9400 1508.0400 ;
        RECT 2662.3400 1513.0000 2663.9400 1513.4800 ;
        RECT 2662.3400 1518.4400 2663.9400 1518.9200 ;
        RECT 2617.3400 1551.0800 2618.9400 1551.5600 ;
        RECT 2617.3400 1556.5200 2618.9400 1557.0000 ;
        RECT 2617.3400 1534.7600 2618.9400 1535.2400 ;
        RECT 2617.3400 1540.2000 2618.9400 1540.6800 ;
        RECT 2617.3400 1545.6400 2618.9400 1546.1200 ;
        RECT 2617.3400 1523.8800 2618.9400 1524.3600 ;
        RECT 2617.3400 1529.3200 2618.9400 1529.8000 ;
        RECT 2617.3400 1507.5600 2618.9400 1508.0400 ;
        RECT 2617.3400 1513.0000 2618.9400 1513.4800 ;
        RECT 2617.3400 1518.4400 2618.9400 1518.9200 ;
        RECT 2673.8800 1496.6800 2676.8800 1497.1600 ;
        RECT 2673.8800 1502.1200 2676.8800 1502.6000 ;
        RECT 2662.3400 1496.6800 2663.9400 1497.1600 ;
        RECT 2662.3400 1502.1200 2663.9400 1502.6000 ;
        RECT 2673.8800 1480.3600 2676.8800 1480.8400 ;
        RECT 2673.8800 1485.8000 2676.8800 1486.2800 ;
        RECT 2673.8800 1491.2400 2676.8800 1491.7200 ;
        RECT 2662.3400 1480.3600 2663.9400 1480.8400 ;
        RECT 2662.3400 1485.8000 2663.9400 1486.2800 ;
        RECT 2662.3400 1491.2400 2663.9400 1491.7200 ;
        RECT 2673.8800 1469.4800 2676.8800 1469.9600 ;
        RECT 2673.8800 1474.9200 2676.8800 1475.4000 ;
        RECT 2662.3400 1469.4800 2663.9400 1469.9600 ;
        RECT 2662.3400 1474.9200 2663.9400 1475.4000 ;
        RECT 2673.8800 1464.0400 2676.8800 1464.5200 ;
        RECT 2662.3400 1464.0400 2663.9400 1464.5200 ;
        RECT 2617.3400 1496.6800 2618.9400 1497.1600 ;
        RECT 2617.3400 1502.1200 2618.9400 1502.6000 ;
        RECT 2617.3400 1480.3600 2618.9400 1480.8400 ;
        RECT 2617.3400 1485.8000 2618.9400 1486.2800 ;
        RECT 2617.3400 1491.2400 2618.9400 1491.7200 ;
        RECT 2617.3400 1469.4800 2618.9400 1469.9600 ;
        RECT 2617.3400 1474.9200 2618.9400 1475.4000 ;
        RECT 2617.3400 1464.0400 2618.9400 1464.5200 ;
        RECT 2572.3400 1551.0800 2573.9400 1551.5600 ;
        RECT 2572.3400 1556.5200 2573.9400 1557.0000 ;
        RECT 2572.3400 1534.7600 2573.9400 1535.2400 ;
        RECT 2572.3400 1540.2000 2573.9400 1540.6800 ;
        RECT 2572.3400 1545.6400 2573.9400 1546.1200 ;
        RECT 2527.3400 1551.0800 2528.9400 1551.5600 ;
        RECT 2527.3400 1556.5200 2528.9400 1557.0000 ;
        RECT 2527.3400 1534.7600 2528.9400 1535.2400 ;
        RECT 2527.3400 1540.2000 2528.9400 1540.6800 ;
        RECT 2527.3400 1545.6400 2528.9400 1546.1200 ;
        RECT 2572.3400 1523.8800 2573.9400 1524.3600 ;
        RECT 2572.3400 1529.3200 2573.9400 1529.8000 ;
        RECT 2572.3400 1507.5600 2573.9400 1508.0400 ;
        RECT 2572.3400 1513.0000 2573.9400 1513.4800 ;
        RECT 2572.3400 1518.4400 2573.9400 1518.9200 ;
        RECT 2527.3400 1523.8800 2528.9400 1524.3600 ;
        RECT 2527.3400 1529.3200 2528.9400 1529.8000 ;
        RECT 2527.3400 1507.5600 2528.9400 1508.0400 ;
        RECT 2527.3400 1513.0000 2528.9400 1513.4800 ;
        RECT 2527.3400 1518.4400 2528.9400 1518.9200 ;
        RECT 2477.7800 1551.0800 2480.7800 1551.5600 ;
        RECT 2477.7800 1556.5200 2480.7800 1557.0000 ;
        RECT 2477.7800 1540.2000 2480.7800 1540.6800 ;
        RECT 2477.7800 1534.7600 2480.7800 1535.2400 ;
        RECT 2477.7800 1545.6400 2480.7800 1546.1200 ;
        RECT 2477.7800 1523.8800 2480.7800 1524.3600 ;
        RECT 2477.7800 1529.3200 2480.7800 1529.8000 ;
        RECT 2477.7800 1513.0000 2480.7800 1513.4800 ;
        RECT 2477.7800 1507.5600 2480.7800 1508.0400 ;
        RECT 2477.7800 1518.4400 2480.7800 1518.9200 ;
        RECT 2572.3400 1496.6800 2573.9400 1497.1600 ;
        RECT 2572.3400 1502.1200 2573.9400 1502.6000 ;
        RECT 2572.3400 1480.3600 2573.9400 1480.8400 ;
        RECT 2572.3400 1485.8000 2573.9400 1486.2800 ;
        RECT 2572.3400 1491.2400 2573.9400 1491.7200 ;
        RECT 2527.3400 1496.6800 2528.9400 1497.1600 ;
        RECT 2527.3400 1502.1200 2528.9400 1502.6000 ;
        RECT 2527.3400 1480.3600 2528.9400 1480.8400 ;
        RECT 2527.3400 1485.8000 2528.9400 1486.2800 ;
        RECT 2527.3400 1491.2400 2528.9400 1491.7200 ;
        RECT 2572.3400 1474.9200 2573.9400 1475.4000 ;
        RECT 2572.3400 1469.4800 2573.9400 1469.9600 ;
        RECT 2572.3400 1464.0400 2573.9400 1464.5200 ;
        RECT 2527.3400 1474.9200 2528.9400 1475.4000 ;
        RECT 2527.3400 1469.4800 2528.9400 1469.9600 ;
        RECT 2527.3400 1464.0400 2528.9400 1464.5200 ;
        RECT 2477.7800 1496.6800 2480.7800 1497.1600 ;
        RECT 2477.7800 1502.1200 2480.7800 1502.6000 ;
        RECT 2477.7800 1485.8000 2480.7800 1486.2800 ;
        RECT 2477.7800 1480.3600 2480.7800 1480.8400 ;
        RECT 2477.7800 1491.2400 2480.7800 1491.7200 ;
        RECT 2477.7800 1469.4800 2480.7800 1469.9600 ;
        RECT 2477.7800 1474.9200 2480.7800 1475.4000 ;
        RECT 2477.7800 1464.0400 2480.7800 1464.5200 ;
        RECT 2477.7800 1662.2300 2676.8800 1665.2300 ;
        RECT 2477.7800 1457.1300 2676.8800 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 1227.4900 2663.9400 1435.5900 ;
        RECT 2617.3400 1227.4900 2618.9400 1435.5900 ;
        RECT 2572.3400 1227.4900 2573.9400 1435.5900 ;
        RECT 2527.3400 1227.4900 2528.9400 1435.5900 ;
        RECT 2673.8800 1227.4900 2676.8800 1435.5900 ;
        RECT 2477.7800 1227.4900 2480.7800 1435.5900 ;
      LAYER met3 ;
        RECT 2673.8800 1430.2400 2676.8800 1430.7200 ;
        RECT 2662.3400 1430.2400 2663.9400 1430.7200 ;
        RECT 2673.8800 1419.3600 2676.8800 1419.8400 ;
        RECT 2673.8800 1424.8000 2676.8800 1425.2800 ;
        RECT 2662.3400 1419.3600 2663.9400 1419.8400 ;
        RECT 2662.3400 1424.8000 2663.9400 1425.2800 ;
        RECT 2673.8800 1403.0400 2676.8800 1403.5200 ;
        RECT 2673.8800 1408.4800 2676.8800 1408.9600 ;
        RECT 2662.3400 1403.0400 2663.9400 1403.5200 ;
        RECT 2662.3400 1408.4800 2663.9400 1408.9600 ;
        RECT 2673.8800 1392.1600 2676.8800 1392.6400 ;
        RECT 2673.8800 1397.6000 2676.8800 1398.0800 ;
        RECT 2662.3400 1392.1600 2663.9400 1392.6400 ;
        RECT 2662.3400 1397.6000 2663.9400 1398.0800 ;
        RECT 2673.8800 1413.9200 2676.8800 1414.4000 ;
        RECT 2662.3400 1413.9200 2663.9400 1414.4000 ;
        RECT 2617.3400 1419.3600 2618.9400 1419.8400 ;
        RECT 2617.3400 1424.8000 2618.9400 1425.2800 ;
        RECT 2617.3400 1430.2400 2618.9400 1430.7200 ;
        RECT 2617.3400 1403.0400 2618.9400 1403.5200 ;
        RECT 2617.3400 1408.4800 2618.9400 1408.9600 ;
        RECT 2617.3400 1397.6000 2618.9400 1398.0800 ;
        RECT 2617.3400 1392.1600 2618.9400 1392.6400 ;
        RECT 2617.3400 1413.9200 2618.9400 1414.4000 ;
        RECT 2673.8800 1375.8400 2676.8800 1376.3200 ;
        RECT 2673.8800 1381.2800 2676.8800 1381.7600 ;
        RECT 2662.3400 1375.8400 2663.9400 1376.3200 ;
        RECT 2662.3400 1381.2800 2663.9400 1381.7600 ;
        RECT 2673.8800 1359.5200 2676.8800 1360.0000 ;
        RECT 2673.8800 1364.9600 2676.8800 1365.4400 ;
        RECT 2673.8800 1370.4000 2676.8800 1370.8800 ;
        RECT 2662.3400 1359.5200 2663.9400 1360.0000 ;
        RECT 2662.3400 1364.9600 2663.9400 1365.4400 ;
        RECT 2662.3400 1370.4000 2663.9400 1370.8800 ;
        RECT 2673.8800 1348.6400 2676.8800 1349.1200 ;
        RECT 2673.8800 1354.0800 2676.8800 1354.5600 ;
        RECT 2662.3400 1348.6400 2663.9400 1349.1200 ;
        RECT 2662.3400 1354.0800 2663.9400 1354.5600 ;
        RECT 2673.8800 1332.3200 2676.8800 1332.8000 ;
        RECT 2673.8800 1337.7600 2676.8800 1338.2400 ;
        RECT 2673.8800 1343.2000 2676.8800 1343.6800 ;
        RECT 2662.3400 1332.3200 2663.9400 1332.8000 ;
        RECT 2662.3400 1337.7600 2663.9400 1338.2400 ;
        RECT 2662.3400 1343.2000 2663.9400 1343.6800 ;
        RECT 2617.3400 1375.8400 2618.9400 1376.3200 ;
        RECT 2617.3400 1381.2800 2618.9400 1381.7600 ;
        RECT 2617.3400 1359.5200 2618.9400 1360.0000 ;
        RECT 2617.3400 1364.9600 2618.9400 1365.4400 ;
        RECT 2617.3400 1370.4000 2618.9400 1370.8800 ;
        RECT 2617.3400 1348.6400 2618.9400 1349.1200 ;
        RECT 2617.3400 1354.0800 2618.9400 1354.5600 ;
        RECT 2617.3400 1332.3200 2618.9400 1332.8000 ;
        RECT 2617.3400 1337.7600 2618.9400 1338.2400 ;
        RECT 2617.3400 1343.2000 2618.9400 1343.6800 ;
        RECT 2673.8800 1386.7200 2676.8800 1387.2000 ;
        RECT 2617.3400 1386.7200 2618.9400 1387.2000 ;
        RECT 2662.3400 1386.7200 2663.9400 1387.2000 ;
        RECT 2572.3400 1419.3600 2573.9400 1419.8400 ;
        RECT 2572.3400 1424.8000 2573.9400 1425.2800 ;
        RECT 2572.3400 1430.2400 2573.9400 1430.7200 ;
        RECT 2527.3400 1419.3600 2528.9400 1419.8400 ;
        RECT 2527.3400 1424.8000 2528.9400 1425.2800 ;
        RECT 2527.3400 1430.2400 2528.9400 1430.7200 ;
        RECT 2572.3400 1403.0400 2573.9400 1403.5200 ;
        RECT 2572.3400 1408.4800 2573.9400 1408.9600 ;
        RECT 2572.3400 1392.1600 2573.9400 1392.6400 ;
        RECT 2572.3400 1397.6000 2573.9400 1398.0800 ;
        RECT 2527.3400 1403.0400 2528.9400 1403.5200 ;
        RECT 2527.3400 1408.4800 2528.9400 1408.9600 ;
        RECT 2527.3400 1392.1600 2528.9400 1392.6400 ;
        RECT 2527.3400 1397.6000 2528.9400 1398.0800 ;
        RECT 2527.3400 1413.9200 2528.9400 1414.4000 ;
        RECT 2572.3400 1413.9200 2573.9400 1414.4000 ;
        RECT 2477.7800 1430.2400 2480.7800 1430.7200 ;
        RECT 2477.7800 1424.8000 2480.7800 1425.2800 ;
        RECT 2477.7800 1419.3600 2480.7800 1419.8400 ;
        RECT 2477.7800 1408.4800 2480.7800 1408.9600 ;
        RECT 2477.7800 1403.0400 2480.7800 1403.5200 ;
        RECT 2477.7800 1397.6000 2480.7800 1398.0800 ;
        RECT 2477.7800 1392.1600 2480.7800 1392.6400 ;
        RECT 2477.7800 1413.9200 2480.7800 1414.4000 ;
        RECT 2572.3400 1375.8400 2573.9400 1376.3200 ;
        RECT 2572.3400 1381.2800 2573.9400 1381.7600 ;
        RECT 2572.3400 1359.5200 2573.9400 1360.0000 ;
        RECT 2572.3400 1364.9600 2573.9400 1365.4400 ;
        RECT 2572.3400 1370.4000 2573.9400 1370.8800 ;
        RECT 2527.3400 1375.8400 2528.9400 1376.3200 ;
        RECT 2527.3400 1381.2800 2528.9400 1381.7600 ;
        RECT 2527.3400 1359.5200 2528.9400 1360.0000 ;
        RECT 2527.3400 1364.9600 2528.9400 1365.4400 ;
        RECT 2527.3400 1370.4000 2528.9400 1370.8800 ;
        RECT 2572.3400 1348.6400 2573.9400 1349.1200 ;
        RECT 2572.3400 1354.0800 2573.9400 1354.5600 ;
        RECT 2572.3400 1332.3200 2573.9400 1332.8000 ;
        RECT 2572.3400 1337.7600 2573.9400 1338.2400 ;
        RECT 2572.3400 1343.2000 2573.9400 1343.6800 ;
        RECT 2527.3400 1348.6400 2528.9400 1349.1200 ;
        RECT 2527.3400 1354.0800 2528.9400 1354.5600 ;
        RECT 2527.3400 1332.3200 2528.9400 1332.8000 ;
        RECT 2527.3400 1337.7600 2528.9400 1338.2400 ;
        RECT 2527.3400 1343.2000 2528.9400 1343.6800 ;
        RECT 2477.7800 1375.8400 2480.7800 1376.3200 ;
        RECT 2477.7800 1381.2800 2480.7800 1381.7600 ;
        RECT 2477.7800 1364.9600 2480.7800 1365.4400 ;
        RECT 2477.7800 1359.5200 2480.7800 1360.0000 ;
        RECT 2477.7800 1370.4000 2480.7800 1370.8800 ;
        RECT 2477.7800 1348.6400 2480.7800 1349.1200 ;
        RECT 2477.7800 1354.0800 2480.7800 1354.5600 ;
        RECT 2477.7800 1337.7600 2480.7800 1338.2400 ;
        RECT 2477.7800 1332.3200 2480.7800 1332.8000 ;
        RECT 2477.7800 1343.2000 2480.7800 1343.6800 ;
        RECT 2477.7800 1386.7200 2480.7800 1387.2000 ;
        RECT 2527.3400 1386.7200 2528.9400 1387.2000 ;
        RECT 2572.3400 1386.7200 2573.9400 1387.2000 ;
        RECT 2673.8800 1321.4400 2676.8800 1321.9200 ;
        RECT 2673.8800 1326.8800 2676.8800 1327.3600 ;
        RECT 2662.3400 1321.4400 2663.9400 1321.9200 ;
        RECT 2662.3400 1326.8800 2663.9400 1327.3600 ;
        RECT 2673.8800 1305.1200 2676.8800 1305.6000 ;
        RECT 2673.8800 1310.5600 2676.8800 1311.0400 ;
        RECT 2673.8800 1316.0000 2676.8800 1316.4800 ;
        RECT 2662.3400 1305.1200 2663.9400 1305.6000 ;
        RECT 2662.3400 1310.5600 2663.9400 1311.0400 ;
        RECT 2662.3400 1316.0000 2663.9400 1316.4800 ;
        RECT 2673.8800 1294.2400 2676.8800 1294.7200 ;
        RECT 2673.8800 1299.6800 2676.8800 1300.1600 ;
        RECT 2662.3400 1294.2400 2663.9400 1294.7200 ;
        RECT 2662.3400 1299.6800 2663.9400 1300.1600 ;
        RECT 2673.8800 1277.9200 2676.8800 1278.4000 ;
        RECT 2673.8800 1283.3600 2676.8800 1283.8400 ;
        RECT 2673.8800 1288.8000 2676.8800 1289.2800 ;
        RECT 2662.3400 1277.9200 2663.9400 1278.4000 ;
        RECT 2662.3400 1283.3600 2663.9400 1283.8400 ;
        RECT 2662.3400 1288.8000 2663.9400 1289.2800 ;
        RECT 2617.3400 1321.4400 2618.9400 1321.9200 ;
        RECT 2617.3400 1326.8800 2618.9400 1327.3600 ;
        RECT 2617.3400 1305.1200 2618.9400 1305.6000 ;
        RECT 2617.3400 1310.5600 2618.9400 1311.0400 ;
        RECT 2617.3400 1316.0000 2618.9400 1316.4800 ;
        RECT 2617.3400 1294.2400 2618.9400 1294.7200 ;
        RECT 2617.3400 1299.6800 2618.9400 1300.1600 ;
        RECT 2617.3400 1277.9200 2618.9400 1278.4000 ;
        RECT 2617.3400 1283.3600 2618.9400 1283.8400 ;
        RECT 2617.3400 1288.8000 2618.9400 1289.2800 ;
        RECT 2673.8800 1267.0400 2676.8800 1267.5200 ;
        RECT 2673.8800 1272.4800 2676.8800 1272.9600 ;
        RECT 2662.3400 1267.0400 2663.9400 1267.5200 ;
        RECT 2662.3400 1272.4800 2663.9400 1272.9600 ;
        RECT 2673.8800 1250.7200 2676.8800 1251.2000 ;
        RECT 2673.8800 1256.1600 2676.8800 1256.6400 ;
        RECT 2673.8800 1261.6000 2676.8800 1262.0800 ;
        RECT 2662.3400 1250.7200 2663.9400 1251.2000 ;
        RECT 2662.3400 1256.1600 2663.9400 1256.6400 ;
        RECT 2662.3400 1261.6000 2663.9400 1262.0800 ;
        RECT 2673.8800 1239.8400 2676.8800 1240.3200 ;
        RECT 2673.8800 1245.2800 2676.8800 1245.7600 ;
        RECT 2662.3400 1239.8400 2663.9400 1240.3200 ;
        RECT 2662.3400 1245.2800 2663.9400 1245.7600 ;
        RECT 2673.8800 1234.4000 2676.8800 1234.8800 ;
        RECT 2662.3400 1234.4000 2663.9400 1234.8800 ;
        RECT 2617.3400 1267.0400 2618.9400 1267.5200 ;
        RECT 2617.3400 1272.4800 2618.9400 1272.9600 ;
        RECT 2617.3400 1250.7200 2618.9400 1251.2000 ;
        RECT 2617.3400 1256.1600 2618.9400 1256.6400 ;
        RECT 2617.3400 1261.6000 2618.9400 1262.0800 ;
        RECT 2617.3400 1239.8400 2618.9400 1240.3200 ;
        RECT 2617.3400 1245.2800 2618.9400 1245.7600 ;
        RECT 2617.3400 1234.4000 2618.9400 1234.8800 ;
        RECT 2572.3400 1321.4400 2573.9400 1321.9200 ;
        RECT 2572.3400 1326.8800 2573.9400 1327.3600 ;
        RECT 2572.3400 1305.1200 2573.9400 1305.6000 ;
        RECT 2572.3400 1310.5600 2573.9400 1311.0400 ;
        RECT 2572.3400 1316.0000 2573.9400 1316.4800 ;
        RECT 2527.3400 1321.4400 2528.9400 1321.9200 ;
        RECT 2527.3400 1326.8800 2528.9400 1327.3600 ;
        RECT 2527.3400 1305.1200 2528.9400 1305.6000 ;
        RECT 2527.3400 1310.5600 2528.9400 1311.0400 ;
        RECT 2527.3400 1316.0000 2528.9400 1316.4800 ;
        RECT 2572.3400 1294.2400 2573.9400 1294.7200 ;
        RECT 2572.3400 1299.6800 2573.9400 1300.1600 ;
        RECT 2572.3400 1277.9200 2573.9400 1278.4000 ;
        RECT 2572.3400 1283.3600 2573.9400 1283.8400 ;
        RECT 2572.3400 1288.8000 2573.9400 1289.2800 ;
        RECT 2527.3400 1294.2400 2528.9400 1294.7200 ;
        RECT 2527.3400 1299.6800 2528.9400 1300.1600 ;
        RECT 2527.3400 1277.9200 2528.9400 1278.4000 ;
        RECT 2527.3400 1283.3600 2528.9400 1283.8400 ;
        RECT 2527.3400 1288.8000 2528.9400 1289.2800 ;
        RECT 2477.7800 1321.4400 2480.7800 1321.9200 ;
        RECT 2477.7800 1326.8800 2480.7800 1327.3600 ;
        RECT 2477.7800 1310.5600 2480.7800 1311.0400 ;
        RECT 2477.7800 1305.1200 2480.7800 1305.6000 ;
        RECT 2477.7800 1316.0000 2480.7800 1316.4800 ;
        RECT 2477.7800 1294.2400 2480.7800 1294.7200 ;
        RECT 2477.7800 1299.6800 2480.7800 1300.1600 ;
        RECT 2477.7800 1283.3600 2480.7800 1283.8400 ;
        RECT 2477.7800 1277.9200 2480.7800 1278.4000 ;
        RECT 2477.7800 1288.8000 2480.7800 1289.2800 ;
        RECT 2572.3400 1267.0400 2573.9400 1267.5200 ;
        RECT 2572.3400 1272.4800 2573.9400 1272.9600 ;
        RECT 2572.3400 1250.7200 2573.9400 1251.2000 ;
        RECT 2572.3400 1256.1600 2573.9400 1256.6400 ;
        RECT 2572.3400 1261.6000 2573.9400 1262.0800 ;
        RECT 2527.3400 1267.0400 2528.9400 1267.5200 ;
        RECT 2527.3400 1272.4800 2528.9400 1272.9600 ;
        RECT 2527.3400 1250.7200 2528.9400 1251.2000 ;
        RECT 2527.3400 1256.1600 2528.9400 1256.6400 ;
        RECT 2527.3400 1261.6000 2528.9400 1262.0800 ;
        RECT 2572.3400 1245.2800 2573.9400 1245.7600 ;
        RECT 2572.3400 1239.8400 2573.9400 1240.3200 ;
        RECT 2572.3400 1234.4000 2573.9400 1234.8800 ;
        RECT 2527.3400 1245.2800 2528.9400 1245.7600 ;
        RECT 2527.3400 1239.8400 2528.9400 1240.3200 ;
        RECT 2527.3400 1234.4000 2528.9400 1234.8800 ;
        RECT 2477.7800 1267.0400 2480.7800 1267.5200 ;
        RECT 2477.7800 1272.4800 2480.7800 1272.9600 ;
        RECT 2477.7800 1256.1600 2480.7800 1256.6400 ;
        RECT 2477.7800 1250.7200 2480.7800 1251.2000 ;
        RECT 2477.7800 1261.6000 2480.7800 1262.0800 ;
        RECT 2477.7800 1239.8400 2480.7800 1240.3200 ;
        RECT 2477.7800 1245.2800 2480.7800 1245.7600 ;
        RECT 2477.7800 1234.4000 2480.7800 1234.8800 ;
        RECT 2477.7800 1432.5900 2676.8800 1435.5900 ;
        RECT 2477.7800 1227.4900 2676.8800 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 997.8500 2663.9400 1205.9500 ;
        RECT 2617.3400 997.8500 2618.9400 1205.9500 ;
        RECT 2572.3400 997.8500 2573.9400 1205.9500 ;
        RECT 2527.3400 997.8500 2528.9400 1205.9500 ;
        RECT 2673.8800 997.8500 2676.8800 1205.9500 ;
        RECT 2477.7800 997.8500 2480.7800 1205.9500 ;
      LAYER met3 ;
        RECT 2673.8800 1200.6000 2676.8800 1201.0800 ;
        RECT 2662.3400 1200.6000 2663.9400 1201.0800 ;
        RECT 2673.8800 1189.7200 2676.8800 1190.2000 ;
        RECT 2673.8800 1195.1600 2676.8800 1195.6400 ;
        RECT 2662.3400 1189.7200 2663.9400 1190.2000 ;
        RECT 2662.3400 1195.1600 2663.9400 1195.6400 ;
        RECT 2673.8800 1173.4000 2676.8800 1173.8800 ;
        RECT 2673.8800 1178.8400 2676.8800 1179.3200 ;
        RECT 2662.3400 1173.4000 2663.9400 1173.8800 ;
        RECT 2662.3400 1178.8400 2663.9400 1179.3200 ;
        RECT 2673.8800 1162.5200 2676.8800 1163.0000 ;
        RECT 2673.8800 1167.9600 2676.8800 1168.4400 ;
        RECT 2662.3400 1162.5200 2663.9400 1163.0000 ;
        RECT 2662.3400 1167.9600 2663.9400 1168.4400 ;
        RECT 2673.8800 1184.2800 2676.8800 1184.7600 ;
        RECT 2662.3400 1184.2800 2663.9400 1184.7600 ;
        RECT 2617.3400 1189.7200 2618.9400 1190.2000 ;
        RECT 2617.3400 1195.1600 2618.9400 1195.6400 ;
        RECT 2617.3400 1200.6000 2618.9400 1201.0800 ;
        RECT 2617.3400 1173.4000 2618.9400 1173.8800 ;
        RECT 2617.3400 1178.8400 2618.9400 1179.3200 ;
        RECT 2617.3400 1167.9600 2618.9400 1168.4400 ;
        RECT 2617.3400 1162.5200 2618.9400 1163.0000 ;
        RECT 2617.3400 1184.2800 2618.9400 1184.7600 ;
        RECT 2673.8800 1146.2000 2676.8800 1146.6800 ;
        RECT 2673.8800 1151.6400 2676.8800 1152.1200 ;
        RECT 2662.3400 1146.2000 2663.9400 1146.6800 ;
        RECT 2662.3400 1151.6400 2663.9400 1152.1200 ;
        RECT 2673.8800 1129.8800 2676.8800 1130.3600 ;
        RECT 2673.8800 1135.3200 2676.8800 1135.8000 ;
        RECT 2673.8800 1140.7600 2676.8800 1141.2400 ;
        RECT 2662.3400 1129.8800 2663.9400 1130.3600 ;
        RECT 2662.3400 1135.3200 2663.9400 1135.8000 ;
        RECT 2662.3400 1140.7600 2663.9400 1141.2400 ;
        RECT 2673.8800 1119.0000 2676.8800 1119.4800 ;
        RECT 2673.8800 1124.4400 2676.8800 1124.9200 ;
        RECT 2662.3400 1119.0000 2663.9400 1119.4800 ;
        RECT 2662.3400 1124.4400 2663.9400 1124.9200 ;
        RECT 2673.8800 1102.6800 2676.8800 1103.1600 ;
        RECT 2673.8800 1108.1200 2676.8800 1108.6000 ;
        RECT 2673.8800 1113.5600 2676.8800 1114.0400 ;
        RECT 2662.3400 1102.6800 2663.9400 1103.1600 ;
        RECT 2662.3400 1108.1200 2663.9400 1108.6000 ;
        RECT 2662.3400 1113.5600 2663.9400 1114.0400 ;
        RECT 2617.3400 1146.2000 2618.9400 1146.6800 ;
        RECT 2617.3400 1151.6400 2618.9400 1152.1200 ;
        RECT 2617.3400 1129.8800 2618.9400 1130.3600 ;
        RECT 2617.3400 1135.3200 2618.9400 1135.8000 ;
        RECT 2617.3400 1140.7600 2618.9400 1141.2400 ;
        RECT 2617.3400 1119.0000 2618.9400 1119.4800 ;
        RECT 2617.3400 1124.4400 2618.9400 1124.9200 ;
        RECT 2617.3400 1102.6800 2618.9400 1103.1600 ;
        RECT 2617.3400 1108.1200 2618.9400 1108.6000 ;
        RECT 2617.3400 1113.5600 2618.9400 1114.0400 ;
        RECT 2673.8800 1157.0800 2676.8800 1157.5600 ;
        RECT 2617.3400 1157.0800 2618.9400 1157.5600 ;
        RECT 2662.3400 1157.0800 2663.9400 1157.5600 ;
        RECT 2572.3400 1189.7200 2573.9400 1190.2000 ;
        RECT 2572.3400 1195.1600 2573.9400 1195.6400 ;
        RECT 2572.3400 1200.6000 2573.9400 1201.0800 ;
        RECT 2527.3400 1189.7200 2528.9400 1190.2000 ;
        RECT 2527.3400 1195.1600 2528.9400 1195.6400 ;
        RECT 2527.3400 1200.6000 2528.9400 1201.0800 ;
        RECT 2572.3400 1173.4000 2573.9400 1173.8800 ;
        RECT 2572.3400 1178.8400 2573.9400 1179.3200 ;
        RECT 2572.3400 1162.5200 2573.9400 1163.0000 ;
        RECT 2572.3400 1167.9600 2573.9400 1168.4400 ;
        RECT 2527.3400 1173.4000 2528.9400 1173.8800 ;
        RECT 2527.3400 1178.8400 2528.9400 1179.3200 ;
        RECT 2527.3400 1162.5200 2528.9400 1163.0000 ;
        RECT 2527.3400 1167.9600 2528.9400 1168.4400 ;
        RECT 2527.3400 1184.2800 2528.9400 1184.7600 ;
        RECT 2572.3400 1184.2800 2573.9400 1184.7600 ;
        RECT 2477.7800 1200.6000 2480.7800 1201.0800 ;
        RECT 2477.7800 1195.1600 2480.7800 1195.6400 ;
        RECT 2477.7800 1189.7200 2480.7800 1190.2000 ;
        RECT 2477.7800 1178.8400 2480.7800 1179.3200 ;
        RECT 2477.7800 1173.4000 2480.7800 1173.8800 ;
        RECT 2477.7800 1167.9600 2480.7800 1168.4400 ;
        RECT 2477.7800 1162.5200 2480.7800 1163.0000 ;
        RECT 2477.7800 1184.2800 2480.7800 1184.7600 ;
        RECT 2572.3400 1146.2000 2573.9400 1146.6800 ;
        RECT 2572.3400 1151.6400 2573.9400 1152.1200 ;
        RECT 2572.3400 1129.8800 2573.9400 1130.3600 ;
        RECT 2572.3400 1135.3200 2573.9400 1135.8000 ;
        RECT 2572.3400 1140.7600 2573.9400 1141.2400 ;
        RECT 2527.3400 1146.2000 2528.9400 1146.6800 ;
        RECT 2527.3400 1151.6400 2528.9400 1152.1200 ;
        RECT 2527.3400 1129.8800 2528.9400 1130.3600 ;
        RECT 2527.3400 1135.3200 2528.9400 1135.8000 ;
        RECT 2527.3400 1140.7600 2528.9400 1141.2400 ;
        RECT 2572.3400 1119.0000 2573.9400 1119.4800 ;
        RECT 2572.3400 1124.4400 2573.9400 1124.9200 ;
        RECT 2572.3400 1102.6800 2573.9400 1103.1600 ;
        RECT 2572.3400 1108.1200 2573.9400 1108.6000 ;
        RECT 2572.3400 1113.5600 2573.9400 1114.0400 ;
        RECT 2527.3400 1119.0000 2528.9400 1119.4800 ;
        RECT 2527.3400 1124.4400 2528.9400 1124.9200 ;
        RECT 2527.3400 1102.6800 2528.9400 1103.1600 ;
        RECT 2527.3400 1108.1200 2528.9400 1108.6000 ;
        RECT 2527.3400 1113.5600 2528.9400 1114.0400 ;
        RECT 2477.7800 1146.2000 2480.7800 1146.6800 ;
        RECT 2477.7800 1151.6400 2480.7800 1152.1200 ;
        RECT 2477.7800 1135.3200 2480.7800 1135.8000 ;
        RECT 2477.7800 1129.8800 2480.7800 1130.3600 ;
        RECT 2477.7800 1140.7600 2480.7800 1141.2400 ;
        RECT 2477.7800 1119.0000 2480.7800 1119.4800 ;
        RECT 2477.7800 1124.4400 2480.7800 1124.9200 ;
        RECT 2477.7800 1108.1200 2480.7800 1108.6000 ;
        RECT 2477.7800 1102.6800 2480.7800 1103.1600 ;
        RECT 2477.7800 1113.5600 2480.7800 1114.0400 ;
        RECT 2477.7800 1157.0800 2480.7800 1157.5600 ;
        RECT 2527.3400 1157.0800 2528.9400 1157.5600 ;
        RECT 2572.3400 1157.0800 2573.9400 1157.5600 ;
        RECT 2673.8800 1091.8000 2676.8800 1092.2800 ;
        RECT 2673.8800 1097.2400 2676.8800 1097.7200 ;
        RECT 2662.3400 1091.8000 2663.9400 1092.2800 ;
        RECT 2662.3400 1097.2400 2663.9400 1097.7200 ;
        RECT 2673.8800 1075.4800 2676.8800 1075.9600 ;
        RECT 2673.8800 1080.9200 2676.8800 1081.4000 ;
        RECT 2673.8800 1086.3600 2676.8800 1086.8400 ;
        RECT 2662.3400 1075.4800 2663.9400 1075.9600 ;
        RECT 2662.3400 1080.9200 2663.9400 1081.4000 ;
        RECT 2662.3400 1086.3600 2663.9400 1086.8400 ;
        RECT 2673.8800 1064.6000 2676.8800 1065.0800 ;
        RECT 2673.8800 1070.0400 2676.8800 1070.5200 ;
        RECT 2662.3400 1064.6000 2663.9400 1065.0800 ;
        RECT 2662.3400 1070.0400 2663.9400 1070.5200 ;
        RECT 2673.8800 1048.2800 2676.8800 1048.7600 ;
        RECT 2673.8800 1053.7200 2676.8800 1054.2000 ;
        RECT 2673.8800 1059.1600 2676.8800 1059.6400 ;
        RECT 2662.3400 1048.2800 2663.9400 1048.7600 ;
        RECT 2662.3400 1053.7200 2663.9400 1054.2000 ;
        RECT 2662.3400 1059.1600 2663.9400 1059.6400 ;
        RECT 2617.3400 1091.8000 2618.9400 1092.2800 ;
        RECT 2617.3400 1097.2400 2618.9400 1097.7200 ;
        RECT 2617.3400 1075.4800 2618.9400 1075.9600 ;
        RECT 2617.3400 1080.9200 2618.9400 1081.4000 ;
        RECT 2617.3400 1086.3600 2618.9400 1086.8400 ;
        RECT 2617.3400 1064.6000 2618.9400 1065.0800 ;
        RECT 2617.3400 1070.0400 2618.9400 1070.5200 ;
        RECT 2617.3400 1048.2800 2618.9400 1048.7600 ;
        RECT 2617.3400 1053.7200 2618.9400 1054.2000 ;
        RECT 2617.3400 1059.1600 2618.9400 1059.6400 ;
        RECT 2673.8800 1037.4000 2676.8800 1037.8800 ;
        RECT 2673.8800 1042.8400 2676.8800 1043.3200 ;
        RECT 2662.3400 1037.4000 2663.9400 1037.8800 ;
        RECT 2662.3400 1042.8400 2663.9400 1043.3200 ;
        RECT 2673.8800 1021.0800 2676.8800 1021.5600 ;
        RECT 2673.8800 1026.5200 2676.8800 1027.0000 ;
        RECT 2673.8800 1031.9600 2676.8800 1032.4400 ;
        RECT 2662.3400 1021.0800 2663.9400 1021.5600 ;
        RECT 2662.3400 1026.5200 2663.9400 1027.0000 ;
        RECT 2662.3400 1031.9600 2663.9400 1032.4400 ;
        RECT 2673.8800 1010.2000 2676.8800 1010.6800 ;
        RECT 2673.8800 1015.6400 2676.8800 1016.1200 ;
        RECT 2662.3400 1010.2000 2663.9400 1010.6800 ;
        RECT 2662.3400 1015.6400 2663.9400 1016.1200 ;
        RECT 2673.8800 1004.7600 2676.8800 1005.2400 ;
        RECT 2662.3400 1004.7600 2663.9400 1005.2400 ;
        RECT 2617.3400 1037.4000 2618.9400 1037.8800 ;
        RECT 2617.3400 1042.8400 2618.9400 1043.3200 ;
        RECT 2617.3400 1021.0800 2618.9400 1021.5600 ;
        RECT 2617.3400 1026.5200 2618.9400 1027.0000 ;
        RECT 2617.3400 1031.9600 2618.9400 1032.4400 ;
        RECT 2617.3400 1010.2000 2618.9400 1010.6800 ;
        RECT 2617.3400 1015.6400 2618.9400 1016.1200 ;
        RECT 2617.3400 1004.7600 2618.9400 1005.2400 ;
        RECT 2572.3400 1091.8000 2573.9400 1092.2800 ;
        RECT 2572.3400 1097.2400 2573.9400 1097.7200 ;
        RECT 2572.3400 1075.4800 2573.9400 1075.9600 ;
        RECT 2572.3400 1080.9200 2573.9400 1081.4000 ;
        RECT 2572.3400 1086.3600 2573.9400 1086.8400 ;
        RECT 2527.3400 1091.8000 2528.9400 1092.2800 ;
        RECT 2527.3400 1097.2400 2528.9400 1097.7200 ;
        RECT 2527.3400 1075.4800 2528.9400 1075.9600 ;
        RECT 2527.3400 1080.9200 2528.9400 1081.4000 ;
        RECT 2527.3400 1086.3600 2528.9400 1086.8400 ;
        RECT 2572.3400 1064.6000 2573.9400 1065.0800 ;
        RECT 2572.3400 1070.0400 2573.9400 1070.5200 ;
        RECT 2572.3400 1048.2800 2573.9400 1048.7600 ;
        RECT 2572.3400 1053.7200 2573.9400 1054.2000 ;
        RECT 2572.3400 1059.1600 2573.9400 1059.6400 ;
        RECT 2527.3400 1064.6000 2528.9400 1065.0800 ;
        RECT 2527.3400 1070.0400 2528.9400 1070.5200 ;
        RECT 2527.3400 1048.2800 2528.9400 1048.7600 ;
        RECT 2527.3400 1053.7200 2528.9400 1054.2000 ;
        RECT 2527.3400 1059.1600 2528.9400 1059.6400 ;
        RECT 2477.7800 1091.8000 2480.7800 1092.2800 ;
        RECT 2477.7800 1097.2400 2480.7800 1097.7200 ;
        RECT 2477.7800 1080.9200 2480.7800 1081.4000 ;
        RECT 2477.7800 1075.4800 2480.7800 1075.9600 ;
        RECT 2477.7800 1086.3600 2480.7800 1086.8400 ;
        RECT 2477.7800 1064.6000 2480.7800 1065.0800 ;
        RECT 2477.7800 1070.0400 2480.7800 1070.5200 ;
        RECT 2477.7800 1053.7200 2480.7800 1054.2000 ;
        RECT 2477.7800 1048.2800 2480.7800 1048.7600 ;
        RECT 2477.7800 1059.1600 2480.7800 1059.6400 ;
        RECT 2572.3400 1037.4000 2573.9400 1037.8800 ;
        RECT 2572.3400 1042.8400 2573.9400 1043.3200 ;
        RECT 2572.3400 1021.0800 2573.9400 1021.5600 ;
        RECT 2572.3400 1026.5200 2573.9400 1027.0000 ;
        RECT 2572.3400 1031.9600 2573.9400 1032.4400 ;
        RECT 2527.3400 1037.4000 2528.9400 1037.8800 ;
        RECT 2527.3400 1042.8400 2528.9400 1043.3200 ;
        RECT 2527.3400 1021.0800 2528.9400 1021.5600 ;
        RECT 2527.3400 1026.5200 2528.9400 1027.0000 ;
        RECT 2527.3400 1031.9600 2528.9400 1032.4400 ;
        RECT 2572.3400 1015.6400 2573.9400 1016.1200 ;
        RECT 2572.3400 1010.2000 2573.9400 1010.6800 ;
        RECT 2572.3400 1004.7600 2573.9400 1005.2400 ;
        RECT 2527.3400 1015.6400 2528.9400 1016.1200 ;
        RECT 2527.3400 1010.2000 2528.9400 1010.6800 ;
        RECT 2527.3400 1004.7600 2528.9400 1005.2400 ;
        RECT 2477.7800 1037.4000 2480.7800 1037.8800 ;
        RECT 2477.7800 1042.8400 2480.7800 1043.3200 ;
        RECT 2477.7800 1026.5200 2480.7800 1027.0000 ;
        RECT 2477.7800 1021.0800 2480.7800 1021.5600 ;
        RECT 2477.7800 1031.9600 2480.7800 1032.4400 ;
        RECT 2477.7800 1010.2000 2480.7800 1010.6800 ;
        RECT 2477.7800 1015.6400 2480.7800 1016.1200 ;
        RECT 2477.7800 1004.7600 2480.7800 1005.2400 ;
        RECT 2477.7800 1202.9500 2676.8800 1205.9500 ;
        RECT 2477.7800 997.8500 2676.8800 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2662.3400 768.2100 2663.9400 976.3100 ;
        RECT 2617.3400 768.2100 2618.9400 976.3100 ;
        RECT 2572.3400 768.2100 2573.9400 976.3100 ;
        RECT 2527.3400 768.2100 2528.9400 976.3100 ;
        RECT 2673.8800 768.2100 2676.8800 976.3100 ;
        RECT 2477.7800 768.2100 2480.7800 976.3100 ;
      LAYER met3 ;
        RECT 2673.8800 970.9600 2676.8800 971.4400 ;
        RECT 2662.3400 970.9600 2663.9400 971.4400 ;
        RECT 2673.8800 960.0800 2676.8800 960.5600 ;
        RECT 2673.8800 965.5200 2676.8800 966.0000 ;
        RECT 2662.3400 960.0800 2663.9400 960.5600 ;
        RECT 2662.3400 965.5200 2663.9400 966.0000 ;
        RECT 2673.8800 943.7600 2676.8800 944.2400 ;
        RECT 2673.8800 949.2000 2676.8800 949.6800 ;
        RECT 2662.3400 943.7600 2663.9400 944.2400 ;
        RECT 2662.3400 949.2000 2663.9400 949.6800 ;
        RECT 2673.8800 932.8800 2676.8800 933.3600 ;
        RECT 2673.8800 938.3200 2676.8800 938.8000 ;
        RECT 2662.3400 932.8800 2663.9400 933.3600 ;
        RECT 2662.3400 938.3200 2663.9400 938.8000 ;
        RECT 2673.8800 954.6400 2676.8800 955.1200 ;
        RECT 2662.3400 954.6400 2663.9400 955.1200 ;
        RECT 2617.3400 960.0800 2618.9400 960.5600 ;
        RECT 2617.3400 965.5200 2618.9400 966.0000 ;
        RECT 2617.3400 970.9600 2618.9400 971.4400 ;
        RECT 2617.3400 943.7600 2618.9400 944.2400 ;
        RECT 2617.3400 949.2000 2618.9400 949.6800 ;
        RECT 2617.3400 938.3200 2618.9400 938.8000 ;
        RECT 2617.3400 932.8800 2618.9400 933.3600 ;
        RECT 2617.3400 954.6400 2618.9400 955.1200 ;
        RECT 2673.8800 916.5600 2676.8800 917.0400 ;
        RECT 2673.8800 922.0000 2676.8800 922.4800 ;
        RECT 2662.3400 916.5600 2663.9400 917.0400 ;
        RECT 2662.3400 922.0000 2663.9400 922.4800 ;
        RECT 2673.8800 900.2400 2676.8800 900.7200 ;
        RECT 2673.8800 905.6800 2676.8800 906.1600 ;
        RECT 2673.8800 911.1200 2676.8800 911.6000 ;
        RECT 2662.3400 900.2400 2663.9400 900.7200 ;
        RECT 2662.3400 905.6800 2663.9400 906.1600 ;
        RECT 2662.3400 911.1200 2663.9400 911.6000 ;
        RECT 2673.8800 889.3600 2676.8800 889.8400 ;
        RECT 2673.8800 894.8000 2676.8800 895.2800 ;
        RECT 2662.3400 889.3600 2663.9400 889.8400 ;
        RECT 2662.3400 894.8000 2663.9400 895.2800 ;
        RECT 2673.8800 873.0400 2676.8800 873.5200 ;
        RECT 2673.8800 878.4800 2676.8800 878.9600 ;
        RECT 2673.8800 883.9200 2676.8800 884.4000 ;
        RECT 2662.3400 873.0400 2663.9400 873.5200 ;
        RECT 2662.3400 878.4800 2663.9400 878.9600 ;
        RECT 2662.3400 883.9200 2663.9400 884.4000 ;
        RECT 2617.3400 916.5600 2618.9400 917.0400 ;
        RECT 2617.3400 922.0000 2618.9400 922.4800 ;
        RECT 2617.3400 900.2400 2618.9400 900.7200 ;
        RECT 2617.3400 905.6800 2618.9400 906.1600 ;
        RECT 2617.3400 911.1200 2618.9400 911.6000 ;
        RECT 2617.3400 889.3600 2618.9400 889.8400 ;
        RECT 2617.3400 894.8000 2618.9400 895.2800 ;
        RECT 2617.3400 873.0400 2618.9400 873.5200 ;
        RECT 2617.3400 878.4800 2618.9400 878.9600 ;
        RECT 2617.3400 883.9200 2618.9400 884.4000 ;
        RECT 2673.8800 927.4400 2676.8800 927.9200 ;
        RECT 2617.3400 927.4400 2618.9400 927.9200 ;
        RECT 2662.3400 927.4400 2663.9400 927.9200 ;
        RECT 2572.3400 960.0800 2573.9400 960.5600 ;
        RECT 2572.3400 965.5200 2573.9400 966.0000 ;
        RECT 2572.3400 970.9600 2573.9400 971.4400 ;
        RECT 2527.3400 960.0800 2528.9400 960.5600 ;
        RECT 2527.3400 965.5200 2528.9400 966.0000 ;
        RECT 2527.3400 970.9600 2528.9400 971.4400 ;
        RECT 2572.3400 943.7600 2573.9400 944.2400 ;
        RECT 2572.3400 949.2000 2573.9400 949.6800 ;
        RECT 2572.3400 932.8800 2573.9400 933.3600 ;
        RECT 2572.3400 938.3200 2573.9400 938.8000 ;
        RECT 2527.3400 943.7600 2528.9400 944.2400 ;
        RECT 2527.3400 949.2000 2528.9400 949.6800 ;
        RECT 2527.3400 932.8800 2528.9400 933.3600 ;
        RECT 2527.3400 938.3200 2528.9400 938.8000 ;
        RECT 2527.3400 954.6400 2528.9400 955.1200 ;
        RECT 2572.3400 954.6400 2573.9400 955.1200 ;
        RECT 2477.7800 970.9600 2480.7800 971.4400 ;
        RECT 2477.7800 965.5200 2480.7800 966.0000 ;
        RECT 2477.7800 960.0800 2480.7800 960.5600 ;
        RECT 2477.7800 949.2000 2480.7800 949.6800 ;
        RECT 2477.7800 943.7600 2480.7800 944.2400 ;
        RECT 2477.7800 938.3200 2480.7800 938.8000 ;
        RECT 2477.7800 932.8800 2480.7800 933.3600 ;
        RECT 2477.7800 954.6400 2480.7800 955.1200 ;
        RECT 2572.3400 916.5600 2573.9400 917.0400 ;
        RECT 2572.3400 922.0000 2573.9400 922.4800 ;
        RECT 2572.3400 900.2400 2573.9400 900.7200 ;
        RECT 2572.3400 905.6800 2573.9400 906.1600 ;
        RECT 2572.3400 911.1200 2573.9400 911.6000 ;
        RECT 2527.3400 916.5600 2528.9400 917.0400 ;
        RECT 2527.3400 922.0000 2528.9400 922.4800 ;
        RECT 2527.3400 900.2400 2528.9400 900.7200 ;
        RECT 2527.3400 905.6800 2528.9400 906.1600 ;
        RECT 2527.3400 911.1200 2528.9400 911.6000 ;
        RECT 2572.3400 889.3600 2573.9400 889.8400 ;
        RECT 2572.3400 894.8000 2573.9400 895.2800 ;
        RECT 2572.3400 873.0400 2573.9400 873.5200 ;
        RECT 2572.3400 878.4800 2573.9400 878.9600 ;
        RECT 2572.3400 883.9200 2573.9400 884.4000 ;
        RECT 2527.3400 889.3600 2528.9400 889.8400 ;
        RECT 2527.3400 894.8000 2528.9400 895.2800 ;
        RECT 2527.3400 873.0400 2528.9400 873.5200 ;
        RECT 2527.3400 878.4800 2528.9400 878.9600 ;
        RECT 2527.3400 883.9200 2528.9400 884.4000 ;
        RECT 2477.7800 916.5600 2480.7800 917.0400 ;
        RECT 2477.7800 922.0000 2480.7800 922.4800 ;
        RECT 2477.7800 905.6800 2480.7800 906.1600 ;
        RECT 2477.7800 900.2400 2480.7800 900.7200 ;
        RECT 2477.7800 911.1200 2480.7800 911.6000 ;
        RECT 2477.7800 889.3600 2480.7800 889.8400 ;
        RECT 2477.7800 894.8000 2480.7800 895.2800 ;
        RECT 2477.7800 878.4800 2480.7800 878.9600 ;
        RECT 2477.7800 873.0400 2480.7800 873.5200 ;
        RECT 2477.7800 883.9200 2480.7800 884.4000 ;
        RECT 2477.7800 927.4400 2480.7800 927.9200 ;
        RECT 2527.3400 927.4400 2528.9400 927.9200 ;
        RECT 2572.3400 927.4400 2573.9400 927.9200 ;
        RECT 2673.8800 862.1600 2676.8800 862.6400 ;
        RECT 2673.8800 867.6000 2676.8800 868.0800 ;
        RECT 2662.3400 862.1600 2663.9400 862.6400 ;
        RECT 2662.3400 867.6000 2663.9400 868.0800 ;
        RECT 2673.8800 845.8400 2676.8800 846.3200 ;
        RECT 2673.8800 851.2800 2676.8800 851.7600 ;
        RECT 2673.8800 856.7200 2676.8800 857.2000 ;
        RECT 2662.3400 845.8400 2663.9400 846.3200 ;
        RECT 2662.3400 851.2800 2663.9400 851.7600 ;
        RECT 2662.3400 856.7200 2663.9400 857.2000 ;
        RECT 2673.8800 834.9600 2676.8800 835.4400 ;
        RECT 2673.8800 840.4000 2676.8800 840.8800 ;
        RECT 2662.3400 834.9600 2663.9400 835.4400 ;
        RECT 2662.3400 840.4000 2663.9400 840.8800 ;
        RECT 2673.8800 818.6400 2676.8800 819.1200 ;
        RECT 2673.8800 824.0800 2676.8800 824.5600 ;
        RECT 2673.8800 829.5200 2676.8800 830.0000 ;
        RECT 2662.3400 818.6400 2663.9400 819.1200 ;
        RECT 2662.3400 824.0800 2663.9400 824.5600 ;
        RECT 2662.3400 829.5200 2663.9400 830.0000 ;
        RECT 2617.3400 862.1600 2618.9400 862.6400 ;
        RECT 2617.3400 867.6000 2618.9400 868.0800 ;
        RECT 2617.3400 845.8400 2618.9400 846.3200 ;
        RECT 2617.3400 851.2800 2618.9400 851.7600 ;
        RECT 2617.3400 856.7200 2618.9400 857.2000 ;
        RECT 2617.3400 834.9600 2618.9400 835.4400 ;
        RECT 2617.3400 840.4000 2618.9400 840.8800 ;
        RECT 2617.3400 818.6400 2618.9400 819.1200 ;
        RECT 2617.3400 824.0800 2618.9400 824.5600 ;
        RECT 2617.3400 829.5200 2618.9400 830.0000 ;
        RECT 2673.8800 807.7600 2676.8800 808.2400 ;
        RECT 2673.8800 813.2000 2676.8800 813.6800 ;
        RECT 2662.3400 807.7600 2663.9400 808.2400 ;
        RECT 2662.3400 813.2000 2663.9400 813.6800 ;
        RECT 2673.8800 791.4400 2676.8800 791.9200 ;
        RECT 2673.8800 796.8800 2676.8800 797.3600 ;
        RECT 2673.8800 802.3200 2676.8800 802.8000 ;
        RECT 2662.3400 791.4400 2663.9400 791.9200 ;
        RECT 2662.3400 796.8800 2663.9400 797.3600 ;
        RECT 2662.3400 802.3200 2663.9400 802.8000 ;
        RECT 2673.8800 780.5600 2676.8800 781.0400 ;
        RECT 2673.8800 786.0000 2676.8800 786.4800 ;
        RECT 2662.3400 780.5600 2663.9400 781.0400 ;
        RECT 2662.3400 786.0000 2663.9400 786.4800 ;
        RECT 2673.8800 775.1200 2676.8800 775.6000 ;
        RECT 2662.3400 775.1200 2663.9400 775.6000 ;
        RECT 2617.3400 807.7600 2618.9400 808.2400 ;
        RECT 2617.3400 813.2000 2618.9400 813.6800 ;
        RECT 2617.3400 791.4400 2618.9400 791.9200 ;
        RECT 2617.3400 796.8800 2618.9400 797.3600 ;
        RECT 2617.3400 802.3200 2618.9400 802.8000 ;
        RECT 2617.3400 780.5600 2618.9400 781.0400 ;
        RECT 2617.3400 786.0000 2618.9400 786.4800 ;
        RECT 2617.3400 775.1200 2618.9400 775.6000 ;
        RECT 2572.3400 862.1600 2573.9400 862.6400 ;
        RECT 2572.3400 867.6000 2573.9400 868.0800 ;
        RECT 2572.3400 845.8400 2573.9400 846.3200 ;
        RECT 2572.3400 851.2800 2573.9400 851.7600 ;
        RECT 2572.3400 856.7200 2573.9400 857.2000 ;
        RECT 2527.3400 862.1600 2528.9400 862.6400 ;
        RECT 2527.3400 867.6000 2528.9400 868.0800 ;
        RECT 2527.3400 845.8400 2528.9400 846.3200 ;
        RECT 2527.3400 851.2800 2528.9400 851.7600 ;
        RECT 2527.3400 856.7200 2528.9400 857.2000 ;
        RECT 2572.3400 834.9600 2573.9400 835.4400 ;
        RECT 2572.3400 840.4000 2573.9400 840.8800 ;
        RECT 2572.3400 818.6400 2573.9400 819.1200 ;
        RECT 2572.3400 824.0800 2573.9400 824.5600 ;
        RECT 2572.3400 829.5200 2573.9400 830.0000 ;
        RECT 2527.3400 834.9600 2528.9400 835.4400 ;
        RECT 2527.3400 840.4000 2528.9400 840.8800 ;
        RECT 2527.3400 818.6400 2528.9400 819.1200 ;
        RECT 2527.3400 824.0800 2528.9400 824.5600 ;
        RECT 2527.3400 829.5200 2528.9400 830.0000 ;
        RECT 2477.7800 862.1600 2480.7800 862.6400 ;
        RECT 2477.7800 867.6000 2480.7800 868.0800 ;
        RECT 2477.7800 851.2800 2480.7800 851.7600 ;
        RECT 2477.7800 845.8400 2480.7800 846.3200 ;
        RECT 2477.7800 856.7200 2480.7800 857.2000 ;
        RECT 2477.7800 834.9600 2480.7800 835.4400 ;
        RECT 2477.7800 840.4000 2480.7800 840.8800 ;
        RECT 2477.7800 824.0800 2480.7800 824.5600 ;
        RECT 2477.7800 818.6400 2480.7800 819.1200 ;
        RECT 2477.7800 829.5200 2480.7800 830.0000 ;
        RECT 2572.3400 807.7600 2573.9400 808.2400 ;
        RECT 2572.3400 813.2000 2573.9400 813.6800 ;
        RECT 2572.3400 791.4400 2573.9400 791.9200 ;
        RECT 2572.3400 796.8800 2573.9400 797.3600 ;
        RECT 2572.3400 802.3200 2573.9400 802.8000 ;
        RECT 2527.3400 807.7600 2528.9400 808.2400 ;
        RECT 2527.3400 813.2000 2528.9400 813.6800 ;
        RECT 2527.3400 791.4400 2528.9400 791.9200 ;
        RECT 2527.3400 796.8800 2528.9400 797.3600 ;
        RECT 2527.3400 802.3200 2528.9400 802.8000 ;
        RECT 2572.3400 786.0000 2573.9400 786.4800 ;
        RECT 2572.3400 780.5600 2573.9400 781.0400 ;
        RECT 2572.3400 775.1200 2573.9400 775.6000 ;
        RECT 2527.3400 786.0000 2528.9400 786.4800 ;
        RECT 2527.3400 780.5600 2528.9400 781.0400 ;
        RECT 2527.3400 775.1200 2528.9400 775.6000 ;
        RECT 2477.7800 807.7600 2480.7800 808.2400 ;
        RECT 2477.7800 813.2000 2480.7800 813.6800 ;
        RECT 2477.7800 796.8800 2480.7800 797.3600 ;
        RECT 2477.7800 791.4400 2480.7800 791.9200 ;
        RECT 2477.7800 802.3200 2480.7800 802.8000 ;
        RECT 2477.7800 780.5600 2480.7800 781.0400 ;
        RECT 2477.7800 786.0000 2480.7800 786.4800 ;
        RECT 2477.7800 775.1200 2480.7800 775.6000 ;
        RECT 2477.7800 973.3100 2676.8800 976.3100 ;
        RECT 2477.7800 768.2100 2676.8800 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2785.1600 2833.6100 2787.1600 2854.5400 ;
        RECT 2698.0000 2833.6100 2700.0000 2854.5400 ;
      LAYER met3 ;
        RECT 2785.1600 2850.0400 2787.1600 2850.5200 ;
        RECT 2698.0000 2850.0400 2700.0000 2850.5200 ;
        RECT 2785.1600 2839.1600 2787.1600 2839.6400 ;
        RECT 2698.0000 2839.1600 2700.0000 2839.6400 ;
        RECT 2698.0000 2844.6000 2700.0000 2845.0800 ;
        RECT 2785.1600 2844.6000 2787.1600 2845.0800 ;
        RECT 2698.0000 2852.5400 2787.1600 2854.5400 ;
        RECT 2698.0000 2833.6100 2787.1600 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 538.5700 2699.5000 746.6700 ;
        RECT 2785.6600 538.5700 2787.1600 746.6700 ;
      LAYER met3 ;
        RECT 2785.6600 741.3200 2787.1600 741.8000 ;
        RECT 2785.6600 735.8800 2787.1600 736.3600 ;
        RECT 2785.6600 730.4400 2787.1600 730.9200 ;
        RECT 2785.6600 719.5600 2787.1600 720.0400 ;
        RECT 2785.6600 714.1200 2787.1600 714.6000 ;
        RECT 2785.6600 708.6800 2787.1600 709.1600 ;
        RECT 2785.6600 703.2400 2787.1600 703.7200 ;
        RECT 2785.6600 725.0000 2787.1600 725.4800 ;
        RECT 2785.6600 692.3600 2787.1600 692.8400 ;
        RECT 2785.6600 686.9200 2787.1600 687.4000 ;
        RECT 2785.6600 681.4800 2787.1600 681.9600 ;
        RECT 2785.6600 676.0400 2787.1600 676.5200 ;
        RECT 2785.6600 670.6000 2787.1600 671.0800 ;
        RECT 2785.6600 665.1600 2787.1600 665.6400 ;
        RECT 2785.6600 659.7200 2787.1600 660.2000 ;
        RECT 2785.6600 654.2800 2787.1600 654.7600 ;
        RECT 2785.6600 648.8400 2787.1600 649.3200 ;
        RECT 2785.6600 643.4000 2787.1600 643.8800 ;
        RECT 2785.6600 697.8000 2787.1600 698.2800 ;
        RECT 2698.0000 741.3200 2699.5000 741.8000 ;
        RECT 2698.0000 735.8800 2699.5000 736.3600 ;
        RECT 2698.0000 730.4400 2699.5000 730.9200 ;
        RECT 2698.0000 719.5600 2699.5000 720.0400 ;
        RECT 2698.0000 714.1200 2699.5000 714.6000 ;
        RECT 2698.0000 708.6800 2699.5000 709.1600 ;
        RECT 2698.0000 703.2400 2699.5000 703.7200 ;
        RECT 2698.0000 725.0000 2699.5000 725.4800 ;
        RECT 2698.0000 692.3600 2699.5000 692.8400 ;
        RECT 2698.0000 686.9200 2699.5000 687.4000 ;
        RECT 2698.0000 681.4800 2699.5000 681.9600 ;
        RECT 2698.0000 676.0400 2699.5000 676.5200 ;
        RECT 2698.0000 670.6000 2699.5000 671.0800 ;
        RECT 2698.0000 665.1600 2699.5000 665.6400 ;
        RECT 2698.0000 659.7200 2699.5000 660.2000 ;
        RECT 2698.0000 654.2800 2699.5000 654.7600 ;
        RECT 2698.0000 648.8400 2699.5000 649.3200 ;
        RECT 2698.0000 643.4000 2699.5000 643.8800 ;
        RECT 2698.0000 697.8000 2699.5000 698.2800 ;
        RECT 2785.6600 637.9600 2787.1600 638.4400 ;
        RECT 2785.6600 632.5200 2787.1600 633.0000 ;
        RECT 2785.6600 627.0800 2787.1600 627.5600 ;
        RECT 2785.6600 621.6400 2787.1600 622.1200 ;
        RECT 2785.6600 616.2000 2787.1600 616.6800 ;
        RECT 2785.6600 610.7600 2787.1600 611.2400 ;
        RECT 2785.6600 605.3200 2787.1600 605.8000 ;
        RECT 2785.6600 599.8800 2787.1600 600.3600 ;
        RECT 2785.6600 594.4400 2787.1600 594.9200 ;
        RECT 2785.6600 589.0000 2787.1600 589.4800 ;
        RECT 2785.6600 583.5600 2787.1600 584.0400 ;
        RECT 2785.6600 578.1200 2787.1600 578.6000 ;
        RECT 2785.6600 572.6800 2787.1600 573.1600 ;
        RECT 2785.6600 567.2400 2787.1600 567.7200 ;
        RECT 2785.6600 561.8000 2787.1600 562.2800 ;
        RECT 2785.6600 556.3600 2787.1600 556.8400 ;
        RECT 2785.6600 550.9200 2787.1600 551.4000 ;
        RECT 2785.6600 545.4800 2787.1600 545.9600 ;
        RECT 2698.0000 637.9600 2699.5000 638.4400 ;
        RECT 2698.0000 632.5200 2699.5000 633.0000 ;
        RECT 2698.0000 627.0800 2699.5000 627.5600 ;
        RECT 2698.0000 621.6400 2699.5000 622.1200 ;
        RECT 2698.0000 616.2000 2699.5000 616.6800 ;
        RECT 2698.0000 610.7600 2699.5000 611.2400 ;
        RECT 2698.0000 605.3200 2699.5000 605.8000 ;
        RECT 2698.0000 599.8800 2699.5000 600.3600 ;
        RECT 2698.0000 594.4400 2699.5000 594.9200 ;
        RECT 2698.0000 589.0000 2699.5000 589.4800 ;
        RECT 2698.0000 583.5600 2699.5000 584.0400 ;
        RECT 2698.0000 578.1200 2699.5000 578.6000 ;
        RECT 2698.0000 572.6800 2699.5000 573.1600 ;
        RECT 2698.0000 567.2400 2699.5000 567.7200 ;
        RECT 2698.0000 561.8000 2699.5000 562.2800 ;
        RECT 2698.0000 556.3600 2699.5000 556.8400 ;
        RECT 2698.0000 550.9200 2699.5000 551.4000 ;
        RECT 2698.0000 545.4800 2699.5000 545.9600 ;
        RECT 2698.0000 745.1700 2787.1600 746.6700 ;
        RECT 2698.0000 538.5700 2787.1600 540.0700 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 308.9300 2699.5000 517.0300 ;
        RECT 2785.6600 308.9300 2787.1600 517.0300 ;
      LAYER met3 ;
        RECT 2785.6600 511.6800 2787.1600 512.1600 ;
        RECT 2785.6600 506.2400 2787.1600 506.7200 ;
        RECT 2785.6600 500.8000 2787.1600 501.2800 ;
        RECT 2785.6600 489.9200 2787.1600 490.4000 ;
        RECT 2785.6600 484.4800 2787.1600 484.9600 ;
        RECT 2785.6600 479.0400 2787.1600 479.5200 ;
        RECT 2785.6600 473.6000 2787.1600 474.0800 ;
        RECT 2785.6600 495.3600 2787.1600 495.8400 ;
        RECT 2785.6600 462.7200 2787.1600 463.2000 ;
        RECT 2785.6600 457.2800 2787.1600 457.7600 ;
        RECT 2785.6600 451.8400 2787.1600 452.3200 ;
        RECT 2785.6600 446.4000 2787.1600 446.8800 ;
        RECT 2785.6600 440.9600 2787.1600 441.4400 ;
        RECT 2785.6600 435.5200 2787.1600 436.0000 ;
        RECT 2785.6600 430.0800 2787.1600 430.5600 ;
        RECT 2785.6600 424.6400 2787.1600 425.1200 ;
        RECT 2785.6600 419.2000 2787.1600 419.6800 ;
        RECT 2785.6600 413.7600 2787.1600 414.2400 ;
        RECT 2785.6600 468.1600 2787.1600 468.6400 ;
        RECT 2698.0000 511.6800 2699.5000 512.1600 ;
        RECT 2698.0000 506.2400 2699.5000 506.7200 ;
        RECT 2698.0000 500.8000 2699.5000 501.2800 ;
        RECT 2698.0000 489.9200 2699.5000 490.4000 ;
        RECT 2698.0000 484.4800 2699.5000 484.9600 ;
        RECT 2698.0000 479.0400 2699.5000 479.5200 ;
        RECT 2698.0000 473.6000 2699.5000 474.0800 ;
        RECT 2698.0000 495.3600 2699.5000 495.8400 ;
        RECT 2698.0000 462.7200 2699.5000 463.2000 ;
        RECT 2698.0000 457.2800 2699.5000 457.7600 ;
        RECT 2698.0000 451.8400 2699.5000 452.3200 ;
        RECT 2698.0000 446.4000 2699.5000 446.8800 ;
        RECT 2698.0000 440.9600 2699.5000 441.4400 ;
        RECT 2698.0000 435.5200 2699.5000 436.0000 ;
        RECT 2698.0000 430.0800 2699.5000 430.5600 ;
        RECT 2698.0000 424.6400 2699.5000 425.1200 ;
        RECT 2698.0000 419.2000 2699.5000 419.6800 ;
        RECT 2698.0000 413.7600 2699.5000 414.2400 ;
        RECT 2698.0000 468.1600 2699.5000 468.6400 ;
        RECT 2785.6600 408.3200 2787.1600 408.8000 ;
        RECT 2785.6600 402.8800 2787.1600 403.3600 ;
        RECT 2785.6600 397.4400 2787.1600 397.9200 ;
        RECT 2785.6600 392.0000 2787.1600 392.4800 ;
        RECT 2785.6600 386.5600 2787.1600 387.0400 ;
        RECT 2785.6600 381.1200 2787.1600 381.6000 ;
        RECT 2785.6600 375.6800 2787.1600 376.1600 ;
        RECT 2785.6600 370.2400 2787.1600 370.7200 ;
        RECT 2785.6600 364.8000 2787.1600 365.2800 ;
        RECT 2785.6600 359.3600 2787.1600 359.8400 ;
        RECT 2785.6600 353.9200 2787.1600 354.4000 ;
        RECT 2785.6600 348.4800 2787.1600 348.9600 ;
        RECT 2785.6600 343.0400 2787.1600 343.5200 ;
        RECT 2785.6600 337.6000 2787.1600 338.0800 ;
        RECT 2785.6600 332.1600 2787.1600 332.6400 ;
        RECT 2785.6600 326.7200 2787.1600 327.2000 ;
        RECT 2785.6600 321.2800 2787.1600 321.7600 ;
        RECT 2785.6600 315.8400 2787.1600 316.3200 ;
        RECT 2698.0000 408.3200 2699.5000 408.8000 ;
        RECT 2698.0000 402.8800 2699.5000 403.3600 ;
        RECT 2698.0000 397.4400 2699.5000 397.9200 ;
        RECT 2698.0000 392.0000 2699.5000 392.4800 ;
        RECT 2698.0000 386.5600 2699.5000 387.0400 ;
        RECT 2698.0000 381.1200 2699.5000 381.6000 ;
        RECT 2698.0000 375.6800 2699.5000 376.1600 ;
        RECT 2698.0000 370.2400 2699.5000 370.7200 ;
        RECT 2698.0000 364.8000 2699.5000 365.2800 ;
        RECT 2698.0000 359.3600 2699.5000 359.8400 ;
        RECT 2698.0000 353.9200 2699.5000 354.4000 ;
        RECT 2698.0000 348.4800 2699.5000 348.9600 ;
        RECT 2698.0000 343.0400 2699.5000 343.5200 ;
        RECT 2698.0000 337.6000 2699.5000 338.0800 ;
        RECT 2698.0000 332.1600 2699.5000 332.6400 ;
        RECT 2698.0000 326.7200 2699.5000 327.2000 ;
        RECT 2698.0000 321.2800 2699.5000 321.7600 ;
        RECT 2698.0000 315.8400 2699.5000 316.3200 ;
        RECT 2698.0000 515.5300 2787.1600 517.0300 ;
        RECT 2698.0000 308.9300 2787.1600 310.4300 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 79.2900 2699.5000 287.3900 ;
        RECT 2785.6600 79.2900 2787.1600 287.3900 ;
      LAYER met3 ;
        RECT 2785.6600 282.0400 2787.1600 282.5200 ;
        RECT 2785.6600 276.6000 2787.1600 277.0800 ;
        RECT 2785.6600 271.1600 2787.1600 271.6400 ;
        RECT 2785.6600 260.2800 2787.1600 260.7600 ;
        RECT 2785.6600 254.8400 2787.1600 255.3200 ;
        RECT 2785.6600 249.4000 2787.1600 249.8800 ;
        RECT 2785.6600 243.9600 2787.1600 244.4400 ;
        RECT 2785.6600 265.7200 2787.1600 266.2000 ;
        RECT 2785.6600 233.0800 2787.1600 233.5600 ;
        RECT 2785.6600 227.6400 2787.1600 228.1200 ;
        RECT 2785.6600 222.2000 2787.1600 222.6800 ;
        RECT 2785.6600 216.7600 2787.1600 217.2400 ;
        RECT 2785.6600 211.3200 2787.1600 211.8000 ;
        RECT 2785.6600 205.8800 2787.1600 206.3600 ;
        RECT 2785.6600 200.4400 2787.1600 200.9200 ;
        RECT 2785.6600 195.0000 2787.1600 195.4800 ;
        RECT 2785.6600 189.5600 2787.1600 190.0400 ;
        RECT 2785.6600 184.1200 2787.1600 184.6000 ;
        RECT 2785.6600 238.5200 2787.1600 239.0000 ;
        RECT 2698.0000 282.0400 2699.5000 282.5200 ;
        RECT 2698.0000 276.6000 2699.5000 277.0800 ;
        RECT 2698.0000 271.1600 2699.5000 271.6400 ;
        RECT 2698.0000 260.2800 2699.5000 260.7600 ;
        RECT 2698.0000 254.8400 2699.5000 255.3200 ;
        RECT 2698.0000 249.4000 2699.5000 249.8800 ;
        RECT 2698.0000 243.9600 2699.5000 244.4400 ;
        RECT 2698.0000 265.7200 2699.5000 266.2000 ;
        RECT 2698.0000 233.0800 2699.5000 233.5600 ;
        RECT 2698.0000 227.6400 2699.5000 228.1200 ;
        RECT 2698.0000 222.2000 2699.5000 222.6800 ;
        RECT 2698.0000 216.7600 2699.5000 217.2400 ;
        RECT 2698.0000 211.3200 2699.5000 211.8000 ;
        RECT 2698.0000 205.8800 2699.5000 206.3600 ;
        RECT 2698.0000 200.4400 2699.5000 200.9200 ;
        RECT 2698.0000 195.0000 2699.5000 195.4800 ;
        RECT 2698.0000 189.5600 2699.5000 190.0400 ;
        RECT 2698.0000 184.1200 2699.5000 184.6000 ;
        RECT 2698.0000 238.5200 2699.5000 239.0000 ;
        RECT 2785.6600 178.6800 2787.1600 179.1600 ;
        RECT 2785.6600 173.2400 2787.1600 173.7200 ;
        RECT 2785.6600 167.8000 2787.1600 168.2800 ;
        RECT 2785.6600 162.3600 2787.1600 162.8400 ;
        RECT 2785.6600 156.9200 2787.1600 157.4000 ;
        RECT 2785.6600 151.4800 2787.1600 151.9600 ;
        RECT 2785.6600 146.0400 2787.1600 146.5200 ;
        RECT 2785.6600 140.6000 2787.1600 141.0800 ;
        RECT 2785.6600 135.1600 2787.1600 135.6400 ;
        RECT 2785.6600 129.7200 2787.1600 130.2000 ;
        RECT 2785.6600 124.2800 2787.1600 124.7600 ;
        RECT 2785.6600 118.8400 2787.1600 119.3200 ;
        RECT 2785.6600 113.4000 2787.1600 113.8800 ;
        RECT 2785.6600 107.9600 2787.1600 108.4400 ;
        RECT 2785.6600 102.5200 2787.1600 103.0000 ;
        RECT 2785.6600 97.0800 2787.1600 97.5600 ;
        RECT 2785.6600 91.6400 2787.1600 92.1200 ;
        RECT 2785.6600 86.2000 2787.1600 86.6800 ;
        RECT 2698.0000 178.6800 2699.5000 179.1600 ;
        RECT 2698.0000 173.2400 2699.5000 173.7200 ;
        RECT 2698.0000 167.8000 2699.5000 168.2800 ;
        RECT 2698.0000 162.3600 2699.5000 162.8400 ;
        RECT 2698.0000 156.9200 2699.5000 157.4000 ;
        RECT 2698.0000 151.4800 2699.5000 151.9600 ;
        RECT 2698.0000 146.0400 2699.5000 146.5200 ;
        RECT 2698.0000 140.6000 2699.5000 141.0800 ;
        RECT 2698.0000 135.1600 2699.5000 135.6400 ;
        RECT 2698.0000 129.7200 2699.5000 130.2000 ;
        RECT 2698.0000 124.2800 2699.5000 124.7600 ;
        RECT 2698.0000 118.8400 2699.5000 119.3200 ;
        RECT 2698.0000 113.4000 2699.5000 113.8800 ;
        RECT 2698.0000 107.9600 2699.5000 108.4400 ;
        RECT 2698.0000 102.5200 2699.5000 103.0000 ;
        RECT 2698.0000 97.0800 2699.5000 97.5600 ;
        RECT 2698.0000 91.6400 2699.5000 92.1200 ;
        RECT 2698.0000 86.2000 2699.5000 86.6800 ;
        RECT 2698.0000 285.8900 2787.1600 287.3900 ;
        RECT 2698.0000 79.2900 2787.1600 80.7900 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'S_term_RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2785.1600 37.6700 2787.1600 58.6000 ;
        RECT 2698.0000 37.6700 2700.0000 58.6000 ;
      LAYER met3 ;
        RECT 2785.1600 54.1000 2787.1600 54.5800 ;
        RECT 2698.0000 54.1000 2700.0000 54.5800 ;
        RECT 2785.1600 43.2200 2787.1600 43.7000 ;
        RECT 2698.0000 43.2200 2700.0000 43.7000 ;
        RECT 2698.0000 48.6600 2700.0000 49.1400 ;
        RECT 2785.1600 48.6600 2787.1600 49.1400 ;
        RECT 2698.0000 56.6000 2787.1600 58.6000 ;
        RECT 2698.0000 37.6700 2787.1600 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 2605.3300 2699.5000 2813.4300 ;
        RECT 2785.6600 2605.3300 2787.1600 2813.4300 ;
      LAYER met3 ;
        RECT 2785.6600 2808.0800 2787.1600 2808.5600 ;
        RECT 2785.6600 2802.6400 2787.1600 2803.1200 ;
        RECT 2785.6600 2797.2000 2787.1600 2797.6800 ;
        RECT 2785.6600 2786.3200 2787.1600 2786.8000 ;
        RECT 2785.6600 2780.8800 2787.1600 2781.3600 ;
        RECT 2785.6600 2775.4400 2787.1600 2775.9200 ;
        RECT 2785.6600 2770.0000 2787.1600 2770.4800 ;
        RECT 2785.6600 2791.7600 2787.1600 2792.2400 ;
        RECT 2785.6600 2759.1200 2787.1600 2759.6000 ;
        RECT 2785.6600 2753.6800 2787.1600 2754.1600 ;
        RECT 2785.6600 2748.2400 2787.1600 2748.7200 ;
        RECT 2785.6600 2742.8000 2787.1600 2743.2800 ;
        RECT 2785.6600 2737.3600 2787.1600 2737.8400 ;
        RECT 2785.6600 2731.9200 2787.1600 2732.4000 ;
        RECT 2785.6600 2726.4800 2787.1600 2726.9600 ;
        RECT 2785.6600 2721.0400 2787.1600 2721.5200 ;
        RECT 2785.6600 2715.6000 2787.1600 2716.0800 ;
        RECT 2785.6600 2710.1600 2787.1600 2710.6400 ;
        RECT 2785.6600 2764.5600 2787.1600 2765.0400 ;
        RECT 2698.0000 2808.0800 2699.5000 2808.5600 ;
        RECT 2698.0000 2802.6400 2699.5000 2803.1200 ;
        RECT 2698.0000 2797.2000 2699.5000 2797.6800 ;
        RECT 2698.0000 2786.3200 2699.5000 2786.8000 ;
        RECT 2698.0000 2780.8800 2699.5000 2781.3600 ;
        RECT 2698.0000 2775.4400 2699.5000 2775.9200 ;
        RECT 2698.0000 2770.0000 2699.5000 2770.4800 ;
        RECT 2698.0000 2791.7600 2699.5000 2792.2400 ;
        RECT 2698.0000 2759.1200 2699.5000 2759.6000 ;
        RECT 2698.0000 2753.6800 2699.5000 2754.1600 ;
        RECT 2698.0000 2748.2400 2699.5000 2748.7200 ;
        RECT 2698.0000 2742.8000 2699.5000 2743.2800 ;
        RECT 2698.0000 2737.3600 2699.5000 2737.8400 ;
        RECT 2698.0000 2731.9200 2699.5000 2732.4000 ;
        RECT 2698.0000 2726.4800 2699.5000 2726.9600 ;
        RECT 2698.0000 2721.0400 2699.5000 2721.5200 ;
        RECT 2698.0000 2715.6000 2699.5000 2716.0800 ;
        RECT 2698.0000 2710.1600 2699.5000 2710.6400 ;
        RECT 2698.0000 2764.5600 2699.5000 2765.0400 ;
        RECT 2785.6600 2704.7200 2787.1600 2705.2000 ;
        RECT 2785.6600 2699.2800 2787.1600 2699.7600 ;
        RECT 2785.6600 2693.8400 2787.1600 2694.3200 ;
        RECT 2785.6600 2688.4000 2787.1600 2688.8800 ;
        RECT 2785.6600 2682.9600 2787.1600 2683.4400 ;
        RECT 2785.6600 2677.5200 2787.1600 2678.0000 ;
        RECT 2785.6600 2672.0800 2787.1600 2672.5600 ;
        RECT 2785.6600 2666.6400 2787.1600 2667.1200 ;
        RECT 2785.6600 2661.2000 2787.1600 2661.6800 ;
        RECT 2785.6600 2655.7600 2787.1600 2656.2400 ;
        RECT 2785.6600 2650.3200 2787.1600 2650.8000 ;
        RECT 2785.6600 2644.8800 2787.1600 2645.3600 ;
        RECT 2785.6600 2639.4400 2787.1600 2639.9200 ;
        RECT 2785.6600 2634.0000 2787.1600 2634.4800 ;
        RECT 2785.6600 2628.5600 2787.1600 2629.0400 ;
        RECT 2785.6600 2623.1200 2787.1600 2623.6000 ;
        RECT 2785.6600 2617.6800 2787.1600 2618.1600 ;
        RECT 2785.6600 2612.2400 2787.1600 2612.7200 ;
        RECT 2698.0000 2704.7200 2699.5000 2705.2000 ;
        RECT 2698.0000 2699.2800 2699.5000 2699.7600 ;
        RECT 2698.0000 2693.8400 2699.5000 2694.3200 ;
        RECT 2698.0000 2688.4000 2699.5000 2688.8800 ;
        RECT 2698.0000 2682.9600 2699.5000 2683.4400 ;
        RECT 2698.0000 2677.5200 2699.5000 2678.0000 ;
        RECT 2698.0000 2672.0800 2699.5000 2672.5600 ;
        RECT 2698.0000 2666.6400 2699.5000 2667.1200 ;
        RECT 2698.0000 2661.2000 2699.5000 2661.6800 ;
        RECT 2698.0000 2655.7600 2699.5000 2656.2400 ;
        RECT 2698.0000 2650.3200 2699.5000 2650.8000 ;
        RECT 2698.0000 2644.8800 2699.5000 2645.3600 ;
        RECT 2698.0000 2639.4400 2699.5000 2639.9200 ;
        RECT 2698.0000 2634.0000 2699.5000 2634.4800 ;
        RECT 2698.0000 2628.5600 2699.5000 2629.0400 ;
        RECT 2698.0000 2623.1200 2699.5000 2623.6000 ;
        RECT 2698.0000 2617.6800 2699.5000 2618.1600 ;
        RECT 2698.0000 2612.2400 2699.5000 2612.7200 ;
        RECT 2698.0000 2811.9300 2787.1600 2813.4300 ;
        RECT 2698.0000 2605.3300 2787.1600 2606.8300 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 2375.6900 2699.5000 2583.7900 ;
        RECT 2785.6600 2375.6900 2787.1600 2583.7900 ;
      LAYER met3 ;
        RECT 2785.6600 2578.4400 2787.1600 2578.9200 ;
        RECT 2785.6600 2573.0000 2787.1600 2573.4800 ;
        RECT 2785.6600 2567.5600 2787.1600 2568.0400 ;
        RECT 2785.6600 2556.6800 2787.1600 2557.1600 ;
        RECT 2785.6600 2551.2400 2787.1600 2551.7200 ;
        RECT 2785.6600 2545.8000 2787.1600 2546.2800 ;
        RECT 2785.6600 2540.3600 2787.1600 2540.8400 ;
        RECT 2785.6600 2562.1200 2787.1600 2562.6000 ;
        RECT 2785.6600 2529.4800 2787.1600 2529.9600 ;
        RECT 2785.6600 2524.0400 2787.1600 2524.5200 ;
        RECT 2785.6600 2518.6000 2787.1600 2519.0800 ;
        RECT 2785.6600 2513.1600 2787.1600 2513.6400 ;
        RECT 2785.6600 2507.7200 2787.1600 2508.2000 ;
        RECT 2785.6600 2502.2800 2787.1600 2502.7600 ;
        RECT 2785.6600 2496.8400 2787.1600 2497.3200 ;
        RECT 2785.6600 2491.4000 2787.1600 2491.8800 ;
        RECT 2785.6600 2485.9600 2787.1600 2486.4400 ;
        RECT 2785.6600 2480.5200 2787.1600 2481.0000 ;
        RECT 2785.6600 2534.9200 2787.1600 2535.4000 ;
        RECT 2698.0000 2578.4400 2699.5000 2578.9200 ;
        RECT 2698.0000 2573.0000 2699.5000 2573.4800 ;
        RECT 2698.0000 2567.5600 2699.5000 2568.0400 ;
        RECT 2698.0000 2556.6800 2699.5000 2557.1600 ;
        RECT 2698.0000 2551.2400 2699.5000 2551.7200 ;
        RECT 2698.0000 2545.8000 2699.5000 2546.2800 ;
        RECT 2698.0000 2540.3600 2699.5000 2540.8400 ;
        RECT 2698.0000 2562.1200 2699.5000 2562.6000 ;
        RECT 2698.0000 2529.4800 2699.5000 2529.9600 ;
        RECT 2698.0000 2524.0400 2699.5000 2524.5200 ;
        RECT 2698.0000 2518.6000 2699.5000 2519.0800 ;
        RECT 2698.0000 2513.1600 2699.5000 2513.6400 ;
        RECT 2698.0000 2507.7200 2699.5000 2508.2000 ;
        RECT 2698.0000 2502.2800 2699.5000 2502.7600 ;
        RECT 2698.0000 2496.8400 2699.5000 2497.3200 ;
        RECT 2698.0000 2491.4000 2699.5000 2491.8800 ;
        RECT 2698.0000 2485.9600 2699.5000 2486.4400 ;
        RECT 2698.0000 2480.5200 2699.5000 2481.0000 ;
        RECT 2698.0000 2534.9200 2699.5000 2535.4000 ;
        RECT 2785.6600 2475.0800 2787.1600 2475.5600 ;
        RECT 2785.6600 2469.6400 2787.1600 2470.1200 ;
        RECT 2785.6600 2464.2000 2787.1600 2464.6800 ;
        RECT 2785.6600 2458.7600 2787.1600 2459.2400 ;
        RECT 2785.6600 2453.3200 2787.1600 2453.8000 ;
        RECT 2785.6600 2447.8800 2787.1600 2448.3600 ;
        RECT 2785.6600 2442.4400 2787.1600 2442.9200 ;
        RECT 2785.6600 2437.0000 2787.1600 2437.4800 ;
        RECT 2785.6600 2431.5600 2787.1600 2432.0400 ;
        RECT 2785.6600 2426.1200 2787.1600 2426.6000 ;
        RECT 2785.6600 2420.6800 2787.1600 2421.1600 ;
        RECT 2785.6600 2415.2400 2787.1600 2415.7200 ;
        RECT 2785.6600 2409.8000 2787.1600 2410.2800 ;
        RECT 2785.6600 2404.3600 2787.1600 2404.8400 ;
        RECT 2785.6600 2398.9200 2787.1600 2399.4000 ;
        RECT 2785.6600 2393.4800 2787.1600 2393.9600 ;
        RECT 2785.6600 2388.0400 2787.1600 2388.5200 ;
        RECT 2785.6600 2382.6000 2787.1600 2383.0800 ;
        RECT 2698.0000 2475.0800 2699.5000 2475.5600 ;
        RECT 2698.0000 2469.6400 2699.5000 2470.1200 ;
        RECT 2698.0000 2464.2000 2699.5000 2464.6800 ;
        RECT 2698.0000 2458.7600 2699.5000 2459.2400 ;
        RECT 2698.0000 2453.3200 2699.5000 2453.8000 ;
        RECT 2698.0000 2447.8800 2699.5000 2448.3600 ;
        RECT 2698.0000 2442.4400 2699.5000 2442.9200 ;
        RECT 2698.0000 2437.0000 2699.5000 2437.4800 ;
        RECT 2698.0000 2431.5600 2699.5000 2432.0400 ;
        RECT 2698.0000 2426.1200 2699.5000 2426.6000 ;
        RECT 2698.0000 2420.6800 2699.5000 2421.1600 ;
        RECT 2698.0000 2415.2400 2699.5000 2415.7200 ;
        RECT 2698.0000 2409.8000 2699.5000 2410.2800 ;
        RECT 2698.0000 2404.3600 2699.5000 2404.8400 ;
        RECT 2698.0000 2398.9200 2699.5000 2399.4000 ;
        RECT 2698.0000 2393.4800 2699.5000 2393.9600 ;
        RECT 2698.0000 2388.0400 2699.5000 2388.5200 ;
        RECT 2698.0000 2382.6000 2699.5000 2383.0800 ;
        RECT 2698.0000 2582.2900 2787.1600 2583.7900 ;
        RECT 2698.0000 2375.6900 2787.1600 2377.1900 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 2146.0500 2699.5000 2354.1500 ;
        RECT 2785.6600 2146.0500 2787.1600 2354.1500 ;
      LAYER met3 ;
        RECT 2785.6600 2348.8000 2787.1600 2349.2800 ;
        RECT 2785.6600 2343.3600 2787.1600 2343.8400 ;
        RECT 2785.6600 2337.9200 2787.1600 2338.4000 ;
        RECT 2785.6600 2327.0400 2787.1600 2327.5200 ;
        RECT 2785.6600 2321.6000 2787.1600 2322.0800 ;
        RECT 2785.6600 2316.1600 2787.1600 2316.6400 ;
        RECT 2785.6600 2310.7200 2787.1600 2311.2000 ;
        RECT 2785.6600 2332.4800 2787.1600 2332.9600 ;
        RECT 2785.6600 2299.8400 2787.1600 2300.3200 ;
        RECT 2785.6600 2294.4000 2787.1600 2294.8800 ;
        RECT 2785.6600 2288.9600 2787.1600 2289.4400 ;
        RECT 2785.6600 2283.5200 2787.1600 2284.0000 ;
        RECT 2785.6600 2278.0800 2787.1600 2278.5600 ;
        RECT 2785.6600 2272.6400 2787.1600 2273.1200 ;
        RECT 2785.6600 2267.2000 2787.1600 2267.6800 ;
        RECT 2785.6600 2261.7600 2787.1600 2262.2400 ;
        RECT 2785.6600 2256.3200 2787.1600 2256.8000 ;
        RECT 2785.6600 2250.8800 2787.1600 2251.3600 ;
        RECT 2785.6600 2305.2800 2787.1600 2305.7600 ;
        RECT 2698.0000 2348.8000 2699.5000 2349.2800 ;
        RECT 2698.0000 2343.3600 2699.5000 2343.8400 ;
        RECT 2698.0000 2337.9200 2699.5000 2338.4000 ;
        RECT 2698.0000 2327.0400 2699.5000 2327.5200 ;
        RECT 2698.0000 2321.6000 2699.5000 2322.0800 ;
        RECT 2698.0000 2316.1600 2699.5000 2316.6400 ;
        RECT 2698.0000 2310.7200 2699.5000 2311.2000 ;
        RECT 2698.0000 2332.4800 2699.5000 2332.9600 ;
        RECT 2698.0000 2299.8400 2699.5000 2300.3200 ;
        RECT 2698.0000 2294.4000 2699.5000 2294.8800 ;
        RECT 2698.0000 2288.9600 2699.5000 2289.4400 ;
        RECT 2698.0000 2283.5200 2699.5000 2284.0000 ;
        RECT 2698.0000 2278.0800 2699.5000 2278.5600 ;
        RECT 2698.0000 2272.6400 2699.5000 2273.1200 ;
        RECT 2698.0000 2267.2000 2699.5000 2267.6800 ;
        RECT 2698.0000 2261.7600 2699.5000 2262.2400 ;
        RECT 2698.0000 2256.3200 2699.5000 2256.8000 ;
        RECT 2698.0000 2250.8800 2699.5000 2251.3600 ;
        RECT 2698.0000 2305.2800 2699.5000 2305.7600 ;
        RECT 2785.6600 2245.4400 2787.1600 2245.9200 ;
        RECT 2785.6600 2240.0000 2787.1600 2240.4800 ;
        RECT 2785.6600 2234.5600 2787.1600 2235.0400 ;
        RECT 2785.6600 2229.1200 2787.1600 2229.6000 ;
        RECT 2785.6600 2223.6800 2787.1600 2224.1600 ;
        RECT 2785.6600 2218.2400 2787.1600 2218.7200 ;
        RECT 2785.6600 2212.8000 2787.1600 2213.2800 ;
        RECT 2785.6600 2207.3600 2787.1600 2207.8400 ;
        RECT 2785.6600 2201.9200 2787.1600 2202.4000 ;
        RECT 2785.6600 2196.4800 2787.1600 2196.9600 ;
        RECT 2785.6600 2191.0400 2787.1600 2191.5200 ;
        RECT 2785.6600 2185.6000 2787.1600 2186.0800 ;
        RECT 2785.6600 2180.1600 2787.1600 2180.6400 ;
        RECT 2785.6600 2174.7200 2787.1600 2175.2000 ;
        RECT 2785.6600 2169.2800 2787.1600 2169.7600 ;
        RECT 2785.6600 2163.8400 2787.1600 2164.3200 ;
        RECT 2785.6600 2158.4000 2787.1600 2158.8800 ;
        RECT 2785.6600 2152.9600 2787.1600 2153.4400 ;
        RECT 2698.0000 2245.4400 2699.5000 2245.9200 ;
        RECT 2698.0000 2240.0000 2699.5000 2240.4800 ;
        RECT 2698.0000 2234.5600 2699.5000 2235.0400 ;
        RECT 2698.0000 2229.1200 2699.5000 2229.6000 ;
        RECT 2698.0000 2223.6800 2699.5000 2224.1600 ;
        RECT 2698.0000 2218.2400 2699.5000 2218.7200 ;
        RECT 2698.0000 2212.8000 2699.5000 2213.2800 ;
        RECT 2698.0000 2207.3600 2699.5000 2207.8400 ;
        RECT 2698.0000 2201.9200 2699.5000 2202.4000 ;
        RECT 2698.0000 2196.4800 2699.5000 2196.9600 ;
        RECT 2698.0000 2191.0400 2699.5000 2191.5200 ;
        RECT 2698.0000 2185.6000 2699.5000 2186.0800 ;
        RECT 2698.0000 2180.1600 2699.5000 2180.6400 ;
        RECT 2698.0000 2174.7200 2699.5000 2175.2000 ;
        RECT 2698.0000 2169.2800 2699.5000 2169.7600 ;
        RECT 2698.0000 2163.8400 2699.5000 2164.3200 ;
        RECT 2698.0000 2158.4000 2699.5000 2158.8800 ;
        RECT 2698.0000 2152.9600 2699.5000 2153.4400 ;
        RECT 2698.0000 2352.6500 2787.1600 2354.1500 ;
        RECT 2698.0000 2146.0500 2787.1600 2147.5500 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 1916.4100 2699.5000 2124.5100 ;
        RECT 2785.6600 1916.4100 2787.1600 2124.5100 ;
      LAYER met3 ;
        RECT 2785.6600 2119.1600 2787.1600 2119.6400 ;
        RECT 2785.6600 2113.7200 2787.1600 2114.2000 ;
        RECT 2785.6600 2108.2800 2787.1600 2108.7600 ;
        RECT 2785.6600 2097.4000 2787.1600 2097.8800 ;
        RECT 2785.6600 2091.9600 2787.1600 2092.4400 ;
        RECT 2785.6600 2086.5200 2787.1600 2087.0000 ;
        RECT 2785.6600 2081.0800 2787.1600 2081.5600 ;
        RECT 2785.6600 2102.8400 2787.1600 2103.3200 ;
        RECT 2785.6600 2070.2000 2787.1600 2070.6800 ;
        RECT 2785.6600 2064.7600 2787.1600 2065.2400 ;
        RECT 2785.6600 2059.3200 2787.1600 2059.8000 ;
        RECT 2785.6600 2053.8800 2787.1600 2054.3600 ;
        RECT 2785.6600 2048.4400 2787.1600 2048.9200 ;
        RECT 2785.6600 2043.0000 2787.1600 2043.4800 ;
        RECT 2785.6600 2037.5600 2787.1600 2038.0400 ;
        RECT 2785.6600 2032.1200 2787.1600 2032.6000 ;
        RECT 2785.6600 2026.6800 2787.1600 2027.1600 ;
        RECT 2785.6600 2021.2400 2787.1600 2021.7200 ;
        RECT 2785.6600 2075.6400 2787.1600 2076.1200 ;
        RECT 2698.0000 2119.1600 2699.5000 2119.6400 ;
        RECT 2698.0000 2113.7200 2699.5000 2114.2000 ;
        RECT 2698.0000 2108.2800 2699.5000 2108.7600 ;
        RECT 2698.0000 2097.4000 2699.5000 2097.8800 ;
        RECT 2698.0000 2091.9600 2699.5000 2092.4400 ;
        RECT 2698.0000 2086.5200 2699.5000 2087.0000 ;
        RECT 2698.0000 2081.0800 2699.5000 2081.5600 ;
        RECT 2698.0000 2102.8400 2699.5000 2103.3200 ;
        RECT 2698.0000 2070.2000 2699.5000 2070.6800 ;
        RECT 2698.0000 2064.7600 2699.5000 2065.2400 ;
        RECT 2698.0000 2059.3200 2699.5000 2059.8000 ;
        RECT 2698.0000 2053.8800 2699.5000 2054.3600 ;
        RECT 2698.0000 2048.4400 2699.5000 2048.9200 ;
        RECT 2698.0000 2043.0000 2699.5000 2043.4800 ;
        RECT 2698.0000 2037.5600 2699.5000 2038.0400 ;
        RECT 2698.0000 2032.1200 2699.5000 2032.6000 ;
        RECT 2698.0000 2026.6800 2699.5000 2027.1600 ;
        RECT 2698.0000 2021.2400 2699.5000 2021.7200 ;
        RECT 2698.0000 2075.6400 2699.5000 2076.1200 ;
        RECT 2785.6600 2015.8000 2787.1600 2016.2800 ;
        RECT 2785.6600 2010.3600 2787.1600 2010.8400 ;
        RECT 2785.6600 2004.9200 2787.1600 2005.4000 ;
        RECT 2785.6600 1999.4800 2787.1600 1999.9600 ;
        RECT 2785.6600 1994.0400 2787.1600 1994.5200 ;
        RECT 2785.6600 1988.6000 2787.1600 1989.0800 ;
        RECT 2785.6600 1983.1600 2787.1600 1983.6400 ;
        RECT 2785.6600 1977.7200 2787.1600 1978.2000 ;
        RECT 2785.6600 1972.2800 2787.1600 1972.7600 ;
        RECT 2785.6600 1966.8400 2787.1600 1967.3200 ;
        RECT 2785.6600 1961.4000 2787.1600 1961.8800 ;
        RECT 2785.6600 1955.9600 2787.1600 1956.4400 ;
        RECT 2785.6600 1950.5200 2787.1600 1951.0000 ;
        RECT 2785.6600 1945.0800 2787.1600 1945.5600 ;
        RECT 2785.6600 1939.6400 2787.1600 1940.1200 ;
        RECT 2785.6600 1934.2000 2787.1600 1934.6800 ;
        RECT 2785.6600 1928.7600 2787.1600 1929.2400 ;
        RECT 2785.6600 1923.3200 2787.1600 1923.8000 ;
        RECT 2698.0000 2015.8000 2699.5000 2016.2800 ;
        RECT 2698.0000 2010.3600 2699.5000 2010.8400 ;
        RECT 2698.0000 2004.9200 2699.5000 2005.4000 ;
        RECT 2698.0000 1999.4800 2699.5000 1999.9600 ;
        RECT 2698.0000 1994.0400 2699.5000 1994.5200 ;
        RECT 2698.0000 1988.6000 2699.5000 1989.0800 ;
        RECT 2698.0000 1983.1600 2699.5000 1983.6400 ;
        RECT 2698.0000 1977.7200 2699.5000 1978.2000 ;
        RECT 2698.0000 1972.2800 2699.5000 1972.7600 ;
        RECT 2698.0000 1966.8400 2699.5000 1967.3200 ;
        RECT 2698.0000 1961.4000 2699.5000 1961.8800 ;
        RECT 2698.0000 1955.9600 2699.5000 1956.4400 ;
        RECT 2698.0000 1950.5200 2699.5000 1951.0000 ;
        RECT 2698.0000 1945.0800 2699.5000 1945.5600 ;
        RECT 2698.0000 1939.6400 2699.5000 1940.1200 ;
        RECT 2698.0000 1934.2000 2699.5000 1934.6800 ;
        RECT 2698.0000 1928.7600 2699.5000 1929.2400 ;
        RECT 2698.0000 1923.3200 2699.5000 1923.8000 ;
        RECT 2698.0000 2123.0100 2787.1600 2124.5100 ;
        RECT 2698.0000 1916.4100 2787.1600 1917.9100 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 1686.7700 2699.5000 1894.8700 ;
        RECT 2785.6600 1686.7700 2787.1600 1894.8700 ;
      LAYER met3 ;
        RECT 2785.6600 1889.5200 2787.1600 1890.0000 ;
        RECT 2785.6600 1884.0800 2787.1600 1884.5600 ;
        RECT 2785.6600 1878.6400 2787.1600 1879.1200 ;
        RECT 2785.6600 1867.7600 2787.1600 1868.2400 ;
        RECT 2785.6600 1862.3200 2787.1600 1862.8000 ;
        RECT 2785.6600 1856.8800 2787.1600 1857.3600 ;
        RECT 2785.6600 1851.4400 2787.1600 1851.9200 ;
        RECT 2785.6600 1873.2000 2787.1600 1873.6800 ;
        RECT 2785.6600 1840.5600 2787.1600 1841.0400 ;
        RECT 2785.6600 1835.1200 2787.1600 1835.6000 ;
        RECT 2785.6600 1829.6800 2787.1600 1830.1600 ;
        RECT 2785.6600 1824.2400 2787.1600 1824.7200 ;
        RECT 2785.6600 1818.8000 2787.1600 1819.2800 ;
        RECT 2785.6600 1813.3600 2787.1600 1813.8400 ;
        RECT 2785.6600 1807.9200 2787.1600 1808.4000 ;
        RECT 2785.6600 1802.4800 2787.1600 1802.9600 ;
        RECT 2785.6600 1797.0400 2787.1600 1797.5200 ;
        RECT 2785.6600 1791.6000 2787.1600 1792.0800 ;
        RECT 2785.6600 1846.0000 2787.1600 1846.4800 ;
        RECT 2698.0000 1889.5200 2699.5000 1890.0000 ;
        RECT 2698.0000 1884.0800 2699.5000 1884.5600 ;
        RECT 2698.0000 1878.6400 2699.5000 1879.1200 ;
        RECT 2698.0000 1867.7600 2699.5000 1868.2400 ;
        RECT 2698.0000 1862.3200 2699.5000 1862.8000 ;
        RECT 2698.0000 1856.8800 2699.5000 1857.3600 ;
        RECT 2698.0000 1851.4400 2699.5000 1851.9200 ;
        RECT 2698.0000 1873.2000 2699.5000 1873.6800 ;
        RECT 2698.0000 1840.5600 2699.5000 1841.0400 ;
        RECT 2698.0000 1835.1200 2699.5000 1835.6000 ;
        RECT 2698.0000 1829.6800 2699.5000 1830.1600 ;
        RECT 2698.0000 1824.2400 2699.5000 1824.7200 ;
        RECT 2698.0000 1818.8000 2699.5000 1819.2800 ;
        RECT 2698.0000 1813.3600 2699.5000 1813.8400 ;
        RECT 2698.0000 1807.9200 2699.5000 1808.4000 ;
        RECT 2698.0000 1802.4800 2699.5000 1802.9600 ;
        RECT 2698.0000 1797.0400 2699.5000 1797.5200 ;
        RECT 2698.0000 1791.6000 2699.5000 1792.0800 ;
        RECT 2698.0000 1846.0000 2699.5000 1846.4800 ;
        RECT 2785.6600 1786.1600 2787.1600 1786.6400 ;
        RECT 2785.6600 1780.7200 2787.1600 1781.2000 ;
        RECT 2785.6600 1775.2800 2787.1600 1775.7600 ;
        RECT 2785.6600 1769.8400 2787.1600 1770.3200 ;
        RECT 2785.6600 1764.4000 2787.1600 1764.8800 ;
        RECT 2785.6600 1758.9600 2787.1600 1759.4400 ;
        RECT 2785.6600 1753.5200 2787.1600 1754.0000 ;
        RECT 2785.6600 1748.0800 2787.1600 1748.5600 ;
        RECT 2785.6600 1742.6400 2787.1600 1743.1200 ;
        RECT 2785.6600 1737.2000 2787.1600 1737.6800 ;
        RECT 2785.6600 1731.7600 2787.1600 1732.2400 ;
        RECT 2785.6600 1726.3200 2787.1600 1726.8000 ;
        RECT 2785.6600 1720.8800 2787.1600 1721.3600 ;
        RECT 2785.6600 1715.4400 2787.1600 1715.9200 ;
        RECT 2785.6600 1710.0000 2787.1600 1710.4800 ;
        RECT 2785.6600 1704.5600 2787.1600 1705.0400 ;
        RECT 2785.6600 1699.1200 2787.1600 1699.6000 ;
        RECT 2785.6600 1693.6800 2787.1600 1694.1600 ;
        RECT 2698.0000 1786.1600 2699.5000 1786.6400 ;
        RECT 2698.0000 1780.7200 2699.5000 1781.2000 ;
        RECT 2698.0000 1775.2800 2699.5000 1775.7600 ;
        RECT 2698.0000 1769.8400 2699.5000 1770.3200 ;
        RECT 2698.0000 1764.4000 2699.5000 1764.8800 ;
        RECT 2698.0000 1758.9600 2699.5000 1759.4400 ;
        RECT 2698.0000 1753.5200 2699.5000 1754.0000 ;
        RECT 2698.0000 1748.0800 2699.5000 1748.5600 ;
        RECT 2698.0000 1742.6400 2699.5000 1743.1200 ;
        RECT 2698.0000 1737.2000 2699.5000 1737.6800 ;
        RECT 2698.0000 1731.7600 2699.5000 1732.2400 ;
        RECT 2698.0000 1726.3200 2699.5000 1726.8000 ;
        RECT 2698.0000 1720.8800 2699.5000 1721.3600 ;
        RECT 2698.0000 1715.4400 2699.5000 1715.9200 ;
        RECT 2698.0000 1710.0000 2699.5000 1710.4800 ;
        RECT 2698.0000 1704.5600 2699.5000 1705.0400 ;
        RECT 2698.0000 1699.1200 2699.5000 1699.6000 ;
        RECT 2698.0000 1693.6800 2699.5000 1694.1600 ;
        RECT 2698.0000 1893.3700 2787.1600 1894.8700 ;
        RECT 2698.0000 1686.7700 2787.1600 1688.2700 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 1457.1300 2699.5000 1665.2300 ;
        RECT 2785.6600 1457.1300 2787.1600 1665.2300 ;
      LAYER met3 ;
        RECT 2785.6600 1659.8800 2787.1600 1660.3600 ;
        RECT 2785.6600 1654.4400 2787.1600 1654.9200 ;
        RECT 2785.6600 1649.0000 2787.1600 1649.4800 ;
        RECT 2785.6600 1638.1200 2787.1600 1638.6000 ;
        RECT 2785.6600 1632.6800 2787.1600 1633.1600 ;
        RECT 2785.6600 1627.2400 2787.1600 1627.7200 ;
        RECT 2785.6600 1621.8000 2787.1600 1622.2800 ;
        RECT 2785.6600 1643.5600 2787.1600 1644.0400 ;
        RECT 2785.6600 1610.9200 2787.1600 1611.4000 ;
        RECT 2785.6600 1605.4800 2787.1600 1605.9600 ;
        RECT 2785.6600 1600.0400 2787.1600 1600.5200 ;
        RECT 2785.6600 1594.6000 2787.1600 1595.0800 ;
        RECT 2785.6600 1589.1600 2787.1600 1589.6400 ;
        RECT 2785.6600 1583.7200 2787.1600 1584.2000 ;
        RECT 2785.6600 1578.2800 2787.1600 1578.7600 ;
        RECT 2785.6600 1572.8400 2787.1600 1573.3200 ;
        RECT 2785.6600 1567.4000 2787.1600 1567.8800 ;
        RECT 2785.6600 1561.9600 2787.1600 1562.4400 ;
        RECT 2785.6600 1616.3600 2787.1600 1616.8400 ;
        RECT 2698.0000 1659.8800 2699.5000 1660.3600 ;
        RECT 2698.0000 1654.4400 2699.5000 1654.9200 ;
        RECT 2698.0000 1649.0000 2699.5000 1649.4800 ;
        RECT 2698.0000 1638.1200 2699.5000 1638.6000 ;
        RECT 2698.0000 1632.6800 2699.5000 1633.1600 ;
        RECT 2698.0000 1627.2400 2699.5000 1627.7200 ;
        RECT 2698.0000 1621.8000 2699.5000 1622.2800 ;
        RECT 2698.0000 1643.5600 2699.5000 1644.0400 ;
        RECT 2698.0000 1610.9200 2699.5000 1611.4000 ;
        RECT 2698.0000 1605.4800 2699.5000 1605.9600 ;
        RECT 2698.0000 1600.0400 2699.5000 1600.5200 ;
        RECT 2698.0000 1594.6000 2699.5000 1595.0800 ;
        RECT 2698.0000 1589.1600 2699.5000 1589.6400 ;
        RECT 2698.0000 1583.7200 2699.5000 1584.2000 ;
        RECT 2698.0000 1578.2800 2699.5000 1578.7600 ;
        RECT 2698.0000 1572.8400 2699.5000 1573.3200 ;
        RECT 2698.0000 1567.4000 2699.5000 1567.8800 ;
        RECT 2698.0000 1561.9600 2699.5000 1562.4400 ;
        RECT 2698.0000 1616.3600 2699.5000 1616.8400 ;
        RECT 2785.6600 1556.5200 2787.1600 1557.0000 ;
        RECT 2785.6600 1551.0800 2787.1600 1551.5600 ;
        RECT 2785.6600 1545.6400 2787.1600 1546.1200 ;
        RECT 2785.6600 1540.2000 2787.1600 1540.6800 ;
        RECT 2785.6600 1534.7600 2787.1600 1535.2400 ;
        RECT 2785.6600 1529.3200 2787.1600 1529.8000 ;
        RECT 2785.6600 1523.8800 2787.1600 1524.3600 ;
        RECT 2785.6600 1518.4400 2787.1600 1518.9200 ;
        RECT 2785.6600 1513.0000 2787.1600 1513.4800 ;
        RECT 2785.6600 1507.5600 2787.1600 1508.0400 ;
        RECT 2785.6600 1502.1200 2787.1600 1502.6000 ;
        RECT 2785.6600 1496.6800 2787.1600 1497.1600 ;
        RECT 2785.6600 1491.2400 2787.1600 1491.7200 ;
        RECT 2785.6600 1485.8000 2787.1600 1486.2800 ;
        RECT 2785.6600 1480.3600 2787.1600 1480.8400 ;
        RECT 2785.6600 1474.9200 2787.1600 1475.4000 ;
        RECT 2785.6600 1469.4800 2787.1600 1469.9600 ;
        RECT 2785.6600 1464.0400 2787.1600 1464.5200 ;
        RECT 2698.0000 1556.5200 2699.5000 1557.0000 ;
        RECT 2698.0000 1551.0800 2699.5000 1551.5600 ;
        RECT 2698.0000 1545.6400 2699.5000 1546.1200 ;
        RECT 2698.0000 1540.2000 2699.5000 1540.6800 ;
        RECT 2698.0000 1534.7600 2699.5000 1535.2400 ;
        RECT 2698.0000 1529.3200 2699.5000 1529.8000 ;
        RECT 2698.0000 1523.8800 2699.5000 1524.3600 ;
        RECT 2698.0000 1518.4400 2699.5000 1518.9200 ;
        RECT 2698.0000 1513.0000 2699.5000 1513.4800 ;
        RECT 2698.0000 1507.5600 2699.5000 1508.0400 ;
        RECT 2698.0000 1502.1200 2699.5000 1502.6000 ;
        RECT 2698.0000 1496.6800 2699.5000 1497.1600 ;
        RECT 2698.0000 1491.2400 2699.5000 1491.7200 ;
        RECT 2698.0000 1485.8000 2699.5000 1486.2800 ;
        RECT 2698.0000 1480.3600 2699.5000 1480.8400 ;
        RECT 2698.0000 1474.9200 2699.5000 1475.4000 ;
        RECT 2698.0000 1469.4800 2699.5000 1469.9600 ;
        RECT 2698.0000 1464.0400 2699.5000 1464.5200 ;
        RECT 2698.0000 1663.7300 2787.1600 1665.2300 ;
        RECT 2698.0000 1457.1300 2787.1600 1458.6300 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 1227.4900 2699.5000 1435.5900 ;
        RECT 2785.6600 1227.4900 2787.1600 1435.5900 ;
      LAYER met3 ;
        RECT 2785.6600 1430.2400 2787.1600 1430.7200 ;
        RECT 2785.6600 1424.8000 2787.1600 1425.2800 ;
        RECT 2785.6600 1419.3600 2787.1600 1419.8400 ;
        RECT 2785.6600 1408.4800 2787.1600 1408.9600 ;
        RECT 2785.6600 1403.0400 2787.1600 1403.5200 ;
        RECT 2785.6600 1397.6000 2787.1600 1398.0800 ;
        RECT 2785.6600 1392.1600 2787.1600 1392.6400 ;
        RECT 2785.6600 1413.9200 2787.1600 1414.4000 ;
        RECT 2785.6600 1381.2800 2787.1600 1381.7600 ;
        RECT 2785.6600 1375.8400 2787.1600 1376.3200 ;
        RECT 2785.6600 1370.4000 2787.1600 1370.8800 ;
        RECT 2785.6600 1364.9600 2787.1600 1365.4400 ;
        RECT 2785.6600 1359.5200 2787.1600 1360.0000 ;
        RECT 2785.6600 1354.0800 2787.1600 1354.5600 ;
        RECT 2785.6600 1348.6400 2787.1600 1349.1200 ;
        RECT 2785.6600 1343.2000 2787.1600 1343.6800 ;
        RECT 2785.6600 1337.7600 2787.1600 1338.2400 ;
        RECT 2785.6600 1332.3200 2787.1600 1332.8000 ;
        RECT 2785.6600 1386.7200 2787.1600 1387.2000 ;
        RECT 2698.0000 1430.2400 2699.5000 1430.7200 ;
        RECT 2698.0000 1424.8000 2699.5000 1425.2800 ;
        RECT 2698.0000 1419.3600 2699.5000 1419.8400 ;
        RECT 2698.0000 1408.4800 2699.5000 1408.9600 ;
        RECT 2698.0000 1403.0400 2699.5000 1403.5200 ;
        RECT 2698.0000 1397.6000 2699.5000 1398.0800 ;
        RECT 2698.0000 1392.1600 2699.5000 1392.6400 ;
        RECT 2698.0000 1413.9200 2699.5000 1414.4000 ;
        RECT 2698.0000 1381.2800 2699.5000 1381.7600 ;
        RECT 2698.0000 1375.8400 2699.5000 1376.3200 ;
        RECT 2698.0000 1370.4000 2699.5000 1370.8800 ;
        RECT 2698.0000 1364.9600 2699.5000 1365.4400 ;
        RECT 2698.0000 1359.5200 2699.5000 1360.0000 ;
        RECT 2698.0000 1354.0800 2699.5000 1354.5600 ;
        RECT 2698.0000 1348.6400 2699.5000 1349.1200 ;
        RECT 2698.0000 1343.2000 2699.5000 1343.6800 ;
        RECT 2698.0000 1337.7600 2699.5000 1338.2400 ;
        RECT 2698.0000 1332.3200 2699.5000 1332.8000 ;
        RECT 2698.0000 1386.7200 2699.5000 1387.2000 ;
        RECT 2785.6600 1326.8800 2787.1600 1327.3600 ;
        RECT 2785.6600 1321.4400 2787.1600 1321.9200 ;
        RECT 2785.6600 1316.0000 2787.1600 1316.4800 ;
        RECT 2785.6600 1310.5600 2787.1600 1311.0400 ;
        RECT 2785.6600 1305.1200 2787.1600 1305.6000 ;
        RECT 2785.6600 1299.6800 2787.1600 1300.1600 ;
        RECT 2785.6600 1294.2400 2787.1600 1294.7200 ;
        RECT 2785.6600 1288.8000 2787.1600 1289.2800 ;
        RECT 2785.6600 1283.3600 2787.1600 1283.8400 ;
        RECT 2785.6600 1277.9200 2787.1600 1278.4000 ;
        RECT 2785.6600 1272.4800 2787.1600 1272.9600 ;
        RECT 2785.6600 1267.0400 2787.1600 1267.5200 ;
        RECT 2785.6600 1261.6000 2787.1600 1262.0800 ;
        RECT 2785.6600 1256.1600 2787.1600 1256.6400 ;
        RECT 2785.6600 1250.7200 2787.1600 1251.2000 ;
        RECT 2785.6600 1245.2800 2787.1600 1245.7600 ;
        RECT 2785.6600 1239.8400 2787.1600 1240.3200 ;
        RECT 2785.6600 1234.4000 2787.1600 1234.8800 ;
        RECT 2698.0000 1326.8800 2699.5000 1327.3600 ;
        RECT 2698.0000 1321.4400 2699.5000 1321.9200 ;
        RECT 2698.0000 1316.0000 2699.5000 1316.4800 ;
        RECT 2698.0000 1310.5600 2699.5000 1311.0400 ;
        RECT 2698.0000 1305.1200 2699.5000 1305.6000 ;
        RECT 2698.0000 1299.6800 2699.5000 1300.1600 ;
        RECT 2698.0000 1294.2400 2699.5000 1294.7200 ;
        RECT 2698.0000 1288.8000 2699.5000 1289.2800 ;
        RECT 2698.0000 1283.3600 2699.5000 1283.8400 ;
        RECT 2698.0000 1277.9200 2699.5000 1278.4000 ;
        RECT 2698.0000 1272.4800 2699.5000 1272.9600 ;
        RECT 2698.0000 1267.0400 2699.5000 1267.5200 ;
        RECT 2698.0000 1261.6000 2699.5000 1262.0800 ;
        RECT 2698.0000 1256.1600 2699.5000 1256.6400 ;
        RECT 2698.0000 1250.7200 2699.5000 1251.2000 ;
        RECT 2698.0000 1245.2800 2699.5000 1245.7600 ;
        RECT 2698.0000 1239.8400 2699.5000 1240.3200 ;
        RECT 2698.0000 1234.4000 2699.5000 1234.8800 ;
        RECT 2698.0000 1434.0900 2787.1600 1435.5900 ;
        RECT 2698.0000 1227.4900 2787.1600 1228.9900 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 997.8500 2699.5000 1205.9500 ;
        RECT 2785.6600 997.8500 2787.1600 1205.9500 ;
      LAYER met3 ;
        RECT 2785.6600 1200.6000 2787.1600 1201.0800 ;
        RECT 2785.6600 1195.1600 2787.1600 1195.6400 ;
        RECT 2785.6600 1189.7200 2787.1600 1190.2000 ;
        RECT 2785.6600 1178.8400 2787.1600 1179.3200 ;
        RECT 2785.6600 1173.4000 2787.1600 1173.8800 ;
        RECT 2785.6600 1167.9600 2787.1600 1168.4400 ;
        RECT 2785.6600 1162.5200 2787.1600 1163.0000 ;
        RECT 2785.6600 1184.2800 2787.1600 1184.7600 ;
        RECT 2785.6600 1151.6400 2787.1600 1152.1200 ;
        RECT 2785.6600 1146.2000 2787.1600 1146.6800 ;
        RECT 2785.6600 1140.7600 2787.1600 1141.2400 ;
        RECT 2785.6600 1135.3200 2787.1600 1135.8000 ;
        RECT 2785.6600 1129.8800 2787.1600 1130.3600 ;
        RECT 2785.6600 1124.4400 2787.1600 1124.9200 ;
        RECT 2785.6600 1119.0000 2787.1600 1119.4800 ;
        RECT 2785.6600 1113.5600 2787.1600 1114.0400 ;
        RECT 2785.6600 1108.1200 2787.1600 1108.6000 ;
        RECT 2785.6600 1102.6800 2787.1600 1103.1600 ;
        RECT 2785.6600 1157.0800 2787.1600 1157.5600 ;
        RECT 2698.0000 1200.6000 2699.5000 1201.0800 ;
        RECT 2698.0000 1195.1600 2699.5000 1195.6400 ;
        RECT 2698.0000 1189.7200 2699.5000 1190.2000 ;
        RECT 2698.0000 1178.8400 2699.5000 1179.3200 ;
        RECT 2698.0000 1173.4000 2699.5000 1173.8800 ;
        RECT 2698.0000 1167.9600 2699.5000 1168.4400 ;
        RECT 2698.0000 1162.5200 2699.5000 1163.0000 ;
        RECT 2698.0000 1184.2800 2699.5000 1184.7600 ;
        RECT 2698.0000 1151.6400 2699.5000 1152.1200 ;
        RECT 2698.0000 1146.2000 2699.5000 1146.6800 ;
        RECT 2698.0000 1140.7600 2699.5000 1141.2400 ;
        RECT 2698.0000 1135.3200 2699.5000 1135.8000 ;
        RECT 2698.0000 1129.8800 2699.5000 1130.3600 ;
        RECT 2698.0000 1124.4400 2699.5000 1124.9200 ;
        RECT 2698.0000 1119.0000 2699.5000 1119.4800 ;
        RECT 2698.0000 1113.5600 2699.5000 1114.0400 ;
        RECT 2698.0000 1108.1200 2699.5000 1108.6000 ;
        RECT 2698.0000 1102.6800 2699.5000 1103.1600 ;
        RECT 2698.0000 1157.0800 2699.5000 1157.5600 ;
        RECT 2785.6600 1097.2400 2787.1600 1097.7200 ;
        RECT 2785.6600 1091.8000 2787.1600 1092.2800 ;
        RECT 2785.6600 1086.3600 2787.1600 1086.8400 ;
        RECT 2785.6600 1080.9200 2787.1600 1081.4000 ;
        RECT 2785.6600 1075.4800 2787.1600 1075.9600 ;
        RECT 2785.6600 1070.0400 2787.1600 1070.5200 ;
        RECT 2785.6600 1064.6000 2787.1600 1065.0800 ;
        RECT 2785.6600 1059.1600 2787.1600 1059.6400 ;
        RECT 2785.6600 1053.7200 2787.1600 1054.2000 ;
        RECT 2785.6600 1048.2800 2787.1600 1048.7600 ;
        RECT 2785.6600 1042.8400 2787.1600 1043.3200 ;
        RECT 2785.6600 1037.4000 2787.1600 1037.8800 ;
        RECT 2785.6600 1031.9600 2787.1600 1032.4400 ;
        RECT 2785.6600 1026.5200 2787.1600 1027.0000 ;
        RECT 2785.6600 1021.0800 2787.1600 1021.5600 ;
        RECT 2785.6600 1015.6400 2787.1600 1016.1200 ;
        RECT 2785.6600 1010.2000 2787.1600 1010.6800 ;
        RECT 2785.6600 1004.7600 2787.1600 1005.2400 ;
        RECT 2698.0000 1097.2400 2699.5000 1097.7200 ;
        RECT 2698.0000 1091.8000 2699.5000 1092.2800 ;
        RECT 2698.0000 1086.3600 2699.5000 1086.8400 ;
        RECT 2698.0000 1080.9200 2699.5000 1081.4000 ;
        RECT 2698.0000 1075.4800 2699.5000 1075.9600 ;
        RECT 2698.0000 1070.0400 2699.5000 1070.5200 ;
        RECT 2698.0000 1064.6000 2699.5000 1065.0800 ;
        RECT 2698.0000 1059.1600 2699.5000 1059.6400 ;
        RECT 2698.0000 1053.7200 2699.5000 1054.2000 ;
        RECT 2698.0000 1048.2800 2699.5000 1048.7600 ;
        RECT 2698.0000 1042.8400 2699.5000 1043.3200 ;
        RECT 2698.0000 1037.4000 2699.5000 1037.8800 ;
        RECT 2698.0000 1031.9600 2699.5000 1032.4400 ;
        RECT 2698.0000 1026.5200 2699.5000 1027.0000 ;
        RECT 2698.0000 1021.0800 2699.5000 1021.5600 ;
        RECT 2698.0000 1015.6400 2699.5000 1016.1200 ;
        RECT 2698.0000 1010.2000 2699.5000 1010.6800 ;
        RECT 2698.0000 1004.7600 2699.5000 1005.2400 ;
        RECT 2698.0000 1204.4500 2787.1600 1205.9500 ;
        RECT 2698.0000 997.8500 2787.1600 999.3500 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2698.0000 768.2100 2699.5000 976.3100 ;
        RECT 2785.6600 768.2100 2787.1600 976.3100 ;
      LAYER met3 ;
        RECT 2785.6600 970.9600 2787.1600 971.4400 ;
        RECT 2785.6600 965.5200 2787.1600 966.0000 ;
        RECT 2785.6600 960.0800 2787.1600 960.5600 ;
        RECT 2785.6600 949.2000 2787.1600 949.6800 ;
        RECT 2785.6600 943.7600 2787.1600 944.2400 ;
        RECT 2785.6600 938.3200 2787.1600 938.8000 ;
        RECT 2785.6600 932.8800 2787.1600 933.3600 ;
        RECT 2785.6600 954.6400 2787.1600 955.1200 ;
        RECT 2785.6600 922.0000 2787.1600 922.4800 ;
        RECT 2785.6600 916.5600 2787.1600 917.0400 ;
        RECT 2785.6600 911.1200 2787.1600 911.6000 ;
        RECT 2785.6600 905.6800 2787.1600 906.1600 ;
        RECT 2785.6600 900.2400 2787.1600 900.7200 ;
        RECT 2785.6600 894.8000 2787.1600 895.2800 ;
        RECT 2785.6600 889.3600 2787.1600 889.8400 ;
        RECT 2785.6600 883.9200 2787.1600 884.4000 ;
        RECT 2785.6600 878.4800 2787.1600 878.9600 ;
        RECT 2785.6600 873.0400 2787.1600 873.5200 ;
        RECT 2785.6600 927.4400 2787.1600 927.9200 ;
        RECT 2698.0000 970.9600 2699.5000 971.4400 ;
        RECT 2698.0000 965.5200 2699.5000 966.0000 ;
        RECT 2698.0000 960.0800 2699.5000 960.5600 ;
        RECT 2698.0000 949.2000 2699.5000 949.6800 ;
        RECT 2698.0000 943.7600 2699.5000 944.2400 ;
        RECT 2698.0000 938.3200 2699.5000 938.8000 ;
        RECT 2698.0000 932.8800 2699.5000 933.3600 ;
        RECT 2698.0000 954.6400 2699.5000 955.1200 ;
        RECT 2698.0000 922.0000 2699.5000 922.4800 ;
        RECT 2698.0000 916.5600 2699.5000 917.0400 ;
        RECT 2698.0000 911.1200 2699.5000 911.6000 ;
        RECT 2698.0000 905.6800 2699.5000 906.1600 ;
        RECT 2698.0000 900.2400 2699.5000 900.7200 ;
        RECT 2698.0000 894.8000 2699.5000 895.2800 ;
        RECT 2698.0000 889.3600 2699.5000 889.8400 ;
        RECT 2698.0000 883.9200 2699.5000 884.4000 ;
        RECT 2698.0000 878.4800 2699.5000 878.9600 ;
        RECT 2698.0000 873.0400 2699.5000 873.5200 ;
        RECT 2698.0000 927.4400 2699.5000 927.9200 ;
        RECT 2785.6600 867.6000 2787.1600 868.0800 ;
        RECT 2785.6600 862.1600 2787.1600 862.6400 ;
        RECT 2785.6600 856.7200 2787.1600 857.2000 ;
        RECT 2785.6600 851.2800 2787.1600 851.7600 ;
        RECT 2785.6600 845.8400 2787.1600 846.3200 ;
        RECT 2785.6600 840.4000 2787.1600 840.8800 ;
        RECT 2785.6600 834.9600 2787.1600 835.4400 ;
        RECT 2785.6600 829.5200 2787.1600 830.0000 ;
        RECT 2785.6600 824.0800 2787.1600 824.5600 ;
        RECT 2785.6600 818.6400 2787.1600 819.1200 ;
        RECT 2785.6600 813.2000 2787.1600 813.6800 ;
        RECT 2785.6600 807.7600 2787.1600 808.2400 ;
        RECT 2785.6600 802.3200 2787.1600 802.8000 ;
        RECT 2785.6600 796.8800 2787.1600 797.3600 ;
        RECT 2785.6600 791.4400 2787.1600 791.9200 ;
        RECT 2785.6600 786.0000 2787.1600 786.4800 ;
        RECT 2785.6600 780.5600 2787.1600 781.0400 ;
        RECT 2785.6600 775.1200 2787.1600 775.6000 ;
        RECT 2698.0000 867.6000 2699.5000 868.0800 ;
        RECT 2698.0000 862.1600 2699.5000 862.6400 ;
        RECT 2698.0000 856.7200 2699.5000 857.2000 ;
        RECT 2698.0000 851.2800 2699.5000 851.7600 ;
        RECT 2698.0000 845.8400 2699.5000 846.3200 ;
        RECT 2698.0000 840.4000 2699.5000 840.8800 ;
        RECT 2698.0000 834.9600 2699.5000 835.4400 ;
        RECT 2698.0000 829.5200 2699.5000 830.0000 ;
        RECT 2698.0000 824.0800 2699.5000 824.5600 ;
        RECT 2698.0000 818.6400 2699.5000 819.1200 ;
        RECT 2698.0000 813.2000 2699.5000 813.6800 ;
        RECT 2698.0000 807.7600 2699.5000 808.2400 ;
        RECT 2698.0000 802.3200 2699.5000 802.8000 ;
        RECT 2698.0000 796.8800 2699.5000 797.3600 ;
        RECT 2698.0000 791.4400 2699.5000 791.9200 ;
        RECT 2698.0000 786.0000 2699.5000 786.4800 ;
        RECT 2698.0000 780.5600 2699.5000 781.0400 ;
        RECT 2698.0000 775.1200 2699.5000 775.6000 ;
        RECT 2698.0000 974.8100 2787.1600 976.3100 ;
        RECT 2698.0000 768.2100 2787.1600 769.7100 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 245.6800 2833.6100 247.6800 2854.5400 ;
        RECT 442.7800 2833.6100 444.7800 2854.5400 ;
      LAYER met3 ;
        RECT 442.7800 2850.0400 444.7800 2850.5200 ;
        RECT 245.6800 2850.0400 247.6800 2850.5200 ;
        RECT 442.7800 2839.1600 444.7800 2839.6400 ;
        RECT 245.6800 2839.1600 247.6800 2839.6400 ;
        RECT 442.7800 2844.6000 444.7800 2845.0800 ;
        RECT 245.6800 2844.6000 247.6800 2845.0800 ;
        RECT 245.6800 2852.5400 444.7800 2854.5400 ;
        RECT 245.6800 2833.6100 444.7800 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 538.5700 431.8400 746.6700 ;
        RECT 385.2400 538.5700 386.8400 746.6700 ;
        RECT 340.2400 538.5700 341.8400 746.6700 ;
        RECT 295.2400 538.5700 296.8400 746.6700 ;
        RECT 441.7800 538.5700 444.7800 746.6700 ;
        RECT 245.6800 538.5700 248.6800 746.6700 ;
      LAYER met3 ;
        RECT 441.7800 741.3200 444.7800 741.8000 ;
        RECT 430.2400 741.3200 431.8400 741.8000 ;
        RECT 441.7800 730.4400 444.7800 730.9200 ;
        RECT 441.7800 735.8800 444.7800 736.3600 ;
        RECT 430.2400 730.4400 431.8400 730.9200 ;
        RECT 430.2400 735.8800 431.8400 736.3600 ;
        RECT 441.7800 714.1200 444.7800 714.6000 ;
        RECT 441.7800 719.5600 444.7800 720.0400 ;
        RECT 430.2400 714.1200 431.8400 714.6000 ;
        RECT 430.2400 719.5600 431.8400 720.0400 ;
        RECT 441.7800 703.2400 444.7800 703.7200 ;
        RECT 441.7800 708.6800 444.7800 709.1600 ;
        RECT 430.2400 703.2400 431.8400 703.7200 ;
        RECT 430.2400 708.6800 431.8400 709.1600 ;
        RECT 441.7800 725.0000 444.7800 725.4800 ;
        RECT 430.2400 725.0000 431.8400 725.4800 ;
        RECT 385.2400 730.4400 386.8400 730.9200 ;
        RECT 385.2400 735.8800 386.8400 736.3600 ;
        RECT 385.2400 741.3200 386.8400 741.8000 ;
        RECT 385.2400 714.1200 386.8400 714.6000 ;
        RECT 385.2400 719.5600 386.8400 720.0400 ;
        RECT 385.2400 708.6800 386.8400 709.1600 ;
        RECT 385.2400 703.2400 386.8400 703.7200 ;
        RECT 385.2400 725.0000 386.8400 725.4800 ;
        RECT 441.7800 686.9200 444.7800 687.4000 ;
        RECT 441.7800 692.3600 444.7800 692.8400 ;
        RECT 430.2400 686.9200 431.8400 687.4000 ;
        RECT 430.2400 692.3600 431.8400 692.8400 ;
        RECT 441.7800 670.6000 444.7800 671.0800 ;
        RECT 441.7800 676.0400 444.7800 676.5200 ;
        RECT 441.7800 681.4800 444.7800 681.9600 ;
        RECT 430.2400 670.6000 431.8400 671.0800 ;
        RECT 430.2400 676.0400 431.8400 676.5200 ;
        RECT 430.2400 681.4800 431.8400 681.9600 ;
        RECT 441.7800 659.7200 444.7800 660.2000 ;
        RECT 441.7800 665.1600 444.7800 665.6400 ;
        RECT 430.2400 659.7200 431.8400 660.2000 ;
        RECT 430.2400 665.1600 431.8400 665.6400 ;
        RECT 441.7800 643.4000 444.7800 643.8800 ;
        RECT 441.7800 648.8400 444.7800 649.3200 ;
        RECT 441.7800 654.2800 444.7800 654.7600 ;
        RECT 430.2400 643.4000 431.8400 643.8800 ;
        RECT 430.2400 648.8400 431.8400 649.3200 ;
        RECT 430.2400 654.2800 431.8400 654.7600 ;
        RECT 385.2400 686.9200 386.8400 687.4000 ;
        RECT 385.2400 692.3600 386.8400 692.8400 ;
        RECT 385.2400 670.6000 386.8400 671.0800 ;
        RECT 385.2400 676.0400 386.8400 676.5200 ;
        RECT 385.2400 681.4800 386.8400 681.9600 ;
        RECT 385.2400 659.7200 386.8400 660.2000 ;
        RECT 385.2400 665.1600 386.8400 665.6400 ;
        RECT 385.2400 643.4000 386.8400 643.8800 ;
        RECT 385.2400 648.8400 386.8400 649.3200 ;
        RECT 385.2400 654.2800 386.8400 654.7600 ;
        RECT 441.7800 697.8000 444.7800 698.2800 ;
        RECT 385.2400 697.8000 386.8400 698.2800 ;
        RECT 430.2400 697.8000 431.8400 698.2800 ;
        RECT 340.2400 730.4400 341.8400 730.9200 ;
        RECT 340.2400 735.8800 341.8400 736.3600 ;
        RECT 340.2400 741.3200 341.8400 741.8000 ;
        RECT 295.2400 730.4400 296.8400 730.9200 ;
        RECT 295.2400 735.8800 296.8400 736.3600 ;
        RECT 295.2400 741.3200 296.8400 741.8000 ;
        RECT 340.2400 714.1200 341.8400 714.6000 ;
        RECT 340.2400 719.5600 341.8400 720.0400 ;
        RECT 340.2400 703.2400 341.8400 703.7200 ;
        RECT 340.2400 708.6800 341.8400 709.1600 ;
        RECT 295.2400 714.1200 296.8400 714.6000 ;
        RECT 295.2400 719.5600 296.8400 720.0400 ;
        RECT 295.2400 703.2400 296.8400 703.7200 ;
        RECT 295.2400 708.6800 296.8400 709.1600 ;
        RECT 295.2400 725.0000 296.8400 725.4800 ;
        RECT 340.2400 725.0000 341.8400 725.4800 ;
        RECT 245.6800 741.3200 248.6800 741.8000 ;
        RECT 245.6800 735.8800 248.6800 736.3600 ;
        RECT 245.6800 730.4400 248.6800 730.9200 ;
        RECT 245.6800 719.5600 248.6800 720.0400 ;
        RECT 245.6800 714.1200 248.6800 714.6000 ;
        RECT 245.6800 708.6800 248.6800 709.1600 ;
        RECT 245.6800 703.2400 248.6800 703.7200 ;
        RECT 245.6800 725.0000 248.6800 725.4800 ;
        RECT 340.2400 686.9200 341.8400 687.4000 ;
        RECT 340.2400 692.3600 341.8400 692.8400 ;
        RECT 340.2400 670.6000 341.8400 671.0800 ;
        RECT 340.2400 676.0400 341.8400 676.5200 ;
        RECT 340.2400 681.4800 341.8400 681.9600 ;
        RECT 295.2400 686.9200 296.8400 687.4000 ;
        RECT 295.2400 692.3600 296.8400 692.8400 ;
        RECT 295.2400 670.6000 296.8400 671.0800 ;
        RECT 295.2400 676.0400 296.8400 676.5200 ;
        RECT 295.2400 681.4800 296.8400 681.9600 ;
        RECT 340.2400 659.7200 341.8400 660.2000 ;
        RECT 340.2400 665.1600 341.8400 665.6400 ;
        RECT 340.2400 643.4000 341.8400 643.8800 ;
        RECT 340.2400 648.8400 341.8400 649.3200 ;
        RECT 340.2400 654.2800 341.8400 654.7600 ;
        RECT 295.2400 659.7200 296.8400 660.2000 ;
        RECT 295.2400 665.1600 296.8400 665.6400 ;
        RECT 295.2400 643.4000 296.8400 643.8800 ;
        RECT 295.2400 648.8400 296.8400 649.3200 ;
        RECT 295.2400 654.2800 296.8400 654.7600 ;
        RECT 245.6800 686.9200 248.6800 687.4000 ;
        RECT 245.6800 692.3600 248.6800 692.8400 ;
        RECT 245.6800 676.0400 248.6800 676.5200 ;
        RECT 245.6800 670.6000 248.6800 671.0800 ;
        RECT 245.6800 681.4800 248.6800 681.9600 ;
        RECT 245.6800 659.7200 248.6800 660.2000 ;
        RECT 245.6800 665.1600 248.6800 665.6400 ;
        RECT 245.6800 648.8400 248.6800 649.3200 ;
        RECT 245.6800 643.4000 248.6800 643.8800 ;
        RECT 245.6800 654.2800 248.6800 654.7600 ;
        RECT 245.6800 697.8000 248.6800 698.2800 ;
        RECT 295.2400 697.8000 296.8400 698.2800 ;
        RECT 340.2400 697.8000 341.8400 698.2800 ;
        RECT 441.7800 632.5200 444.7800 633.0000 ;
        RECT 441.7800 637.9600 444.7800 638.4400 ;
        RECT 430.2400 632.5200 431.8400 633.0000 ;
        RECT 430.2400 637.9600 431.8400 638.4400 ;
        RECT 441.7800 616.2000 444.7800 616.6800 ;
        RECT 441.7800 621.6400 444.7800 622.1200 ;
        RECT 441.7800 627.0800 444.7800 627.5600 ;
        RECT 430.2400 616.2000 431.8400 616.6800 ;
        RECT 430.2400 621.6400 431.8400 622.1200 ;
        RECT 430.2400 627.0800 431.8400 627.5600 ;
        RECT 441.7800 605.3200 444.7800 605.8000 ;
        RECT 441.7800 610.7600 444.7800 611.2400 ;
        RECT 430.2400 605.3200 431.8400 605.8000 ;
        RECT 430.2400 610.7600 431.8400 611.2400 ;
        RECT 441.7800 589.0000 444.7800 589.4800 ;
        RECT 441.7800 594.4400 444.7800 594.9200 ;
        RECT 441.7800 599.8800 444.7800 600.3600 ;
        RECT 430.2400 589.0000 431.8400 589.4800 ;
        RECT 430.2400 594.4400 431.8400 594.9200 ;
        RECT 430.2400 599.8800 431.8400 600.3600 ;
        RECT 385.2400 632.5200 386.8400 633.0000 ;
        RECT 385.2400 637.9600 386.8400 638.4400 ;
        RECT 385.2400 616.2000 386.8400 616.6800 ;
        RECT 385.2400 621.6400 386.8400 622.1200 ;
        RECT 385.2400 627.0800 386.8400 627.5600 ;
        RECT 385.2400 605.3200 386.8400 605.8000 ;
        RECT 385.2400 610.7600 386.8400 611.2400 ;
        RECT 385.2400 589.0000 386.8400 589.4800 ;
        RECT 385.2400 594.4400 386.8400 594.9200 ;
        RECT 385.2400 599.8800 386.8400 600.3600 ;
        RECT 441.7800 578.1200 444.7800 578.6000 ;
        RECT 441.7800 583.5600 444.7800 584.0400 ;
        RECT 430.2400 578.1200 431.8400 578.6000 ;
        RECT 430.2400 583.5600 431.8400 584.0400 ;
        RECT 441.7800 561.8000 444.7800 562.2800 ;
        RECT 441.7800 567.2400 444.7800 567.7200 ;
        RECT 441.7800 572.6800 444.7800 573.1600 ;
        RECT 430.2400 561.8000 431.8400 562.2800 ;
        RECT 430.2400 567.2400 431.8400 567.7200 ;
        RECT 430.2400 572.6800 431.8400 573.1600 ;
        RECT 441.7800 550.9200 444.7800 551.4000 ;
        RECT 441.7800 556.3600 444.7800 556.8400 ;
        RECT 430.2400 550.9200 431.8400 551.4000 ;
        RECT 430.2400 556.3600 431.8400 556.8400 ;
        RECT 441.7800 545.4800 444.7800 545.9600 ;
        RECT 430.2400 545.4800 431.8400 545.9600 ;
        RECT 385.2400 578.1200 386.8400 578.6000 ;
        RECT 385.2400 583.5600 386.8400 584.0400 ;
        RECT 385.2400 561.8000 386.8400 562.2800 ;
        RECT 385.2400 567.2400 386.8400 567.7200 ;
        RECT 385.2400 572.6800 386.8400 573.1600 ;
        RECT 385.2400 550.9200 386.8400 551.4000 ;
        RECT 385.2400 556.3600 386.8400 556.8400 ;
        RECT 385.2400 545.4800 386.8400 545.9600 ;
        RECT 340.2400 632.5200 341.8400 633.0000 ;
        RECT 340.2400 637.9600 341.8400 638.4400 ;
        RECT 340.2400 616.2000 341.8400 616.6800 ;
        RECT 340.2400 621.6400 341.8400 622.1200 ;
        RECT 340.2400 627.0800 341.8400 627.5600 ;
        RECT 295.2400 632.5200 296.8400 633.0000 ;
        RECT 295.2400 637.9600 296.8400 638.4400 ;
        RECT 295.2400 616.2000 296.8400 616.6800 ;
        RECT 295.2400 621.6400 296.8400 622.1200 ;
        RECT 295.2400 627.0800 296.8400 627.5600 ;
        RECT 340.2400 605.3200 341.8400 605.8000 ;
        RECT 340.2400 610.7600 341.8400 611.2400 ;
        RECT 340.2400 589.0000 341.8400 589.4800 ;
        RECT 340.2400 594.4400 341.8400 594.9200 ;
        RECT 340.2400 599.8800 341.8400 600.3600 ;
        RECT 295.2400 605.3200 296.8400 605.8000 ;
        RECT 295.2400 610.7600 296.8400 611.2400 ;
        RECT 295.2400 589.0000 296.8400 589.4800 ;
        RECT 295.2400 594.4400 296.8400 594.9200 ;
        RECT 295.2400 599.8800 296.8400 600.3600 ;
        RECT 245.6800 632.5200 248.6800 633.0000 ;
        RECT 245.6800 637.9600 248.6800 638.4400 ;
        RECT 245.6800 621.6400 248.6800 622.1200 ;
        RECT 245.6800 616.2000 248.6800 616.6800 ;
        RECT 245.6800 627.0800 248.6800 627.5600 ;
        RECT 245.6800 605.3200 248.6800 605.8000 ;
        RECT 245.6800 610.7600 248.6800 611.2400 ;
        RECT 245.6800 594.4400 248.6800 594.9200 ;
        RECT 245.6800 589.0000 248.6800 589.4800 ;
        RECT 245.6800 599.8800 248.6800 600.3600 ;
        RECT 340.2400 578.1200 341.8400 578.6000 ;
        RECT 340.2400 583.5600 341.8400 584.0400 ;
        RECT 340.2400 561.8000 341.8400 562.2800 ;
        RECT 340.2400 567.2400 341.8400 567.7200 ;
        RECT 340.2400 572.6800 341.8400 573.1600 ;
        RECT 295.2400 578.1200 296.8400 578.6000 ;
        RECT 295.2400 583.5600 296.8400 584.0400 ;
        RECT 295.2400 561.8000 296.8400 562.2800 ;
        RECT 295.2400 567.2400 296.8400 567.7200 ;
        RECT 295.2400 572.6800 296.8400 573.1600 ;
        RECT 340.2400 556.3600 341.8400 556.8400 ;
        RECT 340.2400 550.9200 341.8400 551.4000 ;
        RECT 340.2400 545.4800 341.8400 545.9600 ;
        RECT 295.2400 556.3600 296.8400 556.8400 ;
        RECT 295.2400 550.9200 296.8400 551.4000 ;
        RECT 295.2400 545.4800 296.8400 545.9600 ;
        RECT 245.6800 578.1200 248.6800 578.6000 ;
        RECT 245.6800 583.5600 248.6800 584.0400 ;
        RECT 245.6800 567.2400 248.6800 567.7200 ;
        RECT 245.6800 561.8000 248.6800 562.2800 ;
        RECT 245.6800 572.6800 248.6800 573.1600 ;
        RECT 245.6800 550.9200 248.6800 551.4000 ;
        RECT 245.6800 556.3600 248.6800 556.8400 ;
        RECT 245.6800 545.4800 248.6800 545.9600 ;
        RECT 245.6800 743.6700 444.7800 746.6700 ;
        RECT 245.6800 538.5700 444.7800 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 308.9300 431.8400 517.0300 ;
        RECT 385.2400 308.9300 386.8400 517.0300 ;
        RECT 340.2400 308.9300 341.8400 517.0300 ;
        RECT 295.2400 308.9300 296.8400 517.0300 ;
        RECT 441.7800 308.9300 444.7800 517.0300 ;
        RECT 245.6800 308.9300 248.6800 517.0300 ;
      LAYER met3 ;
        RECT 441.7800 511.6800 444.7800 512.1600 ;
        RECT 430.2400 511.6800 431.8400 512.1600 ;
        RECT 441.7800 500.8000 444.7800 501.2800 ;
        RECT 441.7800 506.2400 444.7800 506.7200 ;
        RECT 430.2400 500.8000 431.8400 501.2800 ;
        RECT 430.2400 506.2400 431.8400 506.7200 ;
        RECT 441.7800 484.4800 444.7800 484.9600 ;
        RECT 441.7800 489.9200 444.7800 490.4000 ;
        RECT 430.2400 484.4800 431.8400 484.9600 ;
        RECT 430.2400 489.9200 431.8400 490.4000 ;
        RECT 441.7800 473.6000 444.7800 474.0800 ;
        RECT 441.7800 479.0400 444.7800 479.5200 ;
        RECT 430.2400 473.6000 431.8400 474.0800 ;
        RECT 430.2400 479.0400 431.8400 479.5200 ;
        RECT 441.7800 495.3600 444.7800 495.8400 ;
        RECT 430.2400 495.3600 431.8400 495.8400 ;
        RECT 385.2400 500.8000 386.8400 501.2800 ;
        RECT 385.2400 506.2400 386.8400 506.7200 ;
        RECT 385.2400 511.6800 386.8400 512.1600 ;
        RECT 385.2400 484.4800 386.8400 484.9600 ;
        RECT 385.2400 489.9200 386.8400 490.4000 ;
        RECT 385.2400 479.0400 386.8400 479.5200 ;
        RECT 385.2400 473.6000 386.8400 474.0800 ;
        RECT 385.2400 495.3600 386.8400 495.8400 ;
        RECT 441.7800 457.2800 444.7800 457.7600 ;
        RECT 441.7800 462.7200 444.7800 463.2000 ;
        RECT 430.2400 457.2800 431.8400 457.7600 ;
        RECT 430.2400 462.7200 431.8400 463.2000 ;
        RECT 441.7800 440.9600 444.7800 441.4400 ;
        RECT 441.7800 446.4000 444.7800 446.8800 ;
        RECT 441.7800 451.8400 444.7800 452.3200 ;
        RECT 430.2400 440.9600 431.8400 441.4400 ;
        RECT 430.2400 446.4000 431.8400 446.8800 ;
        RECT 430.2400 451.8400 431.8400 452.3200 ;
        RECT 441.7800 430.0800 444.7800 430.5600 ;
        RECT 441.7800 435.5200 444.7800 436.0000 ;
        RECT 430.2400 430.0800 431.8400 430.5600 ;
        RECT 430.2400 435.5200 431.8400 436.0000 ;
        RECT 441.7800 413.7600 444.7800 414.2400 ;
        RECT 441.7800 419.2000 444.7800 419.6800 ;
        RECT 441.7800 424.6400 444.7800 425.1200 ;
        RECT 430.2400 413.7600 431.8400 414.2400 ;
        RECT 430.2400 419.2000 431.8400 419.6800 ;
        RECT 430.2400 424.6400 431.8400 425.1200 ;
        RECT 385.2400 457.2800 386.8400 457.7600 ;
        RECT 385.2400 462.7200 386.8400 463.2000 ;
        RECT 385.2400 440.9600 386.8400 441.4400 ;
        RECT 385.2400 446.4000 386.8400 446.8800 ;
        RECT 385.2400 451.8400 386.8400 452.3200 ;
        RECT 385.2400 430.0800 386.8400 430.5600 ;
        RECT 385.2400 435.5200 386.8400 436.0000 ;
        RECT 385.2400 413.7600 386.8400 414.2400 ;
        RECT 385.2400 419.2000 386.8400 419.6800 ;
        RECT 385.2400 424.6400 386.8400 425.1200 ;
        RECT 441.7800 468.1600 444.7800 468.6400 ;
        RECT 385.2400 468.1600 386.8400 468.6400 ;
        RECT 430.2400 468.1600 431.8400 468.6400 ;
        RECT 340.2400 500.8000 341.8400 501.2800 ;
        RECT 340.2400 506.2400 341.8400 506.7200 ;
        RECT 340.2400 511.6800 341.8400 512.1600 ;
        RECT 295.2400 500.8000 296.8400 501.2800 ;
        RECT 295.2400 506.2400 296.8400 506.7200 ;
        RECT 295.2400 511.6800 296.8400 512.1600 ;
        RECT 340.2400 484.4800 341.8400 484.9600 ;
        RECT 340.2400 489.9200 341.8400 490.4000 ;
        RECT 340.2400 473.6000 341.8400 474.0800 ;
        RECT 340.2400 479.0400 341.8400 479.5200 ;
        RECT 295.2400 484.4800 296.8400 484.9600 ;
        RECT 295.2400 489.9200 296.8400 490.4000 ;
        RECT 295.2400 473.6000 296.8400 474.0800 ;
        RECT 295.2400 479.0400 296.8400 479.5200 ;
        RECT 295.2400 495.3600 296.8400 495.8400 ;
        RECT 340.2400 495.3600 341.8400 495.8400 ;
        RECT 245.6800 511.6800 248.6800 512.1600 ;
        RECT 245.6800 506.2400 248.6800 506.7200 ;
        RECT 245.6800 500.8000 248.6800 501.2800 ;
        RECT 245.6800 489.9200 248.6800 490.4000 ;
        RECT 245.6800 484.4800 248.6800 484.9600 ;
        RECT 245.6800 479.0400 248.6800 479.5200 ;
        RECT 245.6800 473.6000 248.6800 474.0800 ;
        RECT 245.6800 495.3600 248.6800 495.8400 ;
        RECT 340.2400 457.2800 341.8400 457.7600 ;
        RECT 340.2400 462.7200 341.8400 463.2000 ;
        RECT 340.2400 440.9600 341.8400 441.4400 ;
        RECT 340.2400 446.4000 341.8400 446.8800 ;
        RECT 340.2400 451.8400 341.8400 452.3200 ;
        RECT 295.2400 457.2800 296.8400 457.7600 ;
        RECT 295.2400 462.7200 296.8400 463.2000 ;
        RECT 295.2400 440.9600 296.8400 441.4400 ;
        RECT 295.2400 446.4000 296.8400 446.8800 ;
        RECT 295.2400 451.8400 296.8400 452.3200 ;
        RECT 340.2400 430.0800 341.8400 430.5600 ;
        RECT 340.2400 435.5200 341.8400 436.0000 ;
        RECT 340.2400 413.7600 341.8400 414.2400 ;
        RECT 340.2400 419.2000 341.8400 419.6800 ;
        RECT 340.2400 424.6400 341.8400 425.1200 ;
        RECT 295.2400 430.0800 296.8400 430.5600 ;
        RECT 295.2400 435.5200 296.8400 436.0000 ;
        RECT 295.2400 413.7600 296.8400 414.2400 ;
        RECT 295.2400 419.2000 296.8400 419.6800 ;
        RECT 295.2400 424.6400 296.8400 425.1200 ;
        RECT 245.6800 457.2800 248.6800 457.7600 ;
        RECT 245.6800 462.7200 248.6800 463.2000 ;
        RECT 245.6800 446.4000 248.6800 446.8800 ;
        RECT 245.6800 440.9600 248.6800 441.4400 ;
        RECT 245.6800 451.8400 248.6800 452.3200 ;
        RECT 245.6800 430.0800 248.6800 430.5600 ;
        RECT 245.6800 435.5200 248.6800 436.0000 ;
        RECT 245.6800 419.2000 248.6800 419.6800 ;
        RECT 245.6800 413.7600 248.6800 414.2400 ;
        RECT 245.6800 424.6400 248.6800 425.1200 ;
        RECT 245.6800 468.1600 248.6800 468.6400 ;
        RECT 295.2400 468.1600 296.8400 468.6400 ;
        RECT 340.2400 468.1600 341.8400 468.6400 ;
        RECT 441.7800 402.8800 444.7800 403.3600 ;
        RECT 441.7800 408.3200 444.7800 408.8000 ;
        RECT 430.2400 402.8800 431.8400 403.3600 ;
        RECT 430.2400 408.3200 431.8400 408.8000 ;
        RECT 441.7800 386.5600 444.7800 387.0400 ;
        RECT 441.7800 392.0000 444.7800 392.4800 ;
        RECT 441.7800 397.4400 444.7800 397.9200 ;
        RECT 430.2400 386.5600 431.8400 387.0400 ;
        RECT 430.2400 392.0000 431.8400 392.4800 ;
        RECT 430.2400 397.4400 431.8400 397.9200 ;
        RECT 441.7800 375.6800 444.7800 376.1600 ;
        RECT 441.7800 381.1200 444.7800 381.6000 ;
        RECT 430.2400 375.6800 431.8400 376.1600 ;
        RECT 430.2400 381.1200 431.8400 381.6000 ;
        RECT 441.7800 359.3600 444.7800 359.8400 ;
        RECT 441.7800 364.8000 444.7800 365.2800 ;
        RECT 441.7800 370.2400 444.7800 370.7200 ;
        RECT 430.2400 359.3600 431.8400 359.8400 ;
        RECT 430.2400 364.8000 431.8400 365.2800 ;
        RECT 430.2400 370.2400 431.8400 370.7200 ;
        RECT 385.2400 402.8800 386.8400 403.3600 ;
        RECT 385.2400 408.3200 386.8400 408.8000 ;
        RECT 385.2400 386.5600 386.8400 387.0400 ;
        RECT 385.2400 392.0000 386.8400 392.4800 ;
        RECT 385.2400 397.4400 386.8400 397.9200 ;
        RECT 385.2400 375.6800 386.8400 376.1600 ;
        RECT 385.2400 381.1200 386.8400 381.6000 ;
        RECT 385.2400 359.3600 386.8400 359.8400 ;
        RECT 385.2400 364.8000 386.8400 365.2800 ;
        RECT 385.2400 370.2400 386.8400 370.7200 ;
        RECT 441.7800 348.4800 444.7800 348.9600 ;
        RECT 441.7800 353.9200 444.7800 354.4000 ;
        RECT 430.2400 348.4800 431.8400 348.9600 ;
        RECT 430.2400 353.9200 431.8400 354.4000 ;
        RECT 441.7800 332.1600 444.7800 332.6400 ;
        RECT 441.7800 337.6000 444.7800 338.0800 ;
        RECT 441.7800 343.0400 444.7800 343.5200 ;
        RECT 430.2400 332.1600 431.8400 332.6400 ;
        RECT 430.2400 337.6000 431.8400 338.0800 ;
        RECT 430.2400 343.0400 431.8400 343.5200 ;
        RECT 441.7800 321.2800 444.7800 321.7600 ;
        RECT 441.7800 326.7200 444.7800 327.2000 ;
        RECT 430.2400 321.2800 431.8400 321.7600 ;
        RECT 430.2400 326.7200 431.8400 327.2000 ;
        RECT 441.7800 315.8400 444.7800 316.3200 ;
        RECT 430.2400 315.8400 431.8400 316.3200 ;
        RECT 385.2400 348.4800 386.8400 348.9600 ;
        RECT 385.2400 353.9200 386.8400 354.4000 ;
        RECT 385.2400 332.1600 386.8400 332.6400 ;
        RECT 385.2400 337.6000 386.8400 338.0800 ;
        RECT 385.2400 343.0400 386.8400 343.5200 ;
        RECT 385.2400 321.2800 386.8400 321.7600 ;
        RECT 385.2400 326.7200 386.8400 327.2000 ;
        RECT 385.2400 315.8400 386.8400 316.3200 ;
        RECT 340.2400 402.8800 341.8400 403.3600 ;
        RECT 340.2400 408.3200 341.8400 408.8000 ;
        RECT 340.2400 386.5600 341.8400 387.0400 ;
        RECT 340.2400 392.0000 341.8400 392.4800 ;
        RECT 340.2400 397.4400 341.8400 397.9200 ;
        RECT 295.2400 402.8800 296.8400 403.3600 ;
        RECT 295.2400 408.3200 296.8400 408.8000 ;
        RECT 295.2400 386.5600 296.8400 387.0400 ;
        RECT 295.2400 392.0000 296.8400 392.4800 ;
        RECT 295.2400 397.4400 296.8400 397.9200 ;
        RECT 340.2400 375.6800 341.8400 376.1600 ;
        RECT 340.2400 381.1200 341.8400 381.6000 ;
        RECT 340.2400 359.3600 341.8400 359.8400 ;
        RECT 340.2400 364.8000 341.8400 365.2800 ;
        RECT 340.2400 370.2400 341.8400 370.7200 ;
        RECT 295.2400 375.6800 296.8400 376.1600 ;
        RECT 295.2400 381.1200 296.8400 381.6000 ;
        RECT 295.2400 359.3600 296.8400 359.8400 ;
        RECT 295.2400 364.8000 296.8400 365.2800 ;
        RECT 295.2400 370.2400 296.8400 370.7200 ;
        RECT 245.6800 402.8800 248.6800 403.3600 ;
        RECT 245.6800 408.3200 248.6800 408.8000 ;
        RECT 245.6800 392.0000 248.6800 392.4800 ;
        RECT 245.6800 386.5600 248.6800 387.0400 ;
        RECT 245.6800 397.4400 248.6800 397.9200 ;
        RECT 245.6800 375.6800 248.6800 376.1600 ;
        RECT 245.6800 381.1200 248.6800 381.6000 ;
        RECT 245.6800 364.8000 248.6800 365.2800 ;
        RECT 245.6800 359.3600 248.6800 359.8400 ;
        RECT 245.6800 370.2400 248.6800 370.7200 ;
        RECT 340.2400 348.4800 341.8400 348.9600 ;
        RECT 340.2400 353.9200 341.8400 354.4000 ;
        RECT 340.2400 332.1600 341.8400 332.6400 ;
        RECT 340.2400 337.6000 341.8400 338.0800 ;
        RECT 340.2400 343.0400 341.8400 343.5200 ;
        RECT 295.2400 348.4800 296.8400 348.9600 ;
        RECT 295.2400 353.9200 296.8400 354.4000 ;
        RECT 295.2400 332.1600 296.8400 332.6400 ;
        RECT 295.2400 337.6000 296.8400 338.0800 ;
        RECT 295.2400 343.0400 296.8400 343.5200 ;
        RECT 340.2400 326.7200 341.8400 327.2000 ;
        RECT 340.2400 321.2800 341.8400 321.7600 ;
        RECT 340.2400 315.8400 341.8400 316.3200 ;
        RECT 295.2400 326.7200 296.8400 327.2000 ;
        RECT 295.2400 321.2800 296.8400 321.7600 ;
        RECT 295.2400 315.8400 296.8400 316.3200 ;
        RECT 245.6800 348.4800 248.6800 348.9600 ;
        RECT 245.6800 353.9200 248.6800 354.4000 ;
        RECT 245.6800 337.6000 248.6800 338.0800 ;
        RECT 245.6800 332.1600 248.6800 332.6400 ;
        RECT 245.6800 343.0400 248.6800 343.5200 ;
        RECT 245.6800 321.2800 248.6800 321.7600 ;
        RECT 245.6800 326.7200 248.6800 327.2000 ;
        RECT 245.6800 315.8400 248.6800 316.3200 ;
        RECT 245.6800 514.0300 444.7800 517.0300 ;
        RECT 245.6800 308.9300 444.7800 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 79.2900 431.8400 287.3900 ;
        RECT 385.2400 79.2900 386.8400 287.3900 ;
        RECT 340.2400 79.2900 341.8400 287.3900 ;
        RECT 295.2400 79.2900 296.8400 287.3900 ;
        RECT 441.7800 79.2900 444.7800 287.3900 ;
        RECT 245.6800 79.2900 248.6800 287.3900 ;
      LAYER met3 ;
        RECT 441.7800 282.0400 444.7800 282.5200 ;
        RECT 430.2400 282.0400 431.8400 282.5200 ;
        RECT 441.7800 271.1600 444.7800 271.6400 ;
        RECT 441.7800 276.6000 444.7800 277.0800 ;
        RECT 430.2400 271.1600 431.8400 271.6400 ;
        RECT 430.2400 276.6000 431.8400 277.0800 ;
        RECT 441.7800 254.8400 444.7800 255.3200 ;
        RECT 441.7800 260.2800 444.7800 260.7600 ;
        RECT 430.2400 254.8400 431.8400 255.3200 ;
        RECT 430.2400 260.2800 431.8400 260.7600 ;
        RECT 441.7800 243.9600 444.7800 244.4400 ;
        RECT 441.7800 249.4000 444.7800 249.8800 ;
        RECT 430.2400 243.9600 431.8400 244.4400 ;
        RECT 430.2400 249.4000 431.8400 249.8800 ;
        RECT 441.7800 265.7200 444.7800 266.2000 ;
        RECT 430.2400 265.7200 431.8400 266.2000 ;
        RECT 385.2400 271.1600 386.8400 271.6400 ;
        RECT 385.2400 276.6000 386.8400 277.0800 ;
        RECT 385.2400 282.0400 386.8400 282.5200 ;
        RECT 385.2400 254.8400 386.8400 255.3200 ;
        RECT 385.2400 260.2800 386.8400 260.7600 ;
        RECT 385.2400 249.4000 386.8400 249.8800 ;
        RECT 385.2400 243.9600 386.8400 244.4400 ;
        RECT 385.2400 265.7200 386.8400 266.2000 ;
        RECT 441.7800 227.6400 444.7800 228.1200 ;
        RECT 441.7800 233.0800 444.7800 233.5600 ;
        RECT 430.2400 227.6400 431.8400 228.1200 ;
        RECT 430.2400 233.0800 431.8400 233.5600 ;
        RECT 441.7800 211.3200 444.7800 211.8000 ;
        RECT 441.7800 216.7600 444.7800 217.2400 ;
        RECT 441.7800 222.2000 444.7800 222.6800 ;
        RECT 430.2400 211.3200 431.8400 211.8000 ;
        RECT 430.2400 216.7600 431.8400 217.2400 ;
        RECT 430.2400 222.2000 431.8400 222.6800 ;
        RECT 441.7800 200.4400 444.7800 200.9200 ;
        RECT 441.7800 205.8800 444.7800 206.3600 ;
        RECT 430.2400 200.4400 431.8400 200.9200 ;
        RECT 430.2400 205.8800 431.8400 206.3600 ;
        RECT 441.7800 184.1200 444.7800 184.6000 ;
        RECT 441.7800 189.5600 444.7800 190.0400 ;
        RECT 441.7800 195.0000 444.7800 195.4800 ;
        RECT 430.2400 184.1200 431.8400 184.6000 ;
        RECT 430.2400 189.5600 431.8400 190.0400 ;
        RECT 430.2400 195.0000 431.8400 195.4800 ;
        RECT 385.2400 227.6400 386.8400 228.1200 ;
        RECT 385.2400 233.0800 386.8400 233.5600 ;
        RECT 385.2400 211.3200 386.8400 211.8000 ;
        RECT 385.2400 216.7600 386.8400 217.2400 ;
        RECT 385.2400 222.2000 386.8400 222.6800 ;
        RECT 385.2400 200.4400 386.8400 200.9200 ;
        RECT 385.2400 205.8800 386.8400 206.3600 ;
        RECT 385.2400 184.1200 386.8400 184.6000 ;
        RECT 385.2400 189.5600 386.8400 190.0400 ;
        RECT 385.2400 195.0000 386.8400 195.4800 ;
        RECT 441.7800 238.5200 444.7800 239.0000 ;
        RECT 385.2400 238.5200 386.8400 239.0000 ;
        RECT 430.2400 238.5200 431.8400 239.0000 ;
        RECT 340.2400 271.1600 341.8400 271.6400 ;
        RECT 340.2400 276.6000 341.8400 277.0800 ;
        RECT 340.2400 282.0400 341.8400 282.5200 ;
        RECT 295.2400 271.1600 296.8400 271.6400 ;
        RECT 295.2400 276.6000 296.8400 277.0800 ;
        RECT 295.2400 282.0400 296.8400 282.5200 ;
        RECT 340.2400 254.8400 341.8400 255.3200 ;
        RECT 340.2400 260.2800 341.8400 260.7600 ;
        RECT 340.2400 243.9600 341.8400 244.4400 ;
        RECT 340.2400 249.4000 341.8400 249.8800 ;
        RECT 295.2400 254.8400 296.8400 255.3200 ;
        RECT 295.2400 260.2800 296.8400 260.7600 ;
        RECT 295.2400 243.9600 296.8400 244.4400 ;
        RECT 295.2400 249.4000 296.8400 249.8800 ;
        RECT 295.2400 265.7200 296.8400 266.2000 ;
        RECT 340.2400 265.7200 341.8400 266.2000 ;
        RECT 245.6800 282.0400 248.6800 282.5200 ;
        RECT 245.6800 276.6000 248.6800 277.0800 ;
        RECT 245.6800 271.1600 248.6800 271.6400 ;
        RECT 245.6800 260.2800 248.6800 260.7600 ;
        RECT 245.6800 254.8400 248.6800 255.3200 ;
        RECT 245.6800 249.4000 248.6800 249.8800 ;
        RECT 245.6800 243.9600 248.6800 244.4400 ;
        RECT 245.6800 265.7200 248.6800 266.2000 ;
        RECT 340.2400 227.6400 341.8400 228.1200 ;
        RECT 340.2400 233.0800 341.8400 233.5600 ;
        RECT 340.2400 211.3200 341.8400 211.8000 ;
        RECT 340.2400 216.7600 341.8400 217.2400 ;
        RECT 340.2400 222.2000 341.8400 222.6800 ;
        RECT 295.2400 227.6400 296.8400 228.1200 ;
        RECT 295.2400 233.0800 296.8400 233.5600 ;
        RECT 295.2400 211.3200 296.8400 211.8000 ;
        RECT 295.2400 216.7600 296.8400 217.2400 ;
        RECT 295.2400 222.2000 296.8400 222.6800 ;
        RECT 340.2400 200.4400 341.8400 200.9200 ;
        RECT 340.2400 205.8800 341.8400 206.3600 ;
        RECT 340.2400 184.1200 341.8400 184.6000 ;
        RECT 340.2400 189.5600 341.8400 190.0400 ;
        RECT 340.2400 195.0000 341.8400 195.4800 ;
        RECT 295.2400 200.4400 296.8400 200.9200 ;
        RECT 295.2400 205.8800 296.8400 206.3600 ;
        RECT 295.2400 184.1200 296.8400 184.6000 ;
        RECT 295.2400 189.5600 296.8400 190.0400 ;
        RECT 295.2400 195.0000 296.8400 195.4800 ;
        RECT 245.6800 227.6400 248.6800 228.1200 ;
        RECT 245.6800 233.0800 248.6800 233.5600 ;
        RECT 245.6800 216.7600 248.6800 217.2400 ;
        RECT 245.6800 211.3200 248.6800 211.8000 ;
        RECT 245.6800 222.2000 248.6800 222.6800 ;
        RECT 245.6800 200.4400 248.6800 200.9200 ;
        RECT 245.6800 205.8800 248.6800 206.3600 ;
        RECT 245.6800 189.5600 248.6800 190.0400 ;
        RECT 245.6800 184.1200 248.6800 184.6000 ;
        RECT 245.6800 195.0000 248.6800 195.4800 ;
        RECT 245.6800 238.5200 248.6800 239.0000 ;
        RECT 295.2400 238.5200 296.8400 239.0000 ;
        RECT 340.2400 238.5200 341.8400 239.0000 ;
        RECT 441.7800 173.2400 444.7800 173.7200 ;
        RECT 441.7800 178.6800 444.7800 179.1600 ;
        RECT 430.2400 173.2400 431.8400 173.7200 ;
        RECT 430.2400 178.6800 431.8400 179.1600 ;
        RECT 441.7800 156.9200 444.7800 157.4000 ;
        RECT 441.7800 162.3600 444.7800 162.8400 ;
        RECT 441.7800 167.8000 444.7800 168.2800 ;
        RECT 430.2400 156.9200 431.8400 157.4000 ;
        RECT 430.2400 162.3600 431.8400 162.8400 ;
        RECT 430.2400 167.8000 431.8400 168.2800 ;
        RECT 441.7800 146.0400 444.7800 146.5200 ;
        RECT 441.7800 151.4800 444.7800 151.9600 ;
        RECT 430.2400 146.0400 431.8400 146.5200 ;
        RECT 430.2400 151.4800 431.8400 151.9600 ;
        RECT 441.7800 129.7200 444.7800 130.2000 ;
        RECT 441.7800 135.1600 444.7800 135.6400 ;
        RECT 441.7800 140.6000 444.7800 141.0800 ;
        RECT 430.2400 129.7200 431.8400 130.2000 ;
        RECT 430.2400 135.1600 431.8400 135.6400 ;
        RECT 430.2400 140.6000 431.8400 141.0800 ;
        RECT 385.2400 173.2400 386.8400 173.7200 ;
        RECT 385.2400 178.6800 386.8400 179.1600 ;
        RECT 385.2400 156.9200 386.8400 157.4000 ;
        RECT 385.2400 162.3600 386.8400 162.8400 ;
        RECT 385.2400 167.8000 386.8400 168.2800 ;
        RECT 385.2400 146.0400 386.8400 146.5200 ;
        RECT 385.2400 151.4800 386.8400 151.9600 ;
        RECT 385.2400 129.7200 386.8400 130.2000 ;
        RECT 385.2400 135.1600 386.8400 135.6400 ;
        RECT 385.2400 140.6000 386.8400 141.0800 ;
        RECT 441.7800 118.8400 444.7800 119.3200 ;
        RECT 441.7800 124.2800 444.7800 124.7600 ;
        RECT 430.2400 118.8400 431.8400 119.3200 ;
        RECT 430.2400 124.2800 431.8400 124.7600 ;
        RECT 441.7800 102.5200 444.7800 103.0000 ;
        RECT 441.7800 107.9600 444.7800 108.4400 ;
        RECT 441.7800 113.4000 444.7800 113.8800 ;
        RECT 430.2400 102.5200 431.8400 103.0000 ;
        RECT 430.2400 107.9600 431.8400 108.4400 ;
        RECT 430.2400 113.4000 431.8400 113.8800 ;
        RECT 441.7800 91.6400 444.7800 92.1200 ;
        RECT 441.7800 97.0800 444.7800 97.5600 ;
        RECT 430.2400 91.6400 431.8400 92.1200 ;
        RECT 430.2400 97.0800 431.8400 97.5600 ;
        RECT 441.7800 86.2000 444.7800 86.6800 ;
        RECT 430.2400 86.2000 431.8400 86.6800 ;
        RECT 385.2400 118.8400 386.8400 119.3200 ;
        RECT 385.2400 124.2800 386.8400 124.7600 ;
        RECT 385.2400 102.5200 386.8400 103.0000 ;
        RECT 385.2400 107.9600 386.8400 108.4400 ;
        RECT 385.2400 113.4000 386.8400 113.8800 ;
        RECT 385.2400 91.6400 386.8400 92.1200 ;
        RECT 385.2400 97.0800 386.8400 97.5600 ;
        RECT 385.2400 86.2000 386.8400 86.6800 ;
        RECT 340.2400 173.2400 341.8400 173.7200 ;
        RECT 340.2400 178.6800 341.8400 179.1600 ;
        RECT 340.2400 156.9200 341.8400 157.4000 ;
        RECT 340.2400 162.3600 341.8400 162.8400 ;
        RECT 340.2400 167.8000 341.8400 168.2800 ;
        RECT 295.2400 173.2400 296.8400 173.7200 ;
        RECT 295.2400 178.6800 296.8400 179.1600 ;
        RECT 295.2400 156.9200 296.8400 157.4000 ;
        RECT 295.2400 162.3600 296.8400 162.8400 ;
        RECT 295.2400 167.8000 296.8400 168.2800 ;
        RECT 340.2400 146.0400 341.8400 146.5200 ;
        RECT 340.2400 151.4800 341.8400 151.9600 ;
        RECT 340.2400 129.7200 341.8400 130.2000 ;
        RECT 340.2400 135.1600 341.8400 135.6400 ;
        RECT 340.2400 140.6000 341.8400 141.0800 ;
        RECT 295.2400 146.0400 296.8400 146.5200 ;
        RECT 295.2400 151.4800 296.8400 151.9600 ;
        RECT 295.2400 129.7200 296.8400 130.2000 ;
        RECT 295.2400 135.1600 296.8400 135.6400 ;
        RECT 295.2400 140.6000 296.8400 141.0800 ;
        RECT 245.6800 173.2400 248.6800 173.7200 ;
        RECT 245.6800 178.6800 248.6800 179.1600 ;
        RECT 245.6800 162.3600 248.6800 162.8400 ;
        RECT 245.6800 156.9200 248.6800 157.4000 ;
        RECT 245.6800 167.8000 248.6800 168.2800 ;
        RECT 245.6800 146.0400 248.6800 146.5200 ;
        RECT 245.6800 151.4800 248.6800 151.9600 ;
        RECT 245.6800 135.1600 248.6800 135.6400 ;
        RECT 245.6800 129.7200 248.6800 130.2000 ;
        RECT 245.6800 140.6000 248.6800 141.0800 ;
        RECT 340.2400 118.8400 341.8400 119.3200 ;
        RECT 340.2400 124.2800 341.8400 124.7600 ;
        RECT 340.2400 102.5200 341.8400 103.0000 ;
        RECT 340.2400 107.9600 341.8400 108.4400 ;
        RECT 340.2400 113.4000 341.8400 113.8800 ;
        RECT 295.2400 118.8400 296.8400 119.3200 ;
        RECT 295.2400 124.2800 296.8400 124.7600 ;
        RECT 295.2400 102.5200 296.8400 103.0000 ;
        RECT 295.2400 107.9600 296.8400 108.4400 ;
        RECT 295.2400 113.4000 296.8400 113.8800 ;
        RECT 340.2400 97.0800 341.8400 97.5600 ;
        RECT 340.2400 91.6400 341.8400 92.1200 ;
        RECT 340.2400 86.2000 341.8400 86.6800 ;
        RECT 295.2400 97.0800 296.8400 97.5600 ;
        RECT 295.2400 91.6400 296.8400 92.1200 ;
        RECT 295.2400 86.2000 296.8400 86.6800 ;
        RECT 245.6800 118.8400 248.6800 119.3200 ;
        RECT 245.6800 124.2800 248.6800 124.7600 ;
        RECT 245.6800 107.9600 248.6800 108.4400 ;
        RECT 245.6800 102.5200 248.6800 103.0000 ;
        RECT 245.6800 113.4000 248.6800 113.8800 ;
        RECT 245.6800 91.6400 248.6800 92.1200 ;
        RECT 245.6800 97.0800 248.6800 97.5600 ;
        RECT 245.6800 86.2000 248.6800 86.6800 ;
        RECT 245.6800 284.3900 444.7800 287.3900 ;
        RECT 245.6800 79.2900 444.7800 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 245.6800 37.6700 247.6800 58.6000 ;
        RECT 442.7800 37.6700 444.7800 58.6000 ;
      LAYER met3 ;
        RECT 442.7800 54.1000 444.7800 54.5800 ;
        RECT 245.6800 54.1000 247.6800 54.5800 ;
        RECT 442.7800 43.2200 444.7800 43.7000 ;
        RECT 245.6800 43.2200 247.6800 43.7000 ;
        RECT 442.7800 48.6600 444.7800 49.1400 ;
        RECT 245.6800 48.6600 247.6800 49.1400 ;
        RECT 245.6800 56.6000 444.7800 58.6000 ;
        RECT 245.6800 37.6700 444.7800 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 2605.3300 431.8400 2813.4300 ;
        RECT 385.2400 2605.3300 386.8400 2813.4300 ;
        RECT 340.2400 2605.3300 341.8400 2813.4300 ;
        RECT 295.2400 2605.3300 296.8400 2813.4300 ;
        RECT 441.7800 2605.3300 444.7800 2813.4300 ;
        RECT 245.6800 2605.3300 248.6800 2813.4300 ;
      LAYER met3 ;
        RECT 441.7800 2808.0800 444.7800 2808.5600 ;
        RECT 430.2400 2808.0800 431.8400 2808.5600 ;
        RECT 441.7800 2797.2000 444.7800 2797.6800 ;
        RECT 441.7800 2802.6400 444.7800 2803.1200 ;
        RECT 430.2400 2797.2000 431.8400 2797.6800 ;
        RECT 430.2400 2802.6400 431.8400 2803.1200 ;
        RECT 441.7800 2780.8800 444.7800 2781.3600 ;
        RECT 441.7800 2786.3200 444.7800 2786.8000 ;
        RECT 430.2400 2780.8800 431.8400 2781.3600 ;
        RECT 430.2400 2786.3200 431.8400 2786.8000 ;
        RECT 441.7800 2770.0000 444.7800 2770.4800 ;
        RECT 441.7800 2775.4400 444.7800 2775.9200 ;
        RECT 430.2400 2770.0000 431.8400 2770.4800 ;
        RECT 430.2400 2775.4400 431.8400 2775.9200 ;
        RECT 441.7800 2791.7600 444.7800 2792.2400 ;
        RECT 430.2400 2791.7600 431.8400 2792.2400 ;
        RECT 385.2400 2797.2000 386.8400 2797.6800 ;
        RECT 385.2400 2802.6400 386.8400 2803.1200 ;
        RECT 385.2400 2808.0800 386.8400 2808.5600 ;
        RECT 385.2400 2780.8800 386.8400 2781.3600 ;
        RECT 385.2400 2786.3200 386.8400 2786.8000 ;
        RECT 385.2400 2775.4400 386.8400 2775.9200 ;
        RECT 385.2400 2770.0000 386.8400 2770.4800 ;
        RECT 385.2400 2791.7600 386.8400 2792.2400 ;
        RECT 441.7800 2753.6800 444.7800 2754.1600 ;
        RECT 441.7800 2759.1200 444.7800 2759.6000 ;
        RECT 430.2400 2753.6800 431.8400 2754.1600 ;
        RECT 430.2400 2759.1200 431.8400 2759.6000 ;
        RECT 441.7800 2737.3600 444.7800 2737.8400 ;
        RECT 441.7800 2742.8000 444.7800 2743.2800 ;
        RECT 441.7800 2748.2400 444.7800 2748.7200 ;
        RECT 430.2400 2737.3600 431.8400 2737.8400 ;
        RECT 430.2400 2742.8000 431.8400 2743.2800 ;
        RECT 430.2400 2748.2400 431.8400 2748.7200 ;
        RECT 441.7800 2726.4800 444.7800 2726.9600 ;
        RECT 441.7800 2731.9200 444.7800 2732.4000 ;
        RECT 430.2400 2726.4800 431.8400 2726.9600 ;
        RECT 430.2400 2731.9200 431.8400 2732.4000 ;
        RECT 441.7800 2710.1600 444.7800 2710.6400 ;
        RECT 441.7800 2715.6000 444.7800 2716.0800 ;
        RECT 441.7800 2721.0400 444.7800 2721.5200 ;
        RECT 430.2400 2710.1600 431.8400 2710.6400 ;
        RECT 430.2400 2715.6000 431.8400 2716.0800 ;
        RECT 430.2400 2721.0400 431.8400 2721.5200 ;
        RECT 385.2400 2753.6800 386.8400 2754.1600 ;
        RECT 385.2400 2759.1200 386.8400 2759.6000 ;
        RECT 385.2400 2737.3600 386.8400 2737.8400 ;
        RECT 385.2400 2742.8000 386.8400 2743.2800 ;
        RECT 385.2400 2748.2400 386.8400 2748.7200 ;
        RECT 385.2400 2726.4800 386.8400 2726.9600 ;
        RECT 385.2400 2731.9200 386.8400 2732.4000 ;
        RECT 385.2400 2710.1600 386.8400 2710.6400 ;
        RECT 385.2400 2715.6000 386.8400 2716.0800 ;
        RECT 385.2400 2721.0400 386.8400 2721.5200 ;
        RECT 441.7800 2764.5600 444.7800 2765.0400 ;
        RECT 385.2400 2764.5600 386.8400 2765.0400 ;
        RECT 430.2400 2764.5600 431.8400 2765.0400 ;
        RECT 340.2400 2797.2000 341.8400 2797.6800 ;
        RECT 340.2400 2802.6400 341.8400 2803.1200 ;
        RECT 340.2400 2808.0800 341.8400 2808.5600 ;
        RECT 295.2400 2797.2000 296.8400 2797.6800 ;
        RECT 295.2400 2802.6400 296.8400 2803.1200 ;
        RECT 295.2400 2808.0800 296.8400 2808.5600 ;
        RECT 340.2400 2780.8800 341.8400 2781.3600 ;
        RECT 340.2400 2786.3200 341.8400 2786.8000 ;
        RECT 340.2400 2770.0000 341.8400 2770.4800 ;
        RECT 340.2400 2775.4400 341.8400 2775.9200 ;
        RECT 295.2400 2780.8800 296.8400 2781.3600 ;
        RECT 295.2400 2786.3200 296.8400 2786.8000 ;
        RECT 295.2400 2770.0000 296.8400 2770.4800 ;
        RECT 295.2400 2775.4400 296.8400 2775.9200 ;
        RECT 295.2400 2791.7600 296.8400 2792.2400 ;
        RECT 340.2400 2791.7600 341.8400 2792.2400 ;
        RECT 245.6800 2808.0800 248.6800 2808.5600 ;
        RECT 245.6800 2802.6400 248.6800 2803.1200 ;
        RECT 245.6800 2797.2000 248.6800 2797.6800 ;
        RECT 245.6800 2786.3200 248.6800 2786.8000 ;
        RECT 245.6800 2780.8800 248.6800 2781.3600 ;
        RECT 245.6800 2775.4400 248.6800 2775.9200 ;
        RECT 245.6800 2770.0000 248.6800 2770.4800 ;
        RECT 245.6800 2791.7600 248.6800 2792.2400 ;
        RECT 340.2400 2753.6800 341.8400 2754.1600 ;
        RECT 340.2400 2759.1200 341.8400 2759.6000 ;
        RECT 340.2400 2737.3600 341.8400 2737.8400 ;
        RECT 340.2400 2742.8000 341.8400 2743.2800 ;
        RECT 340.2400 2748.2400 341.8400 2748.7200 ;
        RECT 295.2400 2753.6800 296.8400 2754.1600 ;
        RECT 295.2400 2759.1200 296.8400 2759.6000 ;
        RECT 295.2400 2737.3600 296.8400 2737.8400 ;
        RECT 295.2400 2742.8000 296.8400 2743.2800 ;
        RECT 295.2400 2748.2400 296.8400 2748.7200 ;
        RECT 340.2400 2726.4800 341.8400 2726.9600 ;
        RECT 340.2400 2731.9200 341.8400 2732.4000 ;
        RECT 340.2400 2710.1600 341.8400 2710.6400 ;
        RECT 340.2400 2715.6000 341.8400 2716.0800 ;
        RECT 340.2400 2721.0400 341.8400 2721.5200 ;
        RECT 295.2400 2726.4800 296.8400 2726.9600 ;
        RECT 295.2400 2731.9200 296.8400 2732.4000 ;
        RECT 295.2400 2710.1600 296.8400 2710.6400 ;
        RECT 295.2400 2715.6000 296.8400 2716.0800 ;
        RECT 295.2400 2721.0400 296.8400 2721.5200 ;
        RECT 245.6800 2753.6800 248.6800 2754.1600 ;
        RECT 245.6800 2759.1200 248.6800 2759.6000 ;
        RECT 245.6800 2742.8000 248.6800 2743.2800 ;
        RECT 245.6800 2737.3600 248.6800 2737.8400 ;
        RECT 245.6800 2748.2400 248.6800 2748.7200 ;
        RECT 245.6800 2726.4800 248.6800 2726.9600 ;
        RECT 245.6800 2731.9200 248.6800 2732.4000 ;
        RECT 245.6800 2715.6000 248.6800 2716.0800 ;
        RECT 245.6800 2710.1600 248.6800 2710.6400 ;
        RECT 245.6800 2721.0400 248.6800 2721.5200 ;
        RECT 245.6800 2764.5600 248.6800 2765.0400 ;
        RECT 295.2400 2764.5600 296.8400 2765.0400 ;
        RECT 340.2400 2764.5600 341.8400 2765.0400 ;
        RECT 441.7800 2699.2800 444.7800 2699.7600 ;
        RECT 441.7800 2704.7200 444.7800 2705.2000 ;
        RECT 430.2400 2699.2800 431.8400 2699.7600 ;
        RECT 430.2400 2704.7200 431.8400 2705.2000 ;
        RECT 441.7800 2682.9600 444.7800 2683.4400 ;
        RECT 441.7800 2688.4000 444.7800 2688.8800 ;
        RECT 441.7800 2693.8400 444.7800 2694.3200 ;
        RECT 430.2400 2682.9600 431.8400 2683.4400 ;
        RECT 430.2400 2688.4000 431.8400 2688.8800 ;
        RECT 430.2400 2693.8400 431.8400 2694.3200 ;
        RECT 441.7800 2672.0800 444.7800 2672.5600 ;
        RECT 441.7800 2677.5200 444.7800 2678.0000 ;
        RECT 430.2400 2672.0800 431.8400 2672.5600 ;
        RECT 430.2400 2677.5200 431.8400 2678.0000 ;
        RECT 441.7800 2655.7600 444.7800 2656.2400 ;
        RECT 441.7800 2661.2000 444.7800 2661.6800 ;
        RECT 441.7800 2666.6400 444.7800 2667.1200 ;
        RECT 430.2400 2655.7600 431.8400 2656.2400 ;
        RECT 430.2400 2661.2000 431.8400 2661.6800 ;
        RECT 430.2400 2666.6400 431.8400 2667.1200 ;
        RECT 385.2400 2699.2800 386.8400 2699.7600 ;
        RECT 385.2400 2704.7200 386.8400 2705.2000 ;
        RECT 385.2400 2682.9600 386.8400 2683.4400 ;
        RECT 385.2400 2688.4000 386.8400 2688.8800 ;
        RECT 385.2400 2693.8400 386.8400 2694.3200 ;
        RECT 385.2400 2672.0800 386.8400 2672.5600 ;
        RECT 385.2400 2677.5200 386.8400 2678.0000 ;
        RECT 385.2400 2655.7600 386.8400 2656.2400 ;
        RECT 385.2400 2661.2000 386.8400 2661.6800 ;
        RECT 385.2400 2666.6400 386.8400 2667.1200 ;
        RECT 441.7800 2644.8800 444.7800 2645.3600 ;
        RECT 441.7800 2650.3200 444.7800 2650.8000 ;
        RECT 430.2400 2644.8800 431.8400 2645.3600 ;
        RECT 430.2400 2650.3200 431.8400 2650.8000 ;
        RECT 441.7800 2628.5600 444.7800 2629.0400 ;
        RECT 441.7800 2634.0000 444.7800 2634.4800 ;
        RECT 441.7800 2639.4400 444.7800 2639.9200 ;
        RECT 430.2400 2628.5600 431.8400 2629.0400 ;
        RECT 430.2400 2634.0000 431.8400 2634.4800 ;
        RECT 430.2400 2639.4400 431.8400 2639.9200 ;
        RECT 441.7800 2617.6800 444.7800 2618.1600 ;
        RECT 441.7800 2623.1200 444.7800 2623.6000 ;
        RECT 430.2400 2617.6800 431.8400 2618.1600 ;
        RECT 430.2400 2623.1200 431.8400 2623.6000 ;
        RECT 441.7800 2612.2400 444.7800 2612.7200 ;
        RECT 430.2400 2612.2400 431.8400 2612.7200 ;
        RECT 385.2400 2644.8800 386.8400 2645.3600 ;
        RECT 385.2400 2650.3200 386.8400 2650.8000 ;
        RECT 385.2400 2628.5600 386.8400 2629.0400 ;
        RECT 385.2400 2634.0000 386.8400 2634.4800 ;
        RECT 385.2400 2639.4400 386.8400 2639.9200 ;
        RECT 385.2400 2617.6800 386.8400 2618.1600 ;
        RECT 385.2400 2623.1200 386.8400 2623.6000 ;
        RECT 385.2400 2612.2400 386.8400 2612.7200 ;
        RECT 340.2400 2699.2800 341.8400 2699.7600 ;
        RECT 340.2400 2704.7200 341.8400 2705.2000 ;
        RECT 340.2400 2682.9600 341.8400 2683.4400 ;
        RECT 340.2400 2688.4000 341.8400 2688.8800 ;
        RECT 340.2400 2693.8400 341.8400 2694.3200 ;
        RECT 295.2400 2699.2800 296.8400 2699.7600 ;
        RECT 295.2400 2704.7200 296.8400 2705.2000 ;
        RECT 295.2400 2682.9600 296.8400 2683.4400 ;
        RECT 295.2400 2688.4000 296.8400 2688.8800 ;
        RECT 295.2400 2693.8400 296.8400 2694.3200 ;
        RECT 340.2400 2672.0800 341.8400 2672.5600 ;
        RECT 340.2400 2677.5200 341.8400 2678.0000 ;
        RECT 340.2400 2655.7600 341.8400 2656.2400 ;
        RECT 340.2400 2661.2000 341.8400 2661.6800 ;
        RECT 340.2400 2666.6400 341.8400 2667.1200 ;
        RECT 295.2400 2672.0800 296.8400 2672.5600 ;
        RECT 295.2400 2677.5200 296.8400 2678.0000 ;
        RECT 295.2400 2655.7600 296.8400 2656.2400 ;
        RECT 295.2400 2661.2000 296.8400 2661.6800 ;
        RECT 295.2400 2666.6400 296.8400 2667.1200 ;
        RECT 245.6800 2699.2800 248.6800 2699.7600 ;
        RECT 245.6800 2704.7200 248.6800 2705.2000 ;
        RECT 245.6800 2688.4000 248.6800 2688.8800 ;
        RECT 245.6800 2682.9600 248.6800 2683.4400 ;
        RECT 245.6800 2693.8400 248.6800 2694.3200 ;
        RECT 245.6800 2672.0800 248.6800 2672.5600 ;
        RECT 245.6800 2677.5200 248.6800 2678.0000 ;
        RECT 245.6800 2661.2000 248.6800 2661.6800 ;
        RECT 245.6800 2655.7600 248.6800 2656.2400 ;
        RECT 245.6800 2666.6400 248.6800 2667.1200 ;
        RECT 340.2400 2644.8800 341.8400 2645.3600 ;
        RECT 340.2400 2650.3200 341.8400 2650.8000 ;
        RECT 340.2400 2628.5600 341.8400 2629.0400 ;
        RECT 340.2400 2634.0000 341.8400 2634.4800 ;
        RECT 340.2400 2639.4400 341.8400 2639.9200 ;
        RECT 295.2400 2644.8800 296.8400 2645.3600 ;
        RECT 295.2400 2650.3200 296.8400 2650.8000 ;
        RECT 295.2400 2628.5600 296.8400 2629.0400 ;
        RECT 295.2400 2634.0000 296.8400 2634.4800 ;
        RECT 295.2400 2639.4400 296.8400 2639.9200 ;
        RECT 340.2400 2623.1200 341.8400 2623.6000 ;
        RECT 340.2400 2617.6800 341.8400 2618.1600 ;
        RECT 340.2400 2612.2400 341.8400 2612.7200 ;
        RECT 295.2400 2623.1200 296.8400 2623.6000 ;
        RECT 295.2400 2617.6800 296.8400 2618.1600 ;
        RECT 295.2400 2612.2400 296.8400 2612.7200 ;
        RECT 245.6800 2644.8800 248.6800 2645.3600 ;
        RECT 245.6800 2650.3200 248.6800 2650.8000 ;
        RECT 245.6800 2634.0000 248.6800 2634.4800 ;
        RECT 245.6800 2628.5600 248.6800 2629.0400 ;
        RECT 245.6800 2639.4400 248.6800 2639.9200 ;
        RECT 245.6800 2617.6800 248.6800 2618.1600 ;
        RECT 245.6800 2623.1200 248.6800 2623.6000 ;
        RECT 245.6800 2612.2400 248.6800 2612.7200 ;
        RECT 245.6800 2810.4300 444.7800 2813.4300 ;
        RECT 245.6800 2605.3300 444.7800 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 2375.6900 431.8400 2583.7900 ;
        RECT 385.2400 2375.6900 386.8400 2583.7900 ;
        RECT 340.2400 2375.6900 341.8400 2583.7900 ;
        RECT 295.2400 2375.6900 296.8400 2583.7900 ;
        RECT 441.7800 2375.6900 444.7800 2583.7900 ;
        RECT 245.6800 2375.6900 248.6800 2583.7900 ;
      LAYER met3 ;
        RECT 441.7800 2578.4400 444.7800 2578.9200 ;
        RECT 430.2400 2578.4400 431.8400 2578.9200 ;
        RECT 441.7800 2567.5600 444.7800 2568.0400 ;
        RECT 441.7800 2573.0000 444.7800 2573.4800 ;
        RECT 430.2400 2567.5600 431.8400 2568.0400 ;
        RECT 430.2400 2573.0000 431.8400 2573.4800 ;
        RECT 441.7800 2551.2400 444.7800 2551.7200 ;
        RECT 441.7800 2556.6800 444.7800 2557.1600 ;
        RECT 430.2400 2551.2400 431.8400 2551.7200 ;
        RECT 430.2400 2556.6800 431.8400 2557.1600 ;
        RECT 441.7800 2540.3600 444.7800 2540.8400 ;
        RECT 441.7800 2545.8000 444.7800 2546.2800 ;
        RECT 430.2400 2540.3600 431.8400 2540.8400 ;
        RECT 430.2400 2545.8000 431.8400 2546.2800 ;
        RECT 441.7800 2562.1200 444.7800 2562.6000 ;
        RECT 430.2400 2562.1200 431.8400 2562.6000 ;
        RECT 385.2400 2567.5600 386.8400 2568.0400 ;
        RECT 385.2400 2573.0000 386.8400 2573.4800 ;
        RECT 385.2400 2578.4400 386.8400 2578.9200 ;
        RECT 385.2400 2551.2400 386.8400 2551.7200 ;
        RECT 385.2400 2556.6800 386.8400 2557.1600 ;
        RECT 385.2400 2545.8000 386.8400 2546.2800 ;
        RECT 385.2400 2540.3600 386.8400 2540.8400 ;
        RECT 385.2400 2562.1200 386.8400 2562.6000 ;
        RECT 441.7800 2524.0400 444.7800 2524.5200 ;
        RECT 441.7800 2529.4800 444.7800 2529.9600 ;
        RECT 430.2400 2524.0400 431.8400 2524.5200 ;
        RECT 430.2400 2529.4800 431.8400 2529.9600 ;
        RECT 441.7800 2507.7200 444.7800 2508.2000 ;
        RECT 441.7800 2513.1600 444.7800 2513.6400 ;
        RECT 441.7800 2518.6000 444.7800 2519.0800 ;
        RECT 430.2400 2507.7200 431.8400 2508.2000 ;
        RECT 430.2400 2513.1600 431.8400 2513.6400 ;
        RECT 430.2400 2518.6000 431.8400 2519.0800 ;
        RECT 441.7800 2496.8400 444.7800 2497.3200 ;
        RECT 441.7800 2502.2800 444.7800 2502.7600 ;
        RECT 430.2400 2496.8400 431.8400 2497.3200 ;
        RECT 430.2400 2502.2800 431.8400 2502.7600 ;
        RECT 441.7800 2480.5200 444.7800 2481.0000 ;
        RECT 441.7800 2485.9600 444.7800 2486.4400 ;
        RECT 441.7800 2491.4000 444.7800 2491.8800 ;
        RECT 430.2400 2480.5200 431.8400 2481.0000 ;
        RECT 430.2400 2485.9600 431.8400 2486.4400 ;
        RECT 430.2400 2491.4000 431.8400 2491.8800 ;
        RECT 385.2400 2524.0400 386.8400 2524.5200 ;
        RECT 385.2400 2529.4800 386.8400 2529.9600 ;
        RECT 385.2400 2507.7200 386.8400 2508.2000 ;
        RECT 385.2400 2513.1600 386.8400 2513.6400 ;
        RECT 385.2400 2518.6000 386.8400 2519.0800 ;
        RECT 385.2400 2496.8400 386.8400 2497.3200 ;
        RECT 385.2400 2502.2800 386.8400 2502.7600 ;
        RECT 385.2400 2480.5200 386.8400 2481.0000 ;
        RECT 385.2400 2485.9600 386.8400 2486.4400 ;
        RECT 385.2400 2491.4000 386.8400 2491.8800 ;
        RECT 441.7800 2534.9200 444.7800 2535.4000 ;
        RECT 385.2400 2534.9200 386.8400 2535.4000 ;
        RECT 430.2400 2534.9200 431.8400 2535.4000 ;
        RECT 340.2400 2567.5600 341.8400 2568.0400 ;
        RECT 340.2400 2573.0000 341.8400 2573.4800 ;
        RECT 340.2400 2578.4400 341.8400 2578.9200 ;
        RECT 295.2400 2567.5600 296.8400 2568.0400 ;
        RECT 295.2400 2573.0000 296.8400 2573.4800 ;
        RECT 295.2400 2578.4400 296.8400 2578.9200 ;
        RECT 340.2400 2551.2400 341.8400 2551.7200 ;
        RECT 340.2400 2556.6800 341.8400 2557.1600 ;
        RECT 340.2400 2540.3600 341.8400 2540.8400 ;
        RECT 340.2400 2545.8000 341.8400 2546.2800 ;
        RECT 295.2400 2551.2400 296.8400 2551.7200 ;
        RECT 295.2400 2556.6800 296.8400 2557.1600 ;
        RECT 295.2400 2540.3600 296.8400 2540.8400 ;
        RECT 295.2400 2545.8000 296.8400 2546.2800 ;
        RECT 295.2400 2562.1200 296.8400 2562.6000 ;
        RECT 340.2400 2562.1200 341.8400 2562.6000 ;
        RECT 245.6800 2578.4400 248.6800 2578.9200 ;
        RECT 245.6800 2573.0000 248.6800 2573.4800 ;
        RECT 245.6800 2567.5600 248.6800 2568.0400 ;
        RECT 245.6800 2556.6800 248.6800 2557.1600 ;
        RECT 245.6800 2551.2400 248.6800 2551.7200 ;
        RECT 245.6800 2545.8000 248.6800 2546.2800 ;
        RECT 245.6800 2540.3600 248.6800 2540.8400 ;
        RECT 245.6800 2562.1200 248.6800 2562.6000 ;
        RECT 340.2400 2524.0400 341.8400 2524.5200 ;
        RECT 340.2400 2529.4800 341.8400 2529.9600 ;
        RECT 340.2400 2507.7200 341.8400 2508.2000 ;
        RECT 340.2400 2513.1600 341.8400 2513.6400 ;
        RECT 340.2400 2518.6000 341.8400 2519.0800 ;
        RECT 295.2400 2524.0400 296.8400 2524.5200 ;
        RECT 295.2400 2529.4800 296.8400 2529.9600 ;
        RECT 295.2400 2507.7200 296.8400 2508.2000 ;
        RECT 295.2400 2513.1600 296.8400 2513.6400 ;
        RECT 295.2400 2518.6000 296.8400 2519.0800 ;
        RECT 340.2400 2496.8400 341.8400 2497.3200 ;
        RECT 340.2400 2502.2800 341.8400 2502.7600 ;
        RECT 340.2400 2480.5200 341.8400 2481.0000 ;
        RECT 340.2400 2485.9600 341.8400 2486.4400 ;
        RECT 340.2400 2491.4000 341.8400 2491.8800 ;
        RECT 295.2400 2496.8400 296.8400 2497.3200 ;
        RECT 295.2400 2502.2800 296.8400 2502.7600 ;
        RECT 295.2400 2480.5200 296.8400 2481.0000 ;
        RECT 295.2400 2485.9600 296.8400 2486.4400 ;
        RECT 295.2400 2491.4000 296.8400 2491.8800 ;
        RECT 245.6800 2524.0400 248.6800 2524.5200 ;
        RECT 245.6800 2529.4800 248.6800 2529.9600 ;
        RECT 245.6800 2513.1600 248.6800 2513.6400 ;
        RECT 245.6800 2507.7200 248.6800 2508.2000 ;
        RECT 245.6800 2518.6000 248.6800 2519.0800 ;
        RECT 245.6800 2496.8400 248.6800 2497.3200 ;
        RECT 245.6800 2502.2800 248.6800 2502.7600 ;
        RECT 245.6800 2485.9600 248.6800 2486.4400 ;
        RECT 245.6800 2480.5200 248.6800 2481.0000 ;
        RECT 245.6800 2491.4000 248.6800 2491.8800 ;
        RECT 245.6800 2534.9200 248.6800 2535.4000 ;
        RECT 295.2400 2534.9200 296.8400 2535.4000 ;
        RECT 340.2400 2534.9200 341.8400 2535.4000 ;
        RECT 441.7800 2469.6400 444.7800 2470.1200 ;
        RECT 441.7800 2475.0800 444.7800 2475.5600 ;
        RECT 430.2400 2469.6400 431.8400 2470.1200 ;
        RECT 430.2400 2475.0800 431.8400 2475.5600 ;
        RECT 441.7800 2453.3200 444.7800 2453.8000 ;
        RECT 441.7800 2458.7600 444.7800 2459.2400 ;
        RECT 441.7800 2464.2000 444.7800 2464.6800 ;
        RECT 430.2400 2453.3200 431.8400 2453.8000 ;
        RECT 430.2400 2458.7600 431.8400 2459.2400 ;
        RECT 430.2400 2464.2000 431.8400 2464.6800 ;
        RECT 441.7800 2442.4400 444.7800 2442.9200 ;
        RECT 441.7800 2447.8800 444.7800 2448.3600 ;
        RECT 430.2400 2442.4400 431.8400 2442.9200 ;
        RECT 430.2400 2447.8800 431.8400 2448.3600 ;
        RECT 441.7800 2426.1200 444.7800 2426.6000 ;
        RECT 441.7800 2431.5600 444.7800 2432.0400 ;
        RECT 441.7800 2437.0000 444.7800 2437.4800 ;
        RECT 430.2400 2426.1200 431.8400 2426.6000 ;
        RECT 430.2400 2431.5600 431.8400 2432.0400 ;
        RECT 430.2400 2437.0000 431.8400 2437.4800 ;
        RECT 385.2400 2469.6400 386.8400 2470.1200 ;
        RECT 385.2400 2475.0800 386.8400 2475.5600 ;
        RECT 385.2400 2453.3200 386.8400 2453.8000 ;
        RECT 385.2400 2458.7600 386.8400 2459.2400 ;
        RECT 385.2400 2464.2000 386.8400 2464.6800 ;
        RECT 385.2400 2442.4400 386.8400 2442.9200 ;
        RECT 385.2400 2447.8800 386.8400 2448.3600 ;
        RECT 385.2400 2426.1200 386.8400 2426.6000 ;
        RECT 385.2400 2431.5600 386.8400 2432.0400 ;
        RECT 385.2400 2437.0000 386.8400 2437.4800 ;
        RECT 441.7800 2415.2400 444.7800 2415.7200 ;
        RECT 441.7800 2420.6800 444.7800 2421.1600 ;
        RECT 430.2400 2415.2400 431.8400 2415.7200 ;
        RECT 430.2400 2420.6800 431.8400 2421.1600 ;
        RECT 441.7800 2398.9200 444.7800 2399.4000 ;
        RECT 441.7800 2404.3600 444.7800 2404.8400 ;
        RECT 441.7800 2409.8000 444.7800 2410.2800 ;
        RECT 430.2400 2398.9200 431.8400 2399.4000 ;
        RECT 430.2400 2404.3600 431.8400 2404.8400 ;
        RECT 430.2400 2409.8000 431.8400 2410.2800 ;
        RECT 441.7800 2388.0400 444.7800 2388.5200 ;
        RECT 441.7800 2393.4800 444.7800 2393.9600 ;
        RECT 430.2400 2388.0400 431.8400 2388.5200 ;
        RECT 430.2400 2393.4800 431.8400 2393.9600 ;
        RECT 441.7800 2382.6000 444.7800 2383.0800 ;
        RECT 430.2400 2382.6000 431.8400 2383.0800 ;
        RECT 385.2400 2415.2400 386.8400 2415.7200 ;
        RECT 385.2400 2420.6800 386.8400 2421.1600 ;
        RECT 385.2400 2398.9200 386.8400 2399.4000 ;
        RECT 385.2400 2404.3600 386.8400 2404.8400 ;
        RECT 385.2400 2409.8000 386.8400 2410.2800 ;
        RECT 385.2400 2388.0400 386.8400 2388.5200 ;
        RECT 385.2400 2393.4800 386.8400 2393.9600 ;
        RECT 385.2400 2382.6000 386.8400 2383.0800 ;
        RECT 340.2400 2469.6400 341.8400 2470.1200 ;
        RECT 340.2400 2475.0800 341.8400 2475.5600 ;
        RECT 340.2400 2453.3200 341.8400 2453.8000 ;
        RECT 340.2400 2458.7600 341.8400 2459.2400 ;
        RECT 340.2400 2464.2000 341.8400 2464.6800 ;
        RECT 295.2400 2469.6400 296.8400 2470.1200 ;
        RECT 295.2400 2475.0800 296.8400 2475.5600 ;
        RECT 295.2400 2453.3200 296.8400 2453.8000 ;
        RECT 295.2400 2458.7600 296.8400 2459.2400 ;
        RECT 295.2400 2464.2000 296.8400 2464.6800 ;
        RECT 340.2400 2442.4400 341.8400 2442.9200 ;
        RECT 340.2400 2447.8800 341.8400 2448.3600 ;
        RECT 340.2400 2426.1200 341.8400 2426.6000 ;
        RECT 340.2400 2431.5600 341.8400 2432.0400 ;
        RECT 340.2400 2437.0000 341.8400 2437.4800 ;
        RECT 295.2400 2442.4400 296.8400 2442.9200 ;
        RECT 295.2400 2447.8800 296.8400 2448.3600 ;
        RECT 295.2400 2426.1200 296.8400 2426.6000 ;
        RECT 295.2400 2431.5600 296.8400 2432.0400 ;
        RECT 295.2400 2437.0000 296.8400 2437.4800 ;
        RECT 245.6800 2469.6400 248.6800 2470.1200 ;
        RECT 245.6800 2475.0800 248.6800 2475.5600 ;
        RECT 245.6800 2458.7600 248.6800 2459.2400 ;
        RECT 245.6800 2453.3200 248.6800 2453.8000 ;
        RECT 245.6800 2464.2000 248.6800 2464.6800 ;
        RECT 245.6800 2442.4400 248.6800 2442.9200 ;
        RECT 245.6800 2447.8800 248.6800 2448.3600 ;
        RECT 245.6800 2431.5600 248.6800 2432.0400 ;
        RECT 245.6800 2426.1200 248.6800 2426.6000 ;
        RECT 245.6800 2437.0000 248.6800 2437.4800 ;
        RECT 340.2400 2415.2400 341.8400 2415.7200 ;
        RECT 340.2400 2420.6800 341.8400 2421.1600 ;
        RECT 340.2400 2398.9200 341.8400 2399.4000 ;
        RECT 340.2400 2404.3600 341.8400 2404.8400 ;
        RECT 340.2400 2409.8000 341.8400 2410.2800 ;
        RECT 295.2400 2415.2400 296.8400 2415.7200 ;
        RECT 295.2400 2420.6800 296.8400 2421.1600 ;
        RECT 295.2400 2398.9200 296.8400 2399.4000 ;
        RECT 295.2400 2404.3600 296.8400 2404.8400 ;
        RECT 295.2400 2409.8000 296.8400 2410.2800 ;
        RECT 340.2400 2393.4800 341.8400 2393.9600 ;
        RECT 340.2400 2388.0400 341.8400 2388.5200 ;
        RECT 340.2400 2382.6000 341.8400 2383.0800 ;
        RECT 295.2400 2393.4800 296.8400 2393.9600 ;
        RECT 295.2400 2388.0400 296.8400 2388.5200 ;
        RECT 295.2400 2382.6000 296.8400 2383.0800 ;
        RECT 245.6800 2415.2400 248.6800 2415.7200 ;
        RECT 245.6800 2420.6800 248.6800 2421.1600 ;
        RECT 245.6800 2404.3600 248.6800 2404.8400 ;
        RECT 245.6800 2398.9200 248.6800 2399.4000 ;
        RECT 245.6800 2409.8000 248.6800 2410.2800 ;
        RECT 245.6800 2388.0400 248.6800 2388.5200 ;
        RECT 245.6800 2393.4800 248.6800 2393.9600 ;
        RECT 245.6800 2382.6000 248.6800 2383.0800 ;
        RECT 245.6800 2580.7900 444.7800 2583.7900 ;
        RECT 245.6800 2375.6900 444.7800 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 2146.0500 431.8400 2354.1500 ;
        RECT 385.2400 2146.0500 386.8400 2354.1500 ;
        RECT 340.2400 2146.0500 341.8400 2354.1500 ;
        RECT 295.2400 2146.0500 296.8400 2354.1500 ;
        RECT 441.7800 2146.0500 444.7800 2354.1500 ;
        RECT 245.6800 2146.0500 248.6800 2354.1500 ;
      LAYER met3 ;
        RECT 441.7800 2348.8000 444.7800 2349.2800 ;
        RECT 430.2400 2348.8000 431.8400 2349.2800 ;
        RECT 441.7800 2337.9200 444.7800 2338.4000 ;
        RECT 441.7800 2343.3600 444.7800 2343.8400 ;
        RECT 430.2400 2337.9200 431.8400 2338.4000 ;
        RECT 430.2400 2343.3600 431.8400 2343.8400 ;
        RECT 441.7800 2321.6000 444.7800 2322.0800 ;
        RECT 441.7800 2327.0400 444.7800 2327.5200 ;
        RECT 430.2400 2321.6000 431.8400 2322.0800 ;
        RECT 430.2400 2327.0400 431.8400 2327.5200 ;
        RECT 441.7800 2310.7200 444.7800 2311.2000 ;
        RECT 441.7800 2316.1600 444.7800 2316.6400 ;
        RECT 430.2400 2310.7200 431.8400 2311.2000 ;
        RECT 430.2400 2316.1600 431.8400 2316.6400 ;
        RECT 441.7800 2332.4800 444.7800 2332.9600 ;
        RECT 430.2400 2332.4800 431.8400 2332.9600 ;
        RECT 385.2400 2337.9200 386.8400 2338.4000 ;
        RECT 385.2400 2343.3600 386.8400 2343.8400 ;
        RECT 385.2400 2348.8000 386.8400 2349.2800 ;
        RECT 385.2400 2321.6000 386.8400 2322.0800 ;
        RECT 385.2400 2327.0400 386.8400 2327.5200 ;
        RECT 385.2400 2316.1600 386.8400 2316.6400 ;
        RECT 385.2400 2310.7200 386.8400 2311.2000 ;
        RECT 385.2400 2332.4800 386.8400 2332.9600 ;
        RECT 441.7800 2294.4000 444.7800 2294.8800 ;
        RECT 441.7800 2299.8400 444.7800 2300.3200 ;
        RECT 430.2400 2294.4000 431.8400 2294.8800 ;
        RECT 430.2400 2299.8400 431.8400 2300.3200 ;
        RECT 441.7800 2278.0800 444.7800 2278.5600 ;
        RECT 441.7800 2283.5200 444.7800 2284.0000 ;
        RECT 441.7800 2288.9600 444.7800 2289.4400 ;
        RECT 430.2400 2278.0800 431.8400 2278.5600 ;
        RECT 430.2400 2283.5200 431.8400 2284.0000 ;
        RECT 430.2400 2288.9600 431.8400 2289.4400 ;
        RECT 441.7800 2267.2000 444.7800 2267.6800 ;
        RECT 441.7800 2272.6400 444.7800 2273.1200 ;
        RECT 430.2400 2267.2000 431.8400 2267.6800 ;
        RECT 430.2400 2272.6400 431.8400 2273.1200 ;
        RECT 441.7800 2250.8800 444.7800 2251.3600 ;
        RECT 441.7800 2256.3200 444.7800 2256.8000 ;
        RECT 441.7800 2261.7600 444.7800 2262.2400 ;
        RECT 430.2400 2250.8800 431.8400 2251.3600 ;
        RECT 430.2400 2256.3200 431.8400 2256.8000 ;
        RECT 430.2400 2261.7600 431.8400 2262.2400 ;
        RECT 385.2400 2294.4000 386.8400 2294.8800 ;
        RECT 385.2400 2299.8400 386.8400 2300.3200 ;
        RECT 385.2400 2278.0800 386.8400 2278.5600 ;
        RECT 385.2400 2283.5200 386.8400 2284.0000 ;
        RECT 385.2400 2288.9600 386.8400 2289.4400 ;
        RECT 385.2400 2267.2000 386.8400 2267.6800 ;
        RECT 385.2400 2272.6400 386.8400 2273.1200 ;
        RECT 385.2400 2250.8800 386.8400 2251.3600 ;
        RECT 385.2400 2256.3200 386.8400 2256.8000 ;
        RECT 385.2400 2261.7600 386.8400 2262.2400 ;
        RECT 441.7800 2305.2800 444.7800 2305.7600 ;
        RECT 385.2400 2305.2800 386.8400 2305.7600 ;
        RECT 430.2400 2305.2800 431.8400 2305.7600 ;
        RECT 340.2400 2337.9200 341.8400 2338.4000 ;
        RECT 340.2400 2343.3600 341.8400 2343.8400 ;
        RECT 340.2400 2348.8000 341.8400 2349.2800 ;
        RECT 295.2400 2337.9200 296.8400 2338.4000 ;
        RECT 295.2400 2343.3600 296.8400 2343.8400 ;
        RECT 295.2400 2348.8000 296.8400 2349.2800 ;
        RECT 340.2400 2321.6000 341.8400 2322.0800 ;
        RECT 340.2400 2327.0400 341.8400 2327.5200 ;
        RECT 340.2400 2310.7200 341.8400 2311.2000 ;
        RECT 340.2400 2316.1600 341.8400 2316.6400 ;
        RECT 295.2400 2321.6000 296.8400 2322.0800 ;
        RECT 295.2400 2327.0400 296.8400 2327.5200 ;
        RECT 295.2400 2310.7200 296.8400 2311.2000 ;
        RECT 295.2400 2316.1600 296.8400 2316.6400 ;
        RECT 295.2400 2332.4800 296.8400 2332.9600 ;
        RECT 340.2400 2332.4800 341.8400 2332.9600 ;
        RECT 245.6800 2348.8000 248.6800 2349.2800 ;
        RECT 245.6800 2343.3600 248.6800 2343.8400 ;
        RECT 245.6800 2337.9200 248.6800 2338.4000 ;
        RECT 245.6800 2327.0400 248.6800 2327.5200 ;
        RECT 245.6800 2321.6000 248.6800 2322.0800 ;
        RECT 245.6800 2316.1600 248.6800 2316.6400 ;
        RECT 245.6800 2310.7200 248.6800 2311.2000 ;
        RECT 245.6800 2332.4800 248.6800 2332.9600 ;
        RECT 340.2400 2294.4000 341.8400 2294.8800 ;
        RECT 340.2400 2299.8400 341.8400 2300.3200 ;
        RECT 340.2400 2278.0800 341.8400 2278.5600 ;
        RECT 340.2400 2283.5200 341.8400 2284.0000 ;
        RECT 340.2400 2288.9600 341.8400 2289.4400 ;
        RECT 295.2400 2294.4000 296.8400 2294.8800 ;
        RECT 295.2400 2299.8400 296.8400 2300.3200 ;
        RECT 295.2400 2278.0800 296.8400 2278.5600 ;
        RECT 295.2400 2283.5200 296.8400 2284.0000 ;
        RECT 295.2400 2288.9600 296.8400 2289.4400 ;
        RECT 340.2400 2267.2000 341.8400 2267.6800 ;
        RECT 340.2400 2272.6400 341.8400 2273.1200 ;
        RECT 340.2400 2250.8800 341.8400 2251.3600 ;
        RECT 340.2400 2256.3200 341.8400 2256.8000 ;
        RECT 340.2400 2261.7600 341.8400 2262.2400 ;
        RECT 295.2400 2267.2000 296.8400 2267.6800 ;
        RECT 295.2400 2272.6400 296.8400 2273.1200 ;
        RECT 295.2400 2250.8800 296.8400 2251.3600 ;
        RECT 295.2400 2256.3200 296.8400 2256.8000 ;
        RECT 295.2400 2261.7600 296.8400 2262.2400 ;
        RECT 245.6800 2294.4000 248.6800 2294.8800 ;
        RECT 245.6800 2299.8400 248.6800 2300.3200 ;
        RECT 245.6800 2283.5200 248.6800 2284.0000 ;
        RECT 245.6800 2278.0800 248.6800 2278.5600 ;
        RECT 245.6800 2288.9600 248.6800 2289.4400 ;
        RECT 245.6800 2267.2000 248.6800 2267.6800 ;
        RECT 245.6800 2272.6400 248.6800 2273.1200 ;
        RECT 245.6800 2256.3200 248.6800 2256.8000 ;
        RECT 245.6800 2250.8800 248.6800 2251.3600 ;
        RECT 245.6800 2261.7600 248.6800 2262.2400 ;
        RECT 245.6800 2305.2800 248.6800 2305.7600 ;
        RECT 295.2400 2305.2800 296.8400 2305.7600 ;
        RECT 340.2400 2305.2800 341.8400 2305.7600 ;
        RECT 441.7800 2240.0000 444.7800 2240.4800 ;
        RECT 441.7800 2245.4400 444.7800 2245.9200 ;
        RECT 430.2400 2240.0000 431.8400 2240.4800 ;
        RECT 430.2400 2245.4400 431.8400 2245.9200 ;
        RECT 441.7800 2223.6800 444.7800 2224.1600 ;
        RECT 441.7800 2229.1200 444.7800 2229.6000 ;
        RECT 441.7800 2234.5600 444.7800 2235.0400 ;
        RECT 430.2400 2223.6800 431.8400 2224.1600 ;
        RECT 430.2400 2229.1200 431.8400 2229.6000 ;
        RECT 430.2400 2234.5600 431.8400 2235.0400 ;
        RECT 441.7800 2212.8000 444.7800 2213.2800 ;
        RECT 441.7800 2218.2400 444.7800 2218.7200 ;
        RECT 430.2400 2212.8000 431.8400 2213.2800 ;
        RECT 430.2400 2218.2400 431.8400 2218.7200 ;
        RECT 441.7800 2196.4800 444.7800 2196.9600 ;
        RECT 441.7800 2201.9200 444.7800 2202.4000 ;
        RECT 441.7800 2207.3600 444.7800 2207.8400 ;
        RECT 430.2400 2196.4800 431.8400 2196.9600 ;
        RECT 430.2400 2201.9200 431.8400 2202.4000 ;
        RECT 430.2400 2207.3600 431.8400 2207.8400 ;
        RECT 385.2400 2240.0000 386.8400 2240.4800 ;
        RECT 385.2400 2245.4400 386.8400 2245.9200 ;
        RECT 385.2400 2223.6800 386.8400 2224.1600 ;
        RECT 385.2400 2229.1200 386.8400 2229.6000 ;
        RECT 385.2400 2234.5600 386.8400 2235.0400 ;
        RECT 385.2400 2212.8000 386.8400 2213.2800 ;
        RECT 385.2400 2218.2400 386.8400 2218.7200 ;
        RECT 385.2400 2196.4800 386.8400 2196.9600 ;
        RECT 385.2400 2201.9200 386.8400 2202.4000 ;
        RECT 385.2400 2207.3600 386.8400 2207.8400 ;
        RECT 441.7800 2185.6000 444.7800 2186.0800 ;
        RECT 441.7800 2191.0400 444.7800 2191.5200 ;
        RECT 430.2400 2185.6000 431.8400 2186.0800 ;
        RECT 430.2400 2191.0400 431.8400 2191.5200 ;
        RECT 441.7800 2169.2800 444.7800 2169.7600 ;
        RECT 441.7800 2174.7200 444.7800 2175.2000 ;
        RECT 441.7800 2180.1600 444.7800 2180.6400 ;
        RECT 430.2400 2169.2800 431.8400 2169.7600 ;
        RECT 430.2400 2174.7200 431.8400 2175.2000 ;
        RECT 430.2400 2180.1600 431.8400 2180.6400 ;
        RECT 441.7800 2158.4000 444.7800 2158.8800 ;
        RECT 441.7800 2163.8400 444.7800 2164.3200 ;
        RECT 430.2400 2158.4000 431.8400 2158.8800 ;
        RECT 430.2400 2163.8400 431.8400 2164.3200 ;
        RECT 441.7800 2152.9600 444.7800 2153.4400 ;
        RECT 430.2400 2152.9600 431.8400 2153.4400 ;
        RECT 385.2400 2185.6000 386.8400 2186.0800 ;
        RECT 385.2400 2191.0400 386.8400 2191.5200 ;
        RECT 385.2400 2169.2800 386.8400 2169.7600 ;
        RECT 385.2400 2174.7200 386.8400 2175.2000 ;
        RECT 385.2400 2180.1600 386.8400 2180.6400 ;
        RECT 385.2400 2158.4000 386.8400 2158.8800 ;
        RECT 385.2400 2163.8400 386.8400 2164.3200 ;
        RECT 385.2400 2152.9600 386.8400 2153.4400 ;
        RECT 340.2400 2240.0000 341.8400 2240.4800 ;
        RECT 340.2400 2245.4400 341.8400 2245.9200 ;
        RECT 340.2400 2223.6800 341.8400 2224.1600 ;
        RECT 340.2400 2229.1200 341.8400 2229.6000 ;
        RECT 340.2400 2234.5600 341.8400 2235.0400 ;
        RECT 295.2400 2240.0000 296.8400 2240.4800 ;
        RECT 295.2400 2245.4400 296.8400 2245.9200 ;
        RECT 295.2400 2223.6800 296.8400 2224.1600 ;
        RECT 295.2400 2229.1200 296.8400 2229.6000 ;
        RECT 295.2400 2234.5600 296.8400 2235.0400 ;
        RECT 340.2400 2212.8000 341.8400 2213.2800 ;
        RECT 340.2400 2218.2400 341.8400 2218.7200 ;
        RECT 340.2400 2196.4800 341.8400 2196.9600 ;
        RECT 340.2400 2201.9200 341.8400 2202.4000 ;
        RECT 340.2400 2207.3600 341.8400 2207.8400 ;
        RECT 295.2400 2212.8000 296.8400 2213.2800 ;
        RECT 295.2400 2218.2400 296.8400 2218.7200 ;
        RECT 295.2400 2196.4800 296.8400 2196.9600 ;
        RECT 295.2400 2201.9200 296.8400 2202.4000 ;
        RECT 295.2400 2207.3600 296.8400 2207.8400 ;
        RECT 245.6800 2240.0000 248.6800 2240.4800 ;
        RECT 245.6800 2245.4400 248.6800 2245.9200 ;
        RECT 245.6800 2229.1200 248.6800 2229.6000 ;
        RECT 245.6800 2223.6800 248.6800 2224.1600 ;
        RECT 245.6800 2234.5600 248.6800 2235.0400 ;
        RECT 245.6800 2212.8000 248.6800 2213.2800 ;
        RECT 245.6800 2218.2400 248.6800 2218.7200 ;
        RECT 245.6800 2201.9200 248.6800 2202.4000 ;
        RECT 245.6800 2196.4800 248.6800 2196.9600 ;
        RECT 245.6800 2207.3600 248.6800 2207.8400 ;
        RECT 340.2400 2185.6000 341.8400 2186.0800 ;
        RECT 340.2400 2191.0400 341.8400 2191.5200 ;
        RECT 340.2400 2169.2800 341.8400 2169.7600 ;
        RECT 340.2400 2174.7200 341.8400 2175.2000 ;
        RECT 340.2400 2180.1600 341.8400 2180.6400 ;
        RECT 295.2400 2185.6000 296.8400 2186.0800 ;
        RECT 295.2400 2191.0400 296.8400 2191.5200 ;
        RECT 295.2400 2169.2800 296.8400 2169.7600 ;
        RECT 295.2400 2174.7200 296.8400 2175.2000 ;
        RECT 295.2400 2180.1600 296.8400 2180.6400 ;
        RECT 340.2400 2163.8400 341.8400 2164.3200 ;
        RECT 340.2400 2158.4000 341.8400 2158.8800 ;
        RECT 340.2400 2152.9600 341.8400 2153.4400 ;
        RECT 295.2400 2163.8400 296.8400 2164.3200 ;
        RECT 295.2400 2158.4000 296.8400 2158.8800 ;
        RECT 295.2400 2152.9600 296.8400 2153.4400 ;
        RECT 245.6800 2185.6000 248.6800 2186.0800 ;
        RECT 245.6800 2191.0400 248.6800 2191.5200 ;
        RECT 245.6800 2174.7200 248.6800 2175.2000 ;
        RECT 245.6800 2169.2800 248.6800 2169.7600 ;
        RECT 245.6800 2180.1600 248.6800 2180.6400 ;
        RECT 245.6800 2158.4000 248.6800 2158.8800 ;
        RECT 245.6800 2163.8400 248.6800 2164.3200 ;
        RECT 245.6800 2152.9600 248.6800 2153.4400 ;
        RECT 245.6800 2351.1500 444.7800 2354.1500 ;
        RECT 245.6800 2146.0500 444.7800 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 1916.4100 431.8400 2124.5100 ;
        RECT 385.2400 1916.4100 386.8400 2124.5100 ;
        RECT 340.2400 1916.4100 341.8400 2124.5100 ;
        RECT 295.2400 1916.4100 296.8400 2124.5100 ;
        RECT 441.7800 1916.4100 444.7800 2124.5100 ;
        RECT 245.6800 1916.4100 248.6800 2124.5100 ;
      LAYER met3 ;
        RECT 441.7800 2119.1600 444.7800 2119.6400 ;
        RECT 430.2400 2119.1600 431.8400 2119.6400 ;
        RECT 441.7800 2108.2800 444.7800 2108.7600 ;
        RECT 441.7800 2113.7200 444.7800 2114.2000 ;
        RECT 430.2400 2108.2800 431.8400 2108.7600 ;
        RECT 430.2400 2113.7200 431.8400 2114.2000 ;
        RECT 441.7800 2091.9600 444.7800 2092.4400 ;
        RECT 441.7800 2097.4000 444.7800 2097.8800 ;
        RECT 430.2400 2091.9600 431.8400 2092.4400 ;
        RECT 430.2400 2097.4000 431.8400 2097.8800 ;
        RECT 441.7800 2081.0800 444.7800 2081.5600 ;
        RECT 441.7800 2086.5200 444.7800 2087.0000 ;
        RECT 430.2400 2081.0800 431.8400 2081.5600 ;
        RECT 430.2400 2086.5200 431.8400 2087.0000 ;
        RECT 441.7800 2102.8400 444.7800 2103.3200 ;
        RECT 430.2400 2102.8400 431.8400 2103.3200 ;
        RECT 385.2400 2108.2800 386.8400 2108.7600 ;
        RECT 385.2400 2113.7200 386.8400 2114.2000 ;
        RECT 385.2400 2119.1600 386.8400 2119.6400 ;
        RECT 385.2400 2091.9600 386.8400 2092.4400 ;
        RECT 385.2400 2097.4000 386.8400 2097.8800 ;
        RECT 385.2400 2086.5200 386.8400 2087.0000 ;
        RECT 385.2400 2081.0800 386.8400 2081.5600 ;
        RECT 385.2400 2102.8400 386.8400 2103.3200 ;
        RECT 441.7800 2064.7600 444.7800 2065.2400 ;
        RECT 441.7800 2070.2000 444.7800 2070.6800 ;
        RECT 430.2400 2064.7600 431.8400 2065.2400 ;
        RECT 430.2400 2070.2000 431.8400 2070.6800 ;
        RECT 441.7800 2048.4400 444.7800 2048.9200 ;
        RECT 441.7800 2053.8800 444.7800 2054.3600 ;
        RECT 441.7800 2059.3200 444.7800 2059.8000 ;
        RECT 430.2400 2048.4400 431.8400 2048.9200 ;
        RECT 430.2400 2053.8800 431.8400 2054.3600 ;
        RECT 430.2400 2059.3200 431.8400 2059.8000 ;
        RECT 441.7800 2037.5600 444.7800 2038.0400 ;
        RECT 441.7800 2043.0000 444.7800 2043.4800 ;
        RECT 430.2400 2037.5600 431.8400 2038.0400 ;
        RECT 430.2400 2043.0000 431.8400 2043.4800 ;
        RECT 441.7800 2021.2400 444.7800 2021.7200 ;
        RECT 441.7800 2026.6800 444.7800 2027.1600 ;
        RECT 441.7800 2032.1200 444.7800 2032.6000 ;
        RECT 430.2400 2021.2400 431.8400 2021.7200 ;
        RECT 430.2400 2026.6800 431.8400 2027.1600 ;
        RECT 430.2400 2032.1200 431.8400 2032.6000 ;
        RECT 385.2400 2064.7600 386.8400 2065.2400 ;
        RECT 385.2400 2070.2000 386.8400 2070.6800 ;
        RECT 385.2400 2048.4400 386.8400 2048.9200 ;
        RECT 385.2400 2053.8800 386.8400 2054.3600 ;
        RECT 385.2400 2059.3200 386.8400 2059.8000 ;
        RECT 385.2400 2037.5600 386.8400 2038.0400 ;
        RECT 385.2400 2043.0000 386.8400 2043.4800 ;
        RECT 385.2400 2021.2400 386.8400 2021.7200 ;
        RECT 385.2400 2026.6800 386.8400 2027.1600 ;
        RECT 385.2400 2032.1200 386.8400 2032.6000 ;
        RECT 441.7800 2075.6400 444.7800 2076.1200 ;
        RECT 385.2400 2075.6400 386.8400 2076.1200 ;
        RECT 430.2400 2075.6400 431.8400 2076.1200 ;
        RECT 340.2400 2108.2800 341.8400 2108.7600 ;
        RECT 340.2400 2113.7200 341.8400 2114.2000 ;
        RECT 340.2400 2119.1600 341.8400 2119.6400 ;
        RECT 295.2400 2108.2800 296.8400 2108.7600 ;
        RECT 295.2400 2113.7200 296.8400 2114.2000 ;
        RECT 295.2400 2119.1600 296.8400 2119.6400 ;
        RECT 340.2400 2091.9600 341.8400 2092.4400 ;
        RECT 340.2400 2097.4000 341.8400 2097.8800 ;
        RECT 340.2400 2081.0800 341.8400 2081.5600 ;
        RECT 340.2400 2086.5200 341.8400 2087.0000 ;
        RECT 295.2400 2091.9600 296.8400 2092.4400 ;
        RECT 295.2400 2097.4000 296.8400 2097.8800 ;
        RECT 295.2400 2081.0800 296.8400 2081.5600 ;
        RECT 295.2400 2086.5200 296.8400 2087.0000 ;
        RECT 295.2400 2102.8400 296.8400 2103.3200 ;
        RECT 340.2400 2102.8400 341.8400 2103.3200 ;
        RECT 245.6800 2119.1600 248.6800 2119.6400 ;
        RECT 245.6800 2113.7200 248.6800 2114.2000 ;
        RECT 245.6800 2108.2800 248.6800 2108.7600 ;
        RECT 245.6800 2097.4000 248.6800 2097.8800 ;
        RECT 245.6800 2091.9600 248.6800 2092.4400 ;
        RECT 245.6800 2086.5200 248.6800 2087.0000 ;
        RECT 245.6800 2081.0800 248.6800 2081.5600 ;
        RECT 245.6800 2102.8400 248.6800 2103.3200 ;
        RECT 340.2400 2064.7600 341.8400 2065.2400 ;
        RECT 340.2400 2070.2000 341.8400 2070.6800 ;
        RECT 340.2400 2048.4400 341.8400 2048.9200 ;
        RECT 340.2400 2053.8800 341.8400 2054.3600 ;
        RECT 340.2400 2059.3200 341.8400 2059.8000 ;
        RECT 295.2400 2064.7600 296.8400 2065.2400 ;
        RECT 295.2400 2070.2000 296.8400 2070.6800 ;
        RECT 295.2400 2048.4400 296.8400 2048.9200 ;
        RECT 295.2400 2053.8800 296.8400 2054.3600 ;
        RECT 295.2400 2059.3200 296.8400 2059.8000 ;
        RECT 340.2400 2037.5600 341.8400 2038.0400 ;
        RECT 340.2400 2043.0000 341.8400 2043.4800 ;
        RECT 340.2400 2021.2400 341.8400 2021.7200 ;
        RECT 340.2400 2026.6800 341.8400 2027.1600 ;
        RECT 340.2400 2032.1200 341.8400 2032.6000 ;
        RECT 295.2400 2037.5600 296.8400 2038.0400 ;
        RECT 295.2400 2043.0000 296.8400 2043.4800 ;
        RECT 295.2400 2021.2400 296.8400 2021.7200 ;
        RECT 295.2400 2026.6800 296.8400 2027.1600 ;
        RECT 295.2400 2032.1200 296.8400 2032.6000 ;
        RECT 245.6800 2064.7600 248.6800 2065.2400 ;
        RECT 245.6800 2070.2000 248.6800 2070.6800 ;
        RECT 245.6800 2053.8800 248.6800 2054.3600 ;
        RECT 245.6800 2048.4400 248.6800 2048.9200 ;
        RECT 245.6800 2059.3200 248.6800 2059.8000 ;
        RECT 245.6800 2037.5600 248.6800 2038.0400 ;
        RECT 245.6800 2043.0000 248.6800 2043.4800 ;
        RECT 245.6800 2026.6800 248.6800 2027.1600 ;
        RECT 245.6800 2021.2400 248.6800 2021.7200 ;
        RECT 245.6800 2032.1200 248.6800 2032.6000 ;
        RECT 245.6800 2075.6400 248.6800 2076.1200 ;
        RECT 295.2400 2075.6400 296.8400 2076.1200 ;
        RECT 340.2400 2075.6400 341.8400 2076.1200 ;
        RECT 441.7800 2010.3600 444.7800 2010.8400 ;
        RECT 441.7800 2015.8000 444.7800 2016.2800 ;
        RECT 430.2400 2010.3600 431.8400 2010.8400 ;
        RECT 430.2400 2015.8000 431.8400 2016.2800 ;
        RECT 441.7800 1994.0400 444.7800 1994.5200 ;
        RECT 441.7800 1999.4800 444.7800 1999.9600 ;
        RECT 441.7800 2004.9200 444.7800 2005.4000 ;
        RECT 430.2400 1994.0400 431.8400 1994.5200 ;
        RECT 430.2400 1999.4800 431.8400 1999.9600 ;
        RECT 430.2400 2004.9200 431.8400 2005.4000 ;
        RECT 441.7800 1983.1600 444.7800 1983.6400 ;
        RECT 441.7800 1988.6000 444.7800 1989.0800 ;
        RECT 430.2400 1983.1600 431.8400 1983.6400 ;
        RECT 430.2400 1988.6000 431.8400 1989.0800 ;
        RECT 441.7800 1966.8400 444.7800 1967.3200 ;
        RECT 441.7800 1972.2800 444.7800 1972.7600 ;
        RECT 441.7800 1977.7200 444.7800 1978.2000 ;
        RECT 430.2400 1966.8400 431.8400 1967.3200 ;
        RECT 430.2400 1972.2800 431.8400 1972.7600 ;
        RECT 430.2400 1977.7200 431.8400 1978.2000 ;
        RECT 385.2400 2010.3600 386.8400 2010.8400 ;
        RECT 385.2400 2015.8000 386.8400 2016.2800 ;
        RECT 385.2400 1994.0400 386.8400 1994.5200 ;
        RECT 385.2400 1999.4800 386.8400 1999.9600 ;
        RECT 385.2400 2004.9200 386.8400 2005.4000 ;
        RECT 385.2400 1983.1600 386.8400 1983.6400 ;
        RECT 385.2400 1988.6000 386.8400 1989.0800 ;
        RECT 385.2400 1966.8400 386.8400 1967.3200 ;
        RECT 385.2400 1972.2800 386.8400 1972.7600 ;
        RECT 385.2400 1977.7200 386.8400 1978.2000 ;
        RECT 441.7800 1955.9600 444.7800 1956.4400 ;
        RECT 441.7800 1961.4000 444.7800 1961.8800 ;
        RECT 430.2400 1955.9600 431.8400 1956.4400 ;
        RECT 430.2400 1961.4000 431.8400 1961.8800 ;
        RECT 441.7800 1939.6400 444.7800 1940.1200 ;
        RECT 441.7800 1945.0800 444.7800 1945.5600 ;
        RECT 441.7800 1950.5200 444.7800 1951.0000 ;
        RECT 430.2400 1939.6400 431.8400 1940.1200 ;
        RECT 430.2400 1945.0800 431.8400 1945.5600 ;
        RECT 430.2400 1950.5200 431.8400 1951.0000 ;
        RECT 441.7800 1928.7600 444.7800 1929.2400 ;
        RECT 441.7800 1934.2000 444.7800 1934.6800 ;
        RECT 430.2400 1928.7600 431.8400 1929.2400 ;
        RECT 430.2400 1934.2000 431.8400 1934.6800 ;
        RECT 441.7800 1923.3200 444.7800 1923.8000 ;
        RECT 430.2400 1923.3200 431.8400 1923.8000 ;
        RECT 385.2400 1955.9600 386.8400 1956.4400 ;
        RECT 385.2400 1961.4000 386.8400 1961.8800 ;
        RECT 385.2400 1939.6400 386.8400 1940.1200 ;
        RECT 385.2400 1945.0800 386.8400 1945.5600 ;
        RECT 385.2400 1950.5200 386.8400 1951.0000 ;
        RECT 385.2400 1928.7600 386.8400 1929.2400 ;
        RECT 385.2400 1934.2000 386.8400 1934.6800 ;
        RECT 385.2400 1923.3200 386.8400 1923.8000 ;
        RECT 340.2400 2010.3600 341.8400 2010.8400 ;
        RECT 340.2400 2015.8000 341.8400 2016.2800 ;
        RECT 340.2400 1994.0400 341.8400 1994.5200 ;
        RECT 340.2400 1999.4800 341.8400 1999.9600 ;
        RECT 340.2400 2004.9200 341.8400 2005.4000 ;
        RECT 295.2400 2010.3600 296.8400 2010.8400 ;
        RECT 295.2400 2015.8000 296.8400 2016.2800 ;
        RECT 295.2400 1994.0400 296.8400 1994.5200 ;
        RECT 295.2400 1999.4800 296.8400 1999.9600 ;
        RECT 295.2400 2004.9200 296.8400 2005.4000 ;
        RECT 340.2400 1983.1600 341.8400 1983.6400 ;
        RECT 340.2400 1988.6000 341.8400 1989.0800 ;
        RECT 340.2400 1966.8400 341.8400 1967.3200 ;
        RECT 340.2400 1972.2800 341.8400 1972.7600 ;
        RECT 340.2400 1977.7200 341.8400 1978.2000 ;
        RECT 295.2400 1983.1600 296.8400 1983.6400 ;
        RECT 295.2400 1988.6000 296.8400 1989.0800 ;
        RECT 295.2400 1966.8400 296.8400 1967.3200 ;
        RECT 295.2400 1972.2800 296.8400 1972.7600 ;
        RECT 295.2400 1977.7200 296.8400 1978.2000 ;
        RECT 245.6800 2010.3600 248.6800 2010.8400 ;
        RECT 245.6800 2015.8000 248.6800 2016.2800 ;
        RECT 245.6800 1999.4800 248.6800 1999.9600 ;
        RECT 245.6800 1994.0400 248.6800 1994.5200 ;
        RECT 245.6800 2004.9200 248.6800 2005.4000 ;
        RECT 245.6800 1983.1600 248.6800 1983.6400 ;
        RECT 245.6800 1988.6000 248.6800 1989.0800 ;
        RECT 245.6800 1972.2800 248.6800 1972.7600 ;
        RECT 245.6800 1966.8400 248.6800 1967.3200 ;
        RECT 245.6800 1977.7200 248.6800 1978.2000 ;
        RECT 340.2400 1955.9600 341.8400 1956.4400 ;
        RECT 340.2400 1961.4000 341.8400 1961.8800 ;
        RECT 340.2400 1939.6400 341.8400 1940.1200 ;
        RECT 340.2400 1945.0800 341.8400 1945.5600 ;
        RECT 340.2400 1950.5200 341.8400 1951.0000 ;
        RECT 295.2400 1955.9600 296.8400 1956.4400 ;
        RECT 295.2400 1961.4000 296.8400 1961.8800 ;
        RECT 295.2400 1939.6400 296.8400 1940.1200 ;
        RECT 295.2400 1945.0800 296.8400 1945.5600 ;
        RECT 295.2400 1950.5200 296.8400 1951.0000 ;
        RECT 340.2400 1934.2000 341.8400 1934.6800 ;
        RECT 340.2400 1928.7600 341.8400 1929.2400 ;
        RECT 340.2400 1923.3200 341.8400 1923.8000 ;
        RECT 295.2400 1934.2000 296.8400 1934.6800 ;
        RECT 295.2400 1928.7600 296.8400 1929.2400 ;
        RECT 295.2400 1923.3200 296.8400 1923.8000 ;
        RECT 245.6800 1955.9600 248.6800 1956.4400 ;
        RECT 245.6800 1961.4000 248.6800 1961.8800 ;
        RECT 245.6800 1945.0800 248.6800 1945.5600 ;
        RECT 245.6800 1939.6400 248.6800 1940.1200 ;
        RECT 245.6800 1950.5200 248.6800 1951.0000 ;
        RECT 245.6800 1928.7600 248.6800 1929.2400 ;
        RECT 245.6800 1934.2000 248.6800 1934.6800 ;
        RECT 245.6800 1923.3200 248.6800 1923.8000 ;
        RECT 245.6800 2121.5100 444.7800 2124.5100 ;
        RECT 245.6800 1916.4100 444.7800 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 1686.7700 431.8400 1894.8700 ;
        RECT 385.2400 1686.7700 386.8400 1894.8700 ;
        RECT 340.2400 1686.7700 341.8400 1894.8700 ;
        RECT 295.2400 1686.7700 296.8400 1894.8700 ;
        RECT 441.7800 1686.7700 444.7800 1894.8700 ;
        RECT 245.6800 1686.7700 248.6800 1894.8700 ;
      LAYER met3 ;
        RECT 441.7800 1889.5200 444.7800 1890.0000 ;
        RECT 430.2400 1889.5200 431.8400 1890.0000 ;
        RECT 441.7800 1878.6400 444.7800 1879.1200 ;
        RECT 441.7800 1884.0800 444.7800 1884.5600 ;
        RECT 430.2400 1878.6400 431.8400 1879.1200 ;
        RECT 430.2400 1884.0800 431.8400 1884.5600 ;
        RECT 441.7800 1862.3200 444.7800 1862.8000 ;
        RECT 441.7800 1867.7600 444.7800 1868.2400 ;
        RECT 430.2400 1862.3200 431.8400 1862.8000 ;
        RECT 430.2400 1867.7600 431.8400 1868.2400 ;
        RECT 441.7800 1851.4400 444.7800 1851.9200 ;
        RECT 441.7800 1856.8800 444.7800 1857.3600 ;
        RECT 430.2400 1851.4400 431.8400 1851.9200 ;
        RECT 430.2400 1856.8800 431.8400 1857.3600 ;
        RECT 441.7800 1873.2000 444.7800 1873.6800 ;
        RECT 430.2400 1873.2000 431.8400 1873.6800 ;
        RECT 385.2400 1878.6400 386.8400 1879.1200 ;
        RECT 385.2400 1884.0800 386.8400 1884.5600 ;
        RECT 385.2400 1889.5200 386.8400 1890.0000 ;
        RECT 385.2400 1862.3200 386.8400 1862.8000 ;
        RECT 385.2400 1867.7600 386.8400 1868.2400 ;
        RECT 385.2400 1856.8800 386.8400 1857.3600 ;
        RECT 385.2400 1851.4400 386.8400 1851.9200 ;
        RECT 385.2400 1873.2000 386.8400 1873.6800 ;
        RECT 441.7800 1835.1200 444.7800 1835.6000 ;
        RECT 441.7800 1840.5600 444.7800 1841.0400 ;
        RECT 430.2400 1835.1200 431.8400 1835.6000 ;
        RECT 430.2400 1840.5600 431.8400 1841.0400 ;
        RECT 441.7800 1818.8000 444.7800 1819.2800 ;
        RECT 441.7800 1824.2400 444.7800 1824.7200 ;
        RECT 441.7800 1829.6800 444.7800 1830.1600 ;
        RECT 430.2400 1818.8000 431.8400 1819.2800 ;
        RECT 430.2400 1824.2400 431.8400 1824.7200 ;
        RECT 430.2400 1829.6800 431.8400 1830.1600 ;
        RECT 441.7800 1807.9200 444.7800 1808.4000 ;
        RECT 441.7800 1813.3600 444.7800 1813.8400 ;
        RECT 430.2400 1807.9200 431.8400 1808.4000 ;
        RECT 430.2400 1813.3600 431.8400 1813.8400 ;
        RECT 441.7800 1791.6000 444.7800 1792.0800 ;
        RECT 441.7800 1797.0400 444.7800 1797.5200 ;
        RECT 441.7800 1802.4800 444.7800 1802.9600 ;
        RECT 430.2400 1791.6000 431.8400 1792.0800 ;
        RECT 430.2400 1797.0400 431.8400 1797.5200 ;
        RECT 430.2400 1802.4800 431.8400 1802.9600 ;
        RECT 385.2400 1835.1200 386.8400 1835.6000 ;
        RECT 385.2400 1840.5600 386.8400 1841.0400 ;
        RECT 385.2400 1818.8000 386.8400 1819.2800 ;
        RECT 385.2400 1824.2400 386.8400 1824.7200 ;
        RECT 385.2400 1829.6800 386.8400 1830.1600 ;
        RECT 385.2400 1807.9200 386.8400 1808.4000 ;
        RECT 385.2400 1813.3600 386.8400 1813.8400 ;
        RECT 385.2400 1791.6000 386.8400 1792.0800 ;
        RECT 385.2400 1797.0400 386.8400 1797.5200 ;
        RECT 385.2400 1802.4800 386.8400 1802.9600 ;
        RECT 441.7800 1846.0000 444.7800 1846.4800 ;
        RECT 385.2400 1846.0000 386.8400 1846.4800 ;
        RECT 430.2400 1846.0000 431.8400 1846.4800 ;
        RECT 340.2400 1878.6400 341.8400 1879.1200 ;
        RECT 340.2400 1884.0800 341.8400 1884.5600 ;
        RECT 340.2400 1889.5200 341.8400 1890.0000 ;
        RECT 295.2400 1878.6400 296.8400 1879.1200 ;
        RECT 295.2400 1884.0800 296.8400 1884.5600 ;
        RECT 295.2400 1889.5200 296.8400 1890.0000 ;
        RECT 340.2400 1862.3200 341.8400 1862.8000 ;
        RECT 340.2400 1867.7600 341.8400 1868.2400 ;
        RECT 340.2400 1851.4400 341.8400 1851.9200 ;
        RECT 340.2400 1856.8800 341.8400 1857.3600 ;
        RECT 295.2400 1862.3200 296.8400 1862.8000 ;
        RECT 295.2400 1867.7600 296.8400 1868.2400 ;
        RECT 295.2400 1851.4400 296.8400 1851.9200 ;
        RECT 295.2400 1856.8800 296.8400 1857.3600 ;
        RECT 295.2400 1873.2000 296.8400 1873.6800 ;
        RECT 340.2400 1873.2000 341.8400 1873.6800 ;
        RECT 245.6800 1889.5200 248.6800 1890.0000 ;
        RECT 245.6800 1884.0800 248.6800 1884.5600 ;
        RECT 245.6800 1878.6400 248.6800 1879.1200 ;
        RECT 245.6800 1867.7600 248.6800 1868.2400 ;
        RECT 245.6800 1862.3200 248.6800 1862.8000 ;
        RECT 245.6800 1856.8800 248.6800 1857.3600 ;
        RECT 245.6800 1851.4400 248.6800 1851.9200 ;
        RECT 245.6800 1873.2000 248.6800 1873.6800 ;
        RECT 340.2400 1835.1200 341.8400 1835.6000 ;
        RECT 340.2400 1840.5600 341.8400 1841.0400 ;
        RECT 340.2400 1818.8000 341.8400 1819.2800 ;
        RECT 340.2400 1824.2400 341.8400 1824.7200 ;
        RECT 340.2400 1829.6800 341.8400 1830.1600 ;
        RECT 295.2400 1835.1200 296.8400 1835.6000 ;
        RECT 295.2400 1840.5600 296.8400 1841.0400 ;
        RECT 295.2400 1818.8000 296.8400 1819.2800 ;
        RECT 295.2400 1824.2400 296.8400 1824.7200 ;
        RECT 295.2400 1829.6800 296.8400 1830.1600 ;
        RECT 340.2400 1807.9200 341.8400 1808.4000 ;
        RECT 340.2400 1813.3600 341.8400 1813.8400 ;
        RECT 340.2400 1791.6000 341.8400 1792.0800 ;
        RECT 340.2400 1797.0400 341.8400 1797.5200 ;
        RECT 340.2400 1802.4800 341.8400 1802.9600 ;
        RECT 295.2400 1807.9200 296.8400 1808.4000 ;
        RECT 295.2400 1813.3600 296.8400 1813.8400 ;
        RECT 295.2400 1791.6000 296.8400 1792.0800 ;
        RECT 295.2400 1797.0400 296.8400 1797.5200 ;
        RECT 295.2400 1802.4800 296.8400 1802.9600 ;
        RECT 245.6800 1835.1200 248.6800 1835.6000 ;
        RECT 245.6800 1840.5600 248.6800 1841.0400 ;
        RECT 245.6800 1824.2400 248.6800 1824.7200 ;
        RECT 245.6800 1818.8000 248.6800 1819.2800 ;
        RECT 245.6800 1829.6800 248.6800 1830.1600 ;
        RECT 245.6800 1807.9200 248.6800 1808.4000 ;
        RECT 245.6800 1813.3600 248.6800 1813.8400 ;
        RECT 245.6800 1797.0400 248.6800 1797.5200 ;
        RECT 245.6800 1791.6000 248.6800 1792.0800 ;
        RECT 245.6800 1802.4800 248.6800 1802.9600 ;
        RECT 245.6800 1846.0000 248.6800 1846.4800 ;
        RECT 295.2400 1846.0000 296.8400 1846.4800 ;
        RECT 340.2400 1846.0000 341.8400 1846.4800 ;
        RECT 441.7800 1780.7200 444.7800 1781.2000 ;
        RECT 441.7800 1786.1600 444.7800 1786.6400 ;
        RECT 430.2400 1780.7200 431.8400 1781.2000 ;
        RECT 430.2400 1786.1600 431.8400 1786.6400 ;
        RECT 441.7800 1764.4000 444.7800 1764.8800 ;
        RECT 441.7800 1769.8400 444.7800 1770.3200 ;
        RECT 441.7800 1775.2800 444.7800 1775.7600 ;
        RECT 430.2400 1764.4000 431.8400 1764.8800 ;
        RECT 430.2400 1769.8400 431.8400 1770.3200 ;
        RECT 430.2400 1775.2800 431.8400 1775.7600 ;
        RECT 441.7800 1753.5200 444.7800 1754.0000 ;
        RECT 441.7800 1758.9600 444.7800 1759.4400 ;
        RECT 430.2400 1753.5200 431.8400 1754.0000 ;
        RECT 430.2400 1758.9600 431.8400 1759.4400 ;
        RECT 441.7800 1737.2000 444.7800 1737.6800 ;
        RECT 441.7800 1742.6400 444.7800 1743.1200 ;
        RECT 441.7800 1748.0800 444.7800 1748.5600 ;
        RECT 430.2400 1737.2000 431.8400 1737.6800 ;
        RECT 430.2400 1742.6400 431.8400 1743.1200 ;
        RECT 430.2400 1748.0800 431.8400 1748.5600 ;
        RECT 385.2400 1780.7200 386.8400 1781.2000 ;
        RECT 385.2400 1786.1600 386.8400 1786.6400 ;
        RECT 385.2400 1764.4000 386.8400 1764.8800 ;
        RECT 385.2400 1769.8400 386.8400 1770.3200 ;
        RECT 385.2400 1775.2800 386.8400 1775.7600 ;
        RECT 385.2400 1753.5200 386.8400 1754.0000 ;
        RECT 385.2400 1758.9600 386.8400 1759.4400 ;
        RECT 385.2400 1737.2000 386.8400 1737.6800 ;
        RECT 385.2400 1742.6400 386.8400 1743.1200 ;
        RECT 385.2400 1748.0800 386.8400 1748.5600 ;
        RECT 441.7800 1726.3200 444.7800 1726.8000 ;
        RECT 441.7800 1731.7600 444.7800 1732.2400 ;
        RECT 430.2400 1726.3200 431.8400 1726.8000 ;
        RECT 430.2400 1731.7600 431.8400 1732.2400 ;
        RECT 441.7800 1710.0000 444.7800 1710.4800 ;
        RECT 441.7800 1715.4400 444.7800 1715.9200 ;
        RECT 441.7800 1720.8800 444.7800 1721.3600 ;
        RECT 430.2400 1710.0000 431.8400 1710.4800 ;
        RECT 430.2400 1715.4400 431.8400 1715.9200 ;
        RECT 430.2400 1720.8800 431.8400 1721.3600 ;
        RECT 441.7800 1699.1200 444.7800 1699.6000 ;
        RECT 441.7800 1704.5600 444.7800 1705.0400 ;
        RECT 430.2400 1699.1200 431.8400 1699.6000 ;
        RECT 430.2400 1704.5600 431.8400 1705.0400 ;
        RECT 441.7800 1693.6800 444.7800 1694.1600 ;
        RECT 430.2400 1693.6800 431.8400 1694.1600 ;
        RECT 385.2400 1726.3200 386.8400 1726.8000 ;
        RECT 385.2400 1731.7600 386.8400 1732.2400 ;
        RECT 385.2400 1710.0000 386.8400 1710.4800 ;
        RECT 385.2400 1715.4400 386.8400 1715.9200 ;
        RECT 385.2400 1720.8800 386.8400 1721.3600 ;
        RECT 385.2400 1699.1200 386.8400 1699.6000 ;
        RECT 385.2400 1704.5600 386.8400 1705.0400 ;
        RECT 385.2400 1693.6800 386.8400 1694.1600 ;
        RECT 340.2400 1780.7200 341.8400 1781.2000 ;
        RECT 340.2400 1786.1600 341.8400 1786.6400 ;
        RECT 340.2400 1764.4000 341.8400 1764.8800 ;
        RECT 340.2400 1769.8400 341.8400 1770.3200 ;
        RECT 340.2400 1775.2800 341.8400 1775.7600 ;
        RECT 295.2400 1780.7200 296.8400 1781.2000 ;
        RECT 295.2400 1786.1600 296.8400 1786.6400 ;
        RECT 295.2400 1764.4000 296.8400 1764.8800 ;
        RECT 295.2400 1769.8400 296.8400 1770.3200 ;
        RECT 295.2400 1775.2800 296.8400 1775.7600 ;
        RECT 340.2400 1753.5200 341.8400 1754.0000 ;
        RECT 340.2400 1758.9600 341.8400 1759.4400 ;
        RECT 340.2400 1737.2000 341.8400 1737.6800 ;
        RECT 340.2400 1742.6400 341.8400 1743.1200 ;
        RECT 340.2400 1748.0800 341.8400 1748.5600 ;
        RECT 295.2400 1753.5200 296.8400 1754.0000 ;
        RECT 295.2400 1758.9600 296.8400 1759.4400 ;
        RECT 295.2400 1737.2000 296.8400 1737.6800 ;
        RECT 295.2400 1742.6400 296.8400 1743.1200 ;
        RECT 295.2400 1748.0800 296.8400 1748.5600 ;
        RECT 245.6800 1780.7200 248.6800 1781.2000 ;
        RECT 245.6800 1786.1600 248.6800 1786.6400 ;
        RECT 245.6800 1769.8400 248.6800 1770.3200 ;
        RECT 245.6800 1764.4000 248.6800 1764.8800 ;
        RECT 245.6800 1775.2800 248.6800 1775.7600 ;
        RECT 245.6800 1753.5200 248.6800 1754.0000 ;
        RECT 245.6800 1758.9600 248.6800 1759.4400 ;
        RECT 245.6800 1742.6400 248.6800 1743.1200 ;
        RECT 245.6800 1737.2000 248.6800 1737.6800 ;
        RECT 245.6800 1748.0800 248.6800 1748.5600 ;
        RECT 340.2400 1726.3200 341.8400 1726.8000 ;
        RECT 340.2400 1731.7600 341.8400 1732.2400 ;
        RECT 340.2400 1710.0000 341.8400 1710.4800 ;
        RECT 340.2400 1715.4400 341.8400 1715.9200 ;
        RECT 340.2400 1720.8800 341.8400 1721.3600 ;
        RECT 295.2400 1726.3200 296.8400 1726.8000 ;
        RECT 295.2400 1731.7600 296.8400 1732.2400 ;
        RECT 295.2400 1710.0000 296.8400 1710.4800 ;
        RECT 295.2400 1715.4400 296.8400 1715.9200 ;
        RECT 295.2400 1720.8800 296.8400 1721.3600 ;
        RECT 340.2400 1704.5600 341.8400 1705.0400 ;
        RECT 340.2400 1699.1200 341.8400 1699.6000 ;
        RECT 340.2400 1693.6800 341.8400 1694.1600 ;
        RECT 295.2400 1704.5600 296.8400 1705.0400 ;
        RECT 295.2400 1699.1200 296.8400 1699.6000 ;
        RECT 295.2400 1693.6800 296.8400 1694.1600 ;
        RECT 245.6800 1726.3200 248.6800 1726.8000 ;
        RECT 245.6800 1731.7600 248.6800 1732.2400 ;
        RECT 245.6800 1715.4400 248.6800 1715.9200 ;
        RECT 245.6800 1710.0000 248.6800 1710.4800 ;
        RECT 245.6800 1720.8800 248.6800 1721.3600 ;
        RECT 245.6800 1699.1200 248.6800 1699.6000 ;
        RECT 245.6800 1704.5600 248.6800 1705.0400 ;
        RECT 245.6800 1693.6800 248.6800 1694.1600 ;
        RECT 245.6800 1891.8700 444.7800 1894.8700 ;
        RECT 245.6800 1686.7700 444.7800 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 1457.1300 431.8400 1665.2300 ;
        RECT 385.2400 1457.1300 386.8400 1665.2300 ;
        RECT 340.2400 1457.1300 341.8400 1665.2300 ;
        RECT 295.2400 1457.1300 296.8400 1665.2300 ;
        RECT 441.7800 1457.1300 444.7800 1665.2300 ;
        RECT 245.6800 1457.1300 248.6800 1665.2300 ;
      LAYER met3 ;
        RECT 441.7800 1659.8800 444.7800 1660.3600 ;
        RECT 430.2400 1659.8800 431.8400 1660.3600 ;
        RECT 441.7800 1649.0000 444.7800 1649.4800 ;
        RECT 441.7800 1654.4400 444.7800 1654.9200 ;
        RECT 430.2400 1649.0000 431.8400 1649.4800 ;
        RECT 430.2400 1654.4400 431.8400 1654.9200 ;
        RECT 441.7800 1632.6800 444.7800 1633.1600 ;
        RECT 441.7800 1638.1200 444.7800 1638.6000 ;
        RECT 430.2400 1632.6800 431.8400 1633.1600 ;
        RECT 430.2400 1638.1200 431.8400 1638.6000 ;
        RECT 441.7800 1621.8000 444.7800 1622.2800 ;
        RECT 441.7800 1627.2400 444.7800 1627.7200 ;
        RECT 430.2400 1621.8000 431.8400 1622.2800 ;
        RECT 430.2400 1627.2400 431.8400 1627.7200 ;
        RECT 441.7800 1643.5600 444.7800 1644.0400 ;
        RECT 430.2400 1643.5600 431.8400 1644.0400 ;
        RECT 385.2400 1649.0000 386.8400 1649.4800 ;
        RECT 385.2400 1654.4400 386.8400 1654.9200 ;
        RECT 385.2400 1659.8800 386.8400 1660.3600 ;
        RECT 385.2400 1632.6800 386.8400 1633.1600 ;
        RECT 385.2400 1638.1200 386.8400 1638.6000 ;
        RECT 385.2400 1627.2400 386.8400 1627.7200 ;
        RECT 385.2400 1621.8000 386.8400 1622.2800 ;
        RECT 385.2400 1643.5600 386.8400 1644.0400 ;
        RECT 441.7800 1605.4800 444.7800 1605.9600 ;
        RECT 441.7800 1610.9200 444.7800 1611.4000 ;
        RECT 430.2400 1605.4800 431.8400 1605.9600 ;
        RECT 430.2400 1610.9200 431.8400 1611.4000 ;
        RECT 441.7800 1589.1600 444.7800 1589.6400 ;
        RECT 441.7800 1594.6000 444.7800 1595.0800 ;
        RECT 441.7800 1600.0400 444.7800 1600.5200 ;
        RECT 430.2400 1589.1600 431.8400 1589.6400 ;
        RECT 430.2400 1594.6000 431.8400 1595.0800 ;
        RECT 430.2400 1600.0400 431.8400 1600.5200 ;
        RECT 441.7800 1578.2800 444.7800 1578.7600 ;
        RECT 441.7800 1583.7200 444.7800 1584.2000 ;
        RECT 430.2400 1578.2800 431.8400 1578.7600 ;
        RECT 430.2400 1583.7200 431.8400 1584.2000 ;
        RECT 441.7800 1561.9600 444.7800 1562.4400 ;
        RECT 441.7800 1567.4000 444.7800 1567.8800 ;
        RECT 441.7800 1572.8400 444.7800 1573.3200 ;
        RECT 430.2400 1561.9600 431.8400 1562.4400 ;
        RECT 430.2400 1567.4000 431.8400 1567.8800 ;
        RECT 430.2400 1572.8400 431.8400 1573.3200 ;
        RECT 385.2400 1605.4800 386.8400 1605.9600 ;
        RECT 385.2400 1610.9200 386.8400 1611.4000 ;
        RECT 385.2400 1589.1600 386.8400 1589.6400 ;
        RECT 385.2400 1594.6000 386.8400 1595.0800 ;
        RECT 385.2400 1600.0400 386.8400 1600.5200 ;
        RECT 385.2400 1578.2800 386.8400 1578.7600 ;
        RECT 385.2400 1583.7200 386.8400 1584.2000 ;
        RECT 385.2400 1561.9600 386.8400 1562.4400 ;
        RECT 385.2400 1567.4000 386.8400 1567.8800 ;
        RECT 385.2400 1572.8400 386.8400 1573.3200 ;
        RECT 441.7800 1616.3600 444.7800 1616.8400 ;
        RECT 385.2400 1616.3600 386.8400 1616.8400 ;
        RECT 430.2400 1616.3600 431.8400 1616.8400 ;
        RECT 340.2400 1649.0000 341.8400 1649.4800 ;
        RECT 340.2400 1654.4400 341.8400 1654.9200 ;
        RECT 340.2400 1659.8800 341.8400 1660.3600 ;
        RECT 295.2400 1649.0000 296.8400 1649.4800 ;
        RECT 295.2400 1654.4400 296.8400 1654.9200 ;
        RECT 295.2400 1659.8800 296.8400 1660.3600 ;
        RECT 340.2400 1632.6800 341.8400 1633.1600 ;
        RECT 340.2400 1638.1200 341.8400 1638.6000 ;
        RECT 340.2400 1621.8000 341.8400 1622.2800 ;
        RECT 340.2400 1627.2400 341.8400 1627.7200 ;
        RECT 295.2400 1632.6800 296.8400 1633.1600 ;
        RECT 295.2400 1638.1200 296.8400 1638.6000 ;
        RECT 295.2400 1621.8000 296.8400 1622.2800 ;
        RECT 295.2400 1627.2400 296.8400 1627.7200 ;
        RECT 295.2400 1643.5600 296.8400 1644.0400 ;
        RECT 340.2400 1643.5600 341.8400 1644.0400 ;
        RECT 245.6800 1659.8800 248.6800 1660.3600 ;
        RECT 245.6800 1654.4400 248.6800 1654.9200 ;
        RECT 245.6800 1649.0000 248.6800 1649.4800 ;
        RECT 245.6800 1638.1200 248.6800 1638.6000 ;
        RECT 245.6800 1632.6800 248.6800 1633.1600 ;
        RECT 245.6800 1627.2400 248.6800 1627.7200 ;
        RECT 245.6800 1621.8000 248.6800 1622.2800 ;
        RECT 245.6800 1643.5600 248.6800 1644.0400 ;
        RECT 340.2400 1605.4800 341.8400 1605.9600 ;
        RECT 340.2400 1610.9200 341.8400 1611.4000 ;
        RECT 340.2400 1589.1600 341.8400 1589.6400 ;
        RECT 340.2400 1594.6000 341.8400 1595.0800 ;
        RECT 340.2400 1600.0400 341.8400 1600.5200 ;
        RECT 295.2400 1605.4800 296.8400 1605.9600 ;
        RECT 295.2400 1610.9200 296.8400 1611.4000 ;
        RECT 295.2400 1589.1600 296.8400 1589.6400 ;
        RECT 295.2400 1594.6000 296.8400 1595.0800 ;
        RECT 295.2400 1600.0400 296.8400 1600.5200 ;
        RECT 340.2400 1578.2800 341.8400 1578.7600 ;
        RECT 340.2400 1583.7200 341.8400 1584.2000 ;
        RECT 340.2400 1561.9600 341.8400 1562.4400 ;
        RECT 340.2400 1567.4000 341.8400 1567.8800 ;
        RECT 340.2400 1572.8400 341.8400 1573.3200 ;
        RECT 295.2400 1578.2800 296.8400 1578.7600 ;
        RECT 295.2400 1583.7200 296.8400 1584.2000 ;
        RECT 295.2400 1561.9600 296.8400 1562.4400 ;
        RECT 295.2400 1567.4000 296.8400 1567.8800 ;
        RECT 295.2400 1572.8400 296.8400 1573.3200 ;
        RECT 245.6800 1605.4800 248.6800 1605.9600 ;
        RECT 245.6800 1610.9200 248.6800 1611.4000 ;
        RECT 245.6800 1594.6000 248.6800 1595.0800 ;
        RECT 245.6800 1589.1600 248.6800 1589.6400 ;
        RECT 245.6800 1600.0400 248.6800 1600.5200 ;
        RECT 245.6800 1578.2800 248.6800 1578.7600 ;
        RECT 245.6800 1583.7200 248.6800 1584.2000 ;
        RECT 245.6800 1567.4000 248.6800 1567.8800 ;
        RECT 245.6800 1561.9600 248.6800 1562.4400 ;
        RECT 245.6800 1572.8400 248.6800 1573.3200 ;
        RECT 245.6800 1616.3600 248.6800 1616.8400 ;
        RECT 295.2400 1616.3600 296.8400 1616.8400 ;
        RECT 340.2400 1616.3600 341.8400 1616.8400 ;
        RECT 441.7800 1551.0800 444.7800 1551.5600 ;
        RECT 441.7800 1556.5200 444.7800 1557.0000 ;
        RECT 430.2400 1551.0800 431.8400 1551.5600 ;
        RECT 430.2400 1556.5200 431.8400 1557.0000 ;
        RECT 441.7800 1534.7600 444.7800 1535.2400 ;
        RECT 441.7800 1540.2000 444.7800 1540.6800 ;
        RECT 441.7800 1545.6400 444.7800 1546.1200 ;
        RECT 430.2400 1534.7600 431.8400 1535.2400 ;
        RECT 430.2400 1540.2000 431.8400 1540.6800 ;
        RECT 430.2400 1545.6400 431.8400 1546.1200 ;
        RECT 441.7800 1523.8800 444.7800 1524.3600 ;
        RECT 441.7800 1529.3200 444.7800 1529.8000 ;
        RECT 430.2400 1523.8800 431.8400 1524.3600 ;
        RECT 430.2400 1529.3200 431.8400 1529.8000 ;
        RECT 441.7800 1507.5600 444.7800 1508.0400 ;
        RECT 441.7800 1513.0000 444.7800 1513.4800 ;
        RECT 441.7800 1518.4400 444.7800 1518.9200 ;
        RECT 430.2400 1507.5600 431.8400 1508.0400 ;
        RECT 430.2400 1513.0000 431.8400 1513.4800 ;
        RECT 430.2400 1518.4400 431.8400 1518.9200 ;
        RECT 385.2400 1551.0800 386.8400 1551.5600 ;
        RECT 385.2400 1556.5200 386.8400 1557.0000 ;
        RECT 385.2400 1534.7600 386.8400 1535.2400 ;
        RECT 385.2400 1540.2000 386.8400 1540.6800 ;
        RECT 385.2400 1545.6400 386.8400 1546.1200 ;
        RECT 385.2400 1523.8800 386.8400 1524.3600 ;
        RECT 385.2400 1529.3200 386.8400 1529.8000 ;
        RECT 385.2400 1507.5600 386.8400 1508.0400 ;
        RECT 385.2400 1513.0000 386.8400 1513.4800 ;
        RECT 385.2400 1518.4400 386.8400 1518.9200 ;
        RECT 441.7800 1496.6800 444.7800 1497.1600 ;
        RECT 441.7800 1502.1200 444.7800 1502.6000 ;
        RECT 430.2400 1496.6800 431.8400 1497.1600 ;
        RECT 430.2400 1502.1200 431.8400 1502.6000 ;
        RECT 441.7800 1480.3600 444.7800 1480.8400 ;
        RECT 441.7800 1485.8000 444.7800 1486.2800 ;
        RECT 441.7800 1491.2400 444.7800 1491.7200 ;
        RECT 430.2400 1480.3600 431.8400 1480.8400 ;
        RECT 430.2400 1485.8000 431.8400 1486.2800 ;
        RECT 430.2400 1491.2400 431.8400 1491.7200 ;
        RECT 441.7800 1469.4800 444.7800 1469.9600 ;
        RECT 441.7800 1474.9200 444.7800 1475.4000 ;
        RECT 430.2400 1469.4800 431.8400 1469.9600 ;
        RECT 430.2400 1474.9200 431.8400 1475.4000 ;
        RECT 441.7800 1464.0400 444.7800 1464.5200 ;
        RECT 430.2400 1464.0400 431.8400 1464.5200 ;
        RECT 385.2400 1496.6800 386.8400 1497.1600 ;
        RECT 385.2400 1502.1200 386.8400 1502.6000 ;
        RECT 385.2400 1480.3600 386.8400 1480.8400 ;
        RECT 385.2400 1485.8000 386.8400 1486.2800 ;
        RECT 385.2400 1491.2400 386.8400 1491.7200 ;
        RECT 385.2400 1469.4800 386.8400 1469.9600 ;
        RECT 385.2400 1474.9200 386.8400 1475.4000 ;
        RECT 385.2400 1464.0400 386.8400 1464.5200 ;
        RECT 340.2400 1551.0800 341.8400 1551.5600 ;
        RECT 340.2400 1556.5200 341.8400 1557.0000 ;
        RECT 340.2400 1534.7600 341.8400 1535.2400 ;
        RECT 340.2400 1540.2000 341.8400 1540.6800 ;
        RECT 340.2400 1545.6400 341.8400 1546.1200 ;
        RECT 295.2400 1551.0800 296.8400 1551.5600 ;
        RECT 295.2400 1556.5200 296.8400 1557.0000 ;
        RECT 295.2400 1534.7600 296.8400 1535.2400 ;
        RECT 295.2400 1540.2000 296.8400 1540.6800 ;
        RECT 295.2400 1545.6400 296.8400 1546.1200 ;
        RECT 340.2400 1523.8800 341.8400 1524.3600 ;
        RECT 340.2400 1529.3200 341.8400 1529.8000 ;
        RECT 340.2400 1507.5600 341.8400 1508.0400 ;
        RECT 340.2400 1513.0000 341.8400 1513.4800 ;
        RECT 340.2400 1518.4400 341.8400 1518.9200 ;
        RECT 295.2400 1523.8800 296.8400 1524.3600 ;
        RECT 295.2400 1529.3200 296.8400 1529.8000 ;
        RECT 295.2400 1507.5600 296.8400 1508.0400 ;
        RECT 295.2400 1513.0000 296.8400 1513.4800 ;
        RECT 295.2400 1518.4400 296.8400 1518.9200 ;
        RECT 245.6800 1551.0800 248.6800 1551.5600 ;
        RECT 245.6800 1556.5200 248.6800 1557.0000 ;
        RECT 245.6800 1540.2000 248.6800 1540.6800 ;
        RECT 245.6800 1534.7600 248.6800 1535.2400 ;
        RECT 245.6800 1545.6400 248.6800 1546.1200 ;
        RECT 245.6800 1523.8800 248.6800 1524.3600 ;
        RECT 245.6800 1529.3200 248.6800 1529.8000 ;
        RECT 245.6800 1513.0000 248.6800 1513.4800 ;
        RECT 245.6800 1507.5600 248.6800 1508.0400 ;
        RECT 245.6800 1518.4400 248.6800 1518.9200 ;
        RECT 340.2400 1496.6800 341.8400 1497.1600 ;
        RECT 340.2400 1502.1200 341.8400 1502.6000 ;
        RECT 340.2400 1480.3600 341.8400 1480.8400 ;
        RECT 340.2400 1485.8000 341.8400 1486.2800 ;
        RECT 340.2400 1491.2400 341.8400 1491.7200 ;
        RECT 295.2400 1496.6800 296.8400 1497.1600 ;
        RECT 295.2400 1502.1200 296.8400 1502.6000 ;
        RECT 295.2400 1480.3600 296.8400 1480.8400 ;
        RECT 295.2400 1485.8000 296.8400 1486.2800 ;
        RECT 295.2400 1491.2400 296.8400 1491.7200 ;
        RECT 340.2400 1474.9200 341.8400 1475.4000 ;
        RECT 340.2400 1469.4800 341.8400 1469.9600 ;
        RECT 340.2400 1464.0400 341.8400 1464.5200 ;
        RECT 295.2400 1474.9200 296.8400 1475.4000 ;
        RECT 295.2400 1469.4800 296.8400 1469.9600 ;
        RECT 295.2400 1464.0400 296.8400 1464.5200 ;
        RECT 245.6800 1496.6800 248.6800 1497.1600 ;
        RECT 245.6800 1502.1200 248.6800 1502.6000 ;
        RECT 245.6800 1485.8000 248.6800 1486.2800 ;
        RECT 245.6800 1480.3600 248.6800 1480.8400 ;
        RECT 245.6800 1491.2400 248.6800 1491.7200 ;
        RECT 245.6800 1469.4800 248.6800 1469.9600 ;
        RECT 245.6800 1474.9200 248.6800 1475.4000 ;
        RECT 245.6800 1464.0400 248.6800 1464.5200 ;
        RECT 245.6800 1662.2300 444.7800 1665.2300 ;
        RECT 245.6800 1457.1300 444.7800 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 1227.4900 431.8400 1435.5900 ;
        RECT 385.2400 1227.4900 386.8400 1435.5900 ;
        RECT 340.2400 1227.4900 341.8400 1435.5900 ;
        RECT 295.2400 1227.4900 296.8400 1435.5900 ;
        RECT 441.7800 1227.4900 444.7800 1435.5900 ;
        RECT 245.6800 1227.4900 248.6800 1435.5900 ;
      LAYER met3 ;
        RECT 441.7800 1430.2400 444.7800 1430.7200 ;
        RECT 430.2400 1430.2400 431.8400 1430.7200 ;
        RECT 441.7800 1419.3600 444.7800 1419.8400 ;
        RECT 441.7800 1424.8000 444.7800 1425.2800 ;
        RECT 430.2400 1419.3600 431.8400 1419.8400 ;
        RECT 430.2400 1424.8000 431.8400 1425.2800 ;
        RECT 441.7800 1403.0400 444.7800 1403.5200 ;
        RECT 441.7800 1408.4800 444.7800 1408.9600 ;
        RECT 430.2400 1403.0400 431.8400 1403.5200 ;
        RECT 430.2400 1408.4800 431.8400 1408.9600 ;
        RECT 441.7800 1392.1600 444.7800 1392.6400 ;
        RECT 441.7800 1397.6000 444.7800 1398.0800 ;
        RECT 430.2400 1392.1600 431.8400 1392.6400 ;
        RECT 430.2400 1397.6000 431.8400 1398.0800 ;
        RECT 441.7800 1413.9200 444.7800 1414.4000 ;
        RECT 430.2400 1413.9200 431.8400 1414.4000 ;
        RECT 385.2400 1419.3600 386.8400 1419.8400 ;
        RECT 385.2400 1424.8000 386.8400 1425.2800 ;
        RECT 385.2400 1430.2400 386.8400 1430.7200 ;
        RECT 385.2400 1403.0400 386.8400 1403.5200 ;
        RECT 385.2400 1408.4800 386.8400 1408.9600 ;
        RECT 385.2400 1397.6000 386.8400 1398.0800 ;
        RECT 385.2400 1392.1600 386.8400 1392.6400 ;
        RECT 385.2400 1413.9200 386.8400 1414.4000 ;
        RECT 441.7800 1375.8400 444.7800 1376.3200 ;
        RECT 441.7800 1381.2800 444.7800 1381.7600 ;
        RECT 430.2400 1375.8400 431.8400 1376.3200 ;
        RECT 430.2400 1381.2800 431.8400 1381.7600 ;
        RECT 441.7800 1359.5200 444.7800 1360.0000 ;
        RECT 441.7800 1364.9600 444.7800 1365.4400 ;
        RECT 441.7800 1370.4000 444.7800 1370.8800 ;
        RECT 430.2400 1359.5200 431.8400 1360.0000 ;
        RECT 430.2400 1364.9600 431.8400 1365.4400 ;
        RECT 430.2400 1370.4000 431.8400 1370.8800 ;
        RECT 441.7800 1348.6400 444.7800 1349.1200 ;
        RECT 441.7800 1354.0800 444.7800 1354.5600 ;
        RECT 430.2400 1348.6400 431.8400 1349.1200 ;
        RECT 430.2400 1354.0800 431.8400 1354.5600 ;
        RECT 441.7800 1332.3200 444.7800 1332.8000 ;
        RECT 441.7800 1337.7600 444.7800 1338.2400 ;
        RECT 441.7800 1343.2000 444.7800 1343.6800 ;
        RECT 430.2400 1332.3200 431.8400 1332.8000 ;
        RECT 430.2400 1337.7600 431.8400 1338.2400 ;
        RECT 430.2400 1343.2000 431.8400 1343.6800 ;
        RECT 385.2400 1375.8400 386.8400 1376.3200 ;
        RECT 385.2400 1381.2800 386.8400 1381.7600 ;
        RECT 385.2400 1359.5200 386.8400 1360.0000 ;
        RECT 385.2400 1364.9600 386.8400 1365.4400 ;
        RECT 385.2400 1370.4000 386.8400 1370.8800 ;
        RECT 385.2400 1348.6400 386.8400 1349.1200 ;
        RECT 385.2400 1354.0800 386.8400 1354.5600 ;
        RECT 385.2400 1332.3200 386.8400 1332.8000 ;
        RECT 385.2400 1337.7600 386.8400 1338.2400 ;
        RECT 385.2400 1343.2000 386.8400 1343.6800 ;
        RECT 441.7800 1386.7200 444.7800 1387.2000 ;
        RECT 385.2400 1386.7200 386.8400 1387.2000 ;
        RECT 430.2400 1386.7200 431.8400 1387.2000 ;
        RECT 340.2400 1419.3600 341.8400 1419.8400 ;
        RECT 340.2400 1424.8000 341.8400 1425.2800 ;
        RECT 340.2400 1430.2400 341.8400 1430.7200 ;
        RECT 295.2400 1419.3600 296.8400 1419.8400 ;
        RECT 295.2400 1424.8000 296.8400 1425.2800 ;
        RECT 295.2400 1430.2400 296.8400 1430.7200 ;
        RECT 340.2400 1403.0400 341.8400 1403.5200 ;
        RECT 340.2400 1408.4800 341.8400 1408.9600 ;
        RECT 340.2400 1392.1600 341.8400 1392.6400 ;
        RECT 340.2400 1397.6000 341.8400 1398.0800 ;
        RECT 295.2400 1403.0400 296.8400 1403.5200 ;
        RECT 295.2400 1408.4800 296.8400 1408.9600 ;
        RECT 295.2400 1392.1600 296.8400 1392.6400 ;
        RECT 295.2400 1397.6000 296.8400 1398.0800 ;
        RECT 295.2400 1413.9200 296.8400 1414.4000 ;
        RECT 340.2400 1413.9200 341.8400 1414.4000 ;
        RECT 245.6800 1430.2400 248.6800 1430.7200 ;
        RECT 245.6800 1424.8000 248.6800 1425.2800 ;
        RECT 245.6800 1419.3600 248.6800 1419.8400 ;
        RECT 245.6800 1408.4800 248.6800 1408.9600 ;
        RECT 245.6800 1403.0400 248.6800 1403.5200 ;
        RECT 245.6800 1397.6000 248.6800 1398.0800 ;
        RECT 245.6800 1392.1600 248.6800 1392.6400 ;
        RECT 245.6800 1413.9200 248.6800 1414.4000 ;
        RECT 340.2400 1375.8400 341.8400 1376.3200 ;
        RECT 340.2400 1381.2800 341.8400 1381.7600 ;
        RECT 340.2400 1359.5200 341.8400 1360.0000 ;
        RECT 340.2400 1364.9600 341.8400 1365.4400 ;
        RECT 340.2400 1370.4000 341.8400 1370.8800 ;
        RECT 295.2400 1375.8400 296.8400 1376.3200 ;
        RECT 295.2400 1381.2800 296.8400 1381.7600 ;
        RECT 295.2400 1359.5200 296.8400 1360.0000 ;
        RECT 295.2400 1364.9600 296.8400 1365.4400 ;
        RECT 295.2400 1370.4000 296.8400 1370.8800 ;
        RECT 340.2400 1348.6400 341.8400 1349.1200 ;
        RECT 340.2400 1354.0800 341.8400 1354.5600 ;
        RECT 340.2400 1332.3200 341.8400 1332.8000 ;
        RECT 340.2400 1337.7600 341.8400 1338.2400 ;
        RECT 340.2400 1343.2000 341.8400 1343.6800 ;
        RECT 295.2400 1348.6400 296.8400 1349.1200 ;
        RECT 295.2400 1354.0800 296.8400 1354.5600 ;
        RECT 295.2400 1332.3200 296.8400 1332.8000 ;
        RECT 295.2400 1337.7600 296.8400 1338.2400 ;
        RECT 295.2400 1343.2000 296.8400 1343.6800 ;
        RECT 245.6800 1375.8400 248.6800 1376.3200 ;
        RECT 245.6800 1381.2800 248.6800 1381.7600 ;
        RECT 245.6800 1364.9600 248.6800 1365.4400 ;
        RECT 245.6800 1359.5200 248.6800 1360.0000 ;
        RECT 245.6800 1370.4000 248.6800 1370.8800 ;
        RECT 245.6800 1348.6400 248.6800 1349.1200 ;
        RECT 245.6800 1354.0800 248.6800 1354.5600 ;
        RECT 245.6800 1337.7600 248.6800 1338.2400 ;
        RECT 245.6800 1332.3200 248.6800 1332.8000 ;
        RECT 245.6800 1343.2000 248.6800 1343.6800 ;
        RECT 245.6800 1386.7200 248.6800 1387.2000 ;
        RECT 295.2400 1386.7200 296.8400 1387.2000 ;
        RECT 340.2400 1386.7200 341.8400 1387.2000 ;
        RECT 441.7800 1321.4400 444.7800 1321.9200 ;
        RECT 441.7800 1326.8800 444.7800 1327.3600 ;
        RECT 430.2400 1321.4400 431.8400 1321.9200 ;
        RECT 430.2400 1326.8800 431.8400 1327.3600 ;
        RECT 441.7800 1305.1200 444.7800 1305.6000 ;
        RECT 441.7800 1310.5600 444.7800 1311.0400 ;
        RECT 441.7800 1316.0000 444.7800 1316.4800 ;
        RECT 430.2400 1305.1200 431.8400 1305.6000 ;
        RECT 430.2400 1310.5600 431.8400 1311.0400 ;
        RECT 430.2400 1316.0000 431.8400 1316.4800 ;
        RECT 441.7800 1294.2400 444.7800 1294.7200 ;
        RECT 441.7800 1299.6800 444.7800 1300.1600 ;
        RECT 430.2400 1294.2400 431.8400 1294.7200 ;
        RECT 430.2400 1299.6800 431.8400 1300.1600 ;
        RECT 441.7800 1277.9200 444.7800 1278.4000 ;
        RECT 441.7800 1283.3600 444.7800 1283.8400 ;
        RECT 441.7800 1288.8000 444.7800 1289.2800 ;
        RECT 430.2400 1277.9200 431.8400 1278.4000 ;
        RECT 430.2400 1283.3600 431.8400 1283.8400 ;
        RECT 430.2400 1288.8000 431.8400 1289.2800 ;
        RECT 385.2400 1321.4400 386.8400 1321.9200 ;
        RECT 385.2400 1326.8800 386.8400 1327.3600 ;
        RECT 385.2400 1305.1200 386.8400 1305.6000 ;
        RECT 385.2400 1310.5600 386.8400 1311.0400 ;
        RECT 385.2400 1316.0000 386.8400 1316.4800 ;
        RECT 385.2400 1294.2400 386.8400 1294.7200 ;
        RECT 385.2400 1299.6800 386.8400 1300.1600 ;
        RECT 385.2400 1277.9200 386.8400 1278.4000 ;
        RECT 385.2400 1283.3600 386.8400 1283.8400 ;
        RECT 385.2400 1288.8000 386.8400 1289.2800 ;
        RECT 441.7800 1267.0400 444.7800 1267.5200 ;
        RECT 441.7800 1272.4800 444.7800 1272.9600 ;
        RECT 430.2400 1267.0400 431.8400 1267.5200 ;
        RECT 430.2400 1272.4800 431.8400 1272.9600 ;
        RECT 441.7800 1250.7200 444.7800 1251.2000 ;
        RECT 441.7800 1256.1600 444.7800 1256.6400 ;
        RECT 441.7800 1261.6000 444.7800 1262.0800 ;
        RECT 430.2400 1250.7200 431.8400 1251.2000 ;
        RECT 430.2400 1256.1600 431.8400 1256.6400 ;
        RECT 430.2400 1261.6000 431.8400 1262.0800 ;
        RECT 441.7800 1239.8400 444.7800 1240.3200 ;
        RECT 441.7800 1245.2800 444.7800 1245.7600 ;
        RECT 430.2400 1239.8400 431.8400 1240.3200 ;
        RECT 430.2400 1245.2800 431.8400 1245.7600 ;
        RECT 441.7800 1234.4000 444.7800 1234.8800 ;
        RECT 430.2400 1234.4000 431.8400 1234.8800 ;
        RECT 385.2400 1267.0400 386.8400 1267.5200 ;
        RECT 385.2400 1272.4800 386.8400 1272.9600 ;
        RECT 385.2400 1250.7200 386.8400 1251.2000 ;
        RECT 385.2400 1256.1600 386.8400 1256.6400 ;
        RECT 385.2400 1261.6000 386.8400 1262.0800 ;
        RECT 385.2400 1239.8400 386.8400 1240.3200 ;
        RECT 385.2400 1245.2800 386.8400 1245.7600 ;
        RECT 385.2400 1234.4000 386.8400 1234.8800 ;
        RECT 340.2400 1321.4400 341.8400 1321.9200 ;
        RECT 340.2400 1326.8800 341.8400 1327.3600 ;
        RECT 340.2400 1305.1200 341.8400 1305.6000 ;
        RECT 340.2400 1310.5600 341.8400 1311.0400 ;
        RECT 340.2400 1316.0000 341.8400 1316.4800 ;
        RECT 295.2400 1321.4400 296.8400 1321.9200 ;
        RECT 295.2400 1326.8800 296.8400 1327.3600 ;
        RECT 295.2400 1305.1200 296.8400 1305.6000 ;
        RECT 295.2400 1310.5600 296.8400 1311.0400 ;
        RECT 295.2400 1316.0000 296.8400 1316.4800 ;
        RECT 340.2400 1294.2400 341.8400 1294.7200 ;
        RECT 340.2400 1299.6800 341.8400 1300.1600 ;
        RECT 340.2400 1277.9200 341.8400 1278.4000 ;
        RECT 340.2400 1283.3600 341.8400 1283.8400 ;
        RECT 340.2400 1288.8000 341.8400 1289.2800 ;
        RECT 295.2400 1294.2400 296.8400 1294.7200 ;
        RECT 295.2400 1299.6800 296.8400 1300.1600 ;
        RECT 295.2400 1277.9200 296.8400 1278.4000 ;
        RECT 295.2400 1283.3600 296.8400 1283.8400 ;
        RECT 295.2400 1288.8000 296.8400 1289.2800 ;
        RECT 245.6800 1321.4400 248.6800 1321.9200 ;
        RECT 245.6800 1326.8800 248.6800 1327.3600 ;
        RECT 245.6800 1310.5600 248.6800 1311.0400 ;
        RECT 245.6800 1305.1200 248.6800 1305.6000 ;
        RECT 245.6800 1316.0000 248.6800 1316.4800 ;
        RECT 245.6800 1294.2400 248.6800 1294.7200 ;
        RECT 245.6800 1299.6800 248.6800 1300.1600 ;
        RECT 245.6800 1283.3600 248.6800 1283.8400 ;
        RECT 245.6800 1277.9200 248.6800 1278.4000 ;
        RECT 245.6800 1288.8000 248.6800 1289.2800 ;
        RECT 340.2400 1267.0400 341.8400 1267.5200 ;
        RECT 340.2400 1272.4800 341.8400 1272.9600 ;
        RECT 340.2400 1250.7200 341.8400 1251.2000 ;
        RECT 340.2400 1256.1600 341.8400 1256.6400 ;
        RECT 340.2400 1261.6000 341.8400 1262.0800 ;
        RECT 295.2400 1267.0400 296.8400 1267.5200 ;
        RECT 295.2400 1272.4800 296.8400 1272.9600 ;
        RECT 295.2400 1250.7200 296.8400 1251.2000 ;
        RECT 295.2400 1256.1600 296.8400 1256.6400 ;
        RECT 295.2400 1261.6000 296.8400 1262.0800 ;
        RECT 340.2400 1245.2800 341.8400 1245.7600 ;
        RECT 340.2400 1239.8400 341.8400 1240.3200 ;
        RECT 340.2400 1234.4000 341.8400 1234.8800 ;
        RECT 295.2400 1245.2800 296.8400 1245.7600 ;
        RECT 295.2400 1239.8400 296.8400 1240.3200 ;
        RECT 295.2400 1234.4000 296.8400 1234.8800 ;
        RECT 245.6800 1267.0400 248.6800 1267.5200 ;
        RECT 245.6800 1272.4800 248.6800 1272.9600 ;
        RECT 245.6800 1256.1600 248.6800 1256.6400 ;
        RECT 245.6800 1250.7200 248.6800 1251.2000 ;
        RECT 245.6800 1261.6000 248.6800 1262.0800 ;
        RECT 245.6800 1239.8400 248.6800 1240.3200 ;
        RECT 245.6800 1245.2800 248.6800 1245.7600 ;
        RECT 245.6800 1234.4000 248.6800 1234.8800 ;
        RECT 245.6800 1432.5900 444.7800 1435.5900 ;
        RECT 245.6800 1227.4900 444.7800 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 997.8500 431.8400 1205.9500 ;
        RECT 385.2400 997.8500 386.8400 1205.9500 ;
        RECT 340.2400 997.8500 341.8400 1205.9500 ;
        RECT 295.2400 997.8500 296.8400 1205.9500 ;
        RECT 441.7800 997.8500 444.7800 1205.9500 ;
        RECT 245.6800 997.8500 248.6800 1205.9500 ;
      LAYER met3 ;
        RECT 441.7800 1200.6000 444.7800 1201.0800 ;
        RECT 430.2400 1200.6000 431.8400 1201.0800 ;
        RECT 441.7800 1189.7200 444.7800 1190.2000 ;
        RECT 441.7800 1195.1600 444.7800 1195.6400 ;
        RECT 430.2400 1189.7200 431.8400 1190.2000 ;
        RECT 430.2400 1195.1600 431.8400 1195.6400 ;
        RECT 441.7800 1173.4000 444.7800 1173.8800 ;
        RECT 441.7800 1178.8400 444.7800 1179.3200 ;
        RECT 430.2400 1173.4000 431.8400 1173.8800 ;
        RECT 430.2400 1178.8400 431.8400 1179.3200 ;
        RECT 441.7800 1162.5200 444.7800 1163.0000 ;
        RECT 441.7800 1167.9600 444.7800 1168.4400 ;
        RECT 430.2400 1162.5200 431.8400 1163.0000 ;
        RECT 430.2400 1167.9600 431.8400 1168.4400 ;
        RECT 441.7800 1184.2800 444.7800 1184.7600 ;
        RECT 430.2400 1184.2800 431.8400 1184.7600 ;
        RECT 385.2400 1189.7200 386.8400 1190.2000 ;
        RECT 385.2400 1195.1600 386.8400 1195.6400 ;
        RECT 385.2400 1200.6000 386.8400 1201.0800 ;
        RECT 385.2400 1173.4000 386.8400 1173.8800 ;
        RECT 385.2400 1178.8400 386.8400 1179.3200 ;
        RECT 385.2400 1167.9600 386.8400 1168.4400 ;
        RECT 385.2400 1162.5200 386.8400 1163.0000 ;
        RECT 385.2400 1184.2800 386.8400 1184.7600 ;
        RECT 441.7800 1146.2000 444.7800 1146.6800 ;
        RECT 441.7800 1151.6400 444.7800 1152.1200 ;
        RECT 430.2400 1146.2000 431.8400 1146.6800 ;
        RECT 430.2400 1151.6400 431.8400 1152.1200 ;
        RECT 441.7800 1129.8800 444.7800 1130.3600 ;
        RECT 441.7800 1135.3200 444.7800 1135.8000 ;
        RECT 441.7800 1140.7600 444.7800 1141.2400 ;
        RECT 430.2400 1129.8800 431.8400 1130.3600 ;
        RECT 430.2400 1135.3200 431.8400 1135.8000 ;
        RECT 430.2400 1140.7600 431.8400 1141.2400 ;
        RECT 441.7800 1119.0000 444.7800 1119.4800 ;
        RECT 441.7800 1124.4400 444.7800 1124.9200 ;
        RECT 430.2400 1119.0000 431.8400 1119.4800 ;
        RECT 430.2400 1124.4400 431.8400 1124.9200 ;
        RECT 441.7800 1102.6800 444.7800 1103.1600 ;
        RECT 441.7800 1108.1200 444.7800 1108.6000 ;
        RECT 441.7800 1113.5600 444.7800 1114.0400 ;
        RECT 430.2400 1102.6800 431.8400 1103.1600 ;
        RECT 430.2400 1108.1200 431.8400 1108.6000 ;
        RECT 430.2400 1113.5600 431.8400 1114.0400 ;
        RECT 385.2400 1146.2000 386.8400 1146.6800 ;
        RECT 385.2400 1151.6400 386.8400 1152.1200 ;
        RECT 385.2400 1129.8800 386.8400 1130.3600 ;
        RECT 385.2400 1135.3200 386.8400 1135.8000 ;
        RECT 385.2400 1140.7600 386.8400 1141.2400 ;
        RECT 385.2400 1119.0000 386.8400 1119.4800 ;
        RECT 385.2400 1124.4400 386.8400 1124.9200 ;
        RECT 385.2400 1102.6800 386.8400 1103.1600 ;
        RECT 385.2400 1108.1200 386.8400 1108.6000 ;
        RECT 385.2400 1113.5600 386.8400 1114.0400 ;
        RECT 441.7800 1157.0800 444.7800 1157.5600 ;
        RECT 385.2400 1157.0800 386.8400 1157.5600 ;
        RECT 430.2400 1157.0800 431.8400 1157.5600 ;
        RECT 340.2400 1189.7200 341.8400 1190.2000 ;
        RECT 340.2400 1195.1600 341.8400 1195.6400 ;
        RECT 340.2400 1200.6000 341.8400 1201.0800 ;
        RECT 295.2400 1189.7200 296.8400 1190.2000 ;
        RECT 295.2400 1195.1600 296.8400 1195.6400 ;
        RECT 295.2400 1200.6000 296.8400 1201.0800 ;
        RECT 340.2400 1173.4000 341.8400 1173.8800 ;
        RECT 340.2400 1178.8400 341.8400 1179.3200 ;
        RECT 340.2400 1162.5200 341.8400 1163.0000 ;
        RECT 340.2400 1167.9600 341.8400 1168.4400 ;
        RECT 295.2400 1173.4000 296.8400 1173.8800 ;
        RECT 295.2400 1178.8400 296.8400 1179.3200 ;
        RECT 295.2400 1162.5200 296.8400 1163.0000 ;
        RECT 295.2400 1167.9600 296.8400 1168.4400 ;
        RECT 295.2400 1184.2800 296.8400 1184.7600 ;
        RECT 340.2400 1184.2800 341.8400 1184.7600 ;
        RECT 245.6800 1200.6000 248.6800 1201.0800 ;
        RECT 245.6800 1195.1600 248.6800 1195.6400 ;
        RECT 245.6800 1189.7200 248.6800 1190.2000 ;
        RECT 245.6800 1178.8400 248.6800 1179.3200 ;
        RECT 245.6800 1173.4000 248.6800 1173.8800 ;
        RECT 245.6800 1167.9600 248.6800 1168.4400 ;
        RECT 245.6800 1162.5200 248.6800 1163.0000 ;
        RECT 245.6800 1184.2800 248.6800 1184.7600 ;
        RECT 340.2400 1146.2000 341.8400 1146.6800 ;
        RECT 340.2400 1151.6400 341.8400 1152.1200 ;
        RECT 340.2400 1129.8800 341.8400 1130.3600 ;
        RECT 340.2400 1135.3200 341.8400 1135.8000 ;
        RECT 340.2400 1140.7600 341.8400 1141.2400 ;
        RECT 295.2400 1146.2000 296.8400 1146.6800 ;
        RECT 295.2400 1151.6400 296.8400 1152.1200 ;
        RECT 295.2400 1129.8800 296.8400 1130.3600 ;
        RECT 295.2400 1135.3200 296.8400 1135.8000 ;
        RECT 295.2400 1140.7600 296.8400 1141.2400 ;
        RECT 340.2400 1119.0000 341.8400 1119.4800 ;
        RECT 340.2400 1124.4400 341.8400 1124.9200 ;
        RECT 340.2400 1102.6800 341.8400 1103.1600 ;
        RECT 340.2400 1108.1200 341.8400 1108.6000 ;
        RECT 340.2400 1113.5600 341.8400 1114.0400 ;
        RECT 295.2400 1119.0000 296.8400 1119.4800 ;
        RECT 295.2400 1124.4400 296.8400 1124.9200 ;
        RECT 295.2400 1102.6800 296.8400 1103.1600 ;
        RECT 295.2400 1108.1200 296.8400 1108.6000 ;
        RECT 295.2400 1113.5600 296.8400 1114.0400 ;
        RECT 245.6800 1146.2000 248.6800 1146.6800 ;
        RECT 245.6800 1151.6400 248.6800 1152.1200 ;
        RECT 245.6800 1135.3200 248.6800 1135.8000 ;
        RECT 245.6800 1129.8800 248.6800 1130.3600 ;
        RECT 245.6800 1140.7600 248.6800 1141.2400 ;
        RECT 245.6800 1119.0000 248.6800 1119.4800 ;
        RECT 245.6800 1124.4400 248.6800 1124.9200 ;
        RECT 245.6800 1108.1200 248.6800 1108.6000 ;
        RECT 245.6800 1102.6800 248.6800 1103.1600 ;
        RECT 245.6800 1113.5600 248.6800 1114.0400 ;
        RECT 245.6800 1157.0800 248.6800 1157.5600 ;
        RECT 295.2400 1157.0800 296.8400 1157.5600 ;
        RECT 340.2400 1157.0800 341.8400 1157.5600 ;
        RECT 441.7800 1091.8000 444.7800 1092.2800 ;
        RECT 441.7800 1097.2400 444.7800 1097.7200 ;
        RECT 430.2400 1091.8000 431.8400 1092.2800 ;
        RECT 430.2400 1097.2400 431.8400 1097.7200 ;
        RECT 441.7800 1075.4800 444.7800 1075.9600 ;
        RECT 441.7800 1080.9200 444.7800 1081.4000 ;
        RECT 441.7800 1086.3600 444.7800 1086.8400 ;
        RECT 430.2400 1075.4800 431.8400 1075.9600 ;
        RECT 430.2400 1080.9200 431.8400 1081.4000 ;
        RECT 430.2400 1086.3600 431.8400 1086.8400 ;
        RECT 441.7800 1064.6000 444.7800 1065.0800 ;
        RECT 441.7800 1070.0400 444.7800 1070.5200 ;
        RECT 430.2400 1064.6000 431.8400 1065.0800 ;
        RECT 430.2400 1070.0400 431.8400 1070.5200 ;
        RECT 441.7800 1048.2800 444.7800 1048.7600 ;
        RECT 441.7800 1053.7200 444.7800 1054.2000 ;
        RECT 441.7800 1059.1600 444.7800 1059.6400 ;
        RECT 430.2400 1048.2800 431.8400 1048.7600 ;
        RECT 430.2400 1053.7200 431.8400 1054.2000 ;
        RECT 430.2400 1059.1600 431.8400 1059.6400 ;
        RECT 385.2400 1091.8000 386.8400 1092.2800 ;
        RECT 385.2400 1097.2400 386.8400 1097.7200 ;
        RECT 385.2400 1075.4800 386.8400 1075.9600 ;
        RECT 385.2400 1080.9200 386.8400 1081.4000 ;
        RECT 385.2400 1086.3600 386.8400 1086.8400 ;
        RECT 385.2400 1064.6000 386.8400 1065.0800 ;
        RECT 385.2400 1070.0400 386.8400 1070.5200 ;
        RECT 385.2400 1048.2800 386.8400 1048.7600 ;
        RECT 385.2400 1053.7200 386.8400 1054.2000 ;
        RECT 385.2400 1059.1600 386.8400 1059.6400 ;
        RECT 441.7800 1037.4000 444.7800 1037.8800 ;
        RECT 441.7800 1042.8400 444.7800 1043.3200 ;
        RECT 430.2400 1037.4000 431.8400 1037.8800 ;
        RECT 430.2400 1042.8400 431.8400 1043.3200 ;
        RECT 441.7800 1021.0800 444.7800 1021.5600 ;
        RECT 441.7800 1026.5200 444.7800 1027.0000 ;
        RECT 441.7800 1031.9600 444.7800 1032.4400 ;
        RECT 430.2400 1021.0800 431.8400 1021.5600 ;
        RECT 430.2400 1026.5200 431.8400 1027.0000 ;
        RECT 430.2400 1031.9600 431.8400 1032.4400 ;
        RECT 441.7800 1010.2000 444.7800 1010.6800 ;
        RECT 441.7800 1015.6400 444.7800 1016.1200 ;
        RECT 430.2400 1010.2000 431.8400 1010.6800 ;
        RECT 430.2400 1015.6400 431.8400 1016.1200 ;
        RECT 441.7800 1004.7600 444.7800 1005.2400 ;
        RECT 430.2400 1004.7600 431.8400 1005.2400 ;
        RECT 385.2400 1037.4000 386.8400 1037.8800 ;
        RECT 385.2400 1042.8400 386.8400 1043.3200 ;
        RECT 385.2400 1021.0800 386.8400 1021.5600 ;
        RECT 385.2400 1026.5200 386.8400 1027.0000 ;
        RECT 385.2400 1031.9600 386.8400 1032.4400 ;
        RECT 385.2400 1010.2000 386.8400 1010.6800 ;
        RECT 385.2400 1015.6400 386.8400 1016.1200 ;
        RECT 385.2400 1004.7600 386.8400 1005.2400 ;
        RECT 340.2400 1091.8000 341.8400 1092.2800 ;
        RECT 340.2400 1097.2400 341.8400 1097.7200 ;
        RECT 340.2400 1075.4800 341.8400 1075.9600 ;
        RECT 340.2400 1080.9200 341.8400 1081.4000 ;
        RECT 340.2400 1086.3600 341.8400 1086.8400 ;
        RECT 295.2400 1091.8000 296.8400 1092.2800 ;
        RECT 295.2400 1097.2400 296.8400 1097.7200 ;
        RECT 295.2400 1075.4800 296.8400 1075.9600 ;
        RECT 295.2400 1080.9200 296.8400 1081.4000 ;
        RECT 295.2400 1086.3600 296.8400 1086.8400 ;
        RECT 340.2400 1064.6000 341.8400 1065.0800 ;
        RECT 340.2400 1070.0400 341.8400 1070.5200 ;
        RECT 340.2400 1048.2800 341.8400 1048.7600 ;
        RECT 340.2400 1053.7200 341.8400 1054.2000 ;
        RECT 340.2400 1059.1600 341.8400 1059.6400 ;
        RECT 295.2400 1064.6000 296.8400 1065.0800 ;
        RECT 295.2400 1070.0400 296.8400 1070.5200 ;
        RECT 295.2400 1048.2800 296.8400 1048.7600 ;
        RECT 295.2400 1053.7200 296.8400 1054.2000 ;
        RECT 295.2400 1059.1600 296.8400 1059.6400 ;
        RECT 245.6800 1091.8000 248.6800 1092.2800 ;
        RECT 245.6800 1097.2400 248.6800 1097.7200 ;
        RECT 245.6800 1080.9200 248.6800 1081.4000 ;
        RECT 245.6800 1075.4800 248.6800 1075.9600 ;
        RECT 245.6800 1086.3600 248.6800 1086.8400 ;
        RECT 245.6800 1064.6000 248.6800 1065.0800 ;
        RECT 245.6800 1070.0400 248.6800 1070.5200 ;
        RECT 245.6800 1053.7200 248.6800 1054.2000 ;
        RECT 245.6800 1048.2800 248.6800 1048.7600 ;
        RECT 245.6800 1059.1600 248.6800 1059.6400 ;
        RECT 340.2400 1037.4000 341.8400 1037.8800 ;
        RECT 340.2400 1042.8400 341.8400 1043.3200 ;
        RECT 340.2400 1021.0800 341.8400 1021.5600 ;
        RECT 340.2400 1026.5200 341.8400 1027.0000 ;
        RECT 340.2400 1031.9600 341.8400 1032.4400 ;
        RECT 295.2400 1037.4000 296.8400 1037.8800 ;
        RECT 295.2400 1042.8400 296.8400 1043.3200 ;
        RECT 295.2400 1021.0800 296.8400 1021.5600 ;
        RECT 295.2400 1026.5200 296.8400 1027.0000 ;
        RECT 295.2400 1031.9600 296.8400 1032.4400 ;
        RECT 340.2400 1015.6400 341.8400 1016.1200 ;
        RECT 340.2400 1010.2000 341.8400 1010.6800 ;
        RECT 340.2400 1004.7600 341.8400 1005.2400 ;
        RECT 295.2400 1015.6400 296.8400 1016.1200 ;
        RECT 295.2400 1010.2000 296.8400 1010.6800 ;
        RECT 295.2400 1004.7600 296.8400 1005.2400 ;
        RECT 245.6800 1037.4000 248.6800 1037.8800 ;
        RECT 245.6800 1042.8400 248.6800 1043.3200 ;
        RECT 245.6800 1026.5200 248.6800 1027.0000 ;
        RECT 245.6800 1021.0800 248.6800 1021.5600 ;
        RECT 245.6800 1031.9600 248.6800 1032.4400 ;
        RECT 245.6800 1010.2000 248.6800 1010.6800 ;
        RECT 245.6800 1015.6400 248.6800 1016.1200 ;
        RECT 245.6800 1004.7600 248.6800 1005.2400 ;
        RECT 245.6800 1202.9500 444.7800 1205.9500 ;
        RECT 245.6800 997.8500 444.7800 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 430.2400 768.2100 431.8400 976.3100 ;
        RECT 385.2400 768.2100 386.8400 976.3100 ;
        RECT 340.2400 768.2100 341.8400 976.3100 ;
        RECT 295.2400 768.2100 296.8400 976.3100 ;
        RECT 441.7800 768.2100 444.7800 976.3100 ;
        RECT 245.6800 768.2100 248.6800 976.3100 ;
      LAYER met3 ;
        RECT 441.7800 970.9600 444.7800 971.4400 ;
        RECT 430.2400 970.9600 431.8400 971.4400 ;
        RECT 441.7800 960.0800 444.7800 960.5600 ;
        RECT 441.7800 965.5200 444.7800 966.0000 ;
        RECT 430.2400 960.0800 431.8400 960.5600 ;
        RECT 430.2400 965.5200 431.8400 966.0000 ;
        RECT 441.7800 943.7600 444.7800 944.2400 ;
        RECT 441.7800 949.2000 444.7800 949.6800 ;
        RECT 430.2400 943.7600 431.8400 944.2400 ;
        RECT 430.2400 949.2000 431.8400 949.6800 ;
        RECT 441.7800 932.8800 444.7800 933.3600 ;
        RECT 441.7800 938.3200 444.7800 938.8000 ;
        RECT 430.2400 932.8800 431.8400 933.3600 ;
        RECT 430.2400 938.3200 431.8400 938.8000 ;
        RECT 441.7800 954.6400 444.7800 955.1200 ;
        RECT 430.2400 954.6400 431.8400 955.1200 ;
        RECT 385.2400 960.0800 386.8400 960.5600 ;
        RECT 385.2400 965.5200 386.8400 966.0000 ;
        RECT 385.2400 970.9600 386.8400 971.4400 ;
        RECT 385.2400 943.7600 386.8400 944.2400 ;
        RECT 385.2400 949.2000 386.8400 949.6800 ;
        RECT 385.2400 938.3200 386.8400 938.8000 ;
        RECT 385.2400 932.8800 386.8400 933.3600 ;
        RECT 385.2400 954.6400 386.8400 955.1200 ;
        RECT 441.7800 916.5600 444.7800 917.0400 ;
        RECT 441.7800 922.0000 444.7800 922.4800 ;
        RECT 430.2400 916.5600 431.8400 917.0400 ;
        RECT 430.2400 922.0000 431.8400 922.4800 ;
        RECT 441.7800 900.2400 444.7800 900.7200 ;
        RECT 441.7800 905.6800 444.7800 906.1600 ;
        RECT 441.7800 911.1200 444.7800 911.6000 ;
        RECT 430.2400 900.2400 431.8400 900.7200 ;
        RECT 430.2400 905.6800 431.8400 906.1600 ;
        RECT 430.2400 911.1200 431.8400 911.6000 ;
        RECT 441.7800 889.3600 444.7800 889.8400 ;
        RECT 441.7800 894.8000 444.7800 895.2800 ;
        RECT 430.2400 889.3600 431.8400 889.8400 ;
        RECT 430.2400 894.8000 431.8400 895.2800 ;
        RECT 441.7800 873.0400 444.7800 873.5200 ;
        RECT 441.7800 878.4800 444.7800 878.9600 ;
        RECT 441.7800 883.9200 444.7800 884.4000 ;
        RECT 430.2400 873.0400 431.8400 873.5200 ;
        RECT 430.2400 878.4800 431.8400 878.9600 ;
        RECT 430.2400 883.9200 431.8400 884.4000 ;
        RECT 385.2400 916.5600 386.8400 917.0400 ;
        RECT 385.2400 922.0000 386.8400 922.4800 ;
        RECT 385.2400 900.2400 386.8400 900.7200 ;
        RECT 385.2400 905.6800 386.8400 906.1600 ;
        RECT 385.2400 911.1200 386.8400 911.6000 ;
        RECT 385.2400 889.3600 386.8400 889.8400 ;
        RECT 385.2400 894.8000 386.8400 895.2800 ;
        RECT 385.2400 873.0400 386.8400 873.5200 ;
        RECT 385.2400 878.4800 386.8400 878.9600 ;
        RECT 385.2400 883.9200 386.8400 884.4000 ;
        RECT 441.7800 927.4400 444.7800 927.9200 ;
        RECT 385.2400 927.4400 386.8400 927.9200 ;
        RECT 430.2400 927.4400 431.8400 927.9200 ;
        RECT 340.2400 960.0800 341.8400 960.5600 ;
        RECT 340.2400 965.5200 341.8400 966.0000 ;
        RECT 340.2400 970.9600 341.8400 971.4400 ;
        RECT 295.2400 960.0800 296.8400 960.5600 ;
        RECT 295.2400 965.5200 296.8400 966.0000 ;
        RECT 295.2400 970.9600 296.8400 971.4400 ;
        RECT 340.2400 943.7600 341.8400 944.2400 ;
        RECT 340.2400 949.2000 341.8400 949.6800 ;
        RECT 340.2400 932.8800 341.8400 933.3600 ;
        RECT 340.2400 938.3200 341.8400 938.8000 ;
        RECT 295.2400 943.7600 296.8400 944.2400 ;
        RECT 295.2400 949.2000 296.8400 949.6800 ;
        RECT 295.2400 932.8800 296.8400 933.3600 ;
        RECT 295.2400 938.3200 296.8400 938.8000 ;
        RECT 295.2400 954.6400 296.8400 955.1200 ;
        RECT 340.2400 954.6400 341.8400 955.1200 ;
        RECT 245.6800 970.9600 248.6800 971.4400 ;
        RECT 245.6800 965.5200 248.6800 966.0000 ;
        RECT 245.6800 960.0800 248.6800 960.5600 ;
        RECT 245.6800 949.2000 248.6800 949.6800 ;
        RECT 245.6800 943.7600 248.6800 944.2400 ;
        RECT 245.6800 938.3200 248.6800 938.8000 ;
        RECT 245.6800 932.8800 248.6800 933.3600 ;
        RECT 245.6800 954.6400 248.6800 955.1200 ;
        RECT 340.2400 916.5600 341.8400 917.0400 ;
        RECT 340.2400 922.0000 341.8400 922.4800 ;
        RECT 340.2400 900.2400 341.8400 900.7200 ;
        RECT 340.2400 905.6800 341.8400 906.1600 ;
        RECT 340.2400 911.1200 341.8400 911.6000 ;
        RECT 295.2400 916.5600 296.8400 917.0400 ;
        RECT 295.2400 922.0000 296.8400 922.4800 ;
        RECT 295.2400 900.2400 296.8400 900.7200 ;
        RECT 295.2400 905.6800 296.8400 906.1600 ;
        RECT 295.2400 911.1200 296.8400 911.6000 ;
        RECT 340.2400 889.3600 341.8400 889.8400 ;
        RECT 340.2400 894.8000 341.8400 895.2800 ;
        RECT 340.2400 873.0400 341.8400 873.5200 ;
        RECT 340.2400 878.4800 341.8400 878.9600 ;
        RECT 340.2400 883.9200 341.8400 884.4000 ;
        RECT 295.2400 889.3600 296.8400 889.8400 ;
        RECT 295.2400 894.8000 296.8400 895.2800 ;
        RECT 295.2400 873.0400 296.8400 873.5200 ;
        RECT 295.2400 878.4800 296.8400 878.9600 ;
        RECT 295.2400 883.9200 296.8400 884.4000 ;
        RECT 245.6800 916.5600 248.6800 917.0400 ;
        RECT 245.6800 922.0000 248.6800 922.4800 ;
        RECT 245.6800 905.6800 248.6800 906.1600 ;
        RECT 245.6800 900.2400 248.6800 900.7200 ;
        RECT 245.6800 911.1200 248.6800 911.6000 ;
        RECT 245.6800 889.3600 248.6800 889.8400 ;
        RECT 245.6800 894.8000 248.6800 895.2800 ;
        RECT 245.6800 878.4800 248.6800 878.9600 ;
        RECT 245.6800 873.0400 248.6800 873.5200 ;
        RECT 245.6800 883.9200 248.6800 884.4000 ;
        RECT 245.6800 927.4400 248.6800 927.9200 ;
        RECT 295.2400 927.4400 296.8400 927.9200 ;
        RECT 340.2400 927.4400 341.8400 927.9200 ;
        RECT 441.7800 862.1600 444.7800 862.6400 ;
        RECT 441.7800 867.6000 444.7800 868.0800 ;
        RECT 430.2400 862.1600 431.8400 862.6400 ;
        RECT 430.2400 867.6000 431.8400 868.0800 ;
        RECT 441.7800 845.8400 444.7800 846.3200 ;
        RECT 441.7800 851.2800 444.7800 851.7600 ;
        RECT 441.7800 856.7200 444.7800 857.2000 ;
        RECT 430.2400 845.8400 431.8400 846.3200 ;
        RECT 430.2400 851.2800 431.8400 851.7600 ;
        RECT 430.2400 856.7200 431.8400 857.2000 ;
        RECT 441.7800 834.9600 444.7800 835.4400 ;
        RECT 441.7800 840.4000 444.7800 840.8800 ;
        RECT 430.2400 834.9600 431.8400 835.4400 ;
        RECT 430.2400 840.4000 431.8400 840.8800 ;
        RECT 441.7800 818.6400 444.7800 819.1200 ;
        RECT 441.7800 824.0800 444.7800 824.5600 ;
        RECT 441.7800 829.5200 444.7800 830.0000 ;
        RECT 430.2400 818.6400 431.8400 819.1200 ;
        RECT 430.2400 824.0800 431.8400 824.5600 ;
        RECT 430.2400 829.5200 431.8400 830.0000 ;
        RECT 385.2400 862.1600 386.8400 862.6400 ;
        RECT 385.2400 867.6000 386.8400 868.0800 ;
        RECT 385.2400 845.8400 386.8400 846.3200 ;
        RECT 385.2400 851.2800 386.8400 851.7600 ;
        RECT 385.2400 856.7200 386.8400 857.2000 ;
        RECT 385.2400 834.9600 386.8400 835.4400 ;
        RECT 385.2400 840.4000 386.8400 840.8800 ;
        RECT 385.2400 818.6400 386.8400 819.1200 ;
        RECT 385.2400 824.0800 386.8400 824.5600 ;
        RECT 385.2400 829.5200 386.8400 830.0000 ;
        RECT 441.7800 807.7600 444.7800 808.2400 ;
        RECT 441.7800 813.2000 444.7800 813.6800 ;
        RECT 430.2400 807.7600 431.8400 808.2400 ;
        RECT 430.2400 813.2000 431.8400 813.6800 ;
        RECT 441.7800 791.4400 444.7800 791.9200 ;
        RECT 441.7800 796.8800 444.7800 797.3600 ;
        RECT 441.7800 802.3200 444.7800 802.8000 ;
        RECT 430.2400 791.4400 431.8400 791.9200 ;
        RECT 430.2400 796.8800 431.8400 797.3600 ;
        RECT 430.2400 802.3200 431.8400 802.8000 ;
        RECT 441.7800 780.5600 444.7800 781.0400 ;
        RECT 441.7800 786.0000 444.7800 786.4800 ;
        RECT 430.2400 780.5600 431.8400 781.0400 ;
        RECT 430.2400 786.0000 431.8400 786.4800 ;
        RECT 441.7800 775.1200 444.7800 775.6000 ;
        RECT 430.2400 775.1200 431.8400 775.6000 ;
        RECT 385.2400 807.7600 386.8400 808.2400 ;
        RECT 385.2400 813.2000 386.8400 813.6800 ;
        RECT 385.2400 791.4400 386.8400 791.9200 ;
        RECT 385.2400 796.8800 386.8400 797.3600 ;
        RECT 385.2400 802.3200 386.8400 802.8000 ;
        RECT 385.2400 780.5600 386.8400 781.0400 ;
        RECT 385.2400 786.0000 386.8400 786.4800 ;
        RECT 385.2400 775.1200 386.8400 775.6000 ;
        RECT 340.2400 862.1600 341.8400 862.6400 ;
        RECT 340.2400 867.6000 341.8400 868.0800 ;
        RECT 340.2400 845.8400 341.8400 846.3200 ;
        RECT 340.2400 851.2800 341.8400 851.7600 ;
        RECT 340.2400 856.7200 341.8400 857.2000 ;
        RECT 295.2400 862.1600 296.8400 862.6400 ;
        RECT 295.2400 867.6000 296.8400 868.0800 ;
        RECT 295.2400 845.8400 296.8400 846.3200 ;
        RECT 295.2400 851.2800 296.8400 851.7600 ;
        RECT 295.2400 856.7200 296.8400 857.2000 ;
        RECT 340.2400 834.9600 341.8400 835.4400 ;
        RECT 340.2400 840.4000 341.8400 840.8800 ;
        RECT 340.2400 818.6400 341.8400 819.1200 ;
        RECT 340.2400 824.0800 341.8400 824.5600 ;
        RECT 340.2400 829.5200 341.8400 830.0000 ;
        RECT 295.2400 834.9600 296.8400 835.4400 ;
        RECT 295.2400 840.4000 296.8400 840.8800 ;
        RECT 295.2400 818.6400 296.8400 819.1200 ;
        RECT 295.2400 824.0800 296.8400 824.5600 ;
        RECT 295.2400 829.5200 296.8400 830.0000 ;
        RECT 245.6800 862.1600 248.6800 862.6400 ;
        RECT 245.6800 867.6000 248.6800 868.0800 ;
        RECT 245.6800 851.2800 248.6800 851.7600 ;
        RECT 245.6800 845.8400 248.6800 846.3200 ;
        RECT 245.6800 856.7200 248.6800 857.2000 ;
        RECT 245.6800 834.9600 248.6800 835.4400 ;
        RECT 245.6800 840.4000 248.6800 840.8800 ;
        RECT 245.6800 824.0800 248.6800 824.5600 ;
        RECT 245.6800 818.6400 248.6800 819.1200 ;
        RECT 245.6800 829.5200 248.6800 830.0000 ;
        RECT 340.2400 807.7600 341.8400 808.2400 ;
        RECT 340.2400 813.2000 341.8400 813.6800 ;
        RECT 340.2400 791.4400 341.8400 791.9200 ;
        RECT 340.2400 796.8800 341.8400 797.3600 ;
        RECT 340.2400 802.3200 341.8400 802.8000 ;
        RECT 295.2400 807.7600 296.8400 808.2400 ;
        RECT 295.2400 813.2000 296.8400 813.6800 ;
        RECT 295.2400 791.4400 296.8400 791.9200 ;
        RECT 295.2400 796.8800 296.8400 797.3600 ;
        RECT 295.2400 802.3200 296.8400 802.8000 ;
        RECT 340.2400 786.0000 341.8400 786.4800 ;
        RECT 340.2400 780.5600 341.8400 781.0400 ;
        RECT 340.2400 775.1200 341.8400 775.6000 ;
        RECT 295.2400 786.0000 296.8400 786.4800 ;
        RECT 295.2400 780.5600 296.8400 781.0400 ;
        RECT 295.2400 775.1200 296.8400 775.6000 ;
        RECT 245.6800 807.7600 248.6800 808.2400 ;
        RECT 245.6800 813.2000 248.6800 813.6800 ;
        RECT 245.6800 796.8800 248.6800 797.3600 ;
        RECT 245.6800 791.4400 248.6800 791.9200 ;
        RECT 245.6800 802.3200 248.6800 802.8000 ;
        RECT 245.6800 780.5600 248.6800 781.0400 ;
        RECT 245.6800 786.0000 248.6800 786.4800 ;
        RECT 245.6800 775.1200 248.6800 775.6000 ;
        RECT 245.6800 973.3100 444.7800 976.3100 ;
        RECT 245.6800 768.2100 444.7800 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 465.9000 2833.6100 467.9000 2854.5400 ;
        RECT 663.0000 2833.6100 665.0000 2854.5400 ;
      LAYER met3 ;
        RECT 663.0000 2850.0400 665.0000 2850.5200 ;
        RECT 465.9000 2850.0400 467.9000 2850.5200 ;
        RECT 663.0000 2839.1600 665.0000 2839.6400 ;
        RECT 465.9000 2839.1600 467.9000 2839.6400 ;
        RECT 663.0000 2844.6000 665.0000 2845.0800 ;
        RECT 465.9000 2844.6000 467.9000 2845.0800 ;
        RECT 465.9000 2852.5400 665.0000 2854.5400 ;
        RECT 465.9000 2833.6100 665.0000 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 538.5700 652.0600 746.6700 ;
        RECT 605.4600 538.5700 607.0600 746.6700 ;
        RECT 560.4600 538.5700 562.0600 746.6700 ;
        RECT 515.4600 538.5700 517.0600 746.6700 ;
        RECT 662.0000 538.5700 665.0000 746.6700 ;
        RECT 465.9000 538.5700 468.9000 746.6700 ;
      LAYER met3 ;
        RECT 662.0000 741.3200 665.0000 741.8000 ;
        RECT 650.4600 741.3200 652.0600 741.8000 ;
        RECT 662.0000 730.4400 665.0000 730.9200 ;
        RECT 662.0000 735.8800 665.0000 736.3600 ;
        RECT 650.4600 730.4400 652.0600 730.9200 ;
        RECT 650.4600 735.8800 652.0600 736.3600 ;
        RECT 662.0000 714.1200 665.0000 714.6000 ;
        RECT 662.0000 719.5600 665.0000 720.0400 ;
        RECT 650.4600 714.1200 652.0600 714.6000 ;
        RECT 650.4600 719.5600 652.0600 720.0400 ;
        RECT 662.0000 703.2400 665.0000 703.7200 ;
        RECT 662.0000 708.6800 665.0000 709.1600 ;
        RECT 650.4600 703.2400 652.0600 703.7200 ;
        RECT 650.4600 708.6800 652.0600 709.1600 ;
        RECT 662.0000 725.0000 665.0000 725.4800 ;
        RECT 650.4600 725.0000 652.0600 725.4800 ;
        RECT 605.4600 730.4400 607.0600 730.9200 ;
        RECT 605.4600 735.8800 607.0600 736.3600 ;
        RECT 605.4600 741.3200 607.0600 741.8000 ;
        RECT 605.4600 714.1200 607.0600 714.6000 ;
        RECT 605.4600 719.5600 607.0600 720.0400 ;
        RECT 605.4600 708.6800 607.0600 709.1600 ;
        RECT 605.4600 703.2400 607.0600 703.7200 ;
        RECT 605.4600 725.0000 607.0600 725.4800 ;
        RECT 662.0000 686.9200 665.0000 687.4000 ;
        RECT 662.0000 692.3600 665.0000 692.8400 ;
        RECT 650.4600 686.9200 652.0600 687.4000 ;
        RECT 650.4600 692.3600 652.0600 692.8400 ;
        RECT 662.0000 670.6000 665.0000 671.0800 ;
        RECT 662.0000 676.0400 665.0000 676.5200 ;
        RECT 662.0000 681.4800 665.0000 681.9600 ;
        RECT 650.4600 670.6000 652.0600 671.0800 ;
        RECT 650.4600 676.0400 652.0600 676.5200 ;
        RECT 650.4600 681.4800 652.0600 681.9600 ;
        RECT 662.0000 659.7200 665.0000 660.2000 ;
        RECT 662.0000 665.1600 665.0000 665.6400 ;
        RECT 650.4600 659.7200 652.0600 660.2000 ;
        RECT 650.4600 665.1600 652.0600 665.6400 ;
        RECT 662.0000 643.4000 665.0000 643.8800 ;
        RECT 662.0000 648.8400 665.0000 649.3200 ;
        RECT 662.0000 654.2800 665.0000 654.7600 ;
        RECT 650.4600 643.4000 652.0600 643.8800 ;
        RECT 650.4600 648.8400 652.0600 649.3200 ;
        RECT 650.4600 654.2800 652.0600 654.7600 ;
        RECT 605.4600 686.9200 607.0600 687.4000 ;
        RECT 605.4600 692.3600 607.0600 692.8400 ;
        RECT 605.4600 670.6000 607.0600 671.0800 ;
        RECT 605.4600 676.0400 607.0600 676.5200 ;
        RECT 605.4600 681.4800 607.0600 681.9600 ;
        RECT 605.4600 659.7200 607.0600 660.2000 ;
        RECT 605.4600 665.1600 607.0600 665.6400 ;
        RECT 605.4600 643.4000 607.0600 643.8800 ;
        RECT 605.4600 648.8400 607.0600 649.3200 ;
        RECT 605.4600 654.2800 607.0600 654.7600 ;
        RECT 662.0000 697.8000 665.0000 698.2800 ;
        RECT 605.4600 697.8000 607.0600 698.2800 ;
        RECT 650.4600 697.8000 652.0600 698.2800 ;
        RECT 560.4600 730.4400 562.0600 730.9200 ;
        RECT 560.4600 735.8800 562.0600 736.3600 ;
        RECT 560.4600 741.3200 562.0600 741.8000 ;
        RECT 515.4600 730.4400 517.0600 730.9200 ;
        RECT 515.4600 735.8800 517.0600 736.3600 ;
        RECT 515.4600 741.3200 517.0600 741.8000 ;
        RECT 560.4600 714.1200 562.0600 714.6000 ;
        RECT 560.4600 719.5600 562.0600 720.0400 ;
        RECT 560.4600 703.2400 562.0600 703.7200 ;
        RECT 560.4600 708.6800 562.0600 709.1600 ;
        RECT 515.4600 714.1200 517.0600 714.6000 ;
        RECT 515.4600 719.5600 517.0600 720.0400 ;
        RECT 515.4600 703.2400 517.0600 703.7200 ;
        RECT 515.4600 708.6800 517.0600 709.1600 ;
        RECT 515.4600 725.0000 517.0600 725.4800 ;
        RECT 560.4600 725.0000 562.0600 725.4800 ;
        RECT 465.9000 741.3200 468.9000 741.8000 ;
        RECT 465.9000 735.8800 468.9000 736.3600 ;
        RECT 465.9000 730.4400 468.9000 730.9200 ;
        RECT 465.9000 719.5600 468.9000 720.0400 ;
        RECT 465.9000 714.1200 468.9000 714.6000 ;
        RECT 465.9000 708.6800 468.9000 709.1600 ;
        RECT 465.9000 703.2400 468.9000 703.7200 ;
        RECT 465.9000 725.0000 468.9000 725.4800 ;
        RECT 560.4600 686.9200 562.0600 687.4000 ;
        RECT 560.4600 692.3600 562.0600 692.8400 ;
        RECT 560.4600 670.6000 562.0600 671.0800 ;
        RECT 560.4600 676.0400 562.0600 676.5200 ;
        RECT 560.4600 681.4800 562.0600 681.9600 ;
        RECT 515.4600 686.9200 517.0600 687.4000 ;
        RECT 515.4600 692.3600 517.0600 692.8400 ;
        RECT 515.4600 670.6000 517.0600 671.0800 ;
        RECT 515.4600 676.0400 517.0600 676.5200 ;
        RECT 515.4600 681.4800 517.0600 681.9600 ;
        RECT 560.4600 659.7200 562.0600 660.2000 ;
        RECT 560.4600 665.1600 562.0600 665.6400 ;
        RECT 560.4600 643.4000 562.0600 643.8800 ;
        RECT 560.4600 648.8400 562.0600 649.3200 ;
        RECT 560.4600 654.2800 562.0600 654.7600 ;
        RECT 515.4600 659.7200 517.0600 660.2000 ;
        RECT 515.4600 665.1600 517.0600 665.6400 ;
        RECT 515.4600 643.4000 517.0600 643.8800 ;
        RECT 515.4600 648.8400 517.0600 649.3200 ;
        RECT 515.4600 654.2800 517.0600 654.7600 ;
        RECT 465.9000 686.9200 468.9000 687.4000 ;
        RECT 465.9000 692.3600 468.9000 692.8400 ;
        RECT 465.9000 676.0400 468.9000 676.5200 ;
        RECT 465.9000 670.6000 468.9000 671.0800 ;
        RECT 465.9000 681.4800 468.9000 681.9600 ;
        RECT 465.9000 659.7200 468.9000 660.2000 ;
        RECT 465.9000 665.1600 468.9000 665.6400 ;
        RECT 465.9000 648.8400 468.9000 649.3200 ;
        RECT 465.9000 643.4000 468.9000 643.8800 ;
        RECT 465.9000 654.2800 468.9000 654.7600 ;
        RECT 465.9000 697.8000 468.9000 698.2800 ;
        RECT 515.4600 697.8000 517.0600 698.2800 ;
        RECT 560.4600 697.8000 562.0600 698.2800 ;
        RECT 662.0000 632.5200 665.0000 633.0000 ;
        RECT 662.0000 637.9600 665.0000 638.4400 ;
        RECT 650.4600 632.5200 652.0600 633.0000 ;
        RECT 650.4600 637.9600 652.0600 638.4400 ;
        RECT 662.0000 616.2000 665.0000 616.6800 ;
        RECT 662.0000 621.6400 665.0000 622.1200 ;
        RECT 662.0000 627.0800 665.0000 627.5600 ;
        RECT 650.4600 616.2000 652.0600 616.6800 ;
        RECT 650.4600 621.6400 652.0600 622.1200 ;
        RECT 650.4600 627.0800 652.0600 627.5600 ;
        RECT 662.0000 605.3200 665.0000 605.8000 ;
        RECT 662.0000 610.7600 665.0000 611.2400 ;
        RECT 650.4600 605.3200 652.0600 605.8000 ;
        RECT 650.4600 610.7600 652.0600 611.2400 ;
        RECT 662.0000 589.0000 665.0000 589.4800 ;
        RECT 662.0000 594.4400 665.0000 594.9200 ;
        RECT 662.0000 599.8800 665.0000 600.3600 ;
        RECT 650.4600 589.0000 652.0600 589.4800 ;
        RECT 650.4600 594.4400 652.0600 594.9200 ;
        RECT 650.4600 599.8800 652.0600 600.3600 ;
        RECT 605.4600 632.5200 607.0600 633.0000 ;
        RECT 605.4600 637.9600 607.0600 638.4400 ;
        RECT 605.4600 616.2000 607.0600 616.6800 ;
        RECT 605.4600 621.6400 607.0600 622.1200 ;
        RECT 605.4600 627.0800 607.0600 627.5600 ;
        RECT 605.4600 605.3200 607.0600 605.8000 ;
        RECT 605.4600 610.7600 607.0600 611.2400 ;
        RECT 605.4600 589.0000 607.0600 589.4800 ;
        RECT 605.4600 594.4400 607.0600 594.9200 ;
        RECT 605.4600 599.8800 607.0600 600.3600 ;
        RECT 662.0000 578.1200 665.0000 578.6000 ;
        RECT 662.0000 583.5600 665.0000 584.0400 ;
        RECT 650.4600 578.1200 652.0600 578.6000 ;
        RECT 650.4600 583.5600 652.0600 584.0400 ;
        RECT 662.0000 561.8000 665.0000 562.2800 ;
        RECT 662.0000 567.2400 665.0000 567.7200 ;
        RECT 662.0000 572.6800 665.0000 573.1600 ;
        RECT 650.4600 561.8000 652.0600 562.2800 ;
        RECT 650.4600 567.2400 652.0600 567.7200 ;
        RECT 650.4600 572.6800 652.0600 573.1600 ;
        RECT 662.0000 550.9200 665.0000 551.4000 ;
        RECT 662.0000 556.3600 665.0000 556.8400 ;
        RECT 650.4600 550.9200 652.0600 551.4000 ;
        RECT 650.4600 556.3600 652.0600 556.8400 ;
        RECT 662.0000 545.4800 665.0000 545.9600 ;
        RECT 650.4600 545.4800 652.0600 545.9600 ;
        RECT 605.4600 578.1200 607.0600 578.6000 ;
        RECT 605.4600 583.5600 607.0600 584.0400 ;
        RECT 605.4600 561.8000 607.0600 562.2800 ;
        RECT 605.4600 567.2400 607.0600 567.7200 ;
        RECT 605.4600 572.6800 607.0600 573.1600 ;
        RECT 605.4600 550.9200 607.0600 551.4000 ;
        RECT 605.4600 556.3600 607.0600 556.8400 ;
        RECT 605.4600 545.4800 607.0600 545.9600 ;
        RECT 560.4600 632.5200 562.0600 633.0000 ;
        RECT 560.4600 637.9600 562.0600 638.4400 ;
        RECT 560.4600 616.2000 562.0600 616.6800 ;
        RECT 560.4600 621.6400 562.0600 622.1200 ;
        RECT 560.4600 627.0800 562.0600 627.5600 ;
        RECT 515.4600 632.5200 517.0600 633.0000 ;
        RECT 515.4600 637.9600 517.0600 638.4400 ;
        RECT 515.4600 616.2000 517.0600 616.6800 ;
        RECT 515.4600 621.6400 517.0600 622.1200 ;
        RECT 515.4600 627.0800 517.0600 627.5600 ;
        RECT 560.4600 605.3200 562.0600 605.8000 ;
        RECT 560.4600 610.7600 562.0600 611.2400 ;
        RECT 560.4600 589.0000 562.0600 589.4800 ;
        RECT 560.4600 594.4400 562.0600 594.9200 ;
        RECT 560.4600 599.8800 562.0600 600.3600 ;
        RECT 515.4600 605.3200 517.0600 605.8000 ;
        RECT 515.4600 610.7600 517.0600 611.2400 ;
        RECT 515.4600 589.0000 517.0600 589.4800 ;
        RECT 515.4600 594.4400 517.0600 594.9200 ;
        RECT 515.4600 599.8800 517.0600 600.3600 ;
        RECT 465.9000 632.5200 468.9000 633.0000 ;
        RECT 465.9000 637.9600 468.9000 638.4400 ;
        RECT 465.9000 621.6400 468.9000 622.1200 ;
        RECT 465.9000 616.2000 468.9000 616.6800 ;
        RECT 465.9000 627.0800 468.9000 627.5600 ;
        RECT 465.9000 605.3200 468.9000 605.8000 ;
        RECT 465.9000 610.7600 468.9000 611.2400 ;
        RECT 465.9000 594.4400 468.9000 594.9200 ;
        RECT 465.9000 589.0000 468.9000 589.4800 ;
        RECT 465.9000 599.8800 468.9000 600.3600 ;
        RECT 560.4600 578.1200 562.0600 578.6000 ;
        RECT 560.4600 583.5600 562.0600 584.0400 ;
        RECT 560.4600 561.8000 562.0600 562.2800 ;
        RECT 560.4600 567.2400 562.0600 567.7200 ;
        RECT 560.4600 572.6800 562.0600 573.1600 ;
        RECT 515.4600 578.1200 517.0600 578.6000 ;
        RECT 515.4600 583.5600 517.0600 584.0400 ;
        RECT 515.4600 561.8000 517.0600 562.2800 ;
        RECT 515.4600 567.2400 517.0600 567.7200 ;
        RECT 515.4600 572.6800 517.0600 573.1600 ;
        RECT 560.4600 556.3600 562.0600 556.8400 ;
        RECT 560.4600 550.9200 562.0600 551.4000 ;
        RECT 560.4600 545.4800 562.0600 545.9600 ;
        RECT 515.4600 556.3600 517.0600 556.8400 ;
        RECT 515.4600 550.9200 517.0600 551.4000 ;
        RECT 515.4600 545.4800 517.0600 545.9600 ;
        RECT 465.9000 578.1200 468.9000 578.6000 ;
        RECT 465.9000 583.5600 468.9000 584.0400 ;
        RECT 465.9000 567.2400 468.9000 567.7200 ;
        RECT 465.9000 561.8000 468.9000 562.2800 ;
        RECT 465.9000 572.6800 468.9000 573.1600 ;
        RECT 465.9000 550.9200 468.9000 551.4000 ;
        RECT 465.9000 556.3600 468.9000 556.8400 ;
        RECT 465.9000 545.4800 468.9000 545.9600 ;
        RECT 465.9000 743.6700 665.0000 746.6700 ;
        RECT 465.9000 538.5700 665.0000 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 308.9300 652.0600 517.0300 ;
        RECT 605.4600 308.9300 607.0600 517.0300 ;
        RECT 560.4600 308.9300 562.0600 517.0300 ;
        RECT 515.4600 308.9300 517.0600 517.0300 ;
        RECT 662.0000 308.9300 665.0000 517.0300 ;
        RECT 465.9000 308.9300 468.9000 517.0300 ;
      LAYER met3 ;
        RECT 662.0000 511.6800 665.0000 512.1600 ;
        RECT 650.4600 511.6800 652.0600 512.1600 ;
        RECT 662.0000 500.8000 665.0000 501.2800 ;
        RECT 662.0000 506.2400 665.0000 506.7200 ;
        RECT 650.4600 500.8000 652.0600 501.2800 ;
        RECT 650.4600 506.2400 652.0600 506.7200 ;
        RECT 662.0000 484.4800 665.0000 484.9600 ;
        RECT 662.0000 489.9200 665.0000 490.4000 ;
        RECT 650.4600 484.4800 652.0600 484.9600 ;
        RECT 650.4600 489.9200 652.0600 490.4000 ;
        RECT 662.0000 473.6000 665.0000 474.0800 ;
        RECT 662.0000 479.0400 665.0000 479.5200 ;
        RECT 650.4600 473.6000 652.0600 474.0800 ;
        RECT 650.4600 479.0400 652.0600 479.5200 ;
        RECT 662.0000 495.3600 665.0000 495.8400 ;
        RECT 650.4600 495.3600 652.0600 495.8400 ;
        RECT 605.4600 500.8000 607.0600 501.2800 ;
        RECT 605.4600 506.2400 607.0600 506.7200 ;
        RECT 605.4600 511.6800 607.0600 512.1600 ;
        RECT 605.4600 484.4800 607.0600 484.9600 ;
        RECT 605.4600 489.9200 607.0600 490.4000 ;
        RECT 605.4600 479.0400 607.0600 479.5200 ;
        RECT 605.4600 473.6000 607.0600 474.0800 ;
        RECT 605.4600 495.3600 607.0600 495.8400 ;
        RECT 662.0000 457.2800 665.0000 457.7600 ;
        RECT 662.0000 462.7200 665.0000 463.2000 ;
        RECT 650.4600 457.2800 652.0600 457.7600 ;
        RECT 650.4600 462.7200 652.0600 463.2000 ;
        RECT 662.0000 440.9600 665.0000 441.4400 ;
        RECT 662.0000 446.4000 665.0000 446.8800 ;
        RECT 662.0000 451.8400 665.0000 452.3200 ;
        RECT 650.4600 440.9600 652.0600 441.4400 ;
        RECT 650.4600 446.4000 652.0600 446.8800 ;
        RECT 650.4600 451.8400 652.0600 452.3200 ;
        RECT 662.0000 430.0800 665.0000 430.5600 ;
        RECT 662.0000 435.5200 665.0000 436.0000 ;
        RECT 650.4600 430.0800 652.0600 430.5600 ;
        RECT 650.4600 435.5200 652.0600 436.0000 ;
        RECT 662.0000 413.7600 665.0000 414.2400 ;
        RECT 662.0000 419.2000 665.0000 419.6800 ;
        RECT 662.0000 424.6400 665.0000 425.1200 ;
        RECT 650.4600 413.7600 652.0600 414.2400 ;
        RECT 650.4600 419.2000 652.0600 419.6800 ;
        RECT 650.4600 424.6400 652.0600 425.1200 ;
        RECT 605.4600 457.2800 607.0600 457.7600 ;
        RECT 605.4600 462.7200 607.0600 463.2000 ;
        RECT 605.4600 440.9600 607.0600 441.4400 ;
        RECT 605.4600 446.4000 607.0600 446.8800 ;
        RECT 605.4600 451.8400 607.0600 452.3200 ;
        RECT 605.4600 430.0800 607.0600 430.5600 ;
        RECT 605.4600 435.5200 607.0600 436.0000 ;
        RECT 605.4600 413.7600 607.0600 414.2400 ;
        RECT 605.4600 419.2000 607.0600 419.6800 ;
        RECT 605.4600 424.6400 607.0600 425.1200 ;
        RECT 662.0000 468.1600 665.0000 468.6400 ;
        RECT 605.4600 468.1600 607.0600 468.6400 ;
        RECT 650.4600 468.1600 652.0600 468.6400 ;
        RECT 560.4600 500.8000 562.0600 501.2800 ;
        RECT 560.4600 506.2400 562.0600 506.7200 ;
        RECT 560.4600 511.6800 562.0600 512.1600 ;
        RECT 515.4600 500.8000 517.0600 501.2800 ;
        RECT 515.4600 506.2400 517.0600 506.7200 ;
        RECT 515.4600 511.6800 517.0600 512.1600 ;
        RECT 560.4600 484.4800 562.0600 484.9600 ;
        RECT 560.4600 489.9200 562.0600 490.4000 ;
        RECT 560.4600 473.6000 562.0600 474.0800 ;
        RECT 560.4600 479.0400 562.0600 479.5200 ;
        RECT 515.4600 484.4800 517.0600 484.9600 ;
        RECT 515.4600 489.9200 517.0600 490.4000 ;
        RECT 515.4600 473.6000 517.0600 474.0800 ;
        RECT 515.4600 479.0400 517.0600 479.5200 ;
        RECT 515.4600 495.3600 517.0600 495.8400 ;
        RECT 560.4600 495.3600 562.0600 495.8400 ;
        RECT 465.9000 511.6800 468.9000 512.1600 ;
        RECT 465.9000 506.2400 468.9000 506.7200 ;
        RECT 465.9000 500.8000 468.9000 501.2800 ;
        RECT 465.9000 489.9200 468.9000 490.4000 ;
        RECT 465.9000 484.4800 468.9000 484.9600 ;
        RECT 465.9000 479.0400 468.9000 479.5200 ;
        RECT 465.9000 473.6000 468.9000 474.0800 ;
        RECT 465.9000 495.3600 468.9000 495.8400 ;
        RECT 560.4600 457.2800 562.0600 457.7600 ;
        RECT 560.4600 462.7200 562.0600 463.2000 ;
        RECT 560.4600 440.9600 562.0600 441.4400 ;
        RECT 560.4600 446.4000 562.0600 446.8800 ;
        RECT 560.4600 451.8400 562.0600 452.3200 ;
        RECT 515.4600 457.2800 517.0600 457.7600 ;
        RECT 515.4600 462.7200 517.0600 463.2000 ;
        RECT 515.4600 440.9600 517.0600 441.4400 ;
        RECT 515.4600 446.4000 517.0600 446.8800 ;
        RECT 515.4600 451.8400 517.0600 452.3200 ;
        RECT 560.4600 430.0800 562.0600 430.5600 ;
        RECT 560.4600 435.5200 562.0600 436.0000 ;
        RECT 560.4600 413.7600 562.0600 414.2400 ;
        RECT 560.4600 419.2000 562.0600 419.6800 ;
        RECT 560.4600 424.6400 562.0600 425.1200 ;
        RECT 515.4600 430.0800 517.0600 430.5600 ;
        RECT 515.4600 435.5200 517.0600 436.0000 ;
        RECT 515.4600 413.7600 517.0600 414.2400 ;
        RECT 515.4600 419.2000 517.0600 419.6800 ;
        RECT 515.4600 424.6400 517.0600 425.1200 ;
        RECT 465.9000 457.2800 468.9000 457.7600 ;
        RECT 465.9000 462.7200 468.9000 463.2000 ;
        RECT 465.9000 446.4000 468.9000 446.8800 ;
        RECT 465.9000 440.9600 468.9000 441.4400 ;
        RECT 465.9000 451.8400 468.9000 452.3200 ;
        RECT 465.9000 430.0800 468.9000 430.5600 ;
        RECT 465.9000 435.5200 468.9000 436.0000 ;
        RECT 465.9000 419.2000 468.9000 419.6800 ;
        RECT 465.9000 413.7600 468.9000 414.2400 ;
        RECT 465.9000 424.6400 468.9000 425.1200 ;
        RECT 465.9000 468.1600 468.9000 468.6400 ;
        RECT 515.4600 468.1600 517.0600 468.6400 ;
        RECT 560.4600 468.1600 562.0600 468.6400 ;
        RECT 662.0000 402.8800 665.0000 403.3600 ;
        RECT 662.0000 408.3200 665.0000 408.8000 ;
        RECT 650.4600 402.8800 652.0600 403.3600 ;
        RECT 650.4600 408.3200 652.0600 408.8000 ;
        RECT 662.0000 386.5600 665.0000 387.0400 ;
        RECT 662.0000 392.0000 665.0000 392.4800 ;
        RECT 662.0000 397.4400 665.0000 397.9200 ;
        RECT 650.4600 386.5600 652.0600 387.0400 ;
        RECT 650.4600 392.0000 652.0600 392.4800 ;
        RECT 650.4600 397.4400 652.0600 397.9200 ;
        RECT 662.0000 375.6800 665.0000 376.1600 ;
        RECT 662.0000 381.1200 665.0000 381.6000 ;
        RECT 650.4600 375.6800 652.0600 376.1600 ;
        RECT 650.4600 381.1200 652.0600 381.6000 ;
        RECT 662.0000 359.3600 665.0000 359.8400 ;
        RECT 662.0000 364.8000 665.0000 365.2800 ;
        RECT 662.0000 370.2400 665.0000 370.7200 ;
        RECT 650.4600 359.3600 652.0600 359.8400 ;
        RECT 650.4600 364.8000 652.0600 365.2800 ;
        RECT 650.4600 370.2400 652.0600 370.7200 ;
        RECT 605.4600 402.8800 607.0600 403.3600 ;
        RECT 605.4600 408.3200 607.0600 408.8000 ;
        RECT 605.4600 386.5600 607.0600 387.0400 ;
        RECT 605.4600 392.0000 607.0600 392.4800 ;
        RECT 605.4600 397.4400 607.0600 397.9200 ;
        RECT 605.4600 375.6800 607.0600 376.1600 ;
        RECT 605.4600 381.1200 607.0600 381.6000 ;
        RECT 605.4600 359.3600 607.0600 359.8400 ;
        RECT 605.4600 364.8000 607.0600 365.2800 ;
        RECT 605.4600 370.2400 607.0600 370.7200 ;
        RECT 662.0000 348.4800 665.0000 348.9600 ;
        RECT 662.0000 353.9200 665.0000 354.4000 ;
        RECT 650.4600 348.4800 652.0600 348.9600 ;
        RECT 650.4600 353.9200 652.0600 354.4000 ;
        RECT 662.0000 332.1600 665.0000 332.6400 ;
        RECT 662.0000 337.6000 665.0000 338.0800 ;
        RECT 662.0000 343.0400 665.0000 343.5200 ;
        RECT 650.4600 332.1600 652.0600 332.6400 ;
        RECT 650.4600 337.6000 652.0600 338.0800 ;
        RECT 650.4600 343.0400 652.0600 343.5200 ;
        RECT 662.0000 321.2800 665.0000 321.7600 ;
        RECT 662.0000 326.7200 665.0000 327.2000 ;
        RECT 650.4600 321.2800 652.0600 321.7600 ;
        RECT 650.4600 326.7200 652.0600 327.2000 ;
        RECT 662.0000 315.8400 665.0000 316.3200 ;
        RECT 650.4600 315.8400 652.0600 316.3200 ;
        RECT 605.4600 348.4800 607.0600 348.9600 ;
        RECT 605.4600 353.9200 607.0600 354.4000 ;
        RECT 605.4600 332.1600 607.0600 332.6400 ;
        RECT 605.4600 337.6000 607.0600 338.0800 ;
        RECT 605.4600 343.0400 607.0600 343.5200 ;
        RECT 605.4600 321.2800 607.0600 321.7600 ;
        RECT 605.4600 326.7200 607.0600 327.2000 ;
        RECT 605.4600 315.8400 607.0600 316.3200 ;
        RECT 560.4600 402.8800 562.0600 403.3600 ;
        RECT 560.4600 408.3200 562.0600 408.8000 ;
        RECT 560.4600 386.5600 562.0600 387.0400 ;
        RECT 560.4600 392.0000 562.0600 392.4800 ;
        RECT 560.4600 397.4400 562.0600 397.9200 ;
        RECT 515.4600 402.8800 517.0600 403.3600 ;
        RECT 515.4600 408.3200 517.0600 408.8000 ;
        RECT 515.4600 386.5600 517.0600 387.0400 ;
        RECT 515.4600 392.0000 517.0600 392.4800 ;
        RECT 515.4600 397.4400 517.0600 397.9200 ;
        RECT 560.4600 375.6800 562.0600 376.1600 ;
        RECT 560.4600 381.1200 562.0600 381.6000 ;
        RECT 560.4600 359.3600 562.0600 359.8400 ;
        RECT 560.4600 364.8000 562.0600 365.2800 ;
        RECT 560.4600 370.2400 562.0600 370.7200 ;
        RECT 515.4600 375.6800 517.0600 376.1600 ;
        RECT 515.4600 381.1200 517.0600 381.6000 ;
        RECT 515.4600 359.3600 517.0600 359.8400 ;
        RECT 515.4600 364.8000 517.0600 365.2800 ;
        RECT 515.4600 370.2400 517.0600 370.7200 ;
        RECT 465.9000 402.8800 468.9000 403.3600 ;
        RECT 465.9000 408.3200 468.9000 408.8000 ;
        RECT 465.9000 392.0000 468.9000 392.4800 ;
        RECT 465.9000 386.5600 468.9000 387.0400 ;
        RECT 465.9000 397.4400 468.9000 397.9200 ;
        RECT 465.9000 375.6800 468.9000 376.1600 ;
        RECT 465.9000 381.1200 468.9000 381.6000 ;
        RECT 465.9000 364.8000 468.9000 365.2800 ;
        RECT 465.9000 359.3600 468.9000 359.8400 ;
        RECT 465.9000 370.2400 468.9000 370.7200 ;
        RECT 560.4600 348.4800 562.0600 348.9600 ;
        RECT 560.4600 353.9200 562.0600 354.4000 ;
        RECT 560.4600 332.1600 562.0600 332.6400 ;
        RECT 560.4600 337.6000 562.0600 338.0800 ;
        RECT 560.4600 343.0400 562.0600 343.5200 ;
        RECT 515.4600 348.4800 517.0600 348.9600 ;
        RECT 515.4600 353.9200 517.0600 354.4000 ;
        RECT 515.4600 332.1600 517.0600 332.6400 ;
        RECT 515.4600 337.6000 517.0600 338.0800 ;
        RECT 515.4600 343.0400 517.0600 343.5200 ;
        RECT 560.4600 326.7200 562.0600 327.2000 ;
        RECT 560.4600 321.2800 562.0600 321.7600 ;
        RECT 560.4600 315.8400 562.0600 316.3200 ;
        RECT 515.4600 326.7200 517.0600 327.2000 ;
        RECT 515.4600 321.2800 517.0600 321.7600 ;
        RECT 515.4600 315.8400 517.0600 316.3200 ;
        RECT 465.9000 348.4800 468.9000 348.9600 ;
        RECT 465.9000 353.9200 468.9000 354.4000 ;
        RECT 465.9000 337.6000 468.9000 338.0800 ;
        RECT 465.9000 332.1600 468.9000 332.6400 ;
        RECT 465.9000 343.0400 468.9000 343.5200 ;
        RECT 465.9000 321.2800 468.9000 321.7600 ;
        RECT 465.9000 326.7200 468.9000 327.2000 ;
        RECT 465.9000 315.8400 468.9000 316.3200 ;
        RECT 465.9000 514.0300 665.0000 517.0300 ;
        RECT 465.9000 308.9300 665.0000 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 79.2900 652.0600 287.3900 ;
        RECT 605.4600 79.2900 607.0600 287.3900 ;
        RECT 560.4600 79.2900 562.0600 287.3900 ;
        RECT 515.4600 79.2900 517.0600 287.3900 ;
        RECT 662.0000 79.2900 665.0000 287.3900 ;
        RECT 465.9000 79.2900 468.9000 287.3900 ;
      LAYER met3 ;
        RECT 662.0000 282.0400 665.0000 282.5200 ;
        RECT 650.4600 282.0400 652.0600 282.5200 ;
        RECT 662.0000 271.1600 665.0000 271.6400 ;
        RECT 662.0000 276.6000 665.0000 277.0800 ;
        RECT 650.4600 271.1600 652.0600 271.6400 ;
        RECT 650.4600 276.6000 652.0600 277.0800 ;
        RECT 662.0000 254.8400 665.0000 255.3200 ;
        RECT 662.0000 260.2800 665.0000 260.7600 ;
        RECT 650.4600 254.8400 652.0600 255.3200 ;
        RECT 650.4600 260.2800 652.0600 260.7600 ;
        RECT 662.0000 243.9600 665.0000 244.4400 ;
        RECT 662.0000 249.4000 665.0000 249.8800 ;
        RECT 650.4600 243.9600 652.0600 244.4400 ;
        RECT 650.4600 249.4000 652.0600 249.8800 ;
        RECT 662.0000 265.7200 665.0000 266.2000 ;
        RECT 650.4600 265.7200 652.0600 266.2000 ;
        RECT 605.4600 271.1600 607.0600 271.6400 ;
        RECT 605.4600 276.6000 607.0600 277.0800 ;
        RECT 605.4600 282.0400 607.0600 282.5200 ;
        RECT 605.4600 254.8400 607.0600 255.3200 ;
        RECT 605.4600 260.2800 607.0600 260.7600 ;
        RECT 605.4600 249.4000 607.0600 249.8800 ;
        RECT 605.4600 243.9600 607.0600 244.4400 ;
        RECT 605.4600 265.7200 607.0600 266.2000 ;
        RECT 662.0000 227.6400 665.0000 228.1200 ;
        RECT 662.0000 233.0800 665.0000 233.5600 ;
        RECT 650.4600 227.6400 652.0600 228.1200 ;
        RECT 650.4600 233.0800 652.0600 233.5600 ;
        RECT 662.0000 211.3200 665.0000 211.8000 ;
        RECT 662.0000 216.7600 665.0000 217.2400 ;
        RECT 662.0000 222.2000 665.0000 222.6800 ;
        RECT 650.4600 211.3200 652.0600 211.8000 ;
        RECT 650.4600 216.7600 652.0600 217.2400 ;
        RECT 650.4600 222.2000 652.0600 222.6800 ;
        RECT 662.0000 200.4400 665.0000 200.9200 ;
        RECT 662.0000 205.8800 665.0000 206.3600 ;
        RECT 650.4600 200.4400 652.0600 200.9200 ;
        RECT 650.4600 205.8800 652.0600 206.3600 ;
        RECT 662.0000 184.1200 665.0000 184.6000 ;
        RECT 662.0000 189.5600 665.0000 190.0400 ;
        RECT 662.0000 195.0000 665.0000 195.4800 ;
        RECT 650.4600 184.1200 652.0600 184.6000 ;
        RECT 650.4600 189.5600 652.0600 190.0400 ;
        RECT 650.4600 195.0000 652.0600 195.4800 ;
        RECT 605.4600 227.6400 607.0600 228.1200 ;
        RECT 605.4600 233.0800 607.0600 233.5600 ;
        RECT 605.4600 211.3200 607.0600 211.8000 ;
        RECT 605.4600 216.7600 607.0600 217.2400 ;
        RECT 605.4600 222.2000 607.0600 222.6800 ;
        RECT 605.4600 200.4400 607.0600 200.9200 ;
        RECT 605.4600 205.8800 607.0600 206.3600 ;
        RECT 605.4600 184.1200 607.0600 184.6000 ;
        RECT 605.4600 189.5600 607.0600 190.0400 ;
        RECT 605.4600 195.0000 607.0600 195.4800 ;
        RECT 662.0000 238.5200 665.0000 239.0000 ;
        RECT 605.4600 238.5200 607.0600 239.0000 ;
        RECT 650.4600 238.5200 652.0600 239.0000 ;
        RECT 560.4600 271.1600 562.0600 271.6400 ;
        RECT 560.4600 276.6000 562.0600 277.0800 ;
        RECT 560.4600 282.0400 562.0600 282.5200 ;
        RECT 515.4600 271.1600 517.0600 271.6400 ;
        RECT 515.4600 276.6000 517.0600 277.0800 ;
        RECT 515.4600 282.0400 517.0600 282.5200 ;
        RECT 560.4600 254.8400 562.0600 255.3200 ;
        RECT 560.4600 260.2800 562.0600 260.7600 ;
        RECT 560.4600 243.9600 562.0600 244.4400 ;
        RECT 560.4600 249.4000 562.0600 249.8800 ;
        RECT 515.4600 254.8400 517.0600 255.3200 ;
        RECT 515.4600 260.2800 517.0600 260.7600 ;
        RECT 515.4600 243.9600 517.0600 244.4400 ;
        RECT 515.4600 249.4000 517.0600 249.8800 ;
        RECT 515.4600 265.7200 517.0600 266.2000 ;
        RECT 560.4600 265.7200 562.0600 266.2000 ;
        RECT 465.9000 282.0400 468.9000 282.5200 ;
        RECT 465.9000 276.6000 468.9000 277.0800 ;
        RECT 465.9000 271.1600 468.9000 271.6400 ;
        RECT 465.9000 260.2800 468.9000 260.7600 ;
        RECT 465.9000 254.8400 468.9000 255.3200 ;
        RECT 465.9000 249.4000 468.9000 249.8800 ;
        RECT 465.9000 243.9600 468.9000 244.4400 ;
        RECT 465.9000 265.7200 468.9000 266.2000 ;
        RECT 560.4600 227.6400 562.0600 228.1200 ;
        RECT 560.4600 233.0800 562.0600 233.5600 ;
        RECT 560.4600 211.3200 562.0600 211.8000 ;
        RECT 560.4600 216.7600 562.0600 217.2400 ;
        RECT 560.4600 222.2000 562.0600 222.6800 ;
        RECT 515.4600 227.6400 517.0600 228.1200 ;
        RECT 515.4600 233.0800 517.0600 233.5600 ;
        RECT 515.4600 211.3200 517.0600 211.8000 ;
        RECT 515.4600 216.7600 517.0600 217.2400 ;
        RECT 515.4600 222.2000 517.0600 222.6800 ;
        RECT 560.4600 200.4400 562.0600 200.9200 ;
        RECT 560.4600 205.8800 562.0600 206.3600 ;
        RECT 560.4600 184.1200 562.0600 184.6000 ;
        RECT 560.4600 189.5600 562.0600 190.0400 ;
        RECT 560.4600 195.0000 562.0600 195.4800 ;
        RECT 515.4600 200.4400 517.0600 200.9200 ;
        RECT 515.4600 205.8800 517.0600 206.3600 ;
        RECT 515.4600 184.1200 517.0600 184.6000 ;
        RECT 515.4600 189.5600 517.0600 190.0400 ;
        RECT 515.4600 195.0000 517.0600 195.4800 ;
        RECT 465.9000 227.6400 468.9000 228.1200 ;
        RECT 465.9000 233.0800 468.9000 233.5600 ;
        RECT 465.9000 216.7600 468.9000 217.2400 ;
        RECT 465.9000 211.3200 468.9000 211.8000 ;
        RECT 465.9000 222.2000 468.9000 222.6800 ;
        RECT 465.9000 200.4400 468.9000 200.9200 ;
        RECT 465.9000 205.8800 468.9000 206.3600 ;
        RECT 465.9000 189.5600 468.9000 190.0400 ;
        RECT 465.9000 184.1200 468.9000 184.6000 ;
        RECT 465.9000 195.0000 468.9000 195.4800 ;
        RECT 465.9000 238.5200 468.9000 239.0000 ;
        RECT 515.4600 238.5200 517.0600 239.0000 ;
        RECT 560.4600 238.5200 562.0600 239.0000 ;
        RECT 662.0000 173.2400 665.0000 173.7200 ;
        RECT 662.0000 178.6800 665.0000 179.1600 ;
        RECT 650.4600 173.2400 652.0600 173.7200 ;
        RECT 650.4600 178.6800 652.0600 179.1600 ;
        RECT 662.0000 156.9200 665.0000 157.4000 ;
        RECT 662.0000 162.3600 665.0000 162.8400 ;
        RECT 662.0000 167.8000 665.0000 168.2800 ;
        RECT 650.4600 156.9200 652.0600 157.4000 ;
        RECT 650.4600 162.3600 652.0600 162.8400 ;
        RECT 650.4600 167.8000 652.0600 168.2800 ;
        RECT 662.0000 146.0400 665.0000 146.5200 ;
        RECT 662.0000 151.4800 665.0000 151.9600 ;
        RECT 650.4600 146.0400 652.0600 146.5200 ;
        RECT 650.4600 151.4800 652.0600 151.9600 ;
        RECT 662.0000 129.7200 665.0000 130.2000 ;
        RECT 662.0000 135.1600 665.0000 135.6400 ;
        RECT 662.0000 140.6000 665.0000 141.0800 ;
        RECT 650.4600 129.7200 652.0600 130.2000 ;
        RECT 650.4600 135.1600 652.0600 135.6400 ;
        RECT 650.4600 140.6000 652.0600 141.0800 ;
        RECT 605.4600 173.2400 607.0600 173.7200 ;
        RECT 605.4600 178.6800 607.0600 179.1600 ;
        RECT 605.4600 156.9200 607.0600 157.4000 ;
        RECT 605.4600 162.3600 607.0600 162.8400 ;
        RECT 605.4600 167.8000 607.0600 168.2800 ;
        RECT 605.4600 146.0400 607.0600 146.5200 ;
        RECT 605.4600 151.4800 607.0600 151.9600 ;
        RECT 605.4600 129.7200 607.0600 130.2000 ;
        RECT 605.4600 135.1600 607.0600 135.6400 ;
        RECT 605.4600 140.6000 607.0600 141.0800 ;
        RECT 662.0000 118.8400 665.0000 119.3200 ;
        RECT 662.0000 124.2800 665.0000 124.7600 ;
        RECT 650.4600 118.8400 652.0600 119.3200 ;
        RECT 650.4600 124.2800 652.0600 124.7600 ;
        RECT 662.0000 102.5200 665.0000 103.0000 ;
        RECT 662.0000 107.9600 665.0000 108.4400 ;
        RECT 662.0000 113.4000 665.0000 113.8800 ;
        RECT 650.4600 102.5200 652.0600 103.0000 ;
        RECT 650.4600 107.9600 652.0600 108.4400 ;
        RECT 650.4600 113.4000 652.0600 113.8800 ;
        RECT 662.0000 91.6400 665.0000 92.1200 ;
        RECT 662.0000 97.0800 665.0000 97.5600 ;
        RECT 650.4600 91.6400 652.0600 92.1200 ;
        RECT 650.4600 97.0800 652.0600 97.5600 ;
        RECT 662.0000 86.2000 665.0000 86.6800 ;
        RECT 650.4600 86.2000 652.0600 86.6800 ;
        RECT 605.4600 118.8400 607.0600 119.3200 ;
        RECT 605.4600 124.2800 607.0600 124.7600 ;
        RECT 605.4600 102.5200 607.0600 103.0000 ;
        RECT 605.4600 107.9600 607.0600 108.4400 ;
        RECT 605.4600 113.4000 607.0600 113.8800 ;
        RECT 605.4600 91.6400 607.0600 92.1200 ;
        RECT 605.4600 97.0800 607.0600 97.5600 ;
        RECT 605.4600 86.2000 607.0600 86.6800 ;
        RECT 560.4600 173.2400 562.0600 173.7200 ;
        RECT 560.4600 178.6800 562.0600 179.1600 ;
        RECT 560.4600 156.9200 562.0600 157.4000 ;
        RECT 560.4600 162.3600 562.0600 162.8400 ;
        RECT 560.4600 167.8000 562.0600 168.2800 ;
        RECT 515.4600 173.2400 517.0600 173.7200 ;
        RECT 515.4600 178.6800 517.0600 179.1600 ;
        RECT 515.4600 156.9200 517.0600 157.4000 ;
        RECT 515.4600 162.3600 517.0600 162.8400 ;
        RECT 515.4600 167.8000 517.0600 168.2800 ;
        RECT 560.4600 146.0400 562.0600 146.5200 ;
        RECT 560.4600 151.4800 562.0600 151.9600 ;
        RECT 560.4600 129.7200 562.0600 130.2000 ;
        RECT 560.4600 135.1600 562.0600 135.6400 ;
        RECT 560.4600 140.6000 562.0600 141.0800 ;
        RECT 515.4600 146.0400 517.0600 146.5200 ;
        RECT 515.4600 151.4800 517.0600 151.9600 ;
        RECT 515.4600 129.7200 517.0600 130.2000 ;
        RECT 515.4600 135.1600 517.0600 135.6400 ;
        RECT 515.4600 140.6000 517.0600 141.0800 ;
        RECT 465.9000 173.2400 468.9000 173.7200 ;
        RECT 465.9000 178.6800 468.9000 179.1600 ;
        RECT 465.9000 162.3600 468.9000 162.8400 ;
        RECT 465.9000 156.9200 468.9000 157.4000 ;
        RECT 465.9000 167.8000 468.9000 168.2800 ;
        RECT 465.9000 146.0400 468.9000 146.5200 ;
        RECT 465.9000 151.4800 468.9000 151.9600 ;
        RECT 465.9000 135.1600 468.9000 135.6400 ;
        RECT 465.9000 129.7200 468.9000 130.2000 ;
        RECT 465.9000 140.6000 468.9000 141.0800 ;
        RECT 560.4600 118.8400 562.0600 119.3200 ;
        RECT 560.4600 124.2800 562.0600 124.7600 ;
        RECT 560.4600 102.5200 562.0600 103.0000 ;
        RECT 560.4600 107.9600 562.0600 108.4400 ;
        RECT 560.4600 113.4000 562.0600 113.8800 ;
        RECT 515.4600 118.8400 517.0600 119.3200 ;
        RECT 515.4600 124.2800 517.0600 124.7600 ;
        RECT 515.4600 102.5200 517.0600 103.0000 ;
        RECT 515.4600 107.9600 517.0600 108.4400 ;
        RECT 515.4600 113.4000 517.0600 113.8800 ;
        RECT 560.4600 97.0800 562.0600 97.5600 ;
        RECT 560.4600 91.6400 562.0600 92.1200 ;
        RECT 560.4600 86.2000 562.0600 86.6800 ;
        RECT 515.4600 97.0800 517.0600 97.5600 ;
        RECT 515.4600 91.6400 517.0600 92.1200 ;
        RECT 515.4600 86.2000 517.0600 86.6800 ;
        RECT 465.9000 118.8400 468.9000 119.3200 ;
        RECT 465.9000 124.2800 468.9000 124.7600 ;
        RECT 465.9000 107.9600 468.9000 108.4400 ;
        RECT 465.9000 102.5200 468.9000 103.0000 ;
        RECT 465.9000 113.4000 468.9000 113.8800 ;
        RECT 465.9000 91.6400 468.9000 92.1200 ;
        RECT 465.9000 97.0800 468.9000 97.5600 ;
        RECT 465.9000 86.2000 468.9000 86.6800 ;
        RECT 465.9000 284.3900 665.0000 287.3900 ;
        RECT 465.9000 79.2900 665.0000 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 465.9000 37.6700 467.9000 58.6000 ;
        RECT 663.0000 37.6700 665.0000 58.6000 ;
      LAYER met3 ;
        RECT 663.0000 54.1000 665.0000 54.5800 ;
        RECT 465.9000 54.1000 467.9000 54.5800 ;
        RECT 663.0000 43.2200 665.0000 43.7000 ;
        RECT 465.9000 43.2200 467.9000 43.7000 ;
        RECT 663.0000 48.6600 665.0000 49.1400 ;
        RECT 465.9000 48.6600 467.9000 49.1400 ;
        RECT 465.9000 56.6000 665.0000 58.6000 ;
        RECT 465.9000 37.6700 665.0000 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 2605.3300 652.0600 2813.4300 ;
        RECT 605.4600 2605.3300 607.0600 2813.4300 ;
        RECT 560.4600 2605.3300 562.0600 2813.4300 ;
        RECT 515.4600 2605.3300 517.0600 2813.4300 ;
        RECT 662.0000 2605.3300 665.0000 2813.4300 ;
        RECT 465.9000 2605.3300 468.9000 2813.4300 ;
      LAYER met3 ;
        RECT 662.0000 2808.0800 665.0000 2808.5600 ;
        RECT 650.4600 2808.0800 652.0600 2808.5600 ;
        RECT 662.0000 2797.2000 665.0000 2797.6800 ;
        RECT 662.0000 2802.6400 665.0000 2803.1200 ;
        RECT 650.4600 2797.2000 652.0600 2797.6800 ;
        RECT 650.4600 2802.6400 652.0600 2803.1200 ;
        RECT 662.0000 2780.8800 665.0000 2781.3600 ;
        RECT 662.0000 2786.3200 665.0000 2786.8000 ;
        RECT 650.4600 2780.8800 652.0600 2781.3600 ;
        RECT 650.4600 2786.3200 652.0600 2786.8000 ;
        RECT 662.0000 2770.0000 665.0000 2770.4800 ;
        RECT 662.0000 2775.4400 665.0000 2775.9200 ;
        RECT 650.4600 2770.0000 652.0600 2770.4800 ;
        RECT 650.4600 2775.4400 652.0600 2775.9200 ;
        RECT 662.0000 2791.7600 665.0000 2792.2400 ;
        RECT 650.4600 2791.7600 652.0600 2792.2400 ;
        RECT 605.4600 2797.2000 607.0600 2797.6800 ;
        RECT 605.4600 2802.6400 607.0600 2803.1200 ;
        RECT 605.4600 2808.0800 607.0600 2808.5600 ;
        RECT 605.4600 2780.8800 607.0600 2781.3600 ;
        RECT 605.4600 2786.3200 607.0600 2786.8000 ;
        RECT 605.4600 2775.4400 607.0600 2775.9200 ;
        RECT 605.4600 2770.0000 607.0600 2770.4800 ;
        RECT 605.4600 2791.7600 607.0600 2792.2400 ;
        RECT 662.0000 2753.6800 665.0000 2754.1600 ;
        RECT 662.0000 2759.1200 665.0000 2759.6000 ;
        RECT 650.4600 2753.6800 652.0600 2754.1600 ;
        RECT 650.4600 2759.1200 652.0600 2759.6000 ;
        RECT 662.0000 2737.3600 665.0000 2737.8400 ;
        RECT 662.0000 2742.8000 665.0000 2743.2800 ;
        RECT 662.0000 2748.2400 665.0000 2748.7200 ;
        RECT 650.4600 2737.3600 652.0600 2737.8400 ;
        RECT 650.4600 2742.8000 652.0600 2743.2800 ;
        RECT 650.4600 2748.2400 652.0600 2748.7200 ;
        RECT 662.0000 2726.4800 665.0000 2726.9600 ;
        RECT 662.0000 2731.9200 665.0000 2732.4000 ;
        RECT 650.4600 2726.4800 652.0600 2726.9600 ;
        RECT 650.4600 2731.9200 652.0600 2732.4000 ;
        RECT 662.0000 2710.1600 665.0000 2710.6400 ;
        RECT 662.0000 2715.6000 665.0000 2716.0800 ;
        RECT 662.0000 2721.0400 665.0000 2721.5200 ;
        RECT 650.4600 2710.1600 652.0600 2710.6400 ;
        RECT 650.4600 2715.6000 652.0600 2716.0800 ;
        RECT 650.4600 2721.0400 652.0600 2721.5200 ;
        RECT 605.4600 2753.6800 607.0600 2754.1600 ;
        RECT 605.4600 2759.1200 607.0600 2759.6000 ;
        RECT 605.4600 2737.3600 607.0600 2737.8400 ;
        RECT 605.4600 2742.8000 607.0600 2743.2800 ;
        RECT 605.4600 2748.2400 607.0600 2748.7200 ;
        RECT 605.4600 2726.4800 607.0600 2726.9600 ;
        RECT 605.4600 2731.9200 607.0600 2732.4000 ;
        RECT 605.4600 2710.1600 607.0600 2710.6400 ;
        RECT 605.4600 2715.6000 607.0600 2716.0800 ;
        RECT 605.4600 2721.0400 607.0600 2721.5200 ;
        RECT 662.0000 2764.5600 665.0000 2765.0400 ;
        RECT 605.4600 2764.5600 607.0600 2765.0400 ;
        RECT 650.4600 2764.5600 652.0600 2765.0400 ;
        RECT 560.4600 2797.2000 562.0600 2797.6800 ;
        RECT 560.4600 2802.6400 562.0600 2803.1200 ;
        RECT 560.4600 2808.0800 562.0600 2808.5600 ;
        RECT 515.4600 2797.2000 517.0600 2797.6800 ;
        RECT 515.4600 2802.6400 517.0600 2803.1200 ;
        RECT 515.4600 2808.0800 517.0600 2808.5600 ;
        RECT 560.4600 2780.8800 562.0600 2781.3600 ;
        RECT 560.4600 2786.3200 562.0600 2786.8000 ;
        RECT 560.4600 2770.0000 562.0600 2770.4800 ;
        RECT 560.4600 2775.4400 562.0600 2775.9200 ;
        RECT 515.4600 2780.8800 517.0600 2781.3600 ;
        RECT 515.4600 2786.3200 517.0600 2786.8000 ;
        RECT 515.4600 2770.0000 517.0600 2770.4800 ;
        RECT 515.4600 2775.4400 517.0600 2775.9200 ;
        RECT 515.4600 2791.7600 517.0600 2792.2400 ;
        RECT 560.4600 2791.7600 562.0600 2792.2400 ;
        RECT 465.9000 2808.0800 468.9000 2808.5600 ;
        RECT 465.9000 2802.6400 468.9000 2803.1200 ;
        RECT 465.9000 2797.2000 468.9000 2797.6800 ;
        RECT 465.9000 2786.3200 468.9000 2786.8000 ;
        RECT 465.9000 2780.8800 468.9000 2781.3600 ;
        RECT 465.9000 2775.4400 468.9000 2775.9200 ;
        RECT 465.9000 2770.0000 468.9000 2770.4800 ;
        RECT 465.9000 2791.7600 468.9000 2792.2400 ;
        RECT 560.4600 2753.6800 562.0600 2754.1600 ;
        RECT 560.4600 2759.1200 562.0600 2759.6000 ;
        RECT 560.4600 2737.3600 562.0600 2737.8400 ;
        RECT 560.4600 2742.8000 562.0600 2743.2800 ;
        RECT 560.4600 2748.2400 562.0600 2748.7200 ;
        RECT 515.4600 2753.6800 517.0600 2754.1600 ;
        RECT 515.4600 2759.1200 517.0600 2759.6000 ;
        RECT 515.4600 2737.3600 517.0600 2737.8400 ;
        RECT 515.4600 2742.8000 517.0600 2743.2800 ;
        RECT 515.4600 2748.2400 517.0600 2748.7200 ;
        RECT 560.4600 2726.4800 562.0600 2726.9600 ;
        RECT 560.4600 2731.9200 562.0600 2732.4000 ;
        RECT 560.4600 2710.1600 562.0600 2710.6400 ;
        RECT 560.4600 2715.6000 562.0600 2716.0800 ;
        RECT 560.4600 2721.0400 562.0600 2721.5200 ;
        RECT 515.4600 2726.4800 517.0600 2726.9600 ;
        RECT 515.4600 2731.9200 517.0600 2732.4000 ;
        RECT 515.4600 2710.1600 517.0600 2710.6400 ;
        RECT 515.4600 2715.6000 517.0600 2716.0800 ;
        RECT 515.4600 2721.0400 517.0600 2721.5200 ;
        RECT 465.9000 2753.6800 468.9000 2754.1600 ;
        RECT 465.9000 2759.1200 468.9000 2759.6000 ;
        RECT 465.9000 2742.8000 468.9000 2743.2800 ;
        RECT 465.9000 2737.3600 468.9000 2737.8400 ;
        RECT 465.9000 2748.2400 468.9000 2748.7200 ;
        RECT 465.9000 2726.4800 468.9000 2726.9600 ;
        RECT 465.9000 2731.9200 468.9000 2732.4000 ;
        RECT 465.9000 2715.6000 468.9000 2716.0800 ;
        RECT 465.9000 2710.1600 468.9000 2710.6400 ;
        RECT 465.9000 2721.0400 468.9000 2721.5200 ;
        RECT 465.9000 2764.5600 468.9000 2765.0400 ;
        RECT 515.4600 2764.5600 517.0600 2765.0400 ;
        RECT 560.4600 2764.5600 562.0600 2765.0400 ;
        RECT 662.0000 2699.2800 665.0000 2699.7600 ;
        RECT 662.0000 2704.7200 665.0000 2705.2000 ;
        RECT 650.4600 2699.2800 652.0600 2699.7600 ;
        RECT 650.4600 2704.7200 652.0600 2705.2000 ;
        RECT 662.0000 2682.9600 665.0000 2683.4400 ;
        RECT 662.0000 2688.4000 665.0000 2688.8800 ;
        RECT 662.0000 2693.8400 665.0000 2694.3200 ;
        RECT 650.4600 2682.9600 652.0600 2683.4400 ;
        RECT 650.4600 2688.4000 652.0600 2688.8800 ;
        RECT 650.4600 2693.8400 652.0600 2694.3200 ;
        RECT 662.0000 2672.0800 665.0000 2672.5600 ;
        RECT 662.0000 2677.5200 665.0000 2678.0000 ;
        RECT 650.4600 2672.0800 652.0600 2672.5600 ;
        RECT 650.4600 2677.5200 652.0600 2678.0000 ;
        RECT 662.0000 2655.7600 665.0000 2656.2400 ;
        RECT 662.0000 2661.2000 665.0000 2661.6800 ;
        RECT 662.0000 2666.6400 665.0000 2667.1200 ;
        RECT 650.4600 2655.7600 652.0600 2656.2400 ;
        RECT 650.4600 2661.2000 652.0600 2661.6800 ;
        RECT 650.4600 2666.6400 652.0600 2667.1200 ;
        RECT 605.4600 2699.2800 607.0600 2699.7600 ;
        RECT 605.4600 2704.7200 607.0600 2705.2000 ;
        RECT 605.4600 2682.9600 607.0600 2683.4400 ;
        RECT 605.4600 2688.4000 607.0600 2688.8800 ;
        RECT 605.4600 2693.8400 607.0600 2694.3200 ;
        RECT 605.4600 2672.0800 607.0600 2672.5600 ;
        RECT 605.4600 2677.5200 607.0600 2678.0000 ;
        RECT 605.4600 2655.7600 607.0600 2656.2400 ;
        RECT 605.4600 2661.2000 607.0600 2661.6800 ;
        RECT 605.4600 2666.6400 607.0600 2667.1200 ;
        RECT 662.0000 2644.8800 665.0000 2645.3600 ;
        RECT 662.0000 2650.3200 665.0000 2650.8000 ;
        RECT 650.4600 2644.8800 652.0600 2645.3600 ;
        RECT 650.4600 2650.3200 652.0600 2650.8000 ;
        RECT 662.0000 2628.5600 665.0000 2629.0400 ;
        RECT 662.0000 2634.0000 665.0000 2634.4800 ;
        RECT 662.0000 2639.4400 665.0000 2639.9200 ;
        RECT 650.4600 2628.5600 652.0600 2629.0400 ;
        RECT 650.4600 2634.0000 652.0600 2634.4800 ;
        RECT 650.4600 2639.4400 652.0600 2639.9200 ;
        RECT 662.0000 2617.6800 665.0000 2618.1600 ;
        RECT 662.0000 2623.1200 665.0000 2623.6000 ;
        RECT 650.4600 2617.6800 652.0600 2618.1600 ;
        RECT 650.4600 2623.1200 652.0600 2623.6000 ;
        RECT 662.0000 2612.2400 665.0000 2612.7200 ;
        RECT 650.4600 2612.2400 652.0600 2612.7200 ;
        RECT 605.4600 2644.8800 607.0600 2645.3600 ;
        RECT 605.4600 2650.3200 607.0600 2650.8000 ;
        RECT 605.4600 2628.5600 607.0600 2629.0400 ;
        RECT 605.4600 2634.0000 607.0600 2634.4800 ;
        RECT 605.4600 2639.4400 607.0600 2639.9200 ;
        RECT 605.4600 2617.6800 607.0600 2618.1600 ;
        RECT 605.4600 2623.1200 607.0600 2623.6000 ;
        RECT 605.4600 2612.2400 607.0600 2612.7200 ;
        RECT 560.4600 2699.2800 562.0600 2699.7600 ;
        RECT 560.4600 2704.7200 562.0600 2705.2000 ;
        RECT 560.4600 2682.9600 562.0600 2683.4400 ;
        RECT 560.4600 2688.4000 562.0600 2688.8800 ;
        RECT 560.4600 2693.8400 562.0600 2694.3200 ;
        RECT 515.4600 2699.2800 517.0600 2699.7600 ;
        RECT 515.4600 2704.7200 517.0600 2705.2000 ;
        RECT 515.4600 2682.9600 517.0600 2683.4400 ;
        RECT 515.4600 2688.4000 517.0600 2688.8800 ;
        RECT 515.4600 2693.8400 517.0600 2694.3200 ;
        RECT 560.4600 2672.0800 562.0600 2672.5600 ;
        RECT 560.4600 2677.5200 562.0600 2678.0000 ;
        RECT 560.4600 2655.7600 562.0600 2656.2400 ;
        RECT 560.4600 2661.2000 562.0600 2661.6800 ;
        RECT 560.4600 2666.6400 562.0600 2667.1200 ;
        RECT 515.4600 2672.0800 517.0600 2672.5600 ;
        RECT 515.4600 2677.5200 517.0600 2678.0000 ;
        RECT 515.4600 2655.7600 517.0600 2656.2400 ;
        RECT 515.4600 2661.2000 517.0600 2661.6800 ;
        RECT 515.4600 2666.6400 517.0600 2667.1200 ;
        RECT 465.9000 2699.2800 468.9000 2699.7600 ;
        RECT 465.9000 2704.7200 468.9000 2705.2000 ;
        RECT 465.9000 2688.4000 468.9000 2688.8800 ;
        RECT 465.9000 2682.9600 468.9000 2683.4400 ;
        RECT 465.9000 2693.8400 468.9000 2694.3200 ;
        RECT 465.9000 2672.0800 468.9000 2672.5600 ;
        RECT 465.9000 2677.5200 468.9000 2678.0000 ;
        RECT 465.9000 2661.2000 468.9000 2661.6800 ;
        RECT 465.9000 2655.7600 468.9000 2656.2400 ;
        RECT 465.9000 2666.6400 468.9000 2667.1200 ;
        RECT 560.4600 2644.8800 562.0600 2645.3600 ;
        RECT 560.4600 2650.3200 562.0600 2650.8000 ;
        RECT 560.4600 2628.5600 562.0600 2629.0400 ;
        RECT 560.4600 2634.0000 562.0600 2634.4800 ;
        RECT 560.4600 2639.4400 562.0600 2639.9200 ;
        RECT 515.4600 2644.8800 517.0600 2645.3600 ;
        RECT 515.4600 2650.3200 517.0600 2650.8000 ;
        RECT 515.4600 2628.5600 517.0600 2629.0400 ;
        RECT 515.4600 2634.0000 517.0600 2634.4800 ;
        RECT 515.4600 2639.4400 517.0600 2639.9200 ;
        RECT 560.4600 2623.1200 562.0600 2623.6000 ;
        RECT 560.4600 2617.6800 562.0600 2618.1600 ;
        RECT 560.4600 2612.2400 562.0600 2612.7200 ;
        RECT 515.4600 2623.1200 517.0600 2623.6000 ;
        RECT 515.4600 2617.6800 517.0600 2618.1600 ;
        RECT 515.4600 2612.2400 517.0600 2612.7200 ;
        RECT 465.9000 2644.8800 468.9000 2645.3600 ;
        RECT 465.9000 2650.3200 468.9000 2650.8000 ;
        RECT 465.9000 2634.0000 468.9000 2634.4800 ;
        RECT 465.9000 2628.5600 468.9000 2629.0400 ;
        RECT 465.9000 2639.4400 468.9000 2639.9200 ;
        RECT 465.9000 2617.6800 468.9000 2618.1600 ;
        RECT 465.9000 2623.1200 468.9000 2623.6000 ;
        RECT 465.9000 2612.2400 468.9000 2612.7200 ;
        RECT 465.9000 2810.4300 665.0000 2813.4300 ;
        RECT 465.9000 2605.3300 665.0000 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 2375.6900 652.0600 2583.7900 ;
        RECT 605.4600 2375.6900 607.0600 2583.7900 ;
        RECT 560.4600 2375.6900 562.0600 2583.7900 ;
        RECT 515.4600 2375.6900 517.0600 2583.7900 ;
        RECT 662.0000 2375.6900 665.0000 2583.7900 ;
        RECT 465.9000 2375.6900 468.9000 2583.7900 ;
      LAYER met3 ;
        RECT 662.0000 2578.4400 665.0000 2578.9200 ;
        RECT 650.4600 2578.4400 652.0600 2578.9200 ;
        RECT 662.0000 2567.5600 665.0000 2568.0400 ;
        RECT 662.0000 2573.0000 665.0000 2573.4800 ;
        RECT 650.4600 2567.5600 652.0600 2568.0400 ;
        RECT 650.4600 2573.0000 652.0600 2573.4800 ;
        RECT 662.0000 2551.2400 665.0000 2551.7200 ;
        RECT 662.0000 2556.6800 665.0000 2557.1600 ;
        RECT 650.4600 2551.2400 652.0600 2551.7200 ;
        RECT 650.4600 2556.6800 652.0600 2557.1600 ;
        RECT 662.0000 2540.3600 665.0000 2540.8400 ;
        RECT 662.0000 2545.8000 665.0000 2546.2800 ;
        RECT 650.4600 2540.3600 652.0600 2540.8400 ;
        RECT 650.4600 2545.8000 652.0600 2546.2800 ;
        RECT 662.0000 2562.1200 665.0000 2562.6000 ;
        RECT 650.4600 2562.1200 652.0600 2562.6000 ;
        RECT 605.4600 2567.5600 607.0600 2568.0400 ;
        RECT 605.4600 2573.0000 607.0600 2573.4800 ;
        RECT 605.4600 2578.4400 607.0600 2578.9200 ;
        RECT 605.4600 2551.2400 607.0600 2551.7200 ;
        RECT 605.4600 2556.6800 607.0600 2557.1600 ;
        RECT 605.4600 2545.8000 607.0600 2546.2800 ;
        RECT 605.4600 2540.3600 607.0600 2540.8400 ;
        RECT 605.4600 2562.1200 607.0600 2562.6000 ;
        RECT 662.0000 2524.0400 665.0000 2524.5200 ;
        RECT 662.0000 2529.4800 665.0000 2529.9600 ;
        RECT 650.4600 2524.0400 652.0600 2524.5200 ;
        RECT 650.4600 2529.4800 652.0600 2529.9600 ;
        RECT 662.0000 2507.7200 665.0000 2508.2000 ;
        RECT 662.0000 2513.1600 665.0000 2513.6400 ;
        RECT 662.0000 2518.6000 665.0000 2519.0800 ;
        RECT 650.4600 2507.7200 652.0600 2508.2000 ;
        RECT 650.4600 2513.1600 652.0600 2513.6400 ;
        RECT 650.4600 2518.6000 652.0600 2519.0800 ;
        RECT 662.0000 2496.8400 665.0000 2497.3200 ;
        RECT 662.0000 2502.2800 665.0000 2502.7600 ;
        RECT 650.4600 2496.8400 652.0600 2497.3200 ;
        RECT 650.4600 2502.2800 652.0600 2502.7600 ;
        RECT 662.0000 2480.5200 665.0000 2481.0000 ;
        RECT 662.0000 2485.9600 665.0000 2486.4400 ;
        RECT 662.0000 2491.4000 665.0000 2491.8800 ;
        RECT 650.4600 2480.5200 652.0600 2481.0000 ;
        RECT 650.4600 2485.9600 652.0600 2486.4400 ;
        RECT 650.4600 2491.4000 652.0600 2491.8800 ;
        RECT 605.4600 2524.0400 607.0600 2524.5200 ;
        RECT 605.4600 2529.4800 607.0600 2529.9600 ;
        RECT 605.4600 2507.7200 607.0600 2508.2000 ;
        RECT 605.4600 2513.1600 607.0600 2513.6400 ;
        RECT 605.4600 2518.6000 607.0600 2519.0800 ;
        RECT 605.4600 2496.8400 607.0600 2497.3200 ;
        RECT 605.4600 2502.2800 607.0600 2502.7600 ;
        RECT 605.4600 2480.5200 607.0600 2481.0000 ;
        RECT 605.4600 2485.9600 607.0600 2486.4400 ;
        RECT 605.4600 2491.4000 607.0600 2491.8800 ;
        RECT 662.0000 2534.9200 665.0000 2535.4000 ;
        RECT 605.4600 2534.9200 607.0600 2535.4000 ;
        RECT 650.4600 2534.9200 652.0600 2535.4000 ;
        RECT 560.4600 2567.5600 562.0600 2568.0400 ;
        RECT 560.4600 2573.0000 562.0600 2573.4800 ;
        RECT 560.4600 2578.4400 562.0600 2578.9200 ;
        RECT 515.4600 2567.5600 517.0600 2568.0400 ;
        RECT 515.4600 2573.0000 517.0600 2573.4800 ;
        RECT 515.4600 2578.4400 517.0600 2578.9200 ;
        RECT 560.4600 2551.2400 562.0600 2551.7200 ;
        RECT 560.4600 2556.6800 562.0600 2557.1600 ;
        RECT 560.4600 2540.3600 562.0600 2540.8400 ;
        RECT 560.4600 2545.8000 562.0600 2546.2800 ;
        RECT 515.4600 2551.2400 517.0600 2551.7200 ;
        RECT 515.4600 2556.6800 517.0600 2557.1600 ;
        RECT 515.4600 2540.3600 517.0600 2540.8400 ;
        RECT 515.4600 2545.8000 517.0600 2546.2800 ;
        RECT 515.4600 2562.1200 517.0600 2562.6000 ;
        RECT 560.4600 2562.1200 562.0600 2562.6000 ;
        RECT 465.9000 2578.4400 468.9000 2578.9200 ;
        RECT 465.9000 2573.0000 468.9000 2573.4800 ;
        RECT 465.9000 2567.5600 468.9000 2568.0400 ;
        RECT 465.9000 2556.6800 468.9000 2557.1600 ;
        RECT 465.9000 2551.2400 468.9000 2551.7200 ;
        RECT 465.9000 2545.8000 468.9000 2546.2800 ;
        RECT 465.9000 2540.3600 468.9000 2540.8400 ;
        RECT 465.9000 2562.1200 468.9000 2562.6000 ;
        RECT 560.4600 2524.0400 562.0600 2524.5200 ;
        RECT 560.4600 2529.4800 562.0600 2529.9600 ;
        RECT 560.4600 2507.7200 562.0600 2508.2000 ;
        RECT 560.4600 2513.1600 562.0600 2513.6400 ;
        RECT 560.4600 2518.6000 562.0600 2519.0800 ;
        RECT 515.4600 2524.0400 517.0600 2524.5200 ;
        RECT 515.4600 2529.4800 517.0600 2529.9600 ;
        RECT 515.4600 2507.7200 517.0600 2508.2000 ;
        RECT 515.4600 2513.1600 517.0600 2513.6400 ;
        RECT 515.4600 2518.6000 517.0600 2519.0800 ;
        RECT 560.4600 2496.8400 562.0600 2497.3200 ;
        RECT 560.4600 2502.2800 562.0600 2502.7600 ;
        RECT 560.4600 2480.5200 562.0600 2481.0000 ;
        RECT 560.4600 2485.9600 562.0600 2486.4400 ;
        RECT 560.4600 2491.4000 562.0600 2491.8800 ;
        RECT 515.4600 2496.8400 517.0600 2497.3200 ;
        RECT 515.4600 2502.2800 517.0600 2502.7600 ;
        RECT 515.4600 2480.5200 517.0600 2481.0000 ;
        RECT 515.4600 2485.9600 517.0600 2486.4400 ;
        RECT 515.4600 2491.4000 517.0600 2491.8800 ;
        RECT 465.9000 2524.0400 468.9000 2524.5200 ;
        RECT 465.9000 2529.4800 468.9000 2529.9600 ;
        RECT 465.9000 2513.1600 468.9000 2513.6400 ;
        RECT 465.9000 2507.7200 468.9000 2508.2000 ;
        RECT 465.9000 2518.6000 468.9000 2519.0800 ;
        RECT 465.9000 2496.8400 468.9000 2497.3200 ;
        RECT 465.9000 2502.2800 468.9000 2502.7600 ;
        RECT 465.9000 2485.9600 468.9000 2486.4400 ;
        RECT 465.9000 2480.5200 468.9000 2481.0000 ;
        RECT 465.9000 2491.4000 468.9000 2491.8800 ;
        RECT 465.9000 2534.9200 468.9000 2535.4000 ;
        RECT 515.4600 2534.9200 517.0600 2535.4000 ;
        RECT 560.4600 2534.9200 562.0600 2535.4000 ;
        RECT 662.0000 2469.6400 665.0000 2470.1200 ;
        RECT 662.0000 2475.0800 665.0000 2475.5600 ;
        RECT 650.4600 2469.6400 652.0600 2470.1200 ;
        RECT 650.4600 2475.0800 652.0600 2475.5600 ;
        RECT 662.0000 2453.3200 665.0000 2453.8000 ;
        RECT 662.0000 2458.7600 665.0000 2459.2400 ;
        RECT 662.0000 2464.2000 665.0000 2464.6800 ;
        RECT 650.4600 2453.3200 652.0600 2453.8000 ;
        RECT 650.4600 2458.7600 652.0600 2459.2400 ;
        RECT 650.4600 2464.2000 652.0600 2464.6800 ;
        RECT 662.0000 2442.4400 665.0000 2442.9200 ;
        RECT 662.0000 2447.8800 665.0000 2448.3600 ;
        RECT 650.4600 2442.4400 652.0600 2442.9200 ;
        RECT 650.4600 2447.8800 652.0600 2448.3600 ;
        RECT 662.0000 2426.1200 665.0000 2426.6000 ;
        RECT 662.0000 2431.5600 665.0000 2432.0400 ;
        RECT 662.0000 2437.0000 665.0000 2437.4800 ;
        RECT 650.4600 2426.1200 652.0600 2426.6000 ;
        RECT 650.4600 2431.5600 652.0600 2432.0400 ;
        RECT 650.4600 2437.0000 652.0600 2437.4800 ;
        RECT 605.4600 2469.6400 607.0600 2470.1200 ;
        RECT 605.4600 2475.0800 607.0600 2475.5600 ;
        RECT 605.4600 2453.3200 607.0600 2453.8000 ;
        RECT 605.4600 2458.7600 607.0600 2459.2400 ;
        RECT 605.4600 2464.2000 607.0600 2464.6800 ;
        RECT 605.4600 2442.4400 607.0600 2442.9200 ;
        RECT 605.4600 2447.8800 607.0600 2448.3600 ;
        RECT 605.4600 2426.1200 607.0600 2426.6000 ;
        RECT 605.4600 2431.5600 607.0600 2432.0400 ;
        RECT 605.4600 2437.0000 607.0600 2437.4800 ;
        RECT 662.0000 2415.2400 665.0000 2415.7200 ;
        RECT 662.0000 2420.6800 665.0000 2421.1600 ;
        RECT 650.4600 2415.2400 652.0600 2415.7200 ;
        RECT 650.4600 2420.6800 652.0600 2421.1600 ;
        RECT 662.0000 2398.9200 665.0000 2399.4000 ;
        RECT 662.0000 2404.3600 665.0000 2404.8400 ;
        RECT 662.0000 2409.8000 665.0000 2410.2800 ;
        RECT 650.4600 2398.9200 652.0600 2399.4000 ;
        RECT 650.4600 2404.3600 652.0600 2404.8400 ;
        RECT 650.4600 2409.8000 652.0600 2410.2800 ;
        RECT 662.0000 2388.0400 665.0000 2388.5200 ;
        RECT 662.0000 2393.4800 665.0000 2393.9600 ;
        RECT 650.4600 2388.0400 652.0600 2388.5200 ;
        RECT 650.4600 2393.4800 652.0600 2393.9600 ;
        RECT 662.0000 2382.6000 665.0000 2383.0800 ;
        RECT 650.4600 2382.6000 652.0600 2383.0800 ;
        RECT 605.4600 2415.2400 607.0600 2415.7200 ;
        RECT 605.4600 2420.6800 607.0600 2421.1600 ;
        RECT 605.4600 2398.9200 607.0600 2399.4000 ;
        RECT 605.4600 2404.3600 607.0600 2404.8400 ;
        RECT 605.4600 2409.8000 607.0600 2410.2800 ;
        RECT 605.4600 2388.0400 607.0600 2388.5200 ;
        RECT 605.4600 2393.4800 607.0600 2393.9600 ;
        RECT 605.4600 2382.6000 607.0600 2383.0800 ;
        RECT 560.4600 2469.6400 562.0600 2470.1200 ;
        RECT 560.4600 2475.0800 562.0600 2475.5600 ;
        RECT 560.4600 2453.3200 562.0600 2453.8000 ;
        RECT 560.4600 2458.7600 562.0600 2459.2400 ;
        RECT 560.4600 2464.2000 562.0600 2464.6800 ;
        RECT 515.4600 2469.6400 517.0600 2470.1200 ;
        RECT 515.4600 2475.0800 517.0600 2475.5600 ;
        RECT 515.4600 2453.3200 517.0600 2453.8000 ;
        RECT 515.4600 2458.7600 517.0600 2459.2400 ;
        RECT 515.4600 2464.2000 517.0600 2464.6800 ;
        RECT 560.4600 2442.4400 562.0600 2442.9200 ;
        RECT 560.4600 2447.8800 562.0600 2448.3600 ;
        RECT 560.4600 2426.1200 562.0600 2426.6000 ;
        RECT 560.4600 2431.5600 562.0600 2432.0400 ;
        RECT 560.4600 2437.0000 562.0600 2437.4800 ;
        RECT 515.4600 2442.4400 517.0600 2442.9200 ;
        RECT 515.4600 2447.8800 517.0600 2448.3600 ;
        RECT 515.4600 2426.1200 517.0600 2426.6000 ;
        RECT 515.4600 2431.5600 517.0600 2432.0400 ;
        RECT 515.4600 2437.0000 517.0600 2437.4800 ;
        RECT 465.9000 2469.6400 468.9000 2470.1200 ;
        RECT 465.9000 2475.0800 468.9000 2475.5600 ;
        RECT 465.9000 2458.7600 468.9000 2459.2400 ;
        RECT 465.9000 2453.3200 468.9000 2453.8000 ;
        RECT 465.9000 2464.2000 468.9000 2464.6800 ;
        RECT 465.9000 2442.4400 468.9000 2442.9200 ;
        RECT 465.9000 2447.8800 468.9000 2448.3600 ;
        RECT 465.9000 2431.5600 468.9000 2432.0400 ;
        RECT 465.9000 2426.1200 468.9000 2426.6000 ;
        RECT 465.9000 2437.0000 468.9000 2437.4800 ;
        RECT 560.4600 2415.2400 562.0600 2415.7200 ;
        RECT 560.4600 2420.6800 562.0600 2421.1600 ;
        RECT 560.4600 2398.9200 562.0600 2399.4000 ;
        RECT 560.4600 2404.3600 562.0600 2404.8400 ;
        RECT 560.4600 2409.8000 562.0600 2410.2800 ;
        RECT 515.4600 2415.2400 517.0600 2415.7200 ;
        RECT 515.4600 2420.6800 517.0600 2421.1600 ;
        RECT 515.4600 2398.9200 517.0600 2399.4000 ;
        RECT 515.4600 2404.3600 517.0600 2404.8400 ;
        RECT 515.4600 2409.8000 517.0600 2410.2800 ;
        RECT 560.4600 2393.4800 562.0600 2393.9600 ;
        RECT 560.4600 2388.0400 562.0600 2388.5200 ;
        RECT 560.4600 2382.6000 562.0600 2383.0800 ;
        RECT 515.4600 2393.4800 517.0600 2393.9600 ;
        RECT 515.4600 2388.0400 517.0600 2388.5200 ;
        RECT 515.4600 2382.6000 517.0600 2383.0800 ;
        RECT 465.9000 2415.2400 468.9000 2415.7200 ;
        RECT 465.9000 2420.6800 468.9000 2421.1600 ;
        RECT 465.9000 2404.3600 468.9000 2404.8400 ;
        RECT 465.9000 2398.9200 468.9000 2399.4000 ;
        RECT 465.9000 2409.8000 468.9000 2410.2800 ;
        RECT 465.9000 2388.0400 468.9000 2388.5200 ;
        RECT 465.9000 2393.4800 468.9000 2393.9600 ;
        RECT 465.9000 2382.6000 468.9000 2383.0800 ;
        RECT 465.9000 2580.7900 665.0000 2583.7900 ;
        RECT 465.9000 2375.6900 665.0000 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 2146.0500 652.0600 2354.1500 ;
        RECT 605.4600 2146.0500 607.0600 2354.1500 ;
        RECT 560.4600 2146.0500 562.0600 2354.1500 ;
        RECT 515.4600 2146.0500 517.0600 2354.1500 ;
        RECT 662.0000 2146.0500 665.0000 2354.1500 ;
        RECT 465.9000 2146.0500 468.9000 2354.1500 ;
      LAYER met3 ;
        RECT 662.0000 2348.8000 665.0000 2349.2800 ;
        RECT 650.4600 2348.8000 652.0600 2349.2800 ;
        RECT 662.0000 2337.9200 665.0000 2338.4000 ;
        RECT 662.0000 2343.3600 665.0000 2343.8400 ;
        RECT 650.4600 2337.9200 652.0600 2338.4000 ;
        RECT 650.4600 2343.3600 652.0600 2343.8400 ;
        RECT 662.0000 2321.6000 665.0000 2322.0800 ;
        RECT 662.0000 2327.0400 665.0000 2327.5200 ;
        RECT 650.4600 2321.6000 652.0600 2322.0800 ;
        RECT 650.4600 2327.0400 652.0600 2327.5200 ;
        RECT 662.0000 2310.7200 665.0000 2311.2000 ;
        RECT 662.0000 2316.1600 665.0000 2316.6400 ;
        RECT 650.4600 2310.7200 652.0600 2311.2000 ;
        RECT 650.4600 2316.1600 652.0600 2316.6400 ;
        RECT 662.0000 2332.4800 665.0000 2332.9600 ;
        RECT 650.4600 2332.4800 652.0600 2332.9600 ;
        RECT 605.4600 2337.9200 607.0600 2338.4000 ;
        RECT 605.4600 2343.3600 607.0600 2343.8400 ;
        RECT 605.4600 2348.8000 607.0600 2349.2800 ;
        RECT 605.4600 2321.6000 607.0600 2322.0800 ;
        RECT 605.4600 2327.0400 607.0600 2327.5200 ;
        RECT 605.4600 2316.1600 607.0600 2316.6400 ;
        RECT 605.4600 2310.7200 607.0600 2311.2000 ;
        RECT 605.4600 2332.4800 607.0600 2332.9600 ;
        RECT 662.0000 2294.4000 665.0000 2294.8800 ;
        RECT 662.0000 2299.8400 665.0000 2300.3200 ;
        RECT 650.4600 2294.4000 652.0600 2294.8800 ;
        RECT 650.4600 2299.8400 652.0600 2300.3200 ;
        RECT 662.0000 2278.0800 665.0000 2278.5600 ;
        RECT 662.0000 2283.5200 665.0000 2284.0000 ;
        RECT 662.0000 2288.9600 665.0000 2289.4400 ;
        RECT 650.4600 2278.0800 652.0600 2278.5600 ;
        RECT 650.4600 2283.5200 652.0600 2284.0000 ;
        RECT 650.4600 2288.9600 652.0600 2289.4400 ;
        RECT 662.0000 2267.2000 665.0000 2267.6800 ;
        RECT 662.0000 2272.6400 665.0000 2273.1200 ;
        RECT 650.4600 2267.2000 652.0600 2267.6800 ;
        RECT 650.4600 2272.6400 652.0600 2273.1200 ;
        RECT 662.0000 2250.8800 665.0000 2251.3600 ;
        RECT 662.0000 2256.3200 665.0000 2256.8000 ;
        RECT 662.0000 2261.7600 665.0000 2262.2400 ;
        RECT 650.4600 2250.8800 652.0600 2251.3600 ;
        RECT 650.4600 2256.3200 652.0600 2256.8000 ;
        RECT 650.4600 2261.7600 652.0600 2262.2400 ;
        RECT 605.4600 2294.4000 607.0600 2294.8800 ;
        RECT 605.4600 2299.8400 607.0600 2300.3200 ;
        RECT 605.4600 2278.0800 607.0600 2278.5600 ;
        RECT 605.4600 2283.5200 607.0600 2284.0000 ;
        RECT 605.4600 2288.9600 607.0600 2289.4400 ;
        RECT 605.4600 2267.2000 607.0600 2267.6800 ;
        RECT 605.4600 2272.6400 607.0600 2273.1200 ;
        RECT 605.4600 2250.8800 607.0600 2251.3600 ;
        RECT 605.4600 2256.3200 607.0600 2256.8000 ;
        RECT 605.4600 2261.7600 607.0600 2262.2400 ;
        RECT 662.0000 2305.2800 665.0000 2305.7600 ;
        RECT 605.4600 2305.2800 607.0600 2305.7600 ;
        RECT 650.4600 2305.2800 652.0600 2305.7600 ;
        RECT 560.4600 2337.9200 562.0600 2338.4000 ;
        RECT 560.4600 2343.3600 562.0600 2343.8400 ;
        RECT 560.4600 2348.8000 562.0600 2349.2800 ;
        RECT 515.4600 2337.9200 517.0600 2338.4000 ;
        RECT 515.4600 2343.3600 517.0600 2343.8400 ;
        RECT 515.4600 2348.8000 517.0600 2349.2800 ;
        RECT 560.4600 2321.6000 562.0600 2322.0800 ;
        RECT 560.4600 2327.0400 562.0600 2327.5200 ;
        RECT 560.4600 2310.7200 562.0600 2311.2000 ;
        RECT 560.4600 2316.1600 562.0600 2316.6400 ;
        RECT 515.4600 2321.6000 517.0600 2322.0800 ;
        RECT 515.4600 2327.0400 517.0600 2327.5200 ;
        RECT 515.4600 2310.7200 517.0600 2311.2000 ;
        RECT 515.4600 2316.1600 517.0600 2316.6400 ;
        RECT 515.4600 2332.4800 517.0600 2332.9600 ;
        RECT 560.4600 2332.4800 562.0600 2332.9600 ;
        RECT 465.9000 2348.8000 468.9000 2349.2800 ;
        RECT 465.9000 2343.3600 468.9000 2343.8400 ;
        RECT 465.9000 2337.9200 468.9000 2338.4000 ;
        RECT 465.9000 2327.0400 468.9000 2327.5200 ;
        RECT 465.9000 2321.6000 468.9000 2322.0800 ;
        RECT 465.9000 2316.1600 468.9000 2316.6400 ;
        RECT 465.9000 2310.7200 468.9000 2311.2000 ;
        RECT 465.9000 2332.4800 468.9000 2332.9600 ;
        RECT 560.4600 2294.4000 562.0600 2294.8800 ;
        RECT 560.4600 2299.8400 562.0600 2300.3200 ;
        RECT 560.4600 2278.0800 562.0600 2278.5600 ;
        RECT 560.4600 2283.5200 562.0600 2284.0000 ;
        RECT 560.4600 2288.9600 562.0600 2289.4400 ;
        RECT 515.4600 2294.4000 517.0600 2294.8800 ;
        RECT 515.4600 2299.8400 517.0600 2300.3200 ;
        RECT 515.4600 2278.0800 517.0600 2278.5600 ;
        RECT 515.4600 2283.5200 517.0600 2284.0000 ;
        RECT 515.4600 2288.9600 517.0600 2289.4400 ;
        RECT 560.4600 2267.2000 562.0600 2267.6800 ;
        RECT 560.4600 2272.6400 562.0600 2273.1200 ;
        RECT 560.4600 2250.8800 562.0600 2251.3600 ;
        RECT 560.4600 2256.3200 562.0600 2256.8000 ;
        RECT 560.4600 2261.7600 562.0600 2262.2400 ;
        RECT 515.4600 2267.2000 517.0600 2267.6800 ;
        RECT 515.4600 2272.6400 517.0600 2273.1200 ;
        RECT 515.4600 2250.8800 517.0600 2251.3600 ;
        RECT 515.4600 2256.3200 517.0600 2256.8000 ;
        RECT 515.4600 2261.7600 517.0600 2262.2400 ;
        RECT 465.9000 2294.4000 468.9000 2294.8800 ;
        RECT 465.9000 2299.8400 468.9000 2300.3200 ;
        RECT 465.9000 2283.5200 468.9000 2284.0000 ;
        RECT 465.9000 2278.0800 468.9000 2278.5600 ;
        RECT 465.9000 2288.9600 468.9000 2289.4400 ;
        RECT 465.9000 2267.2000 468.9000 2267.6800 ;
        RECT 465.9000 2272.6400 468.9000 2273.1200 ;
        RECT 465.9000 2256.3200 468.9000 2256.8000 ;
        RECT 465.9000 2250.8800 468.9000 2251.3600 ;
        RECT 465.9000 2261.7600 468.9000 2262.2400 ;
        RECT 465.9000 2305.2800 468.9000 2305.7600 ;
        RECT 515.4600 2305.2800 517.0600 2305.7600 ;
        RECT 560.4600 2305.2800 562.0600 2305.7600 ;
        RECT 662.0000 2240.0000 665.0000 2240.4800 ;
        RECT 662.0000 2245.4400 665.0000 2245.9200 ;
        RECT 650.4600 2240.0000 652.0600 2240.4800 ;
        RECT 650.4600 2245.4400 652.0600 2245.9200 ;
        RECT 662.0000 2223.6800 665.0000 2224.1600 ;
        RECT 662.0000 2229.1200 665.0000 2229.6000 ;
        RECT 662.0000 2234.5600 665.0000 2235.0400 ;
        RECT 650.4600 2223.6800 652.0600 2224.1600 ;
        RECT 650.4600 2229.1200 652.0600 2229.6000 ;
        RECT 650.4600 2234.5600 652.0600 2235.0400 ;
        RECT 662.0000 2212.8000 665.0000 2213.2800 ;
        RECT 662.0000 2218.2400 665.0000 2218.7200 ;
        RECT 650.4600 2212.8000 652.0600 2213.2800 ;
        RECT 650.4600 2218.2400 652.0600 2218.7200 ;
        RECT 662.0000 2196.4800 665.0000 2196.9600 ;
        RECT 662.0000 2201.9200 665.0000 2202.4000 ;
        RECT 662.0000 2207.3600 665.0000 2207.8400 ;
        RECT 650.4600 2196.4800 652.0600 2196.9600 ;
        RECT 650.4600 2201.9200 652.0600 2202.4000 ;
        RECT 650.4600 2207.3600 652.0600 2207.8400 ;
        RECT 605.4600 2240.0000 607.0600 2240.4800 ;
        RECT 605.4600 2245.4400 607.0600 2245.9200 ;
        RECT 605.4600 2223.6800 607.0600 2224.1600 ;
        RECT 605.4600 2229.1200 607.0600 2229.6000 ;
        RECT 605.4600 2234.5600 607.0600 2235.0400 ;
        RECT 605.4600 2212.8000 607.0600 2213.2800 ;
        RECT 605.4600 2218.2400 607.0600 2218.7200 ;
        RECT 605.4600 2196.4800 607.0600 2196.9600 ;
        RECT 605.4600 2201.9200 607.0600 2202.4000 ;
        RECT 605.4600 2207.3600 607.0600 2207.8400 ;
        RECT 662.0000 2185.6000 665.0000 2186.0800 ;
        RECT 662.0000 2191.0400 665.0000 2191.5200 ;
        RECT 650.4600 2185.6000 652.0600 2186.0800 ;
        RECT 650.4600 2191.0400 652.0600 2191.5200 ;
        RECT 662.0000 2169.2800 665.0000 2169.7600 ;
        RECT 662.0000 2174.7200 665.0000 2175.2000 ;
        RECT 662.0000 2180.1600 665.0000 2180.6400 ;
        RECT 650.4600 2169.2800 652.0600 2169.7600 ;
        RECT 650.4600 2174.7200 652.0600 2175.2000 ;
        RECT 650.4600 2180.1600 652.0600 2180.6400 ;
        RECT 662.0000 2158.4000 665.0000 2158.8800 ;
        RECT 662.0000 2163.8400 665.0000 2164.3200 ;
        RECT 650.4600 2158.4000 652.0600 2158.8800 ;
        RECT 650.4600 2163.8400 652.0600 2164.3200 ;
        RECT 662.0000 2152.9600 665.0000 2153.4400 ;
        RECT 650.4600 2152.9600 652.0600 2153.4400 ;
        RECT 605.4600 2185.6000 607.0600 2186.0800 ;
        RECT 605.4600 2191.0400 607.0600 2191.5200 ;
        RECT 605.4600 2169.2800 607.0600 2169.7600 ;
        RECT 605.4600 2174.7200 607.0600 2175.2000 ;
        RECT 605.4600 2180.1600 607.0600 2180.6400 ;
        RECT 605.4600 2158.4000 607.0600 2158.8800 ;
        RECT 605.4600 2163.8400 607.0600 2164.3200 ;
        RECT 605.4600 2152.9600 607.0600 2153.4400 ;
        RECT 560.4600 2240.0000 562.0600 2240.4800 ;
        RECT 560.4600 2245.4400 562.0600 2245.9200 ;
        RECT 560.4600 2223.6800 562.0600 2224.1600 ;
        RECT 560.4600 2229.1200 562.0600 2229.6000 ;
        RECT 560.4600 2234.5600 562.0600 2235.0400 ;
        RECT 515.4600 2240.0000 517.0600 2240.4800 ;
        RECT 515.4600 2245.4400 517.0600 2245.9200 ;
        RECT 515.4600 2223.6800 517.0600 2224.1600 ;
        RECT 515.4600 2229.1200 517.0600 2229.6000 ;
        RECT 515.4600 2234.5600 517.0600 2235.0400 ;
        RECT 560.4600 2212.8000 562.0600 2213.2800 ;
        RECT 560.4600 2218.2400 562.0600 2218.7200 ;
        RECT 560.4600 2196.4800 562.0600 2196.9600 ;
        RECT 560.4600 2201.9200 562.0600 2202.4000 ;
        RECT 560.4600 2207.3600 562.0600 2207.8400 ;
        RECT 515.4600 2212.8000 517.0600 2213.2800 ;
        RECT 515.4600 2218.2400 517.0600 2218.7200 ;
        RECT 515.4600 2196.4800 517.0600 2196.9600 ;
        RECT 515.4600 2201.9200 517.0600 2202.4000 ;
        RECT 515.4600 2207.3600 517.0600 2207.8400 ;
        RECT 465.9000 2240.0000 468.9000 2240.4800 ;
        RECT 465.9000 2245.4400 468.9000 2245.9200 ;
        RECT 465.9000 2229.1200 468.9000 2229.6000 ;
        RECT 465.9000 2223.6800 468.9000 2224.1600 ;
        RECT 465.9000 2234.5600 468.9000 2235.0400 ;
        RECT 465.9000 2212.8000 468.9000 2213.2800 ;
        RECT 465.9000 2218.2400 468.9000 2218.7200 ;
        RECT 465.9000 2201.9200 468.9000 2202.4000 ;
        RECT 465.9000 2196.4800 468.9000 2196.9600 ;
        RECT 465.9000 2207.3600 468.9000 2207.8400 ;
        RECT 560.4600 2185.6000 562.0600 2186.0800 ;
        RECT 560.4600 2191.0400 562.0600 2191.5200 ;
        RECT 560.4600 2169.2800 562.0600 2169.7600 ;
        RECT 560.4600 2174.7200 562.0600 2175.2000 ;
        RECT 560.4600 2180.1600 562.0600 2180.6400 ;
        RECT 515.4600 2185.6000 517.0600 2186.0800 ;
        RECT 515.4600 2191.0400 517.0600 2191.5200 ;
        RECT 515.4600 2169.2800 517.0600 2169.7600 ;
        RECT 515.4600 2174.7200 517.0600 2175.2000 ;
        RECT 515.4600 2180.1600 517.0600 2180.6400 ;
        RECT 560.4600 2163.8400 562.0600 2164.3200 ;
        RECT 560.4600 2158.4000 562.0600 2158.8800 ;
        RECT 560.4600 2152.9600 562.0600 2153.4400 ;
        RECT 515.4600 2163.8400 517.0600 2164.3200 ;
        RECT 515.4600 2158.4000 517.0600 2158.8800 ;
        RECT 515.4600 2152.9600 517.0600 2153.4400 ;
        RECT 465.9000 2185.6000 468.9000 2186.0800 ;
        RECT 465.9000 2191.0400 468.9000 2191.5200 ;
        RECT 465.9000 2174.7200 468.9000 2175.2000 ;
        RECT 465.9000 2169.2800 468.9000 2169.7600 ;
        RECT 465.9000 2180.1600 468.9000 2180.6400 ;
        RECT 465.9000 2158.4000 468.9000 2158.8800 ;
        RECT 465.9000 2163.8400 468.9000 2164.3200 ;
        RECT 465.9000 2152.9600 468.9000 2153.4400 ;
        RECT 465.9000 2351.1500 665.0000 2354.1500 ;
        RECT 465.9000 2146.0500 665.0000 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 1916.4100 652.0600 2124.5100 ;
        RECT 605.4600 1916.4100 607.0600 2124.5100 ;
        RECT 560.4600 1916.4100 562.0600 2124.5100 ;
        RECT 515.4600 1916.4100 517.0600 2124.5100 ;
        RECT 662.0000 1916.4100 665.0000 2124.5100 ;
        RECT 465.9000 1916.4100 468.9000 2124.5100 ;
      LAYER met3 ;
        RECT 662.0000 2119.1600 665.0000 2119.6400 ;
        RECT 650.4600 2119.1600 652.0600 2119.6400 ;
        RECT 662.0000 2108.2800 665.0000 2108.7600 ;
        RECT 662.0000 2113.7200 665.0000 2114.2000 ;
        RECT 650.4600 2108.2800 652.0600 2108.7600 ;
        RECT 650.4600 2113.7200 652.0600 2114.2000 ;
        RECT 662.0000 2091.9600 665.0000 2092.4400 ;
        RECT 662.0000 2097.4000 665.0000 2097.8800 ;
        RECT 650.4600 2091.9600 652.0600 2092.4400 ;
        RECT 650.4600 2097.4000 652.0600 2097.8800 ;
        RECT 662.0000 2081.0800 665.0000 2081.5600 ;
        RECT 662.0000 2086.5200 665.0000 2087.0000 ;
        RECT 650.4600 2081.0800 652.0600 2081.5600 ;
        RECT 650.4600 2086.5200 652.0600 2087.0000 ;
        RECT 662.0000 2102.8400 665.0000 2103.3200 ;
        RECT 650.4600 2102.8400 652.0600 2103.3200 ;
        RECT 605.4600 2108.2800 607.0600 2108.7600 ;
        RECT 605.4600 2113.7200 607.0600 2114.2000 ;
        RECT 605.4600 2119.1600 607.0600 2119.6400 ;
        RECT 605.4600 2091.9600 607.0600 2092.4400 ;
        RECT 605.4600 2097.4000 607.0600 2097.8800 ;
        RECT 605.4600 2086.5200 607.0600 2087.0000 ;
        RECT 605.4600 2081.0800 607.0600 2081.5600 ;
        RECT 605.4600 2102.8400 607.0600 2103.3200 ;
        RECT 662.0000 2064.7600 665.0000 2065.2400 ;
        RECT 662.0000 2070.2000 665.0000 2070.6800 ;
        RECT 650.4600 2064.7600 652.0600 2065.2400 ;
        RECT 650.4600 2070.2000 652.0600 2070.6800 ;
        RECT 662.0000 2048.4400 665.0000 2048.9200 ;
        RECT 662.0000 2053.8800 665.0000 2054.3600 ;
        RECT 662.0000 2059.3200 665.0000 2059.8000 ;
        RECT 650.4600 2048.4400 652.0600 2048.9200 ;
        RECT 650.4600 2053.8800 652.0600 2054.3600 ;
        RECT 650.4600 2059.3200 652.0600 2059.8000 ;
        RECT 662.0000 2037.5600 665.0000 2038.0400 ;
        RECT 662.0000 2043.0000 665.0000 2043.4800 ;
        RECT 650.4600 2037.5600 652.0600 2038.0400 ;
        RECT 650.4600 2043.0000 652.0600 2043.4800 ;
        RECT 662.0000 2021.2400 665.0000 2021.7200 ;
        RECT 662.0000 2026.6800 665.0000 2027.1600 ;
        RECT 662.0000 2032.1200 665.0000 2032.6000 ;
        RECT 650.4600 2021.2400 652.0600 2021.7200 ;
        RECT 650.4600 2026.6800 652.0600 2027.1600 ;
        RECT 650.4600 2032.1200 652.0600 2032.6000 ;
        RECT 605.4600 2064.7600 607.0600 2065.2400 ;
        RECT 605.4600 2070.2000 607.0600 2070.6800 ;
        RECT 605.4600 2048.4400 607.0600 2048.9200 ;
        RECT 605.4600 2053.8800 607.0600 2054.3600 ;
        RECT 605.4600 2059.3200 607.0600 2059.8000 ;
        RECT 605.4600 2037.5600 607.0600 2038.0400 ;
        RECT 605.4600 2043.0000 607.0600 2043.4800 ;
        RECT 605.4600 2021.2400 607.0600 2021.7200 ;
        RECT 605.4600 2026.6800 607.0600 2027.1600 ;
        RECT 605.4600 2032.1200 607.0600 2032.6000 ;
        RECT 662.0000 2075.6400 665.0000 2076.1200 ;
        RECT 605.4600 2075.6400 607.0600 2076.1200 ;
        RECT 650.4600 2075.6400 652.0600 2076.1200 ;
        RECT 560.4600 2108.2800 562.0600 2108.7600 ;
        RECT 560.4600 2113.7200 562.0600 2114.2000 ;
        RECT 560.4600 2119.1600 562.0600 2119.6400 ;
        RECT 515.4600 2108.2800 517.0600 2108.7600 ;
        RECT 515.4600 2113.7200 517.0600 2114.2000 ;
        RECT 515.4600 2119.1600 517.0600 2119.6400 ;
        RECT 560.4600 2091.9600 562.0600 2092.4400 ;
        RECT 560.4600 2097.4000 562.0600 2097.8800 ;
        RECT 560.4600 2081.0800 562.0600 2081.5600 ;
        RECT 560.4600 2086.5200 562.0600 2087.0000 ;
        RECT 515.4600 2091.9600 517.0600 2092.4400 ;
        RECT 515.4600 2097.4000 517.0600 2097.8800 ;
        RECT 515.4600 2081.0800 517.0600 2081.5600 ;
        RECT 515.4600 2086.5200 517.0600 2087.0000 ;
        RECT 515.4600 2102.8400 517.0600 2103.3200 ;
        RECT 560.4600 2102.8400 562.0600 2103.3200 ;
        RECT 465.9000 2119.1600 468.9000 2119.6400 ;
        RECT 465.9000 2113.7200 468.9000 2114.2000 ;
        RECT 465.9000 2108.2800 468.9000 2108.7600 ;
        RECT 465.9000 2097.4000 468.9000 2097.8800 ;
        RECT 465.9000 2091.9600 468.9000 2092.4400 ;
        RECT 465.9000 2086.5200 468.9000 2087.0000 ;
        RECT 465.9000 2081.0800 468.9000 2081.5600 ;
        RECT 465.9000 2102.8400 468.9000 2103.3200 ;
        RECT 560.4600 2064.7600 562.0600 2065.2400 ;
        RECT 560.4600 2070.2000 562.0600 2070.6800 ;
        RECT 560.4600 2048.4400 562.0600 2048.9200 ;
        RECT 560.4600 2053.8800 562.0600 2054.3600 ;
        RECT 560.4600 2059.3200 562.0600 2059.8000 ;
        RECT 515.4600 2064.7600 517.0600 2065.2400 ;
        RECT 515.4600 2070.2000 517.0600 2070.6800 ;
        RECT 515.4600 2048.4400 517.0600 2048.9200 ;
        RECT 515.4600 2053.8800 517.0600 2054.3600 ;
        RECT 515.4600 2059.3200 517.0600 2059.8000 ;
        RECT 560.4600 2037.5600 562.0600 2038.0400 ;
        RECT 560.4600 2043.0000 562.0600 2043.4800 ;
        RECT 560.4600 2021.2400 562.0600 2021.7200 ;
        RECT 560.4600 2026.6800 562.0600 2027.1600 ;
        RECT 560.4600 2032.1200 562.0600 2032.6000 ;
        RECT 515.4600 2037.5600 517.0600 2038.0400 ;
        RECT 515.4600 2043.0000 517.0600 2043.4800 ;
        RECT 515.4600 2021.2400 517.0600 2021.7200 ;
        RECT 515.4600 2026.6800 517.0600 2027.1600 ;
        RECT 515.4600 2032.1200 517.0600 2032.6000 ;
        RECT 465.9000 2064.7600 468.9000 2065.2400 ;
        RECT 465.9000 2070.2000 468.9000 2070.6800 ;
        RECT 465.9000 2053.8800 468.9000 2054.3600 ;
        RECT 465.9000 2048.4400 468.9000 2048.9200 ;
        RECT 465.9000 2059.3200 468.9000 2059.8000 ;
        RECT 465.9000 2037.5600 468.9000 2038.0400 ;
        RECT 465.9000 2043.0000 468.9000 2043.4800 ;
        RECT 465.9000 2026.6800 468.9000 2027.1600 ;
        RECT 465.9000 2021.2400 468.9000 2021.7200 ;
        RECT 465.9000 2032.1200 468.9000 2032.6000 ;
        RECT 465.9000 2075.6400 468.9000 2076.1200 ;
        RECT 515.4600 2075.6400 517.0600 2076.1200 ;
        RECT 560.4600 2075.6400 562.0600 2076.1200 ;
        RECT 662.0000 2010.3600 665.0000 2010.8400 ;
        RECT 662.0000 2015.8000 665.0000 2016.2800 ;
        RECT 650.4600 2010.3600 652.0600 2010.8400 ;
        RECT 650.4600 2015.8000 652.0600 2016.2800 ;
        RECT 662.0000 1994.0400 665.0000 1994.5200 ;
        RECT 662.0000 1999.4800 665.0000 1999.9600 ;
        RECT 662.0000 2004.9200 665.0000 2005.4000 ;
        RECT 650.4600 1994.0400 652.0600 1994.5200 ;
        RECT 650.4600 1999.4800 652.0600 1999.9600 ;
        RECT 650.4600 2004.9200 652.0600 2005.4000 ;
        RECT 662.0000 1983.1600 665.0000 1983.6400 ;
        RECT 662.0000 1988.6000 665.0000 1989.0800 ;
        RECT 650.4600 1983.1600 652.0600 1983.6400 ;
        RECT 650.4600 1988.6000 652.0600 1989.0800 ;
        RECT 662.0000 1966.8400 665.0000 1967.3200 ;
        RECT 662.0000 1972.2800 665.0000 1972.7600 ;
        RECT 662.0000 1977.7200 665.0000 1978.2000 ;
        RECT 650.4600 1966.8400 652.0600 1967.3200 ;
        RECT 650.4600 1972.2800 652.0600 1972.7600 ;
        RECT 650.4600 1977.7200 652.0600 1978.2000 ;
        RECT 605.4600 2010.3600 607.0600 2010.8400 ;
        RECT 605.4600 2015.8000 607.0600 2016.2800 ;
        RECT 605.4600 1994.0400 607.0600 1994.5200 ;
        RECT 605.4600 1999.4800 607.0600 1999.9600 ;
        RECT 605.4600 2004.9200 607.0600 2005.4000 ;
        RECT 605.4600 1983.1600 607.0600 1983.6400 ;
        RECT 605.4600 1988.6000 607.0600 1989.0800 ;
        RECT 605.4600 1966.8400 607.0600 1967.3200 ;
        RECT 605.4600 1972.2800 607.0600 1972.7600 ;
        RECT 605.4600 1977.7200 607.0600 1978.2000 ;
        RECT 662.0000 1955.9600 665.0000 1956.4400 ;
        RECT 662.0000 1961.4000 665.0000 1961.8800 ;
        RECT 650.4600 1955.9600 652.0600 1956.4400 ;
        RECT 650.4600 1961.4000 652.0600 1961.8800 ;
        RECT 662.0000 1939.6400 665.0000 1940.1200 ;
        RECT 662.0000 1945.0800 665.0000 1945.5600 ;
        RECT 662.0000 1950.5200 665.0000 1951.0000 ;
        RECT 650.4600 1939.6400 652.0600 1940.1200 ;
        RECT 650.4600 1945.0800 652.0600 1945.5600 ;
        RECT 650.4600 1950.5200 652.0600 1951.0000 ;
        RECT 662.0000 1928.7600 665.0000 1929.2400 ;
        RECT 662.0000 1934.2000 665.0000 1934.6800 ;
        RECT 650.4600 1928.7600 652.0600 1929.2400 ;
        RECT 650.4600 1934.2000 652.0600 1934.6800 ;
        RECT 662.0000 1923.3200 665.0000 1923.8000 ;
        RECT 650.4600 1923.3200 652.0600 1923.8000 ;
        RECT 605.4600 1955.9600 607.0600 1956.4400 ;
        RECT 605.4600 1961.4000 607.0600 1961.8800 ;
        RECT 605.4600 1939.6400 607.0600 1940.1200 ;
        RECT 605.4600 1945.0800 607.0600 1945.5600 ;
        RECT 605.4600 1950.5200 607.0600 1951.0000 ;
        RECT 605.4600 1928.7600 607.0600 1929.2400 ;
        RECT 605.4600 1934.2000 607.0600 1934.6800 ;
        RECT 605.4600 1923.3200 607.0600 1923.8000 ;
        RECT 560.4600 2010.3600 562.0600 2010.8400 ;
        RECT 560.4600 2015.8000 562.0600 2016.2800 ;
        RECT 560.4600 1994.0400 562.0600 1994.5200 ;
        RECT 560.4600 1999.4800 562.0600 1999.9600 ;
        RECT 560.4600 2004.9200 562.0600 2005.4000 ;
        RECT 515.4600 2010.3600 517.0600 2010.8400 ;
        RECT 515.4600 2015.8000 517.0600 2016.2800 ;
        RECT 515.4600 1994.0400 517.0600 1994.5200 ;
        RECT 515.4600 1999.4800 517.0600 1999.9600 ;
        RECT 515.4600 2004.9200 517.0600 2005.4000 ;
        RECT 560.4600 1983.1600 562.0600 1983.6400 ;
        RECT 560.4600 1988.6000 562.0600 1989.0800 ;
        RECT 560.4600 1966.8400 562.0600 1967.3200 ;
        RECT 560.4600 1972.2800 562.0600 1972.7600 ;
        RECT 560.4600 1977.7200 562.0600 1978.2000 ;
        RECT 515.4600 1983.1600 517.0600 1983.6400 ;
        RECT 515.4600 1988.6000 517.0600 1989.0800 ;
        RECT 515.4600 1966.8400 517.0600 1967.3200 ;
        RECT 515.4600 1972.2800 517.0600 1972.7600 ;
        RECT 515.4600 1977.7200 517.0600 1978.2000 ;
        RECT 465.9000 2010.3600 468.9000 2010.8400 ;
        RECT 465.9000 2015.8000 468.9000 2016.2800 ;
        RECT 465.9000 1999.4800 468.9000 1999.9600 ;
        RECT 465.9000 1994.0400 468.9000 1994.5200 ;
        RECT 465.9000 2004.9200 468.9000 2005.4000 ;
        RECT 465.9000 1983.1600 468.9000 1983.6400 ;
        RECT 465.9000 1988.6000 468.9000 1989.0800 ;
        RECT 465.9000 1972.2800 468.9000 1972.7600 ;
        RECT 465.9000 1966.8400 468.9000 1967.3200 ;
        RECT 465.9000 1977.7200 468.9000 1978.2000 ;
        RECT 560.4600 1955.9600 562.0600 1956.4400 ;
        RECT 560.4600 1961.4000 562.0600 1961.8800 ;
        RECT 560.4600 1939.6400 562.0600 1940.1200 ;
        RECT 560.4600 1945.0800 562.0600 1945.5600 ;
        RECT 560.4600 1950.5200 562.0600 1951.0000 ;
        RECT 515.4600 1955.9600 517.0600 1956.4400 ;
        RECT 515.4600 1961.4000 517.0600 1961.8800 ;
        RECT 515.4600 1939.6400 517.0600 1940.1200 ;
        RECT 515.4600 1945.0800 517.0600 1945.5600 ;
        RECT 515.4600 1950.5200 517.0600 1951.0000 ;
        RECT 560.4600 1934.2000 562.0600 1934.6800 ;
        RECT 560.4600 1928.7600 562.0600 1929.2400 ;
        RECT 560.4600 1923.3200 562.0600 1923.8000 ;
        RECT 515.4600 1934.2000 517.0600 1934.6800 ;
        RECT 515.4600 1928.7600 517.0600 1929.2400 ;
        RECT 515.4600 1923.3200 517.0600 1923.8000 ;
        RECT 465.9000 1955.9600 468.9000 1956.4400 ;
        RECT 465.9000 1961.4000 468.9000 1961.8800 ;
        RECT 465.9000 1945.0800 468.9000 1945.5600 ;
        RECT 465.9000 1939.6400 468.9000 1940.1200 ;
        RECT 465.9000 1950.5200 468.9000 1951.0000 ;
        RECT 465.9000 1928.7600 468.9000 1929.2400 ;
        RECT 465.9000 1934.2000 468.9000 1934.6800 ;
        RECT 465.9000 1923.3200 468.9000 1923.8000 ;
        RECT 465.9000 2121.5100 665.0000 2124.5100 ;
        RECT 465.9000 1916.4100 665.0000 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 1686.7700 652.0600 1894.8700 ;
        RECT 605.4600 1686.7700 607.0600 1894.8700 ;
        RECT 560.4600 1686.7700 562.0600 1894.8700 ;
        RECT 515.4600 1686.7700 517.0600 1894.8700 ;
        RECT 662.0000 1686.7700 665.0000 1894.8700 ;
        RECT 465.9000 1686.7700 468.9000 1894.8700 ;
      LAYER met3 ;
        RECT 662.0000 1889.5200 665.0000 1890.0000 ;
        RECT 650.4600 1889.5200 652.0600 1890.0000 ;
        RECT 662.0000 1878.6400 665.0000 1879.1200 ;
        RECT 662.0000 1884.0800 665.0000 1884.5600 ;
        RECT 650.4600 1878.6400 652.0600 1879.1200 ;
        RECT 650.4600 1884.0800 652.0600 1884.5600 ;
        RECT 662.0000 1862.3200 665.0000 1862.8000 ;
        RECT 662.0000 1867.7600 665.0000 1868.2400 ;
        RECT 650.4600 1862.3200 652.0600 1862.8000 ;
        RECT 650.4600 1867.7600 652.0600 1868.2400 ;
        RECT 662.0000 1851.4400 665.0000 1851.9200 ;
        RECT 662.0000 1856.8800 665.0000 1857.3600 ;
        RECT 650.4600 1851.4400 652.0600 1851.9200 ;
        RECT 650.4600 1856.8800 652.0600 1857.3600 ;
        RECT 662.0000 1873.2000 665.0000 1873.6800 ;
        RECT 650.4600 1873.2000 652.0600 1873.6800 ;
        RECT 605.4600 1878.6400 607.0600 1879.1200 ;
        RECT 605.4600 1884.0800 607.0600 1884.5600 ;
        RECT 605.4600 1889.5200 607.0600 1890.0000 ;
        RECT 605.4600 1862.3200 607.0600 1862.8000 ;
        RECT 605.4600 1867.7600 607.0600 1868.2400 ;
        RECT 605.4600 1856.8800 607.0600 1857.3600 ;
        RECT 605.4600 1851.4400 607.0600 1851.9200 ;
        RECT 605.4600 1873.2000 607.0600 1873.6800 ;
        RECT 662.0000 1835.1200 665.0000 1835.6000 ;
        RECT 662.0000 1840.5600 665.0000 1841.0400 ;
        RECT 650.4600 1835.1200 652.0600 1835.6000 ;
        RECT 650.4600 1840.5600 652.0600 1841.0400 ;
        RECT 662.0000 1818.8000 665.0000 1819.2800 ;
        RECT 662.0000 1824.2400 665.0000 1824.7200 ;
        RECT 662.0000 1829.6800 665.0000 1830.1600 ;
        RECT 650.4600 1818.8000 652.0600 1819.2800 ;
        RECT 650.4600 1824.2400 652.0600 1824.7200 ;
        RECT 650.4600 1829.6800 652.0600 1830.1600 ;
        RECT 662.0000 1807.9200 665.0000 1808.4000 ;
        RECT 662.0000 1813.3600 665.0000 1813.8400 ;
        RECT 650.4600 1807.9200 652.0600 1808.4000 ;
        RECT 650.4600 1813.3600 652.0600 1813.8400 ;
        RECT 662.0000 1791.6000 665.0000 1792.0800 ;
        RECT 662.0000 1797.0400 665.0000 1797.5200 ;
        RECT 662.0000 1802.4800 665.0000 1802.9600 ;
        RECT 650.4600 1791.6000 652.0600 1792.0800 ;
        RECT 650.4600 1797.0400 652.0600 1797.5200 ;
        RECT 650.4600 1802.4800 652.0600 1802.9600 ;
        RECT 605.4600 1835.1200 607.0600 1835.6000 ;
        RECT 605.4600 1840.5600 607.0600 1841.0400 ;
        RECT 605.4600 1818.8000 607.0600 1819.2800 ;
        RECT 605.4600 1824.2400 607.0600 1824.7200 ;
        RECT 605.4600 1829.6800 607.0600 1830.1600 ;
        RECT 605.4600 1807.9200 607.0600 1808.4000 ;
        RECT 605.4600 1813.3600 607.0600 1813.8400 ;
        RECT 605.4600 1791.6000 607.0600 1792.0800 ;
        RECT 605.4600 1797.0400 607.0600 1797.5200 ;
        RECT 605.4600 1802.4800 607.0600 1802.9600 ;
        RECT 662.0000 1846.0000 665.0000 1846.4800 ;
        RECT 605.4600 1846.0000 607.0600 1846.4800 ;
        RECT 650.4600 1846.0000 652.0600 1846.4800 ;
        RECT 560.4600 1878.6400 562.0600 1879.1200 ;
        RECT 560.4600 1884.0800 562.0600 1884.5600 ;
        RECT 560.4600 1889.5200 562.0600 1890.0000 ;
        RECT 515.4600 1878.6400 517.0600 1879.1200 ;
        RECT 515.4600 1884.0800 517.0600 1884.5600 ;
        RECT 515.4600 1889.5200 517.0600 1890.0000 ;
        RECT 560.4600 1862.3200 562.0600 1862.8000 ;
        RECT 560.4600 1867.7600 562.0600 1868.2400 ;
        RECT 560.4600 1851.4400 562.0600 1851.9200 ;
        RECT 560.4600 1856.8800 562.0600 1857.3600 ;
        RECT 515.4600 1862.3200 517.0600 1862.8000 ;
        RECT 515.4600 1867.7600 517.0600 1868.2400 ;
        RECT 515.4600 1851.4400 517.0600 1851.9200 ;
        RECT 515.4600 1856.8800 517.0600 1857.3600 ;
        RECT 515.4600 1873.2000 517.0600 1873.6800 ;
        RECT 560.4600 1873.2000 562.0600 1873.6800 ;
        RECT 465.9000 1889.5200 468.9000 1890.0000 ;
        RECT 465.9000 1884.0800 468.9000 1884.5600 ;
        RECT 465.9000 1878.6400 468.9000 1879.1200 ;
        RECT 465.9000 1867.7600 468.9000 1868.2400 ;
        RECT 465.9000 1862.3200 468.9000 1862.8000 ;
        RECT 465.9000 1856.8800 468.9000 1857.3600 ;
        RECT 465.9000 1851.4400 468.9000 1851.9200 ;
        RECT 465.9000 1873.2000 468.9000 1873.6800 ;
        RECT 560.4600 1835.1200 562.0600 1835.6000 ;
        RECT 560.4600 1840.5600 562.0600 1841.0400 ;
        RECT 560.4600 1818.8000 562.0600 1819.2800 ;
        RECT 560.4600 1824.2400 562.0600 1824.7200 ;
        RECT 560.4600 1829.6800 562.0600 1830.1600 ;
        RECT 515.4600 1835.1200 517.0600 1835.6000 ;
        RECT 515.4600 1840.5600 517.0600 1841.0400 ;
        RECT 515.4600 1818.8000 517.0600 1819.2800 ;
        RECT 515.4600 1824.2400 517.0600 1824.7200 ;
        RECT 515.4600 1829.6800 517.0600 1830.1600 ;
        RECT 560.4600 1807.9200 562.0600 1808.4000 ;
        RECT 560.4600 1813.3600 562.0600 1813.8400 ;
        RECT 560.4600 1791.6000 562.0600 1792.0800 ;
        RECT 560.4600 1797.0400 562.0600 1797.5200 ;
        RECT 560.4600 1802.4800 562.0600 1802.9600 ;
        RECT 515.4600 1807.9200 517.0600 1808.4000 ;
        RECT 515.4600 1813.3600 517.0600 1813.8400 ;
        RECT 515.4600 1791.6000 517.0600 1792.0800 ;
        RECT 515.4600 1797.0400 517.0600 1797.5200 ;
        RECT 515.4600 1802.4800 517.0600 1802.9600 ;
        RECT 465.9000 1835.1200 468.9000 1835.6000 ;
        RECT 465.9000 1840.5600 468.9000 1841.0400 ;
        RECT 465.9000 1824.2400 468.9000 1824.7200 ;
        RECT 465.9000 1818.8000 468.9000 1819.2800 ;
        RECT 465.9000 1829.6800 468.9000 1830.1600 ;
        RECT 465.9000 1807.9200 468.9000 1808.4000 ;
        RECT 465.9000 1813.3600 468.9000 1813.8400 ;
        RECT 465.9000 1797.0400 468.9000 1797.5200 ;
        RECT 465.9000 1791.6000 468.9000 1792.0800 ;
        RECT 465.9000 1802.4800 468.9000 1802.9600 ;
        RECT 465.9000 1846.0000 468.9000 1846.4800 ;
        RECT 515.4600 1846.0000 517.0600 1846.4800 ;
        RECT 560.4600 1846.0000 562.0600 1846.4800 ;
        RECT 662.0000 1780.7200 665.0000 1781.2000 ;
        RECT 662.0000 1786.1600 665.0000 1786.6400 ;
        RECT 650.4600 1780.7200 652.0600 1781.2000 ;
        RECT 650.4600 1786.1600 652.0600 1786.6400 ;
        RECT 662.0000 1764.4000 665.0000 1764.8800 ;
        RECT 662.0000 1769.8400 665.0000 1770.3200 ;
        RECT 662.0000 1775.2800 665.0000 1775.7600 ;
        RECT 650.4600 1764.4000 652.0600 1764.8800 ;
        RECT 650.4600 1769.8400 652.0600 1770.3200 ;
        RECT 650.4600 1775.2800 652.0600 1775.7600 ;
        RECT 662.0000 1753.5200 665.0000 1754.0000 ;
        RECT 662.0000 1758.9600 665.0000 1759.4400 ;
        RECT 650.4600 1753.5200 652.0600 1754.0000 ;
        RECT 650.4600 1758.9600 652.0600 1759.4400 ;
        RECT 662.0000 1737.2000 665.0000 1737.6800 ;
        RECT 662.0000 1742.6400 665.0000 1743.1200 ;
        RECT 662.0000 1748.0800 665.0000 1748.5600 ;
        RECT 650.4600 1737.2000 652.0600 1737.6800 ;
        RECT 650.4600 1742.6400 652.0600 1743.1200 ;
        RECT 650.4600 1748.0800 652.0600 1748.5600 ;
        RECT 605.4600 1780.7200 607.0600 1781.2000 ;
        RECT 605.4600 1786.1600 607.0600 1786.6400 ;
        RECT 605.4600 1764.4000 607.0600 1764.8800 ;
        RECT 605.4600 1769.8400 607.0600 1770.3200 ;
        RECT 605.4600 1775.2800 607.0600 1775.7600 ;
        RECT 605.4600 1753.5200 607.0600 1754.0000 ;
        RECT 605.4600 1758.9600 607.0600 1759.4400 ;
        RECT 605.4600 1737.2000 607.0600 1737.6800 ;
        RECT 605.4600 1742.6400 607.0600 1743.1200 ;
        RECT 605.4600 1748.0800 607.0600 1748.5600 ;
        RECT 662.0000 1726.3200 665.0000 1726.8000 ;
        RECT 662.0000 1731.7600 665.0000 1732.2400 ;
        RECT 650.4600 1726.3200 652.0600 1726.8000 ;
        RECT 650.4600 1731.7600 652.0600 1732.2400 ;
        RECT 662.0000 1710.0000 665.0000 1710.4800 ;
        RECT 662.0000 1715.4400 665.0000 1715.9200 ;
        RECT 662.0000 1720.8800 665.0000 1721.3600 ;
        RECT 650.4600 1710.0000 652.0600 1710.4800 ;
        RECT 650.4600 1715.4400 652.0600 1715.9200 ;
        RECT 650.4600 1720.8800 652.0600 1721.3600 ;
        RECT 662.0000 1699.1200 665.0000 1699.6000 ;
        RECT 662.0000 1704.5600 665.0000 1705.0400 ;
        RECT 650.4600 1699.1200 652.0600 1699.6000 ;
        RECT 650.4600 1704.5600 652.0600 1705.0400 ;
        RECT 662.0000 1693.6800 665.0000 1694.1600 ;
        RECT 650.4600 1693.6800 652.0600 1694.1600 ;
        RECT 605.4600 1726.3200 607.0600 1726.8000 ;
        RECT 605.4600 1731.7600 607.0600 1732.2400 ;
        RECT 605.4600 1710.0000 607.0600 1710.4800 ;
        RECT 605.4600 1715.4400 607.0600 1715.9200 ;
        RECT 605.4600 1720.8800 607.0600 1721.3600 ;
        RECT 605.4600 1699.1200 607.0600 1699.6000 ;
        RECT 605.4600 1704.5600 607.0600 1705.0400 ;
        RECT 605.4600 1693.6800 607.0600 1694.1600 ;
        RECT 560.4600 1780.7200 562.0600 1781.2000 ;
        RECT 560.4600 1786.1600 562.0600 1786.6400 ;
        RECT 560.4600 1764.4000 562.0600 1764.8800 ;
        RECT 560.4600 1769.8400 562.0600 1770.3200 ;
        RECT 560.4600 1775.2800 562.0600 1775.7600 ;
        RECT 515.4600 1780.7200 517.0600 1781.2000 ;
        RECT 515.4600 1786.1600 517.0600 1786.6400 ;
        RECT 515.4600 1764.4000 517.0600 1764.8800 ;
        RECT 515.4600 1769.8400 517.0600 1770.3200 ;
        RECT 515.4600 1775.2800 517.0600 1775.7600 ;
        RECT 560.4600 1753.5200 562.0600 1754.0000 ;
        RECT 560.4600 1758.9600 562.0600 1759.4400 ;
        RECT 560.4600 1737.2000 562.0600 1737.6800 ;
        RECT 560.4600 1742.6400 562.0600 1743.1200 ;
        RECT 560.4600 1748.0800 562.0600 1748.5600 ;
        RECT 515.4600 1753.5200 517.0600 1754.0000 ;
        RECT 515.4600 1758.9600 517.0600 1759.4400 ;
        RECT 515.4600 1737.2000 517.0600 1737.6800 ;
        RECT 515.4600 1742.6400 517.0600 1743.1200 ;
        RECT 515.4600 1748.0800 517.0600 1748.5600 ;
        RECT 465.9000 1780.7200 468.9000 1781.2000 ;
        RECT 465.9000 1786.1600 468.9000 1786.6400 ;
        RECT 465.9000 1769.8400 468.9000 1770.3200 ;
        RECT 465.9000 1764.4000 468.9000 1764.8800 ;
        RECT 465.9000 1775.2800 468.9000 1775.7600 ;
        RECT 465.9000 1753.5200 468.9000 1754.0000 ;
        RECT 465.9000 1758.9600 468.9000 1759.4400 ;
        RECT 465.9000 1742.6400 468.9000 1743.1200 ;
        RECT 465.9000 1737.2000 468.9000 1737.6800 ;
        RECT 465.9000 1748.0800 468.9000 1748.5600 ;
        RECT 560.4600 1726.3200 562.0600 1726.8000 ;
        RECT 560.4600 1731.7600 562.0600 1732.2400 ;
        RECT 560.4600 1710.0000 562.0600 1710.4800 ;
        RECT 560.4600 1715.4400 562.0600 1715.9200 ;
        RECT 560.4600 1720.8800 562.0600 1721.3600 ;
        RECT 515.4600 1726.3200 517.0600 1726.8000 ;
        RECT 515.4600 1731.7600 517.0600 1732.2400 ;
        RECT 515.4600 1710.0000 517.0600 1710.4800 ;
        RECT 515.4600 1715.4400 517.0600 1715.9200 ;
        RECT 515.4600 1720.8800 517.0600 1721.3600 ;
        RECT 560.4600 1704.5600 562.0600 1705.0400 ;
        RECT 560.4600 1699.1200 562.0600 1699.6000 ;
        RECT 560.4600 1693.6800 562.0600 1694.1600 ;
        RECT 515.4600 1704.5600 517.0600 1705.0400 ;
        RECT 515.4600 1699.1200 517.0600 1699.6000 ;
        RECT 515.4600 1693.6800 517.0600 1694.1600 ;
        RECT 465.9000 1726.3200 468.9000 1726.8000 ;
        RECT 465.9000 1731.7600 468.9000 1732.2400 ;
        RECT 465.9000 1715.4400 468.9000 1715.9200 ;
        RECT 465.9000 1710.0000 468.9000 1710.4800 ;
        RECT 465.9000 1720.8800 468.9000 1721.3600 ;
        RECT 465.9000 1699.1200 468.9000 1699.6000 ;
        RECT 465.9000 1704.5600 468.9000 1705.0400 ;
        RECT 465.9000 1693.6800 468.9000 1694.1600 ;
        RECT 465.9000 1891.8700 665.0000 1894.8700 ;
        RECT 465.9000 1686.7700 665.0000 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 1457.1300 652.0600 1665.2300 ;
        RECT 605.4600 1457.1300 607.0600 1665.2300 ;
        RECT 560.4600 1457.1300 562.0600 1665.2300 ;
        RECT 515.4600 1457.1300 517.0600 1665.2300 ;
        RECT 662.0000 1457.1300 665.0000 1665.2300 ;
        RECT 465.9000 1457.1300 468.9000 1665.2300 ;
      LAYER met3 ;
        RECT 662.0000 1659.8800 665.0000 1660.3600 ;
        RECT 650.4600 1659.8800 652.0600 1660.3600 ;
        RECT 662.0000 1649.0000 665.0000 1649.4800 ;
        RECT 662.0000 1654.4400 665.0000 1654.9200 ;
        RECT 650.4600 1649.0000 652.0600 1649.4800 ;
        RECT 650.4600 1654.4400 652.0600 1654.9200 ;
        RECT 662.0000 1632.6800 665.0000 1633.1600 ;
        RECT 662.0000 1638.1200 665.0000 1638.6000 ;
        RECT 650.4600 1632.6800 652.0600 1633.1600 ;
        RECT 650.4600 1638.1200 652.0600 1638.6000 ;
        RECT 662.0000 1621.8000 665.0000 1622.2800 ;
        RECT 662.0000 1627.2400 665.0000 1627.7200 ;
        RECT 650.4600 1621.8000 652.0600 1622.2800 ;
        RECT 650.4600 1627.2400 652.0600 1627.7200 ;
        RECT 662.0000 1643.5600 665.0000 1644.0400 ;
        RECT 650.4600 1643.5600 652.0600 1644.0400 ;
        RECT 605.4600 1649.0000 607.0600 1649.4800 ;
        RECT 605.4600 1654.4400 607.0600 1654.9200 ;
        RECT 605.4600 1659.8800 607.0600 1660.3600 ;
        RECT 605.4600 1632.6800 607.0600 1633.1600 ;
        RECT 605.4600 1638.1200 607.0600 1638.6000 ;
        RECT 605.4600 1627.2400 607.0600 1627.7200 ;
        RECT 605.4600 1621.8000 607.0600 1622.2800 ;
        RECT 605.4600 1643.5600 607.0600 1644.0400 ;
        RECT 662.0000 1605.4800 665.0000 1605.9600 ;
        RECT 662.0000 1610.9200 665.0000 1611.4000 ;
        RECT 650.4600 1605.4800 652.0600 1605.9600 ;
        RECT 650.4600 1610.9200 652.0600 1611.4000 ;
        RECT 662.0000 1589.1600 665.0000 1589.6400 ;
        RECT 662.0000 1594.6000 665.0000 1595.0800 ;
        RECT 662.0000 1600.0400 665.0000 1600.5200 ;
        RECT 650.4600 1589.1600 652.0600 1589.6400 ;
        RECT 650.4600 1594.6000 652.0600 1595.0800 ;
        RECT 650.4600 1600.0400 652.0600 1600.5200 ;
        RECT 662.0000 1578.2800 665.0000 1578.7600 ;
        RECT 662.0000 1583.7200 665.0000 1584.2000 ;
        RECT 650.4600 1578.2800 652.0600 1578.7600 ;
        RECT 650.4600 1583.7200 652.0600 1584.2000 ;
        RECT 662.0000 1561.9600 665.0000 1562.4400 ;
        RECT 662.0000 1567.4000 665.0000 1567.8800 ;
        RECT 662.0000 1572.8400 665.0000 1573.3200 ;
        RECT 650.4600 1561.9600 652.0600 1562.4400 ;
        RECT 650.4600 1567.4000 652.0600 1567.8800 ;
        RECT 650.4600 1572.8400 652.0600 1573.3200 ;
        RECT 605.4600 1605.4800 607.0600 1605.9600 ;
        RECT 605.4600 1610.9200 607.0600 1611.4000 ;
        RECT 605.4600 1589.1600 607.0600 1589.6400 ;
        RECT 605.4600 1594.6000 607.0600 1595.0800 ;
        RECT 605.4600 1600.0400 607.0600 1600.5200 ;
        RECT 605.4600 1578.2800 607.0600 1578.7600 ;
        RECT 605.4600 1583.7200 607.0600 1584.2000 ;
        RECT 605.4600 1561.9600 607.0600 1562.4400 ;
        RECT 605.4600 1567.4000 607.0600 1567.8800 ;
        RECT 605.4600 1572.8400 607.0600 1573.3200 ;
        RECT 662.0000 1616.3600 665.0000 1616.8400 ;
        RECT 605.4600 1616.3600 607.0600 1616.8400 ;
        RECT 650.4600 1616.3600 652.0600 1616.8400 ;
        RECT 560.4600 1649.0000 562.0600 1649.4800 ;
        RECT 560.4600 1654.4400 562.0600 1654.9200 ;
        RECT 560.4600 1659.8800 562.0600 1660.3600 ;
        RECT 515.4600 1649.0000 517.0600 1649.4800 ;
        RECT 515.4600 1654.4400 517.0600 1654.9200 ;
        RECT 515.4600 1659.8800 517.0600 1660.3600 ;
        RECT 560.4600 1632.6800 562.0600 1633.1600 ;
        RECT 560.4600 1638.1200 562.0600 1638.6000 ;
        RECT 560.4600 1621.8000 562.0600 1622.2800 ;
        RECT 560.4600 1627.2400 562.0600 1627.7200 ;
        RECT 515.4600 1632.6800 517.0600 1633.1600 ;
        RECT 515.4600 1638.1200 517.0600 1638.6000 ;
        RECT 515.4600 1621.8000 517.0600 1622.2800 ;
        RECT 515.4600 1627.2400 517.0600 1627.7200 ;
        RECT 515.4600 1643.5600 517.0600 1644.0400 ;
        RECT 560.4600 1643.5600 562.0600 1644.0400 ;
        RECT 465.9000 1659.8800 468.9000 1660.3600 ;
        RECT 465.9000 1654.4400 468.9000 1654.9200 ;
        RECT 465.9000 1649.0000 468.9000 1649.4800 ;
        RECT 465.9000 1638.1200 468.9000 1638.6000 ;
        RECT 465.9000 1632.6800 468.9000 1633.1600 ;
        RECT 465.9000 1627.2400 468.9000 1627.7200 ;
        RECT 465.9000 1621.8000 468.9000 1622.2800 ;
        RECT 465.9000 1643.5600 468.9000 1644.0400 ;
        RECT 560.4600 1605.4800 562.0600 1605.9600 ;
        RECT 560.4600 1610.9200 562.0600 1611.4000 ;
        RECT 560.4600 1589.1600 562.0600 1589.6400 ;
        RECT 560.4600 1594.6000 562.0600 1595.0800 ;
        RECT 560.4600 1600.0400 562.0600 1600.5200 ;
        RECT 515.4600 1605.4800 517.0600 1605.9600 ;
        RECT 515.4600 1610.9200 517.0600 1611.4000 ;
        RECT 515.4600 1589.1600 517.0600 1589.6400 ;
        RECT 515.4600 1594.6000 517.0600 1595.0800 ;
        RECT 515.4600 1600.0400 517.0600 1600.5200 ;
        RECT 560.4600 1578.2800 562.0600 1578.7600 ;
        RECT 560.4600 1583.7200 562.0600 1584.2000 ;
        RECT 560.4600 1561.9600 562.0600 1562.4400 ;
        RECT 560.4600 1567.4000 562.0600 1567.8800 ;
        RECT 560.4600 1572.8400 562.0600 1573.3200 ;
        RECT 515.4600 1578.2800 517.0600 1578.7600 ;
        RECT 515.4600 1583.7200 517.0600 1584.2000 ;
        RECT 515.4600 1561.9600 517.0600 1562.4400 ;
        RECT 515.4600 1567.4000 517.0600 1567.8800 ;
        RECT 515.4600 1572.8400 517.0600 1573.3200 ;
        RECT 465.9000 1605.4800 468.9000 1605.9600 ;
        RECT 465.9000 1610.9200 468.9000 1611.4000 ;
        RECT 465.9000 1594.6000 468.9000 1595.0800 ;
        RECT 465.9000 1589.1600 468.9000 1589.6400 ;
        RECT 465.9000 1600.0400 468.9000 1600.5200 ;
        RECT 465.9000 1578.2800 468.9000 1578.7600 ;
        RECT 465.9000 1583.7200 468.9000 1584.2000 ;
        RECT 465.9000 1567.4000 468.9000 1567.8800 ;
        RECT 465.9000 1561.9600 468.9000 1562.4400 ;
        RECT 465.9000 1572.8400 468.9000 1573.3200 ;
        RECT 465.9000 1616.3600 468.9000 1616.8400 ;
        RECT 515.4600 1616.3600 517.0600 1616.8400 ;
        RECT 560.4600 1616.3600 562.0600 1616.8400 ;
        RECT 662.0000 1551.0800 665.0000 1551.5600 ;
        RECT 662.0000 1556.5200 665.0000 1557.0000 ;
        RECT 650.4600 1551.0800 652.0600 1551.5600 ;
        RECT 650.4600 1556.5200 652.0600 1557.0000 ;
        RECT 662.0000 1534.7600 665.0000 1535.2400 ;
        RECT 662.0000 1540.2000 665.0000 1540.6800 ;
        RECT 662.0000 1545.6400 665.0000 1546.1200 ;
        RECT 650.4600 1534.7600 652.0600 1535.2400 ;
        RECT 650.4600 1540.2000 652.0600 1540.6800 ;
        RECT 650.4600 1545.6400 652.0600 1546.1200 ;
        RECT 662.0000 1523.8800 665.0000 1524.3600 ;
        RECT 662.0000 1529.3200 665.0000 1529.8000 ;
        RECT 650.4600 1523.8800 652.0600 1524.3600 ;
        RECT 650.4600 1529.3200 652.0600 1529.8000 ;
        RECT 662.0000 1507.5600 665.0000 1508.0400 ;
        RECT 662.0000 1513.0000 665.0000 1513.4800 ;
        RECT 662.0000 1518.4400 665.0000 1518.9200 ;
        RECT 650.4600 1507.5600 652.0600 1508.0400 ;
        RECT 650.4600 1513.0000 652.0600 1513.4800 ;
        RECT 650.4600 1518.4400 652.0600 1518.9200 ;
        RECT 605.4600 1551.0800 607.0600 1551.5600 ;
        RECT 605.4600 1556.5200 607.0600 1557.0000 ;
        RECT 605.4600 1534.7600 607.0600 1535.2400 ;
        RECT 605.4600 1540.2000 607.0600 1540.6800 ;
        RECT 605.4600 1545.6400 607.0600 1546.1200 ;
        RECT 605.4600 1523.8800 607.0600 1524.3600 ;
        RECT 605.4600 1529.3200 607.0600 1529.8000 ;
        RECT 605.4600 1507.5600 607.0600 1508.0400 ;
        RECT 605.4600 1513.0000 607.0600 1513.4800 ;
        RECT 605.4600 1518.4400 607.0600 1518.9200 ;
        RECT 662.0000 1496.6800 665.0000 1497.1600 ;
        RECT 662.0000 1502.1200 665.0000 1502.6000 ;
        RECT 650.4600 1496.6800 652.0600 1497.1600 ;
        RECT 650.4600 1502.1200 652.0600 1502.6000 ;
        RECT 662.0000 1480.3600 665.0000 1480.8400 ;
        RECT 662.0000 1485.8000 665.0000 1486.2800 ;
        RECT 662.0000 1491.2400 665.0000 1491.7200 ;
        RECT 650.4600 1480.3600 652.0600 1480.8400 ;
        RECT 650.4600 1485.8000 652.0600 1486.2800 ;
        RECT 650.4600 1491.2400 652.0600 1491.7200 ;
        RECT 662.0000 1469.4800 665.0000 1469.9600 ;
        RECT 662.0000 1474.9200 665.0000 1475.4000 ;
        RECT 650.4600 1469.4800 652.0600 1469.9600 ;
        RECT 650.4600 1474.9200 652.0600 1475.4000 ;
        RECT 662.0000 1464.0400 665.0000 1464.5200 ;
        RECT 650.4600 1464.0400 652.0600 1464.5200 ;
        RECT 605.4600 1496.6800 607.0600 1497.1600 ;
        RECT 605.4600 1502.1200 607.0600 1502.6000 ;
        RECT 605.4600 1480.3600 607.0600 1480.8400 ;
        RECT 605.4600 1485.8000 607.0600 1486.2800 ;
        RECT 605.4600 1491.2400 607.0600 1491.7200 ;
        RECT 605.4600 1469.4800 607.0600 1469.9600 ;
        RECT 605.4600 1474.9200 607.0600 1475.4000 ;
        RECT 605.4600 1464.0400 607.0600 1464.5200 ;
        RECT 560.4600 1551.0800 562.0600 1551.5600 ;
        RECT 560.4600 1556.5200 562.0600 1557.0000 ;
        RECT 560.4600 1534.7600 562.0600 1535.2400 ;
        RECT 560.4600 1540.2000 562.0600 1540.6800 ;
        RECT 560.4600 1545.6400 562.0600 1546.1200 ;
        RECT 515.4600 1551.0800 517.0600 1551.5600 ;
        RECT 515.4600 1556.5200 517.0600 1557.0000 ;
        RECT 515.4600 1534.7600 517.0600 1535.2400 ;
        RECT 515.4600 1540.2000 517.0600 1540.6800 ;
        RECT 515.4600 1545.6400 517.0600 1546.1200 ;
        RECT 560.4600 1523.8800 562.0600 1524.3600 ;
        RECT 560.4600 1529.3200 562.0600 1529.8000 ;
        RECT 560.4600 1507.5600 562.0600 1508.0400 ;
        RECT 560.4600 1513.0000 562.0600 1513.4800 ;
        RECT 560.4600 1518.4400 562.0600 1518.9200 ;
        RECT 515.4600 1523.8800 517.0600 1524.3600 ;
        RECT 515.4600 1529.3200 517.0600 1529.8000 ;
        RECT 515.4600 1507.5600 517.0600 1508.0400 ;
        RECT 515.4600 1513.0000 517.0600 1513.4800 ;
        RECT 515.4600 1518.4400 517.0600 1518.9200 ;
        RECT 465.9000 1551.0800 468.9000 1551.5600 ;
        RECT 465.9000 1556.5200 468.9000 1557.0000 ;
        RECT 465.9000 1540.2000 468.9000 1540.6800 ;
        RECT 465.9000 1534.7600 468.9000 1535.2400 ;
        RECT 465.9000 1545.6400 468.9000 1546.1200 ;
        RECT 465.9000 1523.8800 468.9000 1524.3600 ;
        RECT 465.9000 1529.3200 468.9000 1529.8000 ;
        RECT 465.9000 1513.0000 468.9000 1513.4800 ;
        RECT 465.9000 1507.5600 468.9000 1508.0400 ;
        RECT 465.9000 1518.4400 468.9000 1518.9200 ;
        RECT 560.4600 1496.6800 562.0600 1497.1600 ;
        RECT 560.4600 1502.1200 562.0600 1502.6000 ;
        RECT 560.4600 1480.3600 562.0600 1480.8400 ;
        RECT 560.4600 1485.8000 562.0600 1486.2800 ;
        RECT 560.4600 1491.2400 562.0600 1491.7200 ;
        RECT 515.4600 1496.6800 517.0600 1497.1600 ;
        RECT 515.4600 1502.1200 517.0600 1502.6000 ;
        RECT 515.4600 1480.3600 517.0600 1480.8400 ;
        RECT 515.4600 1485.8000 517.0600 1486.2800 ;
        RECT 515.4600 1491.2400 517.0600 1491.7200 ;
        RECT 560.4600 1474.9200 562.0600 1475.4000 ;
        RECT 560.4600 1469.4800 562.0600 1469.9600 ;
        RECT 560.4600 1464.0400 562.0600 1464.5200 ;
        RECT 515.4600 1474.9200 517.0600 1475.4000 ;
        RECT 515.4600 1469.4800 517.0600 1469.9600 ;
        RECT 515.4600 1464.0400 517.0600 1464.5200 ;
        RECT 465.9000 1496.6800 468.9000 1497.1600 ;
        RECT 465.9000 1502.1200 468.9000 1502.6000 ;
        RECT 465.9000 1485.8000 468.9000 1486.2800 ;
        RECT 465.9000 1480.3600 468.9000 1480.8400 ;
        RECT 465.9000 1491.2400 468.9000 1491.7200 ;
        RECT 465.9000 1469.4800 468.9000 1469.9600 ;
        RECT 465.9000 1474.9200 468.9000 1475.4000 ;
        RECT 465.9000 1464.0400 468.9000 1464.5200 ;
        RECT 465.9000 1662.2300 665.0000 1665.2300 ;
        RECT 465.9000 1457.1300 665.0000 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 1227.4900 652.0600 1435.5900 ;
        RECT 605.4600 1227.4900 607.0600 1435.5900 ;
        RECT 560.4600 1227.4900 562.0600 1435.5900 ;
        RECT 515.4600 1227.4900 517.0600 1435.5900 ;
        RECT 662.0000 1227.4900 665.0000 1435.5900 ;
        RECT 465.9000 1227.4900 468.9000 1435.5900 ;
      LAYER met3 ;
        RECT 662.0000 1430.2400 665.0000 1430.7200 ;
        RECT 650.4600 1430.2400 652.0600 1430.7200 ;
        RECT 662.0000 1419.3600 665.0000 1419.8400 ;
        RECT 662.0000 1424.8000 665.0000 1425.2800 ;
        RECT 650.4600 1419.3600 652.0600 1419.8400 ;
        RECT 650.4600 1424.8000 652.0600 1425.2800 ;
        RECT 662.0000 1403.0400 665.0000 1403.5200 ;
        RECT 662.0000 1408.4800 665.0000 1408.9600 ;
        RECT 650.4600 1403.0400 652.0600 1403.5200 ;
        RECT 650.4600 1408.4800 652.0600 1408.9600 ;
        RECT 662.0000 1392.1600 665.0000 1392.6400 ;
        RECT 662.0000 1397.6000 665.0000 1398.0800 ;
        RECT 650.4600 1392.1600 652.0600 1392.6400 ;
        RECT 650.4600 1397.6000 652.0600 1398.0800 ;
        RECT 662.0000 1413.9200 665.0000 1414.4000 ;
        RECT 650.4600 1413.9200 652.0600 1414.4000 ;
        RECT 605.4600 1419.3600 607.0600 1419.8400 ;
        RECT 605.4600 1424.8000 607.0600 1425.2800 ;
        RECT 605.4600 1430.2400 607.0600 1430.7200 ;
        RECT 605.4600 1403.0400 607.0600 1403.5200 ;
        RECT 605.4600 1408.4800 607.0600 1408.9600 ;
        RECT 605.4600 1397.6000 607.0600 1398.0800 ;
        RECT 605.4600 1392.1600 607.0600 1392.6400 ;
        RECT 605.4600 1413.9200 607.0600 1414.4000 ;
        RECT 662.0000 1375.8400 665.0000 1376.3200 ;
        RECT 662.0000 1381.2800 665.0000 1381.7600 ;
        RECT 650.4600 1375.8400 652.0600 1376.3200 ;
        RECT 650.4600 1381.2800 652.0600 1381.7600 ;
        RECT 662.0000 1359.5200 665.0000 1360.0000 ;
        RECT 662.0000 1364.9600 665.0000 1365.4400 ;
        RECT 662.0000 1370.4000 665.0000 1370.8800 ;
        RECT 650.4600 1359.5200 652.0600 1360.0000 ;
        RECT 650.4600 1364.9600 652.0600 1365.4400 ;
        RECT 650.4600 1370.4000 652.0600 1370.8800 ;
        RECT 662.0000 1348.6400 665.0000 1349.1200 ;
        RECT 662.0000 1354.0800 665.0000 1354.5600 ;
        RECT 650.4600 1348.6400 652.0600 1349.1200 ;
        RECT 650.4600 1354.0800 652.0600 1354.5600 ;
        RECT 662.0000 1332.3200 665.0000 1332.8000 ;
        RECT 662.0000 1337.7600 665.0000 1338.2400 ;
        RECT 662.0000 1343.2000 665.0000 1343.6800 ;
        RECT 650.4600 1332.3200 652.0600 1332.8000 ;
        RECT 650.4600 1337.7600 652.0600 1338.2400 ;
        RECT 650.4600 1343.2000 652.0600 1343.6800 ;
        RECT 605.4600 1375.8400 607.0600 1376.3200 ;
        RECT 605.4600 1381.2800 607.0600 1381.7600 ;
        RECT 605.4600 1359.5200 607.0600 1360.0000 ;
        RECT 605.4600 1364.9600 607.0600 1365.4400 ;
        RECT 605.4600 1370.4000 607.0600 1370.8800 ;
        RECT 605.4600 1348.6400 607.0600 1349.1200 ;
        RECT 605.4600 1354.0800 607.0600 1354.5600 ;
        RECT 605.4600 1332.3200 607.0600 1332.8000 ;
        RECT 605.4600 1337.7600 607.0600 1338.2400 ;
        RECT 605.4600 1343.2000 607.0600 1343.6800 ;
        RECT 662.0000 1386.7200 665.0000 1387.2000 ;
        RECT 605.4600 1386.7200 607.0600 1387.2000 ;
        RECT 650.4600 1386.7200 652.0600 1387.2000 ;
        RECT 560.4600 1419.3600 562.0600 1419.8400 ;
        RECT 560.4600 1424.8000 562.0600 1425.2800 ;
        RECT 560.4600 1430.2400 562.0600 1430.7200 ;
        RECT 515.4600 1419.3600 517.0600 1419.8400 ;
        RECT 515.4600 1424.8000 517.0600 1425.2800 ;
        RECT 515.4600 1430.2400 517.0600 1430.7200 ;
        RECT 560.4600 1403.0400 562.0600 1403.5200 ;
        RECT 560.4600 1408.4800 562.0600 1408.9600 ;
        RECT 560.4600 1392.1600 562.0600 1392.6400 ;
        RECT 560.4600 1397.6000 562.0600 1398.0800 ;
        RECT 515.4600 1403.0400 517.0600 1403.5200 ;
        RECT 515.4600 1408.4800 517.0600 1408.9600 ;
        RECT 515.4600 1392.1600 517.0600 1392.6400 ;
        RECT 515.4600 1397.6000 517.0600 1398.0800 ;
        RECT 515.4600 1413.9200 517.0600 1414.4000 ;
        RECT 560.4600 1413.9200 562.0600 1414.4000 ;
        RECT 465.9000 1430.2400 468.9000 1430.7200 ;
        RECT 465.9000 1424.8000 468.9000 1425.2800 ;
        RECT 465.9000 1419.3600 468.9000 1419.8400 ;
        RECT 465.9000 1408.4800 468.9000 1408.9600 ;
        RECT 465.9000 1403.0400 468.9000 1403.5200 ;
        RECT 465.9000 1397.6000 468.9000 1398.0800 ;
        RECT 465.9000 1392.1600 468.9000 1392.6400 ;
        RECT 465.9000 1413.9200 468.9000 1414.4000 ;
        RECT 560.4600 1375.8400 562.0600 1376.3200 ;
        RECT 560.4600 1381.2800 562.0600 1381.7600 ;
        RECT 560.4600 1359.5200 562.0600 1360.0000 ;
        RECT 560.4600 1364.9600 562.0600 1365.4400 ;
        RECT 560.4600 1370.4000 562.0600 1370.8800 ;
        RECT 515.4600 1375.8400 517.0600 1376.3200 ;
        RECT 515.4600 1381.2800 517.0600 1381.7600 ;
        RECT 515.4600 1359.5200 517.0600 1360.0000 ;
        RECT 515.4600 1364.9600 517.0600 1365.4400 ;
        RECT 515.4600 1370.4000 517.0600 1370.8800 ;
        RECT 560.4600 1348.6400 562.0600 1349.1200 ;
        RECT 560.4600 1354.0800 562.0600 1354.5600 ;
        RECT 560.4600 1332.3200 562.0600 1332.8000 ;
        RECT 560.4600 1337.7600 562.0600 1338.2400 ;
        RECT 560.4600 1343.2000 562.0600 1343.6800 ;
        RECT 515.4600 1348.6400 517.0600 1349.1200 ;
        RECT 515.4600 1354.0800 517.0600 1354.5600 ;
        RECT 515.4600 1332.3200 517.0600 1332.8000 ;
        RECT 515.4600 1337.7600 517.0600 1338.2400 ;
        RECT 515.4600 1343.2000 517.0600 1343.6800 ;
        RECT 465.9000 1375.8400 468.9000 1376.3200 ;
        RECT 465.9000 1381.2800 468.9000 1381.7600 ;
        RECT 465.9000 1364.9600 468.9000 1365.4400 ;
        RECT 465.9000 1359.5200 468.9000 1360.0000 ;
        RECT 465.9000 1370.4000 468.9000 1370.8800 ;
        RECT 465.9000 1348.6400 468.9000 1349.1200 ;
        RECT 465.9000 1354.0800 468.9000 1354.5600 ;
        RECT 465.9000 1337.7600 468.9000 1338.2400 ;
        RECT 465.9000 1332.3200 468.9000 1332.8000 ;
        RECT 465.9000 1343.2000 468.9000 1343.6800 ;
        RECT 465.9000 1386.7200 468.9000 1387.2000 ;
        RECT 515.4600 1386.7200 517.0600 1387.2000 ;
        RECT 560.4600 1386.7200 562.0600 1387.2000 ;
        RECT 662.0000 1321.4400 665.0000 1321.9200 ;
        RECT 662.0000 1326.8800 665.0000 1327.3600 ;
        RECT 650.4600 1321.4400 652.0600 1321.9200 ;
        RECT 650.4600 1326.8800 652.0600 1327.3600 ;
        RECT 662.0000 1305.1200 665.0000 1305.6000 ;
        RECT 662.0000 1310.5600 665.0000 1311.0400 ;
        RECT 662.0000 1316.0000 665.0000 1316.4800 ;
        RECT 650.4600 1305.1200 652.0600 1305.6000 ;
        RECT 650.4600 1310.5600 652.0600 1311.0400 ;
        RECT 650.4600 1316.0000 652.0600 1316.4800 ;
        RECT 662.0000 1294.2400 665.0000 1294.7200 ;
        RECT 662.0000 1299.6800 665.0000 1300.1600 ;
        RECT 650.4600 1294.2400 652.0600 1294.7200 ;
        RECT 650.4600 1299.6800 652.0600 1300.1600 ;
        RECT 662.0000 1277.9200 665.0000 1278.4000 ;
        RECT 662.0000 1283.3600 665.0000 1283.8400 ;
        RECT 662.0000 1288.8000 665.0000 1289.2800 ;
        RECT 650.4600 1277.9200 652.0600 1278.4000 ;
        RECT 650.4600 1283.3600 652.0600 1283.8400 ;
        RECT 650.4600 1288.8000 652.0600 1289.2800 ;
        RECT 605.4600 1321.4400 607.0600 1321.9200 ;
        RECT 605.4600 1326.8800 607.0600 1327.3600 ;
        RECT 605.4600 1305.1200 607.0600 1305.6000 ;
        RECT 605.4600 1310.5600 607.0600 1311.0400 ;
        RECT 605.4600 1316.0000 607.0600 1316.4800 ;
        RECT 605.4600 1294.2400 607.0600 1294.7200 ;
        RECT 605.4600 1299.6800 607.0600 1300.1600 ;
        RECT 605.4600 1277.9200 607.0600 1278.4000 ;
        RECT 605.4600 1283.3600 607.0600 1283.8400 ;
        RECT 605.4600 1288.8000 607.0600 1289.2800 ;
        RECT 662.0000 1267.0400 665.0000 1267.5200 ;
        RECT 662.0000 1272.4800 665.0000 1272.9600 ;
        RECT 650.4600 1267.0400 652.0600 1267.5200 ;
        RECT 650.4600 1272.4800 652.0600 1272.9600 ;
        RECT 662.0000 1250.7200 665.0000 1251.2000 ;
        RECT 662.0000 1256.1600 665.0000 1256.6400 ;
        RECT 662.0000 1261.6000 665.0000 1262.0800 ;
        RECT 650.4600 1250.7200 652.0600 1251.2000 ;
        RECT 650.4600 1256.1600 652.0600 1256.6400 ;
        RECT 650.4600 1261.6000 652.0600 1262.0800 ;
        RECT 662.0000 1239.8400 665.0000 1240.3200 ;
        RECT 662.0000 1245.2800 665.0000 1245.7600 ;
        RECT 650.4600 1239.8400 652.0600 1240.3200 ;
        RECT 650.4600 1245.2800 652.0600 1245.7600 ;
        RECT 662.0000 1234.4000 665.0000 1234.8800 ;
        RECT 650.4600 1234.4000 652.0600 1234.8800 ;
        RECT 605.4600 1267.0400 607.0600 1267.5200 ;
        RECT 605.4600 1272.4800 607.0600 1272.9600 ;
        RECT 605.4600 1250.7200 607.0600 1251.2000 ;
        RECT 605.4600 1256.1600 607.0600 1256.6400 ;
        RECT 605.4600 1261.6000 607.0600 1262.0800 ;
        RECT 605.4600 1239.8400 607.0600 1240.3200 ;
        RECT 605.4600 1245.2800 607.0600 1245.7600 ;
        RECT 605.4600 1234.4000 607.0600 1234.8800 ;
        RECT 560.4600 1321.4400 562.0600 1321.9200 ;
        RECT 560.4600 1326.8800 562.0600 1327.3600 ;
        RECT 560.4600 1305.1200 562.0600 1305.6000 ;
        RECT 560.4600 1310.5600 562.0600 1311.0400 ;
        RECT 560.4600 1316.0000 562.0600 1316.4800 ;
        RECT 515.4600 1321.4400 517.0600 1321.9200 ;
        RECT 515.4600 1326.8800 517.0600 1327.3600 ;
        RECT 515.4600 1305.1200 517.0600 1305.6000 ;
        RECT 515.4600 1310.5600 517.0600 1311.0400 ;
        RECT 515.4600 1316.0000 517.0600 1316.4800 ;
        RECT 560.4600 1294.2400 562.0600 1294.7200 ;
        RECT 560.4600 1299.6800 562.0600 1300.1600 ;
        RECT 560.4600 1277.9200 562.0600 1278.4000 ;
        RECT 560.4600 1283.3600 562.0600 1283.8400 ;
        RECT 560.4600 1288.8000 562.0600 1289.2800 ;
        RECT 515.4600 1294.2400 517.0600 1294.7200 ;
        RECT 515.4600 1299.6800 517.0600 1300.1600 ;
        RECT 515.4600 1277.9200 517.0600 1278.4000 ;
        RECT 515.4600 1283.3600 517.0600 1283.8400 ;
        RECT 515.4600 1288.8000 517.0600 1289.2800 ;
        RECT 465.9000 1321.4400 468.9000 1321.9200 ;
        RECT 465.9000 1326.8800 468.9000 1327.3600 ;
        RECT 465.9000 1310.5600 468.9000 1311.0400 ;
        RECT 465.9000 1305.1200 468.9000 1305.6000 ;
        RECT 465.9000 1316.0000 468.9000 1316.4800 ;
        RECT 465.9000 1294.2400 468.9000 1294.7200 ;
        RECT 465.9000 1299.6800 468.9000 1300.1600 ;
        RECT 465.9000 1283.3600 468.9000 1283.8400 ;
        RECT 465.9000 1277.9200 468.9000 1278.4000 ;
        RECT 465.9000 1288.8000 468.9000 1289.2800 ;
        RECT 560.4600 1267.0400 562.0600 1267.5200 ;
        RECT 560.4600 1272.4800 562.0600 1272.9600 ;
        RECT 560.4600 1250.7200 562.0600 1251.2000 ;
        RECT 560.4600 1256.1600 562.0600 1256.6400 ;
        RECT 560.4600 1261.6000 562.0600 1262.0800 ;
        RECT 515.4600 1267.0400 517.0600 1267.5200 ;
        RECT 515.4600 1272.4800 517.0600 1272.9600 ;
        RECT 515.4600 1250.7200 517.0600 1251.2000 ;
        RECT 515.4600 1256.1600 517.0600 1256.6400 ;
        RECT 515.4600 1261.6000 517.0600 1262.0800 ;
        RECT 560.4600 1245.2800 562.0600 1245.7600 ;
        RECT 560.4600 1239.8400 562.0600 1240.3200 ;
        RECT 560.4600 1234.4000 562.0600 1234.8800 ;
        RECT 515.4600 1245.2800 517.0600 1245.7600 ;
        RECT 515.4600 1239.8400 517.0600 1240.3200 ;
        RECT 515.4600 1234.4000 517.0600 1234.8800 ;
        RECT 465.9000 1267.0400 468.9000 1267.5200 ;
        RECT 465.9000 1272.4800 468.9000 1272.9600 ;
        RECT 465.9000 1256.1600 468.9000 1256.6400 ;
        RECT 465.9000 1250.7200 468.9000 1251.2000 ;
        RECT 465.9000 1261.6000 468.9000 1262.0800 ;
        RECT 465.9000 1239.8400 468.9000 1240.3200 ;
        RECT 465.9000 1245.2800 468.9000 1245.7600 ;
        RECT 465.9000 1234.4000 468.9000 1234.8800 ;
        RECT 465.9000 1432.5900 665.0000 1435.5900 ;
        RECT 465.9000 1227.4900 665.0000 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 997.8500 652.0600 1205.9500 ;
        RECT 605.4600 997.8500 607.0600 1205.9500 ;
        RECT 560.4600 997.8500 562.0600 1205.9500 ;
        RECT 515.4600 997.8500 517.0600 1205.9500 ;
        RECT 662.0000 997.8500 665.0000 1205.9500 ;
        RECT 465.9000 997.8500 468.9000 1205.9500 ;
      LAYER met3 ;
        RECT 662.0000 1200.6000 665.0000 1201.0800 ;
        RECT 650.4600 1200.6000 652.0600 1201.0800 ;
        RECT 662.0000 1189.7200 665.0000 1190.2000 ;
        RECT 662.0000 1195.1600 665.0000 1195.6400 ;
        RECT 650.4600 1189.7200 652.0600 1190.2000 ;
        RECT 650.4600 1195.1600 652.0600 1195.6400 ;
        RECT 662.0000 1173.4000 665.0000 1173.8800 ;
        RECT 662.0000 1178.8400 665.0000 1179.3200 ;
        RECT 650.4600 1173.4000 652.0600 1173.8800 ;
        RECT 650.4600 1178.8400 652.0600 1179.3200 ;
        RECT 662.0000 1162.5200 665.0000 1163.0000 ;
        RECT 662.0000 1167.9600 665.0000 1168.4400 ;
        RECT 650.4600 1162.5200 652.0600 1163.0000 ;
        RECT 650.4600 1167.9600 652.0600 1168.4400 ;
        RECT 662.0000 1184.2800 665.0000 1184.7600 ;
        RECT 650.4600 1184.2800 652.0600 1184.7600 ;
        RECT 605.4600 1189.7200 607.0600 1190.2000 ;
        RECT 605.4600 1195.1600 607.0600 1195.6400 ;
        RECT 605.4600 1200.6000 607.0600 1201.0800 ;
        RECT 605.4600 1173.4000 607.0600 1173.8800 ;
        RECT 605.4600 1178.8400 607.0600 1179.3200 ;
        RECT 605.4600 1167.9600 607.0600 1168.4400 ;
        RECT 605.4600 1162.5200 607.0600 1163.0000 ;
        RECT 605.4600 1184.2800 607.0600 1184.7600 ;
        RECT 662.0000 1146.2000 665.0000 1146.6800 ;
        RECT 662.0000 1151.6400 665.0000 1152.1200 ;
        RECT 650.4600 1146.2000 652.0600 1146.6800 ;
        RECT 650.4600 1151.6400 652.0600 1152.1200 ;
        RECT 662.0000 1129.8800 665.0000 1130.3600 ;
        RECT 662.0000 1135.3200 665.0000 1135.8000 ;
        RECT 662.0000 1140.7600 665.0000 1141.2400 ;
        RECT 650.4600 1129.8800 652.0600 1130.3600 ;
        RECT 650.4600 1135.3200 652.0600 1135.8000 ;
        RECT 650.4600 1140.7600 652.0600 1141.2400 ;
        RECT 662.0000 1119.0000 665.0000 1119.4800 ;
        RECT 662.0000 1124.4400 665.0000 1124.9200 ;
        RECT 650.4600 1119.0000 652.0600 1119.4800 ;
        RECT 650.4600 1124.4400 652.0600 1124.9200 ;
        RECT 662.0000 1102.6800 665.0000 1103.1600 ;
        RECT 662.0000 1108.1200 665.0000 1108.6000 ;
        RECT 662.0000 1113.5600 665.0000 1114.0400 ;
        RECT 650.4600 1102.6800 652.0600 1103.1600 ;
        RECT 650.4600 1108.1200 652.0600 1108.6000 ;
        RECT 650.4600 1113.5600 652.0600 1114.0400 ;
        RECT 605.4600 1146.2000 607.0600 1146.6800 ;
        RECT 605.4600 1151.6400 607.0600 1152.1200 ;
        RECT 605.4600 1129.8800 607.0600 1130.3600 ;
        RECT 605.4600 1135.3200 607.0600 1135.8000 ;
        RECT 605.4600 1140.7600 607.0600 1141.2400 ;
        RECT 605.4600 1119.0000 607.0600 1119.4800 ;
        RECT 605.4600 1124.4400 607.0600 1124.9200 ;
        RECT 605.4600 1102.6800 607.0600 1103.1600 ;
        RECT 605.4600 1108.1200 607.0600 1108.6000 ;
        RECT 605.4600 1113.5600 607.0600 1114.0400 ;
        RECT 662.0000 1157.0800 665.0000 1157.5600 ;
        RECT 605.4600 1157.0800 607.0600 1157.5600 ;
        RECT 650.4600 1157.0800 652.0600 1157.5600 ;
        RECT 560.4600 1189.7200 562.0600 1190.2000 ;
        RECT 560.4600 1195.1600 562.0600 1195.6400 ;
        RECT 560.4600 1200.6000 562.0600 1201.0800 ;
        RECT 515.4600 1189.7200 517.0600 1190.2000 ;
        RECT 515.4600 1195.1600 517.0600 1195.6400 ;
        RECT 515.4600 1200.6000 517.0600 1201.0800 ;
        RECT 560.4600 1173.4000 562.0600 1173.8800 ;
        RECT 560.4600 1178.8400 562.0600 1179.3200 ;
        RECT 560.4600 1162.5200 562.0600 1163.0000 ;
        RECT 560.4600 1167.9600 562.0600 1168.4400 ;
        RECT 515.4600 1173.4000 517.0600 1173.8800 ;
        RECT 515.4600 1178.8400 517.0600 1179.3200 ;
        RECT 515.4600 1162.5200 517.0600 1163.0000 ;
        RECT 515.4600 1167.9600 517.0600 1168.4400 ;
        RECT 515.4600 1184.2800 517.0600 1184.7600 ;
        RECT 560.4600 1184.2800 562.0600 1184.7600 ;
        RECT 465.9000 1200.6000 468.9000 1201.0800 ;
        RECT 465.9000 1195.1600 468.9000 1195.6400 ;
        RECT 465.9000 1189.7200 468.9000 1190.2000 ;
        RECT 465.9000 1178.8400 468.9000 1179.3200 ;
        RECT 465.9000 1173.4000 468.9000 1173.8800 ;
        RECT 465.9000 1167.9600 468.9000 1168.4400 ;
        RECT 465.9000 1162.5200 468.9000 1163.0000 ;
        RECT 465.9000 1184.2800 468.9000 1184.7600 ;
        RECT 560.4600 1146.2000 562.0600 1146.6800 ;
        RECT 560.4600 1151.6400 562.0600 1152.1200 ;
        RECT 560.4600 1129.8800 562.0600 1130.3600 ;
        RECT 560.4600 1135.3200 562.0600 1135.8000 ;
        RECT 560.4600 1140.7600 562.0600 1141.2400 ;
        RECT 515.4600 1146.2000 517.0600 1146.6800 ;
        RECT 515.4600 1151.6400 517.0600 1152.1200 ;
        RECT 515.4600 1129.8800 517.0600 1130.3600 ;
        RECT 515.4600 1135.3200 517.0600 1135.8000 ;
        RECT 515.4600 1140.7600 517.0600 1141.2400 ;
        RECT 560.4600 1119.0000 562.0600 1119.4800 ;
        RECT 560.4600 1124.4400 562.0600 1124.9200 ;
        RECT 560.4600 1102.6800 562.0600 1103.1600 ;
        RECT 560.4600 1108.1200 562.0600 1108.6000 ;
        RECT 560.4600 1113.5600 562.0600 1114.0400 ;
        RECT 515.4600 1119.0000 517.0600 1119.4800 ;
        RECT 515.4600 1124.4400 517.0600 1124.9200 ;
        RECT 515.4600 1102.6800 517.0600 1103.1600 ;
        RECT 515.4600 1108.1200 517.0600 1108.6000 ;
        RECT 515.4600 1113.5600 517.0600 1114.0400 ;
        RECT 465.9000 1146.2000 468.9000 1146.6800 ;
        RECT 465.9000 1151.6400 468.9000 1152.1200 ;
        RECT 465.9000 1135.3200 468.9000 1135.8000 ;
        RECT 465.9000 1129.8800 468.9000 1130.3600 ;
        RECT 465.9000 1140.7600 468.9000 1141.2400 ;
        RECT 465.9000 1119.0000 468.9000 1119.4800 ;
        RECT 465.9000 1124.4400 468.9000 1124.9200 ;
        RECT 465.9000 1108.1200 468.9000 1108.6000 ;
        RECT 465.9000 1102.6800 468.9000 1103.1600 ;
        RECT 465.9000 1113.5600 468.9000 1114.0400 ;
        RECT 465.9000 1157.0800 468.9000 1157.5600 ;
        RECT 515.4600 1157.0800 517.0600 1157.5600 ;
        RECT 560.4600 1157.0800 562.0600 1157.5600 ;
        RECT 662.0000 1091.8000 665.0000 1092.2800 ;
        RECT 662.0000 1097.2400 665.0000 1097.7200 ;
        RECT 650.4600 1091.8000 652.0600 1092.2800 ;
        RECT 650.4600 1097.2400 652.0600 1097.7200 ;
        RECT 662.0000 1075.4800 665.0000 1075.9600 ;
        RECT 662.0000 1080.9200 665.0000 1081.4000 ;
        RECT 662.0000 1086.3600 665.0000 1086.8400 ;
        RECT 650.4600 1075.4800 652.0600 1075.9600 ;
        RECT 650.4600 1080.9200 652.0600 1081.4000 ;
        RECT 650.4600 1086.3600 652.0600 1086.8400 ;
        RECT 662.0000 1064.6000 665.0000 1065.0800 ;
        RECT 662.0000 1070.0400 665.0000 1070.5200 ;
        RECT 650.4600 1064.6000 652.0600 1065.0800 ;
        RECT 650.4600 1070.0400 652.0600 1070.5200 ;
        RECT 662.0000 1048.2800 665.0000 1048.7600 ;
        RECT 662.0000 1053.7200 665.0000 1054.2000 ;
        RECT 662.0000 1059.1600 665.0000 1059.6400 ;
        RECT 650.4600 1048.2800 652.0600 1048.7600 ;
        RECT 650.4600 1053.7200 652.0600 1054.2000 ;
        RECT 650.4600 1059.1600 652.0600 1059.6400 ;
        RECT 605.4600 1091.8000 607.0600 1092.2800 ;
        RECT 605.4600 1097.2400 607.0600 1097.7200 ;
        RECT 605.4600 1075.4800 607.0600 1075.9600 ;
        RECT 605.4600 1080.9200 607.0600 1081.4000 ;
        RECT 605.4600 1086.3600 607.0600 1086.8400 ;
        RECT 605.4600 1064.6000 607.0600 1065.0800 ;
        RECT 605.4600 1070.0400 607.0600 1070.5200 ;
        RECT 605.4600 1048.2800 607.0600 1048.7600 ;
        RECT 605.4600 1053.7200 607.0600 1054.2000 ;
        RECT 605.4600 1059.1600 607.0600 1059.6400 ;
        RECT 662.0000 1037.4000 665.0000 1037.8800 ;
        RECT 662.0000 1042.8400 665.0000 1043.3200 ;
        RECT 650.4600 1037.4000 652.0600 1037.8800 ;
        RECT 650.4600 1042.8400 652.0600 1043.3200 ;
        RECT 662.0000 1021.0800 665.0000 1021.5600 ;
        RECT 662.0000 1026.5200 665.0000 1027.0000 ;
        RECT 662.0000 1031.9600 665.0000 1032.4400 ;
        RECT 650.4600 1021.0800 652.0600 1021.5600 ;
        RECT 650.4600 1026.5200 652.0600 1027.0000 ;
        RECT 650.4600 1031.9600 652.0600 1032.4400 ;
        RECT 662.0000 1010.2000 665.0000 1010.6800 ;
        RECT 662.0000 1015.6400 665.0000 1016.1200 ;
        RECT 650.4600 1010.2000 652.0600 1010.6800 ;
        RECT 650.4600 1015.6400 652.0600 1016.1200 ;
        RECT 662.0000 1004.7600 665.0000 1005.2400 ;
        RECT 650.4600 1004.7600 652.0600 1005.2400 ;
        RECT 605.4600 1037.4000 607.0600 1037.8800 ;
        RECT 605.4600 1042.8400 607.0600 1043.3200 ;
        RECT 605.4600 1021.0800 607.0600 1021.5600 ;
        RECT 605.4600 1026.5200 607.0600 1027.0000 ;
        RECT 605.4600 1031.9600 607.0600 1032.4400 ;
        RECT 605.4600 1010.2000 607.0600 1010.6800 ;
        RECT 605.4600 1015.6400 607.0600 1016.1200 ;
        RECT 605.4600 1004.7600 607.0600 1005.2400 ;
        RECT 560.4600 1091.8000 562.0600 1092.2800 ;
        RECT 560.4600 1097.2400 562.0600 1097.7200 ;
        RECT 560.4600 1075.4800 562.0600 1075.9600 ;
        RECT 560.4600 1080.9200 562.0600 1081.4000 ;
        RECT 560.4600 1086.3600 562.0600 1086.8400 ;
        RECT 515.4600 1091.8000 517.0600 1092.2800 ;
        RECT 515.4600 1097.2400 517.0600 1097.7200 ;
        RECT 515.4600 1075.4800 517.0600 1075.9600 ;
        RECT 515.4600 1080.9200 517.0600 1081.4000 ;
        RECT 515.4600 1086.3600 517.0600 1086.8400 ;
        RECT 560.4600 1064.6000 562.0600 1065.0800 ;
        RECT 560.4600 1070.0400 562.0600 1070.5200 ;
        RECT 560.4600 1048.2800 562.0600 1048.7600 ;
        RECT 560.4600 1053.7200 562.0600 1054.2000 ;
        RECT 560.4600 1059.1600 562.0600 1059.6400 ;
        RECT 515.4600 1064.6000 517.0600 1065.0800 ;
        RECT 515.4600 1070.0400 517.0600 1070.5200 ;
        RECT 515.4600 1048.2800 517.0600 1048.7600 ;
        RECT 515.4600 1053.7200 517.0600 1054.2000 ;
        RECT 515.4600 1059.1600 517.0600 1059.6400 ;
        RECT 465.9000 1091.8000 468.9000 1092.2800 ;
        RECT 465.9000 1097.2400 468.9000 1097.7200 ;
        RECT 465.9000 1080.9200 468.9000 1081.4000 ;
        RECT 465.9000 1075.4800 468.9000 1075.9600 ;
        RECT 465.9000 1086.3600 468.9000 1086.8400 ;
        RECT 465.9000 1064.6000 468.9000 1065.0800 ;
        RECT 465.9000 1070.0400 468.9000 1070.5200 ;
        RECT 465.9000 1053.7200 468.9000 1054.2000 ;
        RECT 465.9000 1048.2800 468.9000 1048.7600 ;
        RECT 465.9000 1059.1600 468.9000 1059.6400 ;
        RECT 560.4600 1037.4000 562.0600 1037.8800 ;
        RECT 560.4600 1042.8400 562.0600 1043.3200 ;
        RECT 560.4600 1021.0800 562.0600 1021.5600 ;
        RECT 560.4600 1026.5200 562.0600 1027.0000 ;
        RECT 560.4600 1031.9600 562.0600 1032.4400 ;
        RECT 515.4600 1037.4000 517.0600 1037.8800 ;
        RECT 515.4600 1042.8400 517.0600 1043.3200 ;
        RECT 515.4600 1021.0800 517.0600 1021.5600 ;
        RECT 515.4600 1026.5200 517.0600 1027.0000 ;
        RECT 515.4600 1031.9600 517.0600 1032.4400 ;
        RECT 560.4600 1015.6400 562.0600 1016.1200 ;
        RECT 560.4600 1010.2000 562.0600 1010.6800 ;
        RECT 560.4600 1004.7600 562.0600 1005.2400 ;
        RECT 515.4600 1015.6400 517.0600 1016.1200 ;
        RECT 515.4600 1010.2000 517.0600 1010.6800 ;
        RECT 515.4600 1004.7600 517.0600 1005.2400 ;
        RECT 465.9000 1037.4000 468.9000 1037.8800 ;
        RECT 465.9000 1042.8400 468.9000 1043.3200 ;
        RECT 465.9000 1026.5200 468.9000 1027.0000 ;
        RECT 465.9000 1021.0800 468.9000 1021.5600 ;
        RECT 465.9000 1031.9600 468.9000 1032.4400 ;
        RECT 465.9000 1010.2000 468.9000 1010.6800 ;
        RECT 465.9000 1015.6400 468.9000 1016.1200 ;
        RECT 465.9000 1004.7600 468.9000 1005.2400 ;
        RECT 465.9000 1202.9500 665.0000 1205.9500 ;
        RECT 465.9000 997.8500 665.0000 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 650.4600 768.2100 652.0600 976.3100 ;
        RECT 605.4600 768.2100 607.0600 976.3100 ;
        RECT 560.4600 768.2100 562.0600 976.3100 ;
        RECT 515.4600 768.2100 517.0600 976.3100 ;
        RECT 662.0000 768.2100 665.0000 976.3100 ;
        RECT 465.9000 768.2100 468.9000 976.3100 ;
      LAYER met3 ;
        RECT 662.0000 970.9600 665.0000 971.4400 ;
        RECT 650.4600 970.9600 652.0600 971.4400 ;
        RECT 662.0000 960.0800 665.0000 960.5600 ;
        RECT 662.0000 965.5200 665.0000 966.0000 ;
        RECT 650.4600 960.0800 652.0600 960.5600 ;
        RECT 650.4600 965.5200 652.0600 966.0000 ;
        RECT 662.0000 943.7600 665.0000 944.2400 ;
        RECT 662.0000 949.2000 665.0000 949.6800 ;
        RECT 650.4600 943.7600 652.0600 944.2400 ;
        RECT 650.4600 949.2000 652.0600 949.6800 ;
        RECT 662.0000 932.8800 665.0000 933.3600 ;
        RECT 662.0000 938.3200 665.0000 938.8000 ;
        RECT 650.4600 932.8800 652.0600 933.3600 ;
        RECT 650.4600 938.3200 652.0600 938.8000 ;
        RECT 662.0000 954.6400 665.0000 955.1200 ;
        RECT 650.4600 954.6400 652.0600 955.1200 ;
        RECT 605.4600 960.0800 607.0600 960.5600 ;
        RECT 605.4600 965.5200 607.0600 966.0000 ;
        RECT 605.4600 970.9600 607.0600 971.4400 ;
        RECT 605.4600 943.7600 607.0600 944.2400 ;
        RECT 605.4600 949.2000 607.0600 949.6800 ;
        RECT 605.4600 938.3200 607.0600 938.8000 ;
        RECT 605.4600 932.8800 607.0600 933.3600 ;
        RECT 605.4600 954.6400 607.0600 955.1200 ;
        RECT 662.0000 916.5600 665.0000 917.0400 ;
        RECT 662.0000 922.0000 665.0000 922.4800 ;
        RECT 650.4600 916.5600 652.0600 917.0400 ;
        RECT 650.4600 922.0000 652.0600 922.4800 ;
        RECT 662.0000 900.2400 665.0000 900.7200 ;
        RECT 662.0000 905.6800 665.0000 906.1600 ;
        RECT 662.0000 911.1200 665.0000 911.6000 ;
        RECT 650.4600 900.2400 652.0600 900.7200 ;
        RECT 650.4600 905.6800 652.0600 906.1600 ;
        RECT 650.4600 911.1200 652.0600 911.6000 ;
        RECT 662.0000 889.3600 665.0000 889.8400 ;
        RECT 662.0000 894.8000 665.0000 895.2800 ;
        RECT 650.4600 889.3600 652.0600 889.8400 ;
        RECT 650.4600 894.8000 652.0600 895.2800 ;
        RECT 662.0000 873.0400 665.0000 873.5200 ;
        RECT 662.0000 878.4800 665.0000 878.9600 ;
        RECT 662.0000 883.9200 665.0000 884.4000 ;
        RECT 650.4600 873.0400 652.0600 873.5200 ;
        RECT 650.4600 878.4800 652.0600 878.9600 ;
        RECT 650.4600 883.9200 652.0600 884.4000 ;
        RECT 605.4600 916.5600 607.0600 917.0400 ;
        RECT 605.4600 922.0000 607.0600 922.4800 ;
        RECT 605.4600 900.2400 607.0600 900.7200 ;
        RECT 605.4600 905.6800 607.0600 906.1600 ;
        RECT 605.4600 911.1200 607.0600 911.6000 ;
        RECT 605.4600 889.3600 607.0600 889.8400 ;
        RECT 605.4600 894.8000 607.0600 895.2800 ;
        RECT 605.4600 873.0400 607.0600 873.5200 ;
        RECT 605.4600 878.4800 607.0600 878.9600 ;
        RECT 605.4600 883.9200 607.0600 884.4000 ;
        RECT 662.0000 927.4400 665.0000 927.9200 ;
        RECT 605.4600 927.4400 607.0600 927.9200 ;
        RECT 650.4600 927.4400 652.0600 927.9200 ;
        RECT 560.4600 960.0800 562.0600 960.5600 ;
        RECT 560.4600 965.5200 562.0600 966.0000 ;
        RECT 560.4600 970.9600 562.0600 971.4400 ;
        RECT 515.4600 960.0800 517.0600 960.5600 ;
        RECT 515.4600 965.5200 517.0600 966.0000 ;
        RECT 515.4600 970.9600 517.0600 971.4400 ;
        RECT 560.4600 943.7600 562.0600 944.2400 ;
        RECT 560.4600 949.2000 562.0600 949.6800 ;
        RECT 560.4600 932.8800 562.0600 933.3600 ;
        RECT 560.4600 938.3200 562.0600 938.8000 ;
        RECT 515.4600 943.7600 517.0600 944.2400 ;
        RECT 515.4600 949.2000 517.0600 949.6800 ;
        RECT 515.4600 932.8800 517.0600 933.3600 ;
        RECT 515.4600 938.3200 517.0600 938.8000 ;
        RECT 515.4600 954.6400 517.0600 955.1200 ;
        RECT 560.4600 954.6400 562.0600 955.1200 ;
        RECT 465.9000 970.9600 468.9000 971.4400 ;
        RECT 465.9000 965.5200 468.9000 966.0000 ;
        RECT 465.9000 960.0800 468.9000 960.5600 ;
        RECT 465.9000 949.2000 468.9000 949.6800 ;
        RECT 465.9000 943.7600 468.9000 944.2400 ;
        RECT 465.9000 938.3200 468.9000 938.8000 ;
        RECT 465.9000 932.8800 468.9000 933.3600 ;
        RECT 465.9000 954.6400 468.9000 955.1200 ;
        RECT 560.4600 916.5600 562.0600 917.0400 ;
        RECT 560.4600 922.0000 562.0600 922.4800 ;
        RECT 560.4600 900.2400 562.0600 900.7200 ;
        RECT 560.4600 905.6800 562.0600 906.1600 ;
        RECT 560.4600 911.1200 562.0600 911.6000 ;
        RECT 515.4600 916.5600 517.0600 917.0400 ;
        RECT 515.4600 922.0000 517.0600 922.4800 ;
        RECT 515.4600 900.2400 517.0600 900.7200 ;
        RECT 515.4600 905.6800 517.0600 906.1600 ;
        RECT 515.4600 911.1200 517.0600 911.6000 ;
        RECT 560.4600 889.3600 562.0600 889.8400 ;
        RECT 560.4600 894.8000 562.0600 895.2800 ;
        RECT 560.4600 873.0400 562.0600 873.5200 ;
        RECT 560.4600 878.4800 562.0600 878.9600 ;
        RECT 560.4600 883.9200 562.0600 884.4000 ;
        RECT 515.4600 889.3600 517.0600 889.8400 ;
        RECT 515.4600 894.8000 517.0600 895.2800 ;
        RECT 515.4600 873.0400 517.0600 873.5200 ;
        RECT 515.4600 878.4800 517.0600 878.9600 ;
        RECT 515.4600 883.9200 517.0600 884.4000 ;
        RECT 465.9000 916.5600 468.9000 917.0400 ;
        RECT 465.9000 922.0000 468.9000 922.4800 ;
        RECT 465.9000 905.6800 468.9000 906.1600 ;
        RECT 465.9000 900.2400 468.9000 900.7200 ;
        RECT 465.9000 911.1200 468.9000 911.6000 ;
        RECT 465.9000 889.3600 468.9000 889.8400 ;
        RECT 465.9000 894.8000 468.9000 895.2800 ;
        RECT 465.9000 878.4800 468.9000 878.9600 ;
        RECT 465.9000 873.0400 468.9000 873.5200 ;
        RECT 465.9000 883.9200 468.9000 884.4000 ;
        RECT 465.9000 927.4400 468.9000 927.9200 ;
        RECT 515.4600 927.4400 517.0600 927.9200 ;
        RECT 560.4600 927.4400 562.0600 927.9200 ;
        RECT 662.0000 862.1600 665.0000 862.6400 ;
        RECT 662.0000 867.6000 665.0000 868.0800 ;
        RECT 650.4600 862.1600 652.0600 862.6400 ;
        RECT 650.4600 867.6000 652.0600 868.0800 ;
        RECT 662.0000 845.8400 665.0000 846.3200 ;
        RECT 662.0000 851.2800 665.0000 851.7600 ;
        RECT 662.0000 856.7200 665.0000 857.2000 ;
        RECT 650.4600 845.8400 652.0600 846.3200 ;
        RECT 650.4600 851.2800 652.0600 851.7600 ;
        RECT 650.4600 856.7200 652.0600 857.2000 ;
        RECT 662.0000 834.9600 665.0000 835.4400 ;
        RECT 662.0000 840.4000 665.0000 840.8800 ;
        RECT 650.4600 834.9600 652.0600 835.4400 ;
        RECT 650.4600 840.4000 652.0600 840.8800 ;
        RECT 662.0000 818.6400 665.0000 819.1200 ;
        RECT 662.0000 824.0800 665.0000 824.5600 ;
        RECT 662.0000 829.5200 665.0000 830.0000 ;
        RECT 650.4600 818.6400 652.0600 819.1200 ;
        RECT 650.4600 824.0800 652.0600 824.5600 ;
        RECT 650.4600 829.5200 652.0600 830.0000 ;
        RECT 605.4600 862.1600 607.0600 862.6400 ;
        RECT 605.4600 867.6000 607.0600 868.0800 ;
        RECT 605.4600 845.8400 607.0600 846.3200 ;
        RECT 605.4600 851.2800 607.0600 851.7600 ;
        RECT 605.4600 856.7200 607.0600 857.2000 ;
        RECT 605.4600 834.9600 607.0600 835.4400 ;
        RECT 605.4600 840.4000 607.0600 840.8800 ;
        RECT 605.4600 818.6400 607.0600 819.1200 ;
        RECT 605.4600 824.0800 607.0600 824.5600 ;
        RECT 605.4600 829.5200 607.0600 830.0000 ;
        RECT 662.0000 807.7600 665.0000 808.2400 ;
        RECT 662.0000 813.2000 665.0000 813.6800 ;
        RECT 650.4600 807.7600 652.0600 808.2400 ;
        RECT 650.4600 813.2000 652.0600 813.6800 ;
        RECT 662.0000 791.4400 665.0000 791.9200 ;
        RECT 662.0000 796.8800 665.0000 797.3600 ;
        RECT 662.0000 802.3200 665.0000 802.8000 ;
        RECT 650.4600 791.4400 652.0600 791.9200 ;
        RECT 650.4600 796.8800 652.0600 797.3600 ;
        RECT 650.4600 802.3200 652.0600 802.8000 ;
        RECT 662.0000 780.5600 665.0000 781.0400 ;
        RECT 662.0000 786.0000 665.0000 786.4800 ;
        RECT 650.4600 780.5600 652.0600 781.0400 ;
        RECT 650.4600 786.0000 652.0600 786.4800 ;
        RECT 662.0000 775.1200 665.0000 775.6000 ;
        RECT 650.4600 775.1200 652.0600 775.6000 ;
        RECT 605.4600 807.7600 607.0600 808.2400 ;
        RECT 605.4600 813.2000 607.0600 813.6800 ;
        RECT 605.4600 791.4400 607.0600 791.9200 ;
        RECT 605.4600 796.8800 607.0600 797.3600 ;
        RECT 605.4600 802.3200 607.0600 802.8000 ;
        RECT 605.4600 780.5600 607.0600 781.0400 ;
        RECT 605.4600 786.0000 607.0600 786.4800 ;
        RECT 605.4600 775.1200 607.0600 775.6000 ;
        RECT 560.4600 862.1600 562.0600 862.6400 ;
        RECT 560.4600 867.6000 562.0600 868.0800 ;
        RECT 560.4600 845.8400 562.0600 846.3200 ;
        RECT 560.4600 851.2800 562.0600 851.7600 ;
        RECT 560.4600 856.7200 562.0600 857.2000 ;
        RECT 515.4600 862.1600 517.0600 862.6400 ;
        RECT 515.4600 867.6000 517.0600 868.0800 ;
        RECT 515.4600 845.8400 517.0600 846.3200 ;
        RECT 515.4600 851.2800 517.0600 851.7600 ;
        RECT 515.4600 856.7200 517.0600 857.2000 ;
        RECT 560.4600 834.9600 562.0600 835.4400 ;
        RECT 560.4600 840.4000 562.0600 840.8800 ;
        RECT 560.4600 818.6400 562.0600 819.1200 ;
        RECT 560.4600 824.0800 562.0600 824.5600 ;
        RECT 560.4600 829.5200 562.0600 830.0000 ;
        RECT 515.4600 834.9600 517.0600 835.4400 ;
        RECT 515.4600 840.4000 517.0600 840.8800 ;
        RECT 515.4600 818.6400 517.0600 819.1200 ;
        RECT 515.4600 824.0800 517.0600 824.5600 ;
        RECT 515.4600 829.5200 517.0600 830.0000 ;
        RECT 465.9000 862.1600 468.9000 862.6400 ;
        RECT 465.9000 867.6000 468.9000 868.0800 ;
        RECT 465.9000 851.2800 468.9000 851.7600 ;
        RECT 465.9000 845.8400 468.9000 846.3200 ;
        RECT 465.9000 856.7200 468.9000 857.2000 ;
        RECT 465.9000 834.9600 468.9000 835.4400 ;
        RECT 465.9000 840.4000 468.9000 840.8800 ;
        RECT 465.9000 824.0800 468.9000 824.5600 ;
        RECT 465.9000 818.6400 468.9000 819.1200 ;
        RECT 465.9000 829.5200 468.9000 830.0000 ;
        RECT 560.4600 807.7600 562.0600 808.2400 ;
        RECT 560.4600 813.2000 562.0600 813.6800 ;
        RECT 560.4600 791.4400 562.0600 791.9200 ;
        RECT 560.4600 796.8800 562.0600 797.3600 ;
        RECT 560.4600 802.3200 562.0600 802.8000 ;
        RECT 515.4600 807.7600 517.0600 808.2400 ;
        RECT 515.4600 813.2000 517.0600 813.6800 ;
        RECT 515.4600 791.4400 517.0600 791.9200 ;
        RECT 515.4600 796.8800 517.0600 797.3600 ;
        RECT 515.4600 802.3200 517.0600 802.8000 ;
        RECT 560.4600 786.0000 562.0600 786.4800 ;
        RECT 560.4600 780.5600 562.0600 781.0400 ;
        RECT 560.4600 775.1200 562.0600 775.6000 ;
        RECT 515.4600 786.0000 517.0600 786.4800 ;
        RECT 515.4600 780.5600 517.0600 781.0400 ;
        RECT 515.4600 775.1200 517.0600 775.6000 ;
        RECT 465.9000 807.7600 468.9000 808.2400 ;
        RECT 465.9000 813.2000 468.9000 813.6800 ;
        RECT 465.9000 796.8800 468.9000 797.3600 ;
        RECT 465.9000 791.4400 468.9000 791.9200 ;
        RECT 465.9000 802.3200 468.9000 802.8000 ;
        RECT 465.9000 780.5600 468.9000 781.0400 ;
        RECT 465.9000 786.0000 468.9000 786.4800 ;
        RECT 465.9000 775.1200 468.9000 775.6000 ;
        RECT 465.9000 973.3100 665.0000 976.3100 ;
        RECT 465.9000 768.2100 665.0000 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 686.1200 2833.6100 688.1200 2854.5400 ;
        RECT 883.2200 2833.6100 885.2200 2854.5400 ;
      LAYER met3 ;
        RECT 883.2200 2850.0400 885.2200 2850.5200 ;
        RECT 686.1200 2850.0400 688.1200 2850.5200 ;
        RECT 883.2200 2839.1600 885.2200 2839.6400 ;
        RECT 686.1200 2839.1600 688.1200 2839.6400 ;
        RECT 883.2200 2844.6000 885.2200 2845.0800 ;
        RECT 686.1200 2844.6000 688.1200 2845.0800 ;
        RECT 686.1200 2852.5400 885.2200 2854.5400 ;
        RECT 686.1200 2833.6100 885.2200 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 538.5700 872.2800 746.6700 ;
        RECT 825.6800 538.5700 827.2800 746.6700 ;
        RECT 780.6800 538.5700 782.2800 746.6700 ;
        RECT 735.6800 538.5700 737.2800 746.6700 ;
        RECT 882.2200 538.5700 885.2200 746.6700 ;
        RECT 686.1200 538.5700 689.1200 746.6700 ;
      LAYER met3 ;
        RECT 882.2200 741.3200 885.2200 741.8000 ;
        RECT 870.6800 741.3200 872.2800 741.8000 ;
        RECT 882.2200 730.4400 885.2200 730.9200 ;
        RECT 882.2200 735.8800 885.2200 736.3600 ;
        RECT 870.6800 730.4400 872.2800 730.9200 ;
        RECT 870.6800 735.8800 872.2800 736.3600 ;
        RECT 882.2200 714.1200 885.2200 714.6000 ;
        RECT 882.2200 719.5600 885.2200 720.0400 ;
        RECT 870.6800 714.1200 872.2800 714.6000 ;
        RECT 870.6800 719.5600 872.2800 720.0400 ;
        RECT 882.2200 703.2400 885.2200 703.7200 ;
        RECT 882.2200 708.6800 885.2200 709.1600 ;
        RECT 870.6800 703.2400 872.2800 703.7200 ;
        RECT 870.6800 708.6800 872.2800 709.1600 ;
        RECT 882.2200 725.0000 885.2200 725.4800 ;
        RECT 870.6800 725.0000 872.2800 725.4800 ;
        RECT 825.6800 730.4400 827.2800 730.9200 ;
        RECT 825.6800 735.8800 827.2800 736.3600 ;
        RECT 825.6800 741.3200 827.2800 741.8000 ;
        RECT 825.6800 714.1200 827.2800 714.6000 ;
        RECT 825.6800 719.5600 827.2800 720.0400 ;
        RECT 825.6800 708.6800 827.2800 709.1600 ;
        RECT 825.6800 703.2400 827.2800 703.7200 ;
        RECT 825.6800 725.0000 827.2800 725.4800 ;
        RECT 882.2200 686.9200 885.2200 687.4000 ;
        RECT 882.2200 692.3600 885.2200 692.8400 ;
        RECT 870.6800 686.9200 872.2800 687.4000 ;
        RECT 870.6800 692.3600 872.2800 692.8400 ;
        RECT 882.2200 670.6000 885.2200 671.0800 ;
        RECT 882.2200 676.0400 885.2200 676.5200 ;
        RECT 882.2200 681.4800 885.2200 681.9600 ;
        RECT 870.6800 670.6000 872.2800 671.0800 ;
        RECT 870.6800 676.0400 872.2800 676.5200 ;
        RECT 870.6800 681.4800 872.2800 681.9600 ;
        RECT 882.2200 659.7200 885.2200 660.2000 ;
        RECT 882.2200 665.1600 885.2200 665.6400 ;
        RECT 870.6800 659.7200 872.2800 660.2000 ;
        RECT 870.6800 665.1600 872.2800 665.6400 ;
        RECT 882.2200 643.4000 885.2200 643.8800 ;
        RECT 882.2200 648.8400 885.2200 649.3200 ;
        RECT 882.2200 654.2800 885.2200 654.7600 ;
        RECT 870.6800 643.4000 872.2800 643.8800 ;
        RECT 870.6800 648.8400 872.2800 649.3200 ;
        RECT 870.6800 654.2800 872.2800 654.7600 ;
        RECT 825.6800 686.9200 827.2800 687.4000 ;
        RECT 825.6800 692.3600 827.2800 692.8400 ;
        RECT 825.6800 670.6000 827.2800 671.0800 ;
        RECT 825.6800 676.0400 827.2800 676.5200 ;
        RECT 825.6800 681.4800 827.2800 681.9600 ;
        RECT 825.6800 659.7200 827.2800 660.2000 ;
        RECT 825.6800 665.1600 827.2800 665.6400 ;
        RECT 825.6800 643.4000 827.2800 643.8800 ;
        RECT 825.6800 648.8400 827.2800 649.3200 ;
        RECT 825.6800 654.2800 827.2800 654.7600 ;
        RECT 882.2200 697.8000 885.2200 698.2800 ;
        RECT 825.6800 697.8000 827.2800 698.2800 ;
        RECT 870.6800 697.8000 872.2800 698.2800 ;
        RECT 780.6800 730.4400 782.2800 730.9200 ;
        RECT 780.6800 735.8800 782.2800 736.3600 ;
        RECT 780.6800 741.3200 782.2800 741.8000 ;
        RECT 735.6800 730.4400 737.2800 730.9200 ;
        RECT 735.6800 735.8800 737.2800 736.3600 ;
        RECT 735.6800 741.3200 737.2800 741.8000 ;
        RECT 780.6800 714.1200 782.2800 714.6000 ;
        RECT 780.6800 719.5600 782.2800 720.0400 ;
        RECT 780.6800 703.2400 782.2800 703.7200 ;
        RECT 780.6800 708.6800 782.2800 709.1600 ;
        RECT 735.6800 714.1200 737.2800 714.6000 ;
        RECT 735.6800 719.5600 737.2800 720.0400 ;
        RECT 735.6800 703.2400 737.2800 703.7200 ;
        RECT 735.6800 708.6800 737.2800 709.1600 ;
        RECT 735.6800 725.0000 737.2800 725.4800 ;
        RECT 780.6800 725.0000 782.2800 725.4800 ;
        RECT 686.1200 741.3200 689.1200 741.8000 ;
        RECT 686.1200 735.8800 689.1200 736.3600 ;
        RECT 686.1200 730.4400 689.1200 730.9200 ;
        RECT 686.1200 719.5600 689.1200 720.0400 ;
        RECT 686.1200 714.1200 689.1200 714.6000 ;
        RECT 686.1200 708.6800 689.1200 709.1600 ;
        RECT 686.1200 703.2400 689.1200 703.7200 ;
        RECT 686.1200 725.0000 689.1200 725.4800 ;
        RECT 780.6800 686.9200 782.2800 687.4000 ;
        RECT 780.6800 692.3600 782.2800 692.8400 ;
        RECT 780.6800 670.6000 782.2800 671.0800 ;
        RECT 780.6800 676.0400 782.2800 676.5200 ;
        RECT 780.6800 681.4800 782.2800 681.9600 ;
        RECT 735.6800 686.9200 737.2800 687.4000 ;
        RECT 735.6800 692.3600 737.2800 692.8400 ;
        RECT 735.6800 670.6000 737.2800 671.0800 ;
        RECT 735.6800 676.0400 737.2800 676.5200 ;
        RECT 735.6800 681.4800 737.2800 681.9600 ;
        RECT 780.6800 659.7200 782.2800 660.2000 ;
        RECT 780.6800 665.1600 782.2800 665.6400 ;
        RECT 780.6800 643.4000 782.2800 643.8800 ;
        RECT 780.6800 648.8400 782.2800 649.3200 ;
        RECT 780.6800 654.2800 782.2800 654.7600 ;
        RECT 735.6800 659.7200 737.2800 660.2000 ;
        RECT 735.6800 665.1600 737.2800 665.6400 ;
        RECT 735.6800 643.4000 737.2800 643.8800 ;
        RECT 735.6800 648.8400 737.2800 649.3200 ;
        RECT 735.6800 654.2800 737.2800 654.7600 ;
        RECT 686.1200 686.9200 689.1200 687.4000 ;
        RECT 686.1200 692.3600 689.1200 692.8400 ;
        RECT 686.1200 676.0400 689.1200 676.5200 ;
        RECT 686.1200 670.6000 689.1200 671.0800 ;
        RECT 686.1200 681.4800 689.1200 681.9600 ;
        RECT 686.1200 659.7200 689.1200 660.2000 ;
        RECT 686.1200 665.1600 689.1200 665.6400 ;
        RECT 686.1200 648.8400 689.1200 649.3200 ;
        RECT 686.1200 643.4000 689.1200 643.8800 ;
        RECT 686.1200 654.2800 689.1200 654.7600 ;
        RECT 686.1200 697.8000 689.1200 698.2800 ;
        RECT 735.6800 697.8000 737.2800 698.2800 ;
        RECT 780.6800 697.8000 782.2800 698.2800 ;
        RECT 882.2200 632.5200 885.2200 633.0000 ;
        RECT 882.2200 637.9600 885.2200 638.4400 ;
        RECT 870.6800 632.5200 872.2800 633.0000 ;
        RECT 870.6800 637.9600 872.2800 638.4400 ;
        RECT 882.2200 616.2000 885.2200 616.6800 ;
        RECT 882.2200 621.6400 885.2200 622.1200 ;
        RECT 882.2200 627.0800 885.2200 627.5600 ;
        RECT 870.6800 616.2000 872.2800 616.6800 ;
        RECT 870.6800 621.6400 872.2800 622.1200 ;
        RECT 870.6800 627.0800 872.2800 627.5600 ;
        RECT 882.2200 605.3200 885.2200 605.8000 ;
        RECT 882.2200 610.7600 885.2200 611.2400 ;
        RECT 870.6800 605.3200 872.2800 605.8000 ;
        RECT 870.6800 610.7600 872.2800 611.2400 ;
        RECT 882.2200 589.0000 885.2200 589.4800 ;
        RECT 882.2200 594.4400 885.2200 594.9200 ;
        RECT 882.2200 599.8800 885.2200 600.3600 ;
        RECT 870.6800 589.0000 872.2800 589.4800 ;
        RECT 870.6800 594.4400 872.2800 594.9200 ;
        RECT 870.6800 599.8800 872.2800 600.3600 ;
        RECT 825.6800 632.5200 827.2800 633.0000 ;
        RECT 825.6800 637.9600 827.2800 638.4400 ;
        RECT 825.6800 616.2000 827.2800 616.6800 ;
        RECT 825.6800 621.6400 827.2800 622.1200 ;
        RECT 825.6800 627.0800 827.2800 627.5600 ;
        RECT 825.6800 605.3200 827.2800 605.8000 ;
        RECT 825.6800 610.7600 827.2800 611.2400 ;
        RECT 825.6800 589.0000 827.2800 589.4800 ;
        RECT 825.6800 594.4400 827.2800 594.9200 ;
        RECT 825.6800 599.8800 827.2800 600.3600 ;
        RECT 882.2200 578.1200 885.2200 578.6000 ;
        RECT 882.2200 583.5600 885.2200 584.0400 ;
        RECT 870.6800 578.1200 872.2800 578.6000 ;
        RECT 870.6800 583.5600 872.2800 584.0400 ;
        RECT 882.2200 561.8000 885.2200 562.2800 ;
        RECT 882.2200 567.2400 885.2200 567.7200 ;
        RECT 882.2200 572.6800 885.2200 573.1600 ;
        RECT 870.6800 561.8000 872.2800 562.2800 ;
        RECT 870.6800 567.2400 872.2800 567.7200 ;
        RECT 870.6800 572.6800 872.2800 573.1600 ;
        RECT 882.2200 550.9200 885.2200 551.4000 ;
        RECT 882.2200 556.3600 885.2200 556.8400 ;
        RECT 870.6800 550.9200 872.2800 551.4000 ;
        RECT 870.6800 556.3600 872.2800 556.8400 ;
        RECT 882.2200 545.4800 885.2200 545.9600 ;
        RECT 870.6800 545.4800 872.2800 545.9600 ;
        RECT 825.6800 578.1200 827.2800 578.6000 ;
        RECT 825.6800 583.5600 827.2800 584.0400 ;
        RECT 825.6800 561.8000 827.2800 562.2800 ;
        RECT 825.6800 567.2400 827.2800 567.7200 ;
        RECT 825.6800 572.6800 827.2800 573.1600 ;
        RECT 825.6800 550.9200 827.2800 551.4000 ;
        RECT 825.6800 556.3600 827.2800 556.8400 ;
        RECT 825.6800 545.4800 827.2800 545.9600 ;
        RECT 780.6800 632.5200 782.2800 633.0000 ;
        RECT 780.6800 637.9600 782.2800 638.4400 ;
        RECT 780.6800 616.2000 782.2800 616.6800 ;
        RECT 780.6800 621.6400 782.2800 622.1200 ;
        RECT 780.6800 627.0800 782.2800 627.5600 ;
        RECT 735.6800 632.5200 737.2800 633.0000 ;
        RECT 735.6800 637.9600 737.2800 638.4400 ;
        RECT 735.6800 616.2000 737.2800 616.6800 ;
        RECT 735.6800 621.6400 737.2800 622.1200 ;
        RECT 735.6800 627.0800 737.2800 627.5600 ;
        RECT 780.6800 605.3200 782.2800 605.8000 ;
        RECT 780.6800 610.7600 782.2800 611.2400 ;
        RECT 780.6800 589.0000 782.2800 589.4800 ;
        RECT 780.6800 594.4400 782.2800 594.9200 ;
        RECT 780.6800 599.8800 782.2800 600.3600 ;
        RECT 735.6800 605.3200 737.2800 605.8000 ;
        RECT 735.6800 610.7600 737.2800 611.2400 ;
        RECT 735.6800 589.0000 737.2800 589.4800 ;
        RECT 735.6800 594.4400 737.2800 594.9200 ;
        RECT 735.6800 599.8800 737.2800 600.3600 ;
        RECT 686.1200 632.5200 689.1200 633.0000 ;
        RECT 686.1200 637.9600 689.1200 638.4400 ;
        RECT 686.1200 621.6400 689.1200 622.1200 ;
        RECT 686.1200 616.2000 689.1200 616.6800 ;
        RECT 686.1200 627.0800 689.1200 627.5600 ;
        RECT 686.1200 605.3200 689.1200 605.8000 ;
        RECT 686.1200 610.7600 689.1200 611.2400 ;
        RECT 686.1200 594.4400 689.1200 594.9200 ;
        RECT 686.1200 589.0000 689.1200 589.4800 ;
        RECT 686.1200 599.8800 689.1200 600.3600 ;
        RECT 780.6800 578.1200 782.2800 578.6000 ;
        RECT 780.6800 583.5600 782.2800 584.0400 ;
        RECT 780.6800 561.8000 782.2800 562.2800 ;
        RECT 780.6800 567.2400 782.2800 567.7200 ;
        RECT 780.6800 572.6800 782.2800 573.1600 ;
        RECT 735.6800 578.1200 737.2800 578.6000 ;
        RECT 735.6800 583.5600 737.2800 584.0400 ;
        RECT 735.6800 561.8000 737.2800 562.2800 ;
        RECT 735.6800 567.2400 737.2800 567.7200 ;
        RECT 735.6800 572.6800 737.2800 573.1600 ;
        RECT 780.6800 556.3600 782.2800 556.8400 ;
        RECT 780.6800 550.9200 782.2800 551.4000 ;
        RECT 780.6800 545.4800 782.2800 545.9600 ;
        RECT 735.6800 556.3600 737.2800 556.8400 ;
        RECT 735.6800 550.9200 737.2800 551.4000 ;
        RECT 735.6800 545.4800 737.2800 545.9600 ;
        RECT 686.1200 578.1200 689.1200 578.6000 ;
        RECT 686.1200 583.5600 689.1200 584.0400 ;
        RECT 686.1200 567.2400 689.1200 567.7200 ;
        RECT 686.1200 561.8000 689.1200 562.2800 ;
        RECT 686.1200 572.6800 689.1200 573.1600 ;
        RECT 686.1200 550.9200 689.1200 551.4000 ;
        RECT 686.1200 556.3600 689.1200 556.8400 ;
        RECT 686.1200 545.4800 689.1200 545.9600 ;
        RECT 686.1200 743.6700 885.2200 746.6700 ;
        RECT 686.1200 538.5700 885.2200 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 308.9300 872.2800 517.0300 ;
        RECT 825.6800 308.9300 827.2800 517.0300 ;
        RECT 780.6800 308.9300 782.2800 517.0300 ;
        RECT 735.6800 308.9300 737.2800 517.0300 ;
        RECT 882.2200 308.9300 885.2200 517.0300 ;
        RECT 686.1200 308.9300 689.1200 517.0300 ;
      LAYER met3 ;
        RECT 882.2200 511.6800 885.2200 512.1600 ;
        RECT 870.6800 511.6800 872.2800 512.1600 ;
        RECT 882.2200 500.8000 885.2200 501.2800 ;
        RECT 882.2200 506.2400 885.2200 506.7200 ;
        RECT 870.6800 500.8000 872.2800 501.2800 ;
        RECT 870.6800 506.2400 872.2800 506.7200 ;
        RECT 882.2200 484.4800 885.2200 484.9600 ;
        RECT 882.2200 489.9200 885.2200 490.4000 ;
        RECT 870.6800 484.4800 872.2800 484.9600 ;
        RECT 870.6800 489.9200 872.2800 490.4000 ;
        RECT 882.2200 473.6000 885.2200 474.0800 ;
        RECT 882.2200 479.0400 885.2200 479.5200 ;
        RECT 870.6800 473.6000 872.2800 474.0800 ;
        RECT 870.6800 479.0400 872.2800 479.5200 ;
        RECT 882.2200 495.3600 885.2200 495.8400 ;
        RECT 870.6800 495.3600 872.2800 495.8400 ;
        RECT 825.6800 500.8000 827.2800 501.2800 ;
        RECT 825.6800 506.2400 827.2800 506.7200 ;
        RECT 825.6800 511.6800 827.2800 512.1600 ;
        RECT 825.6800 484.4800 827.2800 484.9600 ;
        RECT 825.6800 489.9200 827.2800 490.4000 ;
        RECT 825.6800 479.0400 827.2800 479.5200 ;
        RECT 825.6800 473.6000 827.2800 474.0800 ;
        RECT 825.6800 495.3600 827.2800 495.8400 ;
        RECT 882.2200 457.2800 885.2200 457.7600 ;
        RECT 882.2200 462.7200 885.2200 463.2000 ;
        RECT 870.6800 457.2800 872.2800 457.7600 ;
        RECT 870.6800 462.7200 872.2800 463.2000 ;
        RECT 882.2200 440.9600 885.2200 441.4400 ;
        RECT 882.2200 446.4000 885.2200 446.8800 ;
        RECT 882.2200 451.8400 885.2200 452.3200 ;
        RECT 870.6800 440.9600 872.2800 441.4400 ;
        RECT 870.6800 446.4000 872.2800 446.8800 ;
        RECT 870.6800 451.8400 872.2800 452.3200 ;
        RECT 882.2200 430.0800 885.2200 430.5600 ;
        RECT 882.2200 435.5200 885.2200 436.0000 ;
        RECT 870.6800 430.0800 872.2800 430.5600 ;
        RECT 870.6800 435.5200 872.2800 436.0000 ;
        RECT 882.2200 413.7600 885.2200 414.2400 ;
        RECT 882.2200 419.2000 885.2200 419.6800 ;
        RECT 882.2200 424.6400 885.2200 425.1200 ;
        RECT 870.6800 413.7600 872.2800 414.2400 ;
        RECT 870.6800 419.2000 872.2800 419.6800 ;
        RECT 870.6800 424.6400 872.2800 425.1200 ;
        RECT 825.6800 457.2800 827.2800 457.7600 ;
        RECT 825.6800 462.7200 827.2800 463.2000 ;
        RECT 825.6800 440.9600 827.2800 441.4400 ;
        RECT 825.6800 446.4000 827.2800 446.8800 ;
        RECT 825.6800 451.8400 827.2800 452.3200 ;
        RECT 825.6800 430.0800 827.2800 430.5600 ;
        RECT 825.6800 435.5200 827.2800 436.0000 ;
        RECT 825.6800 413.7600 827.2800 414.2400 ;
        RECT 825.6800 419.2000 827.2800 419.6800 ;
        RECT 825.6800 424.6400 827.2800 425.1200 ;
        RECT 882.2200 468.1600 885.2200 468.6400 ;
        RECT 825.6800 468.1600 827.2800 468.6400 ;
        RECT 870.6800 468.1600 872.2800 468.6400 ;
        RECT 780.6800 500.8000 782.2800 501.2800 ;
        RECT 780.6800 506.2400 782.2800 506.7200 ;
        RECT 780.6800 511.6800 782.2800 512.1600 ;
        RECT 735.6800 500.8000 737.2800 501.2800 ;
        RECT 735.6800 506.2400 737.2800 506.7200 ;
        RECT 735.6800 511.6800 737.2800 512.1600 ;
        RECT 780.6800 484.4800 782.2800 484.9600 ;
        RECT 780.6800 489.9200 782.2800 490.4000 ;
        RECT 780.6800 473.6000 782.2800 474.0800 ;
        RECT 780.6800 479.0400 782.2800 479.5200 ;
        RECT 735.6800 484.4800 737.2800 484.9600 ;
        RECT 735.6800 489.9200 737.2800 490.4000 ;
        RECT 735.6800 473.6000 737.2800 474.0800 ;
        RECT 735.6800 479.0400 737.2800 479.5200 ;
        RECT 735.6800 495.3600 737.2800 495.8400 ;
        RECT 780.6800 495.3600 782.2800 495.8400 ;
        RECT 686.1200 511.6800 689.1200 512.1600 ;
        RECT 686.1200 506.2400 689.1200 506.7200 ;
        RECT 686.1200 500.8000 689.1200 501.2800 ;
        RECT 686.1200 489.9200 689.1200 490.4000 ;
        RECT 686.1200 484.4800 689.1200 484.9600 ;
        RECT 686.1200 479.0400 689.1200 479.5200 ;
        RECT 686.1200 473.6000 689.1200 474.0800 ;
        RECT 686.1200 495.3600 689.1200 495.8400 ;
        RECT 780.6800 457.2800 782.2800 457.7600 ;
        RECT 780.6800 462.7200 782.2800 463.2000 ;
        RECT 780.6800 440.9600 782.2800 441.4400 ;
        RECT 780.6800 446.4000 782.2800 446.8800 ;
        RECT 780.6800 451.8400 782.2800 452.3200 ;
        RECT 735.6800 457.2800 737.2800 457.7600 ;
        RECT 735.6800 462.7200 737.2800 463.2000 ;
        RECT 735.6800 440.9600 737.2800 441.4400 ;
        RECT 735.6800 446.4000 737.2800 446.8800 ;
        RECT 735.6800 451.8400 737.2800 452.3200 ;
        RECT 780.6800 430.0800 782.2800 430.5600 ;
        RECT 780.6800 435.5200 782.2800 436.0000 ;
        RECT 780.6800 413.7600 782.2800 414.2400 ;
        RECT 780.6800 419.2000 782.2800 419.6800 ;
        RECT 780.6800 424.6400 782.2800 425.1200 ;
        RECT 735.6800 430.0800 737.2800 430.5600 ;
        RECT 735.6800 435.5200 737.2800 436.0000 ;
        RECT 735.6800 413.7600 737.2800 414.2400 ;
        RECT 735.6800 419.2000 737.2800 419.6800 ;
        RECT 735.6800 424.6400 737.2800 425.1200 ;
        RECT 686.1200 457.2800 689.1200 457.7600 ;
        RECT 686.1200 462.7200 689.1200 463.2000 ;
        RECT 686.1200 446.4000 689.1200 446.8800 ;
        RECT 686.1200 440.9600 689.1200 441.4400 ;
        RECT 686.1200 451.8400 689.1200 452.3200 ;
        RECT 686.1200 430.0800 689.1200 430.5600 ;
        RECT 686.1200 435.5200 689.1200 436.0000 ;
        RECT 686.1200 419.2000 689.1200 419.6800 ;
        RECT 686.1200 413.7600 689.1200 414.2400 ;
        RECT 686.1200 424.6400 689.1200 425.1200 ;
        RECT 686.1200 468.1600 689.1200 468.6400 ;
        RECT 735.6800 468.1600 737.2800 468.6400 ;
        RECT 780.6800 468.1600 782.2800 468.6400 ;
        RECT 882.2200 402.8800 885.2200 403.3600 ;
        RECT 882.2200 408.3200 885.2200 408.8000 ;
        RECT 870.6800 402.8800 872.2800 403.3600 ;
        RECT 870.6800 408.3200 872.2800 408.8000 ;
        RECT 882.2200 386.5600 885.2200 387.0400 ;
        RECT 882.2200 392.0000 885.2200 392.4800 ;
        RECT 882.2200 397.4400 885.2200 397.9200 ;
        RECT 870.6800 386.5600 872.2800 387.0400 ;
        RECT 870.6800 392.0000 872.2800 392.4800 ;
        RECT 870.6800 397.4400 872.2800 397.9200 ;
        RECT 882.2200 375.6800 885.2200 376.1600 ;
        RECT 882.2200 381.1200 885.2200 381.6000 ;
        RECT 870.6800 375.6800 872.2800 376.1600 ;
        RECT 870.6800 381.1200 872.2800 381.6000 ;
        RECT 882.2200 359.3600 885.2200 359.8400 ;
        RECT 882.2200 364.8000 885.2200 365.2800 ;
        RECT 882.2200 370.2400 885.2200 370.7200 ;
        RECT 870.6800 359.3600 872.2800 359.8400 ;
        RECT 870.6800 364.8000 872.2800 365.2800 ;
        RECT 870.6800 370.2400 872.2800 370.7200 ;
        RECT 825.6800 402.8800 827.2800 403.3600 ;
        RECT 825.6800 408.3200 827.2800 408.8000 ;
        RECT 825.6800 386.5600 827.2800 387.0400 ;
        RECT 825.6800 392.0000 827.2800 392.4800 ;
        RECT 825.6800 397.4400 827.2800 397.9200 ;
        RECT 825.6800 375.6800 827.2800 376.1600 ;
        RECT 825.6800 381.1200 827.2800 381.6000 ;
        RECT 825.6800 359.3600 827.2800 359.8400 ;
        RECT 825.6800 364.8000 827.2800 365.2800 ;
        RECT 825.6800 370.2400 827.2800 370.7200 ;
        RECT 882.2200 348.4800 885.2200 348.9600 ;
        RECT 882.2200 353.9200 885.2200 354.4000 ;
        RECT 870.6800 348.4800 872.2800 348.9600 ;
        RECT 870.6800 353.9200 872.2800 354.4000 ;
        RECT 882.2200 332.1600 885.2200 332.6400 ;
        RECT 882.2200 337.6000 885.2200 338.0800 ;
        RECT 882.2200 343.0400 885.2200 343.5200 ;
        RECT 870.6800 332.1600 872.2800 332.6400 ;
        RECT 870.6800 337.6000 872.2800 338.0800 ;
        RECT 870.6800 343.0400 872.2800 343.5200 ;
        RECT 882.2200 321.2800 885.2200 321.7600 ;
        RECT 882.2200 326.7200 885.2200 327.2000 ;
        RECT 870.6800 321.2800 872.2800 321.7600 ;
        RECT 870.6800 326.7200 872.2800 327.2000 ;
        RECT 882.2200 315.8400 885.2200 316.3200 ;
        RECT 870.6800 315.8400 872.2800 316.3200 ;
        RECT 825.6800 348.4800 827.2800 348.9600 ;
        RECT 825.6800 353.9200 827.2800 354.4000 ;
        RECT 825.6800 332.1600 827.2800 332.6400 ;
        RECT 825.6800 337.6000 827.2800 338.0800 ;
        RECT 825.6800 343.0400 827.2800 343.5200 ;
        RECT 825.6800 321.2800 827.2800 321.7600 ;
        RECT 825.6800 326.7200 827.2800 327.2000 ;
        RECT 825.6800 315.8400 827.2800 316.3200 ;
        RECT 780.6800 402.8800 782.2800 403.3600 ;
        RECT 780.6800 408.3200 782.2800 408.8000 ;
        RECT 780.6800 386.5600 782.2800 387.0400 ;
        RECT 780.6800 392.0000 782.2800 392.4800 ;
        RECT 780.6800 397.4400 782.2800 397.9200 ;
        RECT 735.6800 402.8800 737.2800 403.3600 ;
        RECT 735.6800 408.3200 737.2800 408.8000 ;
        RECT 735.6800 386.5600 737.2800 387.0400 ;
        RECT 735.6800 392.0000 737.2800 392.4800 ;
        RECT 735.6800 397.4400 737.2800 397.9200 ;
        RECT 780.6800 375.6800 782.2800 376.1600 ;
        RECT 780.6800 381.1200 782.2800 381.6000 ;
        RECT 780.6800 359.3600 782.2800 359.8400 ;
        RECT 780.6800 364.8000 782.2800 365.2800 ;
        RECT 780.6800 370.2400 782.2800 370.7200 ;
        RECT 735.6800 375.6800 737.2800 376.1600 ;
        RECT 735.6800 381.1200 737.2800 381.6000 ;
        RECT 735.6800 359.3600 737.2800 359.8400 ;
        RECT 735.6800 364.8000 737.2800 365.2800 ;
        RECT 735.6800 370.2400 737.2800 370.7200 ;
        RECT 686.1200 402.8800 689.1200 403.3600 ;
        RECT 686.1200 408.3200 689.1200 408.8000 ;
        RECT 686.1200 392.0000 689.1200 392.4800 ;
        RECT 686.1200 386.5600 689.1200 387.0400 ;
        RECT 686.1200 397.4400 689.1200 397.9200 ;
        RECT 686.1200 375.6800 689.1200 376.1600 ;
        RECT 686.1200 381.1200 689.1200 381.6000 ;
        RECT 686.1200 364.8000 689.1200 365.2800 ;
        RECT 686.1200 359.3600 689.1200 359.8400 ;
        RECT 686.1200 370.2400 689.1200 370.7200 ;
        RECT 780.6800 348.4800 782.2800 348.9600 ;
        RECT 780.6800 353.9200 782.2800 354.4000 ;
        RECT 780.6800 332.1600 782.2800 332.6400 ;
        RECT 780.6800 337.6000 782.2800 338.0800 ;
        RECT 780.6800 343.0400 782.2800 343.5200 ;
        RECT 735.6800 348.4800 737.2800 348.9600 ;
        RECT 735.6800 353.9200 737.2800 354.4000 ;
        RECT 735.6800 332.1600 737.2800 332.6400 ;
        RECT 735.6800 337.6000 737.2800 338.0800 ;
        RECT 735.6800 343.0400 737.2800 343.5200 ;
        RECT 780.6800 326.7200 782.2800 327.2000 ;
        RECT 780.6800 321.2800 782.2800 321.7600 ;
        RECT 780.6800 315.8400 782.2800 316.3200 ;
        RECT 735.6800 326.7200 737.2800 327.2000 ;
        RECT 735.6800 321.2800 737.2800 321.7600 ;
        RECT 735.6800 315.8400 737.2800 316.3200 ;
        RECT 686.1200 348.4800 689.1200 348.9600 ;
        RECT 686.1200 353.9200 689.1200 354.4000 ;
        RECT 686.1200 337.6000 689.1200 338.0800 ;
        RECT 686.1200 332.1600 689.1200 332.6400 ;
        RECT 686.1200 343.0400 689.1200 343.5200 ;
        RECT 686.1200 321.2800 689.1200 321.7600 ;
        RECT 686.1200 326.7200 689.1200 327.2000 ;
        RECT 686.1200 315.8400 689.1200 316.3200 ;
        RECT 686.1200 514.0300 885.2200 517.0300 ;
        RECT 686.1200 308.9300 885.2200 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 79.2900 872.2800 287.3900 ;
        RECT 825.6800 79.2900 827.2800 287.3900 ;
        RECT 780.6800 79.2900 782.2800 287.3900 ;
        RECT 735.6800 79.2900 737.2800 287.3900 ;
        RECT 882.2200 79.2900 885.2200 287.3900 ;
        RECT 686.1200 79.2900 689.1200 287.3900 ;
      LAYER met3 ;
        RECT 882.2200 282.0400 885.2200 282.5200 ;
        RECT 870.6800 282.0400 872.2800 282.5200 ;
        RECT 882.2200 271.1600 885.2200 271.6400 ;
        RECT 882.2200 276.6000 885.2200 277.0800 ;
        RECT 870.6800 271.1600 872.2800 271.6400 ;
        RECT 870.6800 276.6000 872.2800 277.0800 ;
        RECT 882.2200 254.8400 885.2200 255.3200 ;
        RECT 882.2200 260.2800 885.2200 260.7600 ;
        RECT 870.6800 254.8400 872.2800 255.3200 ;
        RECT 870.6800 260.2800 872.2800 260.7600 ;
        RECT 882.2200 243.9600 885.2200 244.4400 ;
        RECT 882.2200 249.4000 885.2200 249.8800 ;
        RECT 870.6800 243.9600 872.2800 244.4400 ;
        RECT 870.6800 249.4000 872.2800 249.8800 ;
        RECT 882.2200 265.7200 885.2200 266.2000 ;
        RECT 870.6800 265.7200 872.2800 266.2000 ;
        RECT 825.6800 271.1600 827.2800 271.6400 ;
        RECT 825.6800 276.6000 827.2800 277.0800 ;
        RECT 825.6800 282.0400 827.2800 282.5200 ;
        RECT 825.6800 254.8400 827.2800 255.3200 ;
        RECT 825.6800 260.2800 827.2800 260.7600 ;
        RECT 825.6800 249.4000 827.2800 249.8800 ;
        RECT 825.6800 243.9600 827.2800 244.4400 ;
        RECT 825.6800 265.7200 827.2800 266.2000 ;
        RECT 882.2200 227.6400 885.2200 228.1200 ;
        RECT 882.2200 233.0800 885.2200 233.5600 ;
        RECT 870.6800 227.6400 872.2800 228.1200 ;
        RECT 870.6800 233.0800 872.2800 233.5600 ;
        RECT 882.2200 211.3200 885.2200 211.8000 ;
        RECT 882.2200 216.7600 885.2200 217.2400 ;
        RECT 882.2200 222.2000 885.2200 222.6800 ;
        RECT 870.6800 211.3200 872.2800 211.8000 ;
        RECT 870.6800 216.7600 872.2800 217.2400 ;
        RECT 870.6800 222.2000 872.2800 222.6800 ;
        RECT 882.2200 200.4400 885.2200 200.9200 ;
        RECT 882.2200 205.8800 885.2200 206.3600 ;
        RECT 870.6800 200.4400 872.2800 200.9200 ;
        RECT 870.6800 205.8800 872.2800 206.3600 ;
        RECT 882.2200 184.1200 885.2200 184.6000 ;
        RECT 882.2200 189.5600 885.2200 190.0400 ;
        RECT 882.2200 195.0000 885.2200 195.4800 ;
        RECT 870.6800 184.1200 872.2800 184.6000 ;
        RECT 870.6800 189.5600 872.2800 190.0400 ;
        RECT 870.6800 195.0000 872.2800 195.4800 ;
        RECT 825.6800 227.6400 827.2800 228.1200 ;
        RECT 825.6800 233.0800 827.2800 233.5600 ;
        RECT 825.6800 211.3200 827.2800 211.8000 ;
        RECT 825.6800 216.7600 827.2800 217.2400 ;
        RECT 825.6800 222.2000 827.2800 222.6800 ;
        RECT 825.6800 200.4400 827.2800 200.9200 ;
        RECT 825.6800 205.8800 827.2800 206.3600 ;
        RECT 825.6800 184.1200 827.2800 184.6000 ;
        RECT 825.6800 189.5600 827.2800 190.0400 ;
        RECT 825.6800 195.0000 827.2800 195.4800 ;
        RECT 882.2200 238.5200 885.2200 239.0000 ;
        RECT 825.6800 238.5200 827.2800 239.0000 ;
        RECT 870.6800 238.5200 872.2800 239.0000 ;
        RECT 780.6800 271.1600 782.2800 271.6400 ;
        RECT 780.6800 276.6000 782.2800 277.0800 ;
        RECT 780.6800 282.0400 782.2800 282.5200 ;
        RECT 735.6800 271.1600 737.2800 271.6400 ;
        RECT 735.6800 276.6000 737.2800 277.0800 ;
        RECT 735.6800 282.0400 737.2800 282.5200 ;
        RECT 780.6800 254.8400 782.2800 255.3200 ;
        RECT 780.6800 260.2800 782.2800 260.7600 ;
        RECT 780.6800 243.9600 782.2800 244.4400 ;
        RECT 780.6800 249.4000 782.2800 249.8800 ;
        RECT 735.6800 254.8400 737.2800 255.3200 ;
        RECT 735.6800 260.2800 737.2800 260.7600 ;
        RECT 735.6800 243.9600 737.2800 244.4400 ;
        RECT 735.6800 249.4000 737.2800 249.8800 ;
        RECT 735.6800 265.7200 737.2800 266.2000 ;
        RECT 780.6800 265.7200 782.2800 266.2000 ;
        RECT 686.1200 282.0400 689.1200 282.5200 ;
        RECT 686.1200 276.6000 689.1200 277.0800 ;
        RECT 686.1200 271.1600 689.1200 271.6400 ;
        RECT 686.1200 260.2800 689.1200 260.7600 ;
        RECT 686.1200 254.8400 689.1200 255.3200 ;
        RECT 686.1200 249.4000 689.1200 249.8800 ;
        RECT 686.1200 243.9600 689.1200 244.4400 ;
        RECT 686.1200 265.7200 689.1200 266.2000 ;
        RECT 780.6800 227.6400 782.2800 228.1200 ;
        RECT 780.6800 233.0800 782.2800 233.5600 ;
        RECT 780.6800 211.3200 782.2800 211.8000 ;
        RECT 780.6800 216.7600 782.2800 217.2400 ;
        RECT 780.6800 222.2000 782.2800 222.6800 ;
        RECT 735.6800 227.6400 737.2800 228.1200 ;
        RECT 735.6800 233.0800 737.2800 233.5600 ;
        RECT 735.6800 211.3200 737.2800 211.8000 ;
        RECT 735.6800 216.7600 737.2800 217.2400 ;
        RECT 735.6800 222.2000 737.2800 222.6800 ;
        RECT 780.6800 200.4400 782.2800 200.9200 ;
        RECT 780.6800 205.8800 782.2800 206.3600 ;
        RECT 780.6800 184.1200 782.2800 184.6000 ;
        RECT 780.6800 189.5600 782.2800 190.0400 ;
        RECT 780.6800 195.0000 782.2800 195.4800 ;
        RECT 735.6800 200.4400 737.2800 200.9200 ;
        RECT 735.6800 205.8800 737.2800 206.3600 ;
        RECT 735.6800 184.1200 737.2800 184.6000 ;
        RECT 735.6800 189.5600 737.2800 190.0400 ;
        RECT 735.6800 195.0000 737.2800 195.4800 ;
        RECT 686.1200 227.6400 689.1200 228.1200 ;
        RECT 686.1200 233.0800 689.1200 233.5600 ;
        RECT 686.1200 216.7600 689.1200 217.2400 ;
        RECT 686.1200 211.3200 689.1200 211.8000 ;
        RECT 686.1200 222.2000 689.1200 222.6800 ;
        RECT 686.1200 200.4400 689.1200 200.9200 ;
        RECT 686.1200 205.8800 689.1200 206.3600 ;
        RECT 686.1200 189.5600 689.1200 190.0400 ;
        RECT 686.1200 184.1200 689.1200 184.6000 ;
        RECT 686.1200 195.0000 689.1200 195.4800 ;
        RECT 686.1200 238.5200 689.1200 239.0000 ;
        RECT 735.6800 238.5200 737.2800 239.0000 ;
        RECT 780.6800 238.5200 782.2800 239.0000 ;
        RECT 882.2200 173.2400 885.2200 173.7200 ;
        RECT 882.2200 178.6800 885.2200 179.1600 ;
        RECT 870.6800 173.2400 872.2800 173.7200 ;
        RECT 870.6800 178.6800 872.2800 179.1600 ;
        RECT 882.2200 156.9200 885.2200 157.4000 ;
        RECT 882.2200 162.3600 885.2200 162.8400 ;
        RECT 882.2200 167.8000 885.2200 168.2800 ;
        RECT 870.6800 156.9200 872.2800 157.4000 ;
        RECT 870.6800 162.3600 872.2800 162.8400 ;
        RECT 870.6800 167.8000 872.2800 168.2800 ;
        RECT 882.2200 146.0400 885.2200 146.5200 ;
        RECT 882.2200 151.4800 885.2200 151.9600 ;
        RECT 870.6800 146.0400 872.2800 146.5200 ;
        RECT 870.6800 151.4800 872.2800 151.9600 ;
        RECT 882.2200 129.7200 885.2200 130.2000 ;
        RECT 882.2200 135.1600 885.2200 135.6400 ;
        RECT 882.2200 140.6000 885.2200 141.0800 ;
        RECT 870.6800 129.7200 872.2800 130.2000 ;
        RECT 870.6800 135.1600 872.2800 135.6400 ;
        RECT 870.6800 140.6000 872.2800 141.0800 ;
        RECT 825.6800 173.2400 827.2800 173.7200 ;
        RECT 825.6800 178.6800 827.2800 179.1600 ;
        RECT 825.6800 156.9200 827.2800 157.4000 ;
        RECT 825.6800 162.3600 827.2800 162.8400 ;
        RECT 825.6800 167.8000 827.2800 168.2800 ;
        RECT 825.6800 146.0400 827.2800 146.5200 ;
        RECT 825.6800 151.4800 827.2800 151.9600 ;
        RECT 825.6800 129.7200 827.2800 130.2000 ;
        RECT 825.6800 135.1600 827.2800 135.6400 ;
        RECT 825.6800 140.6000 827.2800 141.0800 ;
        RECT 882.2200 118.8400 885.2200 119.3200 ;
        RECT 882.2200 124.2800 885.2200 124.7600 ;
        RECT 870.6800 118.8400 872.2800 119.3200 ;
        RECT 870.6800 124.2800 872.2800 124.7600 ;
        RECT 882.2200 102.5200 885.2200 103.0000 ;
        RECT 882.2200 107.9600 885.2200 108.4400 ;
        RECT 882.2200 113.4000 885.2200 113.8800 ;
        RECT 870.6800 102.5200 872.2800 103.0000 ;
        RECT 870.6800 107.9600 872.2800 108.4400 ;
        RECT 870.6800 113.4000 872.2800 113.8800 ;
        RECT 882.2200 91.6400 885.2200 92.1200 ;
        RECT 882.2200 97.0800 885.2200 97.5600 ;
        RECT 870.6800 91.6400 872.2800 92.1200 ;
        RECT 870.6800 97.0800 872.2800 97.5600 ;
        RECT 882.2200 86.2000 885.2200 86.6800 ;
        RECT 870.6800 86.2000 872.2800 86.6800 ;
        RECT 825.6800 118.8400 827.2800 119.3200 ;
        RECT 825.6800 124.2800 827.2800 124.7600 ;
        RECT 825.6800 102.5200 827.2800 103.0000 ;
        RECT 825.6800 107.9600 827.2800 108.4400 ;
        RECT 825.6800 113.4000 827.2800 113.8800 ;
        RECT 825.6800 91.6400 827.2800 92.1200 ;
        RECT 825.6800 97.0800 827.2800 97.5600 ;
        RECT 825.6800 86.2000 827.2800 86.6800 ;
        RECT 780.6800 173.2400 782.2800 173.7200 ;
        RECT 780.6800 178.6800 782.2800 179.1600 ;
        RECT 780.6800 156.9200 782.2800 157.4000 ;
        RECT 780.6800 162.3600 782.2800 162.8400 ;
        RECT 780.6800 167.8000 782.2800 168.2800 ;
        RECT 735.6800 173.2400 737.2800 173.7200 ;
        RECT 735.6800 178.6800 737.2800 179.1600 ;
        RECT 735.6800 156.9200 737.2800 157.4000 ;
        RECT 735.6800 162.3600 737.2800 162.8400 ;
        RECT 735.6800 167.8000 737.2800 168.2800 ;
        RECT 780.6800 146.0400 782.2800 146.5200 ;
        RECT 780.6800 151.4800 782.2800 151.9600 ;
        RECT 780.6800 129.7200 782.2800 130.2000 ;
        RECT 780.6800 135.1600 782.2800 135.6400 ;
        RECT 780.6800 140.6000 782.2800 141.0800 ;
        RECT 735.6800 146.0400 737.2800 146.5200 ;
        RECT 735.6800 151.4800 737.2800 151.9600 ;
        RECT 735.6800 129.7200 737.2800 130.2000 ;
        RECT 735.6800 135.1600 737.2800 135.6400 ;
        RECT 735.6800 140.6000 737.2800 141.0800 ;
        RECT 686.1200 173.2400 689.1200 173.7200 ;
        RECT 686.1200 178.6800 689.1200 179.1600 ;
        RECT 686.1200 162.3600 689.1200 162.8400 ;
        RECT 686.1200 156.9200 689.1200 157.4000 ;
        RECT 686.1200 167.8000 689.1200 168.2800 ;
        RECT 686.1200 146.0400 689.1200 146.5200 ;
        RECT 686.1200 151.4800 689.1200 151.9600 ;
        RECT 686.1200 135.1600 689.1200 135.6400 ;
        RECT 686.1200 129.7200 689.1200 130.2000 ;
        RECT 686.1200 140.6000 689.1200 141.0800 ;
        RECT 780.6800 118.8400 782.2800 119.3200 ;
        RECT 780.6800 124.2800 782.2800 124.7600 ;
        RECT 780.6800 102.5200 782.2800 103.0000 ;
        RECT 780.6800 107.9600 782.2800 108.4400 ;
        RECT 780.6800 113.4000 782.2800 113.8800 ;
        RECT 735.6800 118.8400 737.2800 119.3200 ;
        RECT 735.6800 124.2800 737.2800 124.7600 ;
        RECT 735.6800 102.5200 737.2800 103.0000 ;
        RECT 735.6800 107.9600 737.2800 108.4400 ;
        RECT 735.6800 113.4000 737.2800 113.8800 ;
        RECT 780.6800 97.0800 782.2800 97.5600 ;
        RECT 780.6800 91.6400 782.2800 92.1200 ;
        RECT 780.6800 86.2000 782.2800 86.6800 ;
        RECT 735.6800 97.0800 737.2800 97.5600 ;
        RECT 735.6800 91.6400 737.2800 92.1200 ;
        RECT 735.6800 86.2000 737.2800 86.6800 ;
        RECT 686.1200 118.8400 689.1200 119.3200 ;
        RECT 686.1200 124.2800 689.1200 124.7600 ;
        RECT 686.1200 107.9600 689.1200 108.4400 ;
        RECT 686.1200 102.5200 689.1200 103.0000 ;
        RECT 686.1200 113.4000 689.1200 113.8800 ;
        RECT 686.1200 91.6400 689.1200 92.1200 ;
        RECT 686.1200 97.0800 689.1200 97.5600 ;
        RECT 686.1200 86.2000 689.1200 86.6800 ;
        RECT 686.1200 284.3900 885.2200 287.3900 ;
        RECT 686.1200 79.2900 885.2200 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 686.1200 37.6700 688.1200 58.6000 ;
        RECT 883.2200 37.6700 885.2200 58.6000 ;
      LAYER met3 ;
        RECT 883.2200 54.1000 885.2200 54.5800 ;
        RECT 686.1200 54.1000 688.1200 54.5800 ;
        RECT 883.2200 43.2200 885.2200 43.7000 ;
        RECT 686.1200 43.2200 688.1200 43.7000 ;
        RECT 883.2200 48.6600 885.2200 49.1400 ;
        RECT 686.1200 48.6600 688.1200 49.1400 ;
        RECT 686.1200 56.6000 885.2200 58.6000 ;
        RECT 686.1200 37.6700 885.2200 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 2605.3300 872.2800 2813.4300 ;
        RECT 825.6800 2605.3300 827.2800 2813.4300 ;
        RECT 780.6800 2605.3300 782.2800 2813.4300 ;
        RECT 735.6800 2605.3300 737.2800 2813.4300 ;
        RECT 882.2200 2605.3300 885.2200 2813.4300 ;
        RECT 686.1200 2605.3300 689.1200 2813.4300 ;
      LAYER met3 ;
        RECT 882.2200 2808.0800 885.2200 2808.5600 ;
        RECT 870.6800 2808.0800 872.2800 2808.5600 ;
        RECT 882.2200 2797.2000 885.2200 2797.6800 ;
        RECT 882.2200 2802.6400 885.2200 2803.1200 ;
        RECT 870.6800 2797.2000 872.2800 2797.6800 ;
        RECT 870.6800 2802.6400 872.2800 2803.1200 ;
        RECT 882.2200 2780.8800 885.2200 2781.3600 ;
        RECT 882.2200 2786.3200 885.2200 2786.8000 ;
        RECT 870.6800 2780.8800 872.2800 2781.3600 ;
        RECT 870.6800 2786.3200 872.2800 2786.8000 ;
        RECT 882.2200 2770.0000 885.2200 2770.4800 ;
        RECT 882.2200 2775.4400 885.2200 2775.9200 ;
        RECT 870.6800 2770.0000 872.2800 2770.4800 ;
        RECT 870.6800 2775.4400 872.2800 2775.9200 ;
        RECT 882.2200 2791.7600 885.2200 2792.2400 ;
        RECT 870.6800 2791.7600 872.2800 2792.2400 ;
        RECT 825.6800 2797.2000 827.2800 2797.6800 ;
        RECT 825.6800 2802.6400 827.2800 2803.1200 ;
        RECT 825.6800 2808.0800 827.2800 2808.5600 ;
        RECT 825.6800 2780.8800 827.2800 2781.3600 ;
        RECT 825.6800 2786.3200 827.2800 2786.8000 ;
        RECT 825.6800 2775.4400 827.2800 2775.9200 ;
        RECT 825.6800 2770.0000 827.2800 2770.4800 ;
        RECT 825.6800 2791.7600 827.2800 2792.2400 ;
        RECT 882.2200 2753.6800 885.2200 2754.1600 ;
        RECT 882.2200 2759.1200 885.2200 2759.6000 ;
        RECT 870.6800 2753.6800 872.2800 2754.1600 ;
        RECT 870.6800 2759.1200 872.2800 2759.6000 ;
        RECT 882.2200 2737.3600 885.2200 2737.8400 ;
        RECT 882.2200 2742.8000 885.2200 2743.2800 ;
        RECT 882.2200 2748.2400 885.2200 2748.7200 ;
        RECT 870.6800 2737.3600 872.2800 2737.8400 ;
        RECT 870.6800 2742.8000 872.2800 2743.2800 ;
        RECT 870.6800 2748.2400 872.2800 2748.7200 ;
        RECT 882.2200 2726.4800 885.2200 2726.9600 ;
        RECT 882.2200 2731.9200 885.2200 2732.4000 ;
        RECT 870.6800 2726.4800 872.2800 2726.9600 ;
        RECT 870.6800 2731.9200 872.2800 2732.4000 ;
        RECT 882.2200 2710.1600 885.2200 2710.6400 ;
        RECT 882.2200 2715.6000 885.2200 2716.0800 ;
        RECT 882.2200 2721.0400 885.2200 2721.5200 ;
        RECT 870.6800 2710.1600 872.2800 2710.6400 ;
        RECT 870.6800 2715.6000 872.2800 2716.0800 ;
        RECT 870.6800 2721.0400 872.2800 2721.5200 ;
        RECT 825.6800 2753.6800 827.2800 2754.1600 ;
        RECT 825.6800 2759.1200 827.2800 2759.6000 ;
        RECT 825.6800 2737.3600 827.2800 2737.8400 ;
        RECT 825.6800 2742.8000 827.2800 2743.2800 ;
        RECT 825.6800 2748.2400 827.2800 2748.7200 ;
        RECT 825.6800 2726.4800 827.2800 2726.9600 ;
        RECT 825.6800 2731.9200 827.2800 2732.4000 ;
        RECT 825.6800 2710.1600 827.2800 2710.6400 ;
        RECT 825.6800 2715.6000 827.2800 2716.0800 ;
        RECT 825.6800 2721.0400 827.2800 2721.5200 ;
        RECT 882.2200 2764.5600 885.2200 2765.0400 ;
        RECT 825.6800 2764.5600 827.2800 2765.0400 ;
        RECT 870.6800 2764.5600 872.2800 2765.0400 ;
        RECT 780.6800 2797.2000 782.2800 2797.6800 ;
        RECT 780.6800 2802.6400 782.2800 2803.1200 ;
        RECT 780.6800 2808.0800 782.2800 2808.5600 ;
        RECT 735.6800 2797.2000 737.2800 2797.6800 ;
        RECT 735.6800 2802.6400 737.2800 2803.1200 ;
        RECT 735.6800 2808.0800 737.2800 2808.5600 ;
        RECT 780.6800 2780.8800 782.2800 2781.3600 ;
        RECT 780.6800 2786.3200 782.2800 2786.8000 ;
        RECT 780.6800 2770.0000 782.2800 2770.4800 ;
        RECT 780.6800 2775.4400 782.2800 2775.9200 ;
        RECT 735.6800 2780.8800 737.2800 2781.3600 ;
        RECT 735.6800 2786.3200 737.2800 2786.8000 ;
        RECT 735.6800 2770.0000 737.2800 2770.4800 ;
        RECT 735.6800 2775.4400 737.2800 2775.9200 ;
        RECT 735.6800 2791.7600 737.2800 2792.2400 ;
        RECT 780.6800 2791.7600 782.2800 2792.2400 ;
        RECT 686.1200 2808.0800 689.1200 2808.5600 ;
        RECT 686.1200 2802.6400 689.1200 2803.1200 ;
        RECT 686.1200 2797.2000 689.1200 2797.6800 ;
        RECT 686.1200 2786.3200 689.1200 2786.8000 ;
        RECT 686.1200 2780.8800 689.1200 2781.3600 ;
        RECT 686.1200 2775.4400 689.1200 2775.9200 ;
        RECT 686.1200 2770.0000 689.1200 2770.4800 ;
        RECT 686.1200 2791.7600 689.1200 2792.2400 ;
        RECT 780.6800 2753.6800 782.2800 2754.1600 ;
        RECT 780.6800 2759.1200 782.2800 2759.6000 ;
        RECT 780.6800 2737.3600 782.2800 2737.8400 ;
        RECT 780.6800 2742.8000 782.2800 2743.2800 ;
        RECT 780.6800 2748.2400 782.2800 2748.7200 ;
        RECT 735.6800 2753.6800 737.2800 2754.1600 ;
        RECT 735.6800 2759.1200 737.2800 2759.6000 ;
        RECT 735.6800 2737.3600 737.2800 2737.8400 ;
        RECT 735.6800 2742.8000 737.2800 2743.2800 ;
        RECT 735.6800 2748.2400 737.2800 2748.7200 ;
        RECT 780.6800 2726.4800 782.2800 2726.9600 ;
        RECT 780.6800 2731.9200 782.2800 2732.4000 ;
        RECT 780.6800 2710.1600 782.2800 2710.6400 ;
        RECT 780.6800 2715.6000 782.2800 2716.0800 ;
        RECT 780.6800 2721.0400 782.2800 2721.5200 ;
        RECT 735.6800 2726.4800 737.2800 2726.9600 ;
        RECT 735.6800 2731.9200 737.2800 2732.4000 ;
        RECT 735.6800 2710.1600 737.2800 2710.6400 ;
        RECT 735.6800 2715.6000 737.2800 2716.0800 ;
        RECT 735.6800 2721.0400 737.2800 2721.5200 ;
        RECT 686.1200 2753.6800 689.1200 2754.1600 ;
        RECT 686.1200 2759.1200 689.1200 2759.6000 ;
        RECT 686.1200 2742.8000 689.1200 2743.2800 ;
        RECT 686.1200 2737.3600 689.1200 2737.8400 ;
        RECT 686.1200 2748.2400 689.1200 2748.7200 ;
        RECT 686.1200 2726.4800 689.1200 2726.9600 ;
        RECT 686.1200 2731.9200 689.1200 2732.4000 ;
        RECT 686.1200 2715.6000 689.1200 2716.0800 ;
        RECT 686.1200 2710.1600 689.1200 2710.6400 ;
        RECT 686.1200 2721.0400 689.1200 2721.5200 ;
        RECT 686.1200 2764.5600 689.1200 2765.0400 ;
        RECT 735.6800 2764.5600 737.2800 2765.0400 ;
        RECT 780.6800 2764.5600 782.2800 2765.0400 ;
        RECT 882.2200 2699.2800 885.2200 2699.7600 ;
        RECT 882.2200 2704.7200 885.2200 2705.2000 ;
        RECT 870.6800 2699.2800 872.2800 2699.7600 ;
        RECT 870.6800 2704.7200 872.2800 2705.2000 ;
        RECT 882.2200 2682.9600 885.2200 2683.4400 ;
        RECT 882.2200 2688.4000 885.2200 2688.8800 ;
        RECT 882.2200 2693.8400 885.2200 2694.3200 ;
        RECT 870.6800 2682.9600 872.2800 2683.4400 ;
        RECT 870.6800 2688.4000 872.2800 2688.8800 ;
        RECT 870.6800 2693.8400 872.2800 2694.3200 ;
        RECT 882.2200 2672.0800 885.2200 2672.5600 ;
        RECT 882.2200 2677.5200 885.2200 2678.0000 ;
        RECT 870.6800 2672.0800 872.2800 2672.5600 ;
        RECT 870.6800 2677.5200 872.2800 2678.0000 ;
        RECT 882.2200 2655.7600 885.2200 2656.2400 ;
        RECT 882.2200 2661.2000 885.2200 2661.6800 ;
        RECT 882.2200 2666.6400 885.2200 2667.1200 ;
        RECT 870.6800 2655.7600 872.2800 2656.2400 ;
        RECT 870.6800 2661.2000 872.2800 2661.6800 ;
        RECT 870.6800 2666.6400 872.2800 2667.1200 ;
        RECT 825.6800 2699.2800 827.2800 2699.7600 ;
        RECT 825.6800 2704.7200 827.2800 2705.2000 ;
        RECT 825.6800 2682.9600 827.2800 2683.4400 ;
        RECT 825.6800 2688.4000 827.2800 2688.8800 ;
        RECT 825.6800 2693.8400 827.2800 2694.3200 ;
        RECT 825.6800 2672.0800 827.2800 2672.5600 ;
        RECT 825.6800 2677.5200 827.2800 2678.0000 ;
        RECT 825.6800 2655.7600 827.2800 2656.2400 ;
        RECT 825.6800 2661.2000 827.2800 2661.6800 ;
        RECT 825.6800 2666.6400 827.2800 2667.1200 ;
        RECT 882.2200 2644.8800 885.2200 2645.3600 ;
        RECT 882.2200 2650.3200 885.2200 2650.8000 ;
        RECT 870.6800 2644.8800 872.2800 2645.3600 ;
        RECT 870.6800 2650.3200 872.2800 2650.8000 ;
        RECT 882.2200 2628.5600 885.2200 2629.0400 ;
        RECT 882.2200 2634.0000 885.2200 2634.4800 ;
        RECT 882.2200 2639.4400 885.2200 2639.9200 ;
        RECT 870.6800 2628.5600 872.2800 2629.0400 ;
        RECT 870.6800 2634.0000 872.2800 2634.4800 ;
        RECT 870.6800 2639.4400 872.2800 2639.9200 ;
        RECT 882.2200 2617.6800 885.2200 2618.1600 ;
        RECT 882.2200 2623.1200 885.2200 2623.6000 ;
        RECT 870.6800 2617.6800 872.2800 2618.1600 ;
        RECT 870.6800 2623.1200 872.2800 2623.6000 ;
        RECT 882.2200 2612.2400 885.2200 2612.7200 ;
        RECT 870.6800 2612.2400 872.2800 2612.7200 ;
        RECT 825.6800 2644.8800 827.2800 2645.3600 ;
        RECT 825.6800 2650.3200 827.2800 2650.8000 ;
        RECT 825.6800 2628.5600 827.2800 2629.0400 ;
        RECT 825.6800 2634.0000 827.2800 2634.4800 ;
        RECT 825.6800 2639.4400 827.2800 2639.9200 ;
        RECT 825.6800 2617.6800 827.2800 2618.1600 ;
        RECT 825.6800 2623.1200 827.2800 2623.6000 ;
        RECT 825.6800 2612.2400 827.2800 2612.7200 ;
        RECT 780.6800 2699.2800 782.2800 2699.7600 ;
        RECT 780.6800 2704.7200 782.2800 2705.2000 ;
        RECT 780.6800 2682.9600 782.2800 2683.4400 ;
        RECT 780.6800 2688.4000 782.2800 2688.8800 ;
        RECT 780.6800 2693.8400 782.2800 2694.3200 ;
        RECT 735.6800 2699.2800 737.2800 2699.7600 ;
        RECT 735.6800 2704.7200 737.2800 2705.2000 ;
        RECT 735.6800 2682.9600 737.2800 2683.4400 ;
        RECT 735.6800 2688.4000 737.2800 2688.8800 ;
        RECT 735.6800 2693.8400 737.2800 2694.3200 ;
        RECT 780.6800 2672.0800 782.2800 2672.5600 ;
        RECT 780.6800 2677.5200 782.2800 2678.0000 ;
        RECT 780.6800 2655.7600 782.2800 2656.2400 ;
        RECT 780.6800 2661.2000 782.2800 2661.6800 ;
        RECT 780.6800 2666.6400 782.2800 2667.1200 ;
        RECT 735.6800 2672.0800 737.2800 2672.5600 ;
        RECT 735.6800 2677.5200 737.2800 2678.0000 ;
        RECT 735.6800 2655.7600 737.2800 2656.2400 ;
        RECT 735.6800 2661.2000 737.2800 2661.6800 ;
        RECT 735.6800 2666.6400 737.2800 2667.1200 ;
        RECT 686.1200 2699.2800 689.1200 2699.7600 ;
        RECT 686.1200 2704.7200 689.1200 2705.2000 ;
        RECT 686.1200 2688.4000 689.1200 2688.8800 ;
        RECT 686.1200 2682.9600 689.1200 2683.4400 ;
        RECT 686.1200 2693.8400 689.1200 2694.3200 ;
        RECT 686.1200 2672.0800 689.1200 2672.5600 ;
        RECT 686.1200 2677.5200 689.1200 2678.0000 ;
        RECT 686.1200 2661.2000 689.1200 2661.6800 ;
        RECT 686.1200 2655.7600 689.1200 2656.2400 ;
        RECT 686.1200 2666.6400 689.1200 2667.1200 ;
        RECT 780.6800 2644.8800 782.2800 2645.3600 ;
        RECT 780.6800 2650.3200 782.2800 2650.8000 ;
        RECT 780.6800 2628.5600 782.2800 2629.0400 ;
        RECT 780.6800 2634.0000 782.2800 2634.4800 ;
        RECT 780.6800 2639.4400 782.2800 2639.9200 ;
        RECT 735.6800 2644.8800 737.2800 2645.3600 ;
        RECT 735.6800 2650.3200 737.2800 2650.8000 ;
        RECT 735.6800 2628.5600 737.2800 2629.0400 ;
        RECT 735.6800 2634.0000 737.2800 2634.4800 ;
        RECT 735.6800 2639.4400 737.2800 2639.9200 ;
        RECT 780.6800 2623.1200 782.2800 2623.6000 ;
        RECT 780.6800 2617.6800 782.2800 2618.1600 ;
        RECT 780.6800 2612.2400 782.2800 2612.7200 ;
        RECT 735.6800 2623.1200 737.2800 2623.6000 ;
        RECT 735.6800 2617.6800 737.2800 2618.1600 ;
        RECT 735.6800 2612.2400 737.2800 2612.7200 ;
        RECT 686.1200 2644.8800 689.1200 2645.3600 ;
        RECT 686.1200 2650.3200 689.1200 2650.8000 ;
        RECT 686.1200 2634.0000 689.1200 2634.4800 ;
        RECT 686.1200 2628.5600 689.1200 2629.0400 ;
        RECT 686.1200 2639.4400 689.1200 2639.9200 ;
        RECT 686.1200 2617.6800 689.1200 2618.1600 ;
        RECT 686.1200 2623.1200 689.1200 2623.6000 ;
        RECT 686.1200 2612.2400 689.1200 2612.7200 ;
        RECT 686.1200 2810.4300 885.2200 2813.4300 ;
        RECT 686.1200 2605.3300 885.2200 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 2375.6900 872.2800 2583.7900 ;
        RECT 825.6800 2375.6900 827.2800 2583.7900 ;
        RECT 780.6800 2375.6900 782.2800 2583.7900 ;
        RECT 735.6800 2375.6900 737.2800 2583.7900 ;
        RECT 882.2200 2375.6900 885.2200 2583.7900 ;
        RECT 686.1200 2375.6900 689.1200 2583.7900 ;
      LAYER met3 ;
        RECT 882.2200 2578.4400 885.2200 2578.9200 ;
        RECT 870.6800 2578.4400 872.2800 2578.9200 ;
        RECT 882.2200 2567.5600 885.2200 2568.0400 ;
        RECT 882.2200 2573.0000 885.2200 2573.4800 ;
        RECT 870.6800 2567.5600 872.2800 2568.0400 ;
        RECT 870.6800 2573.0000 872.2800 2573.4800 ;
        RECT 882.2200 2551.2400 885.2200 2551.7200 ;
        RECT 882.2200 2556.6800 885.2200 2557.1600 ;
        RECT 870.6800 2551.2400 872.2800 2551.7200 ;
        RECT 870.6800 2556.6800 872.2800 2557.1600 ;
        RECT 882.2200 2540.3600 885.2200 2540.8400 ;
        RECT 882.2200 2545.8000 885.2200 2546.2800 ;
        RECT 870.6800 2540.3600 872.2800 2540.8400 ;
        RECT 870.6800 2545.8000 872.2800 2546.2800 ;
        RECT 882.2200 2562.1200 885.2200 2562.6000 ;
        RECT 870.6800 2562.1200 872.2800 2562.6000 ;
        RECT 825.6800 2567.5600 827.2800 2568.0400 ;
        RECT 825.6800 2573.0000 827.2800 2573.4800 ;
        RECT 825.6800 2578.4400 827.2800 2578.9200 ;
        RECT 825.6800 2551.2400 827.2800 2551.7200 ;
        RECT 825.6800 2556.6800 827.2800 2557.1600 ;
        RECT 825.6800 2545.8000 827.2800 2546.2800 ;
        RECT 825.6800 2540.3600 827.2800 2540.8400 ;
        RECT 825.6800 2562.1200 827.2800 2562.6000 ;
        RECT 882.2200 2524.0400 885.2200 2524.5200 ;
        RECT 882.2200 2529.4800 885.2200 2529.9600 ;
        RECT 870.6800 2524.0400 872.2800 2524.5200 ;
        RECT 870.6800 2529.4800 872.2800 2529.9600 ;
        RECT 882.2200 2507.7200 885.2200 2508.2000 ;
        RECT 882.2200 2513.1600 885.2200 2513.6400 ;
        RECT 882.2200 2518.6000 885.2200 2519.0800 ;
        RECT 870.6800 2507.7200 872.2800 2508.2000 ;
        RECT 870.6800 2513.1600 872.2800 2513.6400 ;
        RECT 870.6800 2518.6000 872.2800 2519.0800 ;
        RECT 882.2200 2496.8400 885.2200 2497.3200 ;
        RECT 882.2200 2502.2800 885.2200 2502.7600 ;
        RECT 870.6800 2496.8400 872.2800 2497.3200 ;
        RECT 870.6800 2502.2800 872.2800 2502.7600 ;
        RECT 882.2200 2480.5200 885.2200 2481.0000 ;
        RECT 882.2200 2485.9600 885.2200 2486.4400 ;
        RECT 882.2200 2491.4000 885.2200 2491.8800 ;
        RECT 870.6800 2480.5200 872.2800 2481.0000 ;
        RECT 870.6800 2485.9600 872.2800 2486.4400 ;
        RECT 870.6800 2491.4000 872.2800 2491.8800 ;
        RECT 825.6800 2524.0400 827.2800 2524.5200 ;
        RECT 825.6800 2529.4800 827.2800 2529.9600 ;
        RECT 825.6800 2507.7200 827.2800 2508.2000 ;
        RECT 825.6800 2513.1600 827.2800 2513.6400 ;
        RECT 825.6800 2518.6000 827.2800 2519.0800 ;
        RECT 825.6800 2496.8400 827.2800 2497.3200 ;
        RECT 825.6800 2502.2800 827.2800 2502.7600 ;
        RECT 825.6800 2480.5200 827.2800 2481.0000 ;
        RECT 825.6800 2485.9600 827.2800 2486.4400 ;
        RECT 825.6800 2491.4000 827.2800 2491.8800 ;
        RECT 882.2200 2534.9200 885.2200 2535.4000 ;
        RECT 825.6800 2534.9200 827.2800 2535.4000 ;
        RECT 870.6800 2534.9200 872.2800 2535.4000 ;
        RECT 780.6800 2567.5600 782.2800 2568.0400 ;
        RECT 780.6800 2573.0000 782.2800 2573.4800 ;
        RECT 780.6800 2578.4400 782.2800 2578.9200 ;
        RECT 735.6800 2567.5600 737.2800 2568.0400 ;
        RECT 735.6800 2573.0000 737.2800 2573.4800 ;
        RECT 735.6800 2578.4400 737.2800 2578.9200 ;
        RECT 780.6800 2551.2400 782.2800 2551.7200 ;
        RECT 780.6800 2556.6800 782.2800 2557.1600 ;
        RECT 780.6800 2540.3600 782.2800 2540.8400 ;
        RECT 780.6800 2545.8000 782.2800 2546.2800 ;
        RECT 735.6800 2551.2400 737.2800 2551.7200 ;
        RECT 735.6800 2556.6800 737.2800 2557.1600 ;
        RECT 735.6800 2540.3600 737.2800 2540.8400 ;
        RECT 735.6800 2545.8000 737.2800 2546.2800 ;
        RECT 735.6800 2562.1200 737.2800 2562.6000 ;
        RECT 780.6800 2562.1200 782.2800 2562.6000 ;
        RECT 686.1200 2578.4400 689.1200 2578.9200 ;
        RECT 686.1200 2573.0000 689.1200 2573.4800 ;
        RECT 686.1200 2567.5600 689.1200 2568.0400 ;
        RECT 686.1200 2556.6800 689.1200 2557.1600 ;
        RECT 686.1200 2551.2400 689.1200 2551.7200 ;
        RECT 686.1200 2545.8000 689.1200 2546.2800 ;
        RECT 686.1200 2540.3600 689.1200 2540.8400 ;
        RECT 686.1200 2562.1200 689.1200 2562.6000 ;
        RECT 780.6800 2524.0400 782.2800 2524.5200 ;
        RECT 780.6800 2529.4800 782.2800 2529.9600 ;
        RECT 780.6800 2507.7200 782.2800 2508.2000 ;
        RECT 780.6800 2513.1600 782.2800 2513.6400 ;
        RECT 780.6800 2518.6000 782.2800 2519.0800 ;
        RECT 735.6800 2524.0400 737.2800 2524.5200 ;
        RECT 735.6800 2529.4800 737.2800 2529.9600 ;
        RECT 735.6800 2507.7200 737.2800 2508.2000 ;
        RECT 735.6800 2513.1600 737.2800 2513.6400 ;
        RECT 735.6800 2518.6000 737.2800 2519.0800 ;
        RECT 780.6800 2496.8400 782.2800 2497.3200 ;
        RECT 780.6800 2502.2800 782.2800 2502.7600 ;
        RECT 780.6800 2480.5200 782.2800 2481.0000 ;
        RECT 780.6800 2485.9600 782.2800 2486.4400 ;
        RECT 780.6800 2491.4000 782.2800 2491.8800 ;
        RECT 735.6800 2496.8400 737.2800 2497.3200 ;
        RECT 735.6800 2502.2800 737.2800 2502.7600 ;
        RECT 735.6800 2480.5200 737.2800 2481.0000 ;
        RECT 735.6800 2485.9600 737.2800 2486.4400 ;
        RECT 735.6800 2491.4000 737.2800 2491.8800 ;
        RECT 686.1200 2524.0400 689.1200 2524.5200 ;
        RECT 686.1200 2529.4800 689.1200 2529.9600 ;
        RECT 686.1200 2513.1600 689.1200 2513.6400 ;
        RECT 686.1200 2507.7200 689.1200 2508.2000 ;
        RECT 686.1200 2518.6000 689.1200 2519.0800 ;
        RECT 686.1200 2496.8400 689.1200 2497.3200 ;
        RECT 686.1200 2502.2800 689.1200 2502.7600 ;
        RECT 686.1200 2485.9600 689.1200 2486.4400 ;
        RECT 686.1200 2480.5200 689.1200 2481.0000 ;
        RECT 686.1200 2491.4000 689.1200 2491.8800 ;
        RECT 686.1200 2534.9200 689.1200 2535.4000 ;
        RECT 735.6800 2534.9200 737.2800 2535.4000 ;
        RECT 780.6800 2534.9200 782.2800 2535.4000 ;
        RECT 882.2200 2469.6400 885.2200 2470.1200 ;
        RECT 882.2200 2475.0800 885.2200 2475.5600 ;
        RECT 870.6800 2469.6400 872.2800 2470.1200 ;
        RECT 870.6800 2475.0800 872.2800 2475.5600 ;
        RECT 882.2200 2453.3200 885.2200 2453.8000 ;
        RECT 882.2200 2458.7600 885.2200 2459.2400 ;
        RECT 882.2200 2464.2000 885.2200 2464.6800 ;
        RECT 870.6800 2453.3200 872.2800 2453.8000 ;
        RECT 870.6800 2458.7600 872.2800 2459.2400 ;
        RECT 870.6800 2464.2000 872.2800 2464.6800 ;
        RECT 882.2200 2442.4400 885.2200 2442.9200 ;
        RECT 882.2200 2447.8800 885.2200 2448.3600 ;
        RECT 870.6800 2442.4400 872.2800 2442.9200 ;
        RECT 870.6800 2447.8800 872.2800 2448.3600 ;
        RECT 882.2200 2426.1200 885.2200 2426.6000 ;
        RECT 882.2200 2431.5600 885.2200 2432.0400 ;
        RECT 882.2200 2437.0000 885.2200 2437.4800 ;
        RECT 870.6800 2426.1200 872.2800 2426.6000 ;
        RECT 870.6800 2431.5600 872.2800 2432.0400 ;
        RECT 870.6800 2437.0000 872.2800 2437.4800 ;
        RECT 825.6800 2469.6400 827.2800 2470.1200 ;
        RECT 825.6800 2475.0800 827.2800 2475.5600 ;
        RECT 825.6800 2453.3200 827.2800 2453.8000 ;
        RECT 825.6800 2458.7600 827.2800 2459.2400 ;
        RECT 825.6800 2464.2000 827.2800 2464.6800 ;
        RECT 825.6800 2442.4400 827.2800 2442.9200 ;
        RECT 825.6800 2447.8800 827.2800 2448.3600 ;
        RECT 825.6800 2426.1200 827.2800 2426.6000 ;
        RECT 825.6800 2431.5600 827.2800 2432.0400 ;
        RECT 825.6800 2437.0000 827.2800 2437.4800 ;
        RECT 882.2200 2415.2400 885.2200 2415.7200 ;
        RECT 882.2200 2420.6800 885.2200 2421.1600 ;
        RECT 870.6800 2415.2400 872.2800 2415.7200 ;
        RECT 870.6800 2420.6800 872.2800 2421.1600 ;
        RECT 882.2200 2398.9200 885.2200 2399.4000 ;
        RECT 882.2200 2404.3600 885.2200 2404.8400 ;
        RECT 882.2200 2409.8000 885.2200 2410.2800 ;
        RECT 870.6800 2398.9200 872.2800 2399.4000 ;
        RECT 870.6800 2404.3600 872.2800 2404.8400 ;
        RECT 870.6800 2409.8000 872.2800 2410.2800 ;
        RECT 882.2200 2388.0400 885.2200 2388.5200 ;
        RECT 882.2200 2393.4800 885.2200 2393.9600 ;
        RECT 870.6800 2388.0400 872.2800 2388.5200 ;
        RECT 870.6800 2393.4800 872.2800 2393.9600 ;
        RECT 882.2200 2382.6000 885.2200 2383.0800 ;
        RECT 870.6800 2382.6000 872.2800 2383.0800 ;
        RECT 825.6800 2415.2400 827.2800 2415.7200 ;
        RECT 825.6800 2420.6800 827.2800 2421.1600 ;
        RECT 825.6800 2398.9200 827.2800 2399.4000 ;
        RECT 825.6800 2404.3600 827.2800 2404.8400 ;
        RECT 825.6800 2409.8000 827.2800 2410.2800 ;
        RECT 825.6800 2388.0400 827.2800 2388.5200 ;
        RECT 825.6800 2393.4800 827.2800 2393.9600 ;
        RECT 825.6800 2382.6000 827.2800 2383.0800 ;
        RECT 780.6800 2469.6400 782.2800 2470.1200 ;
        RECT 780.6800 2475.0800 782.2800 2475.5600 ;
        RECT 780.6800 2453.3200 782.2800 2453.8000 ;
        RECT 780.6800 2458.7600 782.2800 2459.2400 ;
        RECT 780.6800 2464.2000 782.2800 2464.6800 ;
        RECT 735.6800 2469.6400 737.2800 2470.1200 ;
        RECT 735.6800 2475.0800 737.2800 2475.5600 ;
        RECT 735.6800 2453.3200 737.2800 2453.8000 ;
        RECT 735.6800 2458.7600 737.2800 2459.2400 ;
        RECT 735.6800 2464.2000 737.2800 2464.6800 ;
        RECT 780.6800 2442.4400 782.2800 2442.9200 ;
        RECT 780.6800 2447.8800 782.2800 2448.3600 ;
        RECT 780.6800 2426.1200 782.2800 2426.6000 ;
        RECT 780.6800 2431.5600 782.2800 2432.0400 ;
        RECT 780.6800 2437.0000 782.2800 2437.4800 ;
        RECT 735.6800 2442.4400 737.2800 2442.9200 ;
        RECT 735.6800 2447.8800 737.2800 2448.3600 ;
        RECT 735.6800 2426.1200 737.2800 2426.6000 ;
        RECT 735.6800 2431.5600 737.2800 2432.0400 ;
        RECT 735.6800 2437.0000 737.2800 2437.4800 ;
        RECT 686.1200 2469.6400 689.1200 2470.1200 ;
        RECT 686.1200 2475.0800 689.1200 2475.5600 ;
        RECT 686.1200 2458.7600 689.1200 2459.2400 ;
        RECT 686.1200 2453.3200 689.1200 2453.8000 ;
        RECT 686.1200 2464.2000 689.1200 2464.6800 ;
        RECT 686.1200 2442.4400 689.1200 2442.9200 ;
        RECT 686.1200 2447.8800 689.1200 2448.3600 ;
        RECT 686.1200 2431.5600 689.1200 2432.0400 ;
        RECT 686.1200 2426.1200 689.1200 2426.6000 ;
        RECT 686.1200 2437.0000 689.1200 2437.4800 ;
        RECT 780.6800 2415.2400 782.2800 2415.7200 ;
        RECT 780.6800 2420.6800 782.2800 2421.1600 ;
        RECT 780.6800 2398.9200 782.2800 2399.4000 ;
        RECT 780.6800 2404.3600 782.2800 2404.8400 ;
        RECT 780.6800 2409.8000 782.2800 2410.2800 ;
        RECT 735.6800 2415.2400 737.2800 2415.7200 ;
        RECT 735.6800 2420.6800 737.2800 2421.1600 ;
        RECT 735.6800 2398.9200 737.2800 2399.4000 ;
        RECT 735.6800 2404.3600 737.2800 2404.8400 ;
        RECT 735.6800 2409.8000 737.2800 2410.2800 ;
        RECT 780.6800 2393.4800 782.2800 2393.9600 ;
        RECT 780.6800 2388.0400 782.2800 2388.5200 ;
        RECT 780.6800 2382.6000 782.2800 2383.0800 ;
        RECT 735.6800 2393.4800 737.2800 2393.9600 ;
        RECT 735.6800 2388.0400 737.2800 2388.5200 ;
        RECT 735.6800 2382.6000 737.2800 2383.0800 ;
        RECT 686.1200 2415.2400 689.1200 2415.7200 ;
        RECT 686.1200 2420.6800 689.1200 2421.1600 ;
        RECT 686.1200 2404.3600 689.1200 2404.8400 ;
        RECT 686.1200 2398.9200 689.1200 2399.4000 ;
        RECT 686.1200 2409.8000 689.1200 2410.2800 ;
        RECT 686.1200 2388.0400 689.1200 2388.5200 ;
        RECT 686.1200 2393.4800 689.1200 2393.9600 ;
        RECT 686.1200 2382.6000 689.1200 2383.0800 ;
        RECT 686.1200 2580.7900 885.2200 2583.7900 ;
        RECT 686.1200 2375.6900 885.2200 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 2146.0500 872.2800 2354.1500 ;
        RECT 825.6800 2146.0500 827.2800 2354.1500 ;
        RECT 780.6800 2146.0500 782.2800 2354.1500 ;
        RECT 735.6800 2146.0500 737.2800 2354.1500 ;
        RECT 882.2200 2146.0500 885.2200 2354.1500 ;
        RECT 686.1200 2146.0500 689.1200 2354.1500 ;
      LAYER met3 ;
        RECT 882.2200 2348.8000 885.2200 2349.2800 ;
        RECT 870.6800 2348.8000 872.2800 2349.2800 ;
        RECT 882.2200 2337.9200 885.2200 2338.4000 ;
        RECT 882.2200 2343.3600 885.2200 2343.8400 ;
        RECT 870.6800 2337.9200 872.2800 2338.4000 ;
        RECT 870.6800 2343.3600 872.2800 2343.8400 ;
        RECT 882.2200 2321.6000 885.2200 2322.0800 ;
        RECT 882.2200 2327.0400 885.2200 2327.5200 ;
        RECT 870.6800 2321.6000 872.2800 2322.0800 ;
        RECT 870.6800 2327.0400 872.2800 2327.5200 ;
        RECT 882.2200 2310.7200 885.2200 2311.2000 ;
        RECT 882.2200 2316.1600 885.2200 2316.6400 ;
        RECT 870.6800 2310.7200 872.2800 2311.2000 ;
        RECT 870.6800 2316.1600 872.2800 2316.6400 ;
        RECT 882.2200 2332.4800 885.2200 2332.9600 ;
        RECT 870.6800 2332.4800 872.2800 2332.9600 ;
        RECT 825.6800 2337.9200 827.2800 2338.4000 ;
        RECT 825.6800 2343.3600 827.2800 2343.8400 ;
        RECT 825.6800 2348.8000 827.2800 2349.2800 ;
        RECT 825.6800 2321.6000 827.2800 2322.0800 ;
        RECT 825.6800 2327.0400 827.2800 2327.5200 ;
        RECT 825.6800 2316.1600 827.2800 2316.6400 ;
        RECT 825.6800 2310.7200 827.2800 2311.2000 ;
        RECT 825.6800 2332.4800 827.2800 2332.9600 ;
        RECT 882.2200 2294.4000 885.2200 2294.8800 ;
        RECT 882.2200 2299.8400 885.2200 2300.3200 ;
        RECT 870.6800 2294.4000 872.2800 2294.8800 ;
        RECT 870.6800 2299.8400 872.2800 2300.3200 ;
        RECT 882.2200 2278.0800 885.2200 2278.5600 ;
        RECT 882.2200 2283.5200 885.2200 2284.0000 ;
        RECT 882.2200 2288.9600 885.2200 2289.4400 ;
        RECT 870.6800 2278.0800 872.2800 2278.5600 ;
        RECT 870.6800 2283.5200 872.2800 2284.0000 ;
        RECT 870.6800 2288.9600 872.2800 2289.4400 ;
        RECT 882.2200 2267.2000 885.2200 2267.6800 ;
        RECT 882.2200 2272.6400 885.2200 2273.1200 ;
        RECT 870.6800 2267.2000 872.2800 2267.6800 ;
        RECT 870.6800 2272.6400 872.2800 2273.1200 ;
        RECT 882.2200 2250.8800 885.2200 2251.3600 ;
        RECT 882.2200 2256.3200 885.2200 2256.8000 ;
        RECT 882.2200 2261.7600 885.2200 2262.2400 ;
        RECT 870.6800 2250.8800 872.2800 2251.3600 ;
        RECT 870.6800 2256.3200 872.2800 2256.8000 ;
        RECT 870.6800 2261.7600 872.2800 2262.2400 ;
        RECT 825.6800 2294.4000 827.2800 2294.8800 ;
        RECT 825.6800 2299.8400 827.2800 2300.3200 ;
        RECT 825.6800 2278.0800 827.2800 2278.5600 ;
        RECT 825.6800 2283.5200 827.2800 2284.0000 ;
        RECT 825.6800 2288.9600 827.2800 2289.4400 ;
        RECT 825.6800 2267.2000 827.2800 2267.6800 ;
        RECT 825.6800 2272.6400 827.2800 2273.1200 ;
        RECT 825.6800 2250.8800 827.2800 2251.3600 ;
        RECT 825.6800 2256.3200 827.2800 2256.8000 ;
        RECT 825.6800 2261.7600 827.2800 2262.2400 ;
        RECT 882.2200 2305.2800 885.2200 2305.7600 ;
        RECT 825.6800 2305.2800 827.2800 2305.7600 ;
        RECT 870.6800 2305.2800 872.2800 2305.7600 ;
        RECT 780.6800 2337.9200 782.2800 2338.4000 ;
        RECT 780.6800 2343.3600 782.2800 2343.8400 ;
        RECT 780.6800 2348.8000 782.2800 2349.2800 ;
        RECT 735.6800 2337.9200 737.2800 2338.4000 ;
        RECT 735.6800 2343.3600 737.2800 2343.8400 ;
        RECT 735.6800 2348.8000 737.2800 2349.2800 ;
        RECT 780.6800 2321.6000 782.2800 2322.0800 ;
        RECT 780.6800 2327.0400 782.2800 2327.5200 ;
        RECT 780.6800 2310.7200 782.2800 2311.2000 ;
        RECT 780.6800 2316.1600 782.2800 2316.6400 ;
        RECT 735.6800 2321.6000 737.2800 2322.0800 ;
        RECT 735.6800 2327.0400 737.2800 2327.5200 ;
        RECT 735.6800 2310.7200 737.2800 2311.2000 ;
        RECT 735.6800 2316.1600 737.2800 2316.6400 ;
        RECT 735.6800 2332.4800 737.2800 2332.9600 ;
        RECT 780.6800 2332.4800 782.2800 2332.9600 ;
        RECT 686.1200 2348.8000 689.1200 2349.2800 ;
        RECT 686.1200 2343.3600 689.1200 2343.8400 ;
        RECT 686.1200 2337.9200 689.1200 2338.4000 ;
        RECT 686.1200 2327.0400 689.1200 2327.5200 ;
        RECT 686.1200 2321.6000 689.1200 2322.0800 ;
        RECT 686.1200 2316.1600 689.1200 2316.6400 ;
        RECT 686.1200 2310.7200 689.1200 2311.2000 ;
        RECT 686.1200 2332.4800 689.1200 2332.9600 ;
        RECT 780.6800 2294.4000 782.2800 2294.8800 ;
        RECT 780.6800 2299.8400 782.2800 2300.3200 ;
        RECT 780.6800 2278.0800 782.2800 2278.5600 ;
        RECT 780.6800 2283.5200 782.2800 2284.0000 ;
        RECT 780.6800 2288.9600 782.2800 2289.4400 ;
        RECT 735.6800 2294.4000 737.2800 2294.8800 ;
        RECT 735.6800 2299.8400 737.2800 2300.3200 ;
        RECT 735.6800 2278.0800 737.2800 2278.5600 ;
        RECT 735.6800 2283.5200 737.2800 2284.0000 ;
        RECT 735.6800 2288.9600 737.2800 2289.4400 ;
        RECT 780.6800 2267.2000 782.2800 2267.6800 ;
        RECT 780.6800 2272.6400 782.2800 2273.1200 ;
        RECT 780.6800 2250.8800 782.2800 2251.3600 ;
        RECT 780.6800 2256.3200 782.2800 2256.8000 ;
        RECT 780.6800 2261.7600 782.2800 2262.2400 ;
        RECT 735.6800 2267.2000 737.2800 2267.6800 ;
        RECT 735.6800 2272.6400 737.2800 2273.1200 ;
        RECT 735.6800 2250.8800 737.2800 2251.3600 ;
        RECT 735.6800 2256.3200 737.2800 2256.8000 ;
        RECT 735.6800 2261.7600 737.2800 2262.2400 ;
        RECT 686.1200 2294.4000 689.1200 2294.8800 ;
        RECT 686.1200 2299.8400 689.1200 2300.3200 ;
        RECT 686.1200 2283.5200 689.1200 2284.0000 ;
        RECT 686.1200 2278.0800 689.1200 2278.5600 ;
        RECT 686.1200 2288.9600 689.1200 2289.4400 ;
        RECT 686.1200 2267.2000 689.1200 2267.6800 ;
        RECT 686.1200 2272.6400 689.1200 2273.1200 ;
        RECT 686.1200 2256.3200 689.1200 2256.8000 ;
        RECT 686.1200 2250.8800 689.1200 2251.3600 ;
        RECT 686.1200 2261.7600 689.1200 2262.2400 ;
        RECT 686.1200 2305.2800 689.1200 2305.7600 ;
        RECT 735.6800 2305.2800 737.2800 2305.7600 ;
        RECT 780.6800 2305.2800 782.2800 2305.7600 ;
        RECT 882.2200 2240.0000 885.2200 2240.4800 ;
        RECT 882.2200 2245.4400 885.2200 2245.9200 ;
        RECT 870.6800 2240.0000 872.2800 2240.4800 ;
        RECT 870.6800 2245.4400 872.2800 2245.9200 ;
        RECT 882.2200 2223.6800 885.2200 2224.1600 ;
        RECT 882.2200 2229.1200 885.2200 2229.6000 ;
        RECT 882.2200 2234.5600 885.2200 2235.0400 ;
        RECT 870.6800 2223.6800 872.2800 2224.1600 ;
        RECT 870.6800 2229.1200 872.2800 2229.6000 ;
        RECT 870.6800 2234.5600 872.2800 2235.0400 ;
        RECT 882.2200 2212.8000 885.2200 2213.2800 ;
        RECT 882.2200 2218.2400 885.2200 2218.7200 ;
        RECT 870.6800 2212.8000 872.2800 2213.2800 ;
        RECT 870.6800 2218.2400 872.2800 2218.7200 ;
        RECT 882.2200 2196.4800 885.2200 2196.9600 ;
        RECT 882.2200 2201.9200 885.2200 2202.4000 ;
        RECT 882.2200 2207.3600 885.2200 2207.8400 ;
        RECT 870.6800 2196.4800 872.2800 2196.9600 ;
        RECT 870.6800 2201.9200 872.2800 2202.4000 ;
        RECT 870.6800 2207.3600 872.2800 2207.8400 ;
        RECT 825.6800 2240.0000 827.2800 2240.4800 ;
        RECT 825.6800 2245.4400 827.2800 2245.9200 ;
        RECT 825.6800 2223.6800 827.2800 2224.1600 ;
        RECT 825.6800 2229.1200 827.2800 2229.6000 ;
        RECT 825.6800 2234.5600 827.2800 2235.0400 ;
        RECT 825.6800 2212.8000 827.2800 2213.2800 ;
        RECT 825.6800 2218.2400 827.2800 2218.7200 ;
        RECT 825.6800 2196.4800 827.2800 2196.9600 ;
        RECT 825.6800 2201.9200 827.2800 2202.4000 ;
        RECT 825.6800 2207.3600 827.2800 2207.8400 ;
        RECT 882.2200 2185.6000 885.2200 2186.0800 ;
        RECT 882.2200 2191.0400 885.2200 2191.5200 ;
        RECT 870.6800 2185.6000 872.2800 2186.0800 ;
        RECT 870.6800 2191.0400 872.2800 2191.5200 ;
        RECT 882.2200 2169.2800 885.2200 2169.7600 ;
        RECT 882.2200 2174.7200 885.2200 2175.2000 ;
        RECT 882.2200 2180.1600 885.2200 2180.6400 ;
        RECT 870.6800 2169.2800 872.2800 2169.7600 ;
        RECT 870.6800 2174.7200 872.2800 2175.2000 ;
        RECT 870.6800 2180.1600 872.2800 2180.6400 ;
        RECT 882.2200 2158.4000 885.2200 2158.8800 ;
        RECT 882.2200 2163.8400 885.2200 2164.3200 ;
        RECT 870.6800 2158.4000 872.2800 2158.8800 ;
        RECT 870.6800 2163.8400 872.2800 2164.3200 ;
        RECT 882.2200 2152.9600 885.2200 2153.4400 ;
        RECT 870.6800 2152.9600 872.2800 2153.4400 ;
        RECT 825.6800 2185.6000 827.2800 2186.0800 ;
        RECT 825.6800 2191.0400 827.2800 2191.5200 ;
        RECT 825.6800 2169.2800 827.2800 2169.7600 ;
        RECT 825.6800 2174.7200 827.2800 2175.2000 ;
        RECT 825.6800 2180.1600 827.2800 2180.6400 ;
        RECT 825.6800 2158.4000 827.2800 2158.8800 ;
        RECT 825.6800 2163.8400 827.2800 2164.3200 ;
        RECT 825.6800 2152.9600 827.2800 2153.4400 ;
        RECT 780.6800 2240.0000 782.2800 2240.4800 ;
        RECT 780.6800 2245.4400 782.2800 2245.9200 ;
        RECT 780.6800 2223.6800 782.2800 2224.1600 ;
        RECT 780.6800 2229.1200 782.2800 2229.6000 ;
        RECT 780.6800 2234.5600 782.2800 2235.0400 ;
        RECT 735.6800 2240.0000 737.2800 2240.4800 ;
        RECT 735.6800 2245.4400 737.2800 2245.9200 ;
        RECT 735.6800 2223.6800 737.2800 2224.1600 ;
        RECT 735.6800 2229.1200 737.2800 2229.6000 ;
        RECT 735.6800 2234.5600 737.2800 2235.0400 ;
        RECT 780.6800 2212.8000 782.2800 2213.2800 ;
        RECT 780.6800 2218.2400 782.2800 2218.7200 ;
        RECT 780.6800 2196.4800 782.2800 2196.9600 ;
        RECT 780.6800 2201.9200 782.2800 2202.4000 ;
        RECT 780.6800 2207.3600 782.2800 2207.8400 ;
        RECT 735.6800 2212.8000 737.2800 2213.2800 ;
        RECT 735.6800 2218.2400 737.2800 2218.7200 ;
        RECT 735.6800 2196.4800 737.2800 2196.9600 ;
        RECT 735.6800 2201.9200 737.2800 2202.4000 ;
        RECT 735.6800 2207.3600 737.2800 2207.8400 ;
        RECT 686.1200 2240.0000 689.1200 2240.4800 ;
        RECT 686.1200 2245.4400 689.1200 2245.9200 ;
        RECT 686.1200 2229.1200 689.1200 2229.6000 ;
        RECT 686.1200 2223.6800 689.1200 2224.1600 ;
        RECT 686.1200 2234.5600 689.1200 2235.0400 ;
        RECT 686.1200 2212.8000 689.1200 2213.2800 ;
        RECT 686.1200 2218.2400 689.1200 2218.7200 ;
        RECT 686.1200 2201.9200 689.1200 2202.4000 ;
        RECT 686.1200 2196.4800 689.1200 2196.9600 ;
        RECT 686.1200 2207.3600 689.1200 2207.8400 ;
        RECT 780.6800 2185.6000 782.2800 2186.0800 ;
        RECT 780.6800 2191.0400 782.2800 2191.5200 ;
        RECT 780.6800 2169.2800 782.2800 2169.7600 ;
        RECT 780.6800 2174.7200 782.2800 2175.2000 ;
        RECT 780.6800 2180.1600 782.2800 2180.6400 ;
        RECT 735.6800 2185.6000 737.2800 2186.0800 ;
        RECT 735.6800 2191.0400 737.2800 2191.5200 ;
        RECT 735.6800 2169.2800 737.2800 2169.7600 ;
        RECT 735.6800 2174.7200 737.2800 2175.2000 ;
        RECT 735.6800 2180.1600 737.2800 2180.6400 ;
        RECT 780.6800 2163.8400 782.2800 2164.3200 ;
        RECT 780.6800 2158.4000 782.2800 2158.8800 ;
        RECT 780.6800 2152.9600 782.2800 2153.4400 ;
        RECT 735.6800 2163.8400 737.2800 2164.3200 ;
        RECT 735.6800 2158.4000 737.2800 2158.8800 ;
        RECT 735.6800 2152.9600 737.2800 2153.4400 ;
        RECT 686.1200 2185.6000 689.1200 2186.0800 ;
        RECT 686.1200 2191.0400 689.1200 2191.5200 ;
        RECT 686.1200 2174.7200 689.1200 2175.2000 ;
        RECT 686.1200 2169.2800 689.1200 2169.7600 ;
        RECT 686.1200 2180.1600 689.1200 2180.6400 ;
        RECT 686.1200 2158.4000 689.1200 2158.8800 ;
        RECT 686.1200 2163.8400 689.1200 2164.3200 ;
        RECT 686.1200 2152.9600 689.1200 2153.4400 ;
        RECT 686.1200 2351.1500 885.2200 2354.1500 ;
        RECT 686.1200 2146.0500 885.2200 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 1916.4100 872.2800 2124.5100 ;
        RECT 825.6800 1916.4100 827.2800 2124.5100 ;
        RECT 780.6800 1916.4100 782.2800 2124.5100 ;
        RECT 735.6800 1916.4100 737.2800 2124.5100 ;
        RECT 882.2200 1916.4100 885.2200 2124.5100 ;
        RECT 686.1200 1916.4100 689.1200 2124.5100 ;
      LAYER met3 ;
        RECT 882.2200 2119.1600 885.2200 2119.6400 ;
        RECT 870.6800 2119.1600 872.2800 2119.6400 ;
        RECT 882.2200 2108.2800 885.2200 2108.7600 ;
        RECT 882.2200 2113.7200 885.2200 2114.2000 ;
        RECT 870.6800 2108.2800 872.2800 2108.7600 ;
        RECT 870.6800 2113.7200 872.2800 2114.2000 ;
        RECT 882.2200 2091.9600 885.2200 2092.4400 ;
        RECT 882.2200 2097.4000 885.2200 2097.8800 ;
        RECT 870.6800 2091.9600 872.2800 2092.4400 ;
        RECT 870.6800 2097.4000 872.2800 2097.8800 ;
        RECT 882.2200 2081.0800 885.2200 2081.5600 ;
        RECT 882.2200 2086.5200 885.2200 2087.0000 ;
        RECT 870.6800 2081.0800 872.2800 2081.5600 ;
        RECT 870.6800 2086.5200 872.2800 2087.0000 ;
        RECT 882.2200 2102.8400 885.2200 2103.3200 ;
        RECT 870.6800 2102.8400 872.2800 2103.3200 ;
        RECT 825.6800 2108.2800 827.2800 2108.7600 ;
        RECT 825.6800 2113.7200 827.2800 2114.2000 ;
        RECT 825.6800 2119.1600 827.2800 2119.6400 ;
        RECT 825.6800 2091.9600 827.2800 2092.4400 ;
        RECT 825.6800 2097.4000 827.2800 2097.8800 ;
        RECT 825.6800 2086.5200 827.2800 2087.0000 ;
        RECT 825.6800 2081.0800 827.2800 2081.5600 ;
        RECT 825.6800 2102.8400 827.2800 2103.3200 ;
        RECT 882.2200 2064.7600 885.2200 2065.2400 ;
        RECT 882.2200 2070.2000 885.2200 2070.6800 ;
        RECT 870.6800 2064.7600 872.2800 2065.2400 ;
        RECT 870.6800 2070.2000 872.2800 2070.6800 ;
        RECT 882.2200 2048.4400 885.2200 2048.9200 ;
        RECT 882.2200 2053.8800 885.2200 2054.3600 ;
        RECT 882.2200 2059.3200 885.2200 2059.8000 ;
        RECT 870.6800 2048.4400 872.2800 2048.9200 ;
        RECT 870.6800 2053.8800 872.2800 2054.3600 ;
        RECT 870.6800 2059.3200 872.2800 2059.8000 ;
        RECT 882.2200 2037.5600 885.2200 2038.0400 ;
        RECT 882.2200 2043.0000 885.2200 2043.4800 ;
        RECT 870.6800 2037.5600 872.2800 2038.0400 ;
        RECT 870.6800 2043.0000 872.2800 2043.4800 ;
        RECT 882.2200 2021.2400 885.2200 2021.7200 ;
        RECT 882.2200 2026.6800 885.2200 2027.1600 ;
        RECT 882.2200 2032.1200 885.2200 2032.6000 ;
        RECT 870.6800 2021.2400 872.2800 2021.7200 ;
        RECT 870.6800 2026.6800 872.2800 2027.1600 ;
        RECT 870.6800 2032.1200 872.2800 2032.6000 ;
        RECT 825.6800 2064.7600 827.2800 2065.2400 ;
        RECT 825.6800 2070.2000 827.2800 2070.6800 ;
        RECT 825.6800 2048.4400 827.2800 2048.9200 ;
        RECT 825.6800 2053.8800 827.2800 2054.3600 ;
        RECT 825.6800 2059.3200 827.2800 2059.8000 ;
        RECT 825.6800 2037.5600 827.2800 2038.0400 ;
        RECT 825.6800 2043.0000 827.2800 2043.4800 ;
        RECT 825.6800 2021.2400 827.2800 2021.7200 ;
        RECT 825.6800 2026.6800 827.2800 2027.1600 ;
        RECT 825.6800 2032.1200 827.2800 2032.6000 ;
        RECT 882.2200 2075.6400 885.2200 2076.1200 ;
        RECT 825.6800 2075.6400 827.2800 2076.1200 ;
        RECT 870.6800 2075.6400 872.2800 2076.1200 ;
        RECT 780.6800 2108.2800 782.2800 2108.7600 ;
        RECT 780.6800 2113.7200 782.2800 2114.2000 ;
        RECT 780.6800 2119.1600 782.2800 2119.6400 ;
        RECT 735.6800 2108.2800 737.2800 2108.7600 ;
        RECT 735.6800 2113.7200 737.2800 2114.2000 ;
        RECT 735.6800 2119.1600 737.2800 2119.6400 ;
        RECT 780.6800 2091.9600 782.2800 2092.4400 ;
        RECT 780.6800 2097.4000 782.2800 2097.8800 ;
        RECT 780.6800 2081.0800 782.2800 2081.5600 ;
        RECT 780.6800 2086.5200 782.2800 2087.0000 ;
        RECT 735.6800 2091.9600 737.2800 2092.4400 ;
        RECT 735.6800 2097.4000 737.2800 2097.8800 ;
        RECT 735.6800 2081.0800 737.2800 2081.5600 ;
        RECT 735.6800 2086.5200 737.2800 2087.0000 ;
        RECT 735.6800 2102.8400 737.2800 2103.3200 ;
        RECT 780.6800 2102.8400 782.2800 2103.3200 ;
        RECT 686.1200 2119.1600 689.1200 2119.6400 ;
        RECT 686.1200 2113.7200 689.1200 2114.2000 ;
        RECT 686.1200 2108.2800 689.1200 2108.7600 ;
        RECT 686.1200 2097.4000 689.1200 2097.8800 ;
        RECT 686.1200 2091.9600 689.1200 2092.4400 ;
        RECT 686.1200 2086.5200 689.1200 2087.0000 ;
        RECT 686.1200 2081.0800 689.1200 2081.5600 ;
        RECT 686.1200 2102.8400 689.1200 2103.3200 ;
        RECT 780.6800 2064.7600 782.2800 2065.2400 ;
        RECT 780.6800 2070.2000 782.2800 2070.6800 ;
        RECT 780.6800 2048.4400 782.2800 2048.9200 ;
        RECT 780.6800 2053.8800 782.2800 2054.3600 ;
        RECT 780.6800 2059.3200 782.2800 2059.8000 ;
        RECT 735.6800 2064.7600 737.2800 2065.2400 ;
        RECT 735.6800 2070.2000 737.2800 2070.6800 ;
        RECT 735.6800 2048.4400 737.2800 2048.9200 ;
        RECT 735.6800 2053.8800 737.2800 2054.3600 ;
        RECT 735.6800 2059.3200 737.2800 2059.8000 ;
        RECT 780.6800 2037.5600 782.2800 2038.0400 ;
        RECT 780.6800 2043.0000 782.2800 2043.4800 ;
        RECT 780.6800 2021.2400 782.2800 2021.7200 ;
        RECT 780.6800 2026.6800 782.2800 2027.1600 ;
        RECT 780.6800 2032.1200 782.2800 2032.6000 ;
        RECT 735.6800 2037.5600 737.2800 2038.0400 ;
        RECT 735.6800 2043.0000 737.2800 2043.4800 ;
        RECT 735.6800 2021.2400 737.2800 2021.7200 ;
        RECT 735.6800 2026.6800 737.2800 2027.1600 ;
        RECT 735.6800 2032.1200 737.2800 2032.6000 ;
        RECT 686.1200 2064.7600 689.1200 2065.2400 ;
        RECT 686.1200 2070.2000 689.1200 2070.6800 ;
        RECT 686.1200 2053.8800 689.1200 2054.3600 ;
        RECT 686.1200 2048.4400 689.1200 2048.9200 ;
        RECT 686.1200 2059.3200 689.1200 2059.8000 ;
        RECT 686.1200 2037.5600 689.1200 2038.0400 ;
        RECT 686.1200 2043.0000 689.1200 2043.4800 ;
        RECT 686.1200 2026.6800 689.1200 2027.1600 ;
        RECT 686.1200 2021.2400 689.1200 2021.7200 ;
        RECT 686.1200 2032.1200 689.1200 2032.6000 ;
        RECT 686.1200 2075.6400 689.1200 2076.1200 ;
        RECT 735.6800 2075.6400 737.2800 2076.1200 ;
        RECT 780.6800 2075.6400 782.2800 2076.1200 ;
        RECT 882.2200 2010.3600 885.2200 2010.8400 ;
        RECT 882.2200 2015.8000 885.2200 2016.2800 ;
        RECT 870.6800 2010.3600 872.2800 2010.8400 ;
        RECT 870.6800 2015.8000 872.2800 2016.2800 ;
        RECT 882.2200 1994.0400 885.2200 1994.5200 ;
        RECT 882.2200 1999.4800 885.2200 1999.9600 ;
        RECT 882.2200 2004.9200 885.2200 2005.4000 ;
        RECT 870.6800 1994.0400 872.2800 1994.5200 ;
        RECT 870.6800 1999.4800 872.2800 1999.9600 ;
        RECT 870.6800 2004.9200 872.2800 2005.4000 ;
        RECT 882.2200 1983.1600 885.2200 1983.6400 ;
        RECT 882.2200 1988.6000 885.2200 1989.0800 ;
        RECT 870.6800 1983.1600 872.2800 1983.6400 ;
        RECT 870.6800 1988.6000 872.2800 1989.0800 ;
        RECT 882.2200 1966.8400 885.2200 1967.3200 ;
        RECT 882.2200 1972.2800 885.2200 1972.7600 ;
        RECT 882.2200 1977.7200 885.2200 1978.2000 ;
        RECT 870.6800 1966.8400 872.2800 1967.3200 ;
        RECT 870.6800 1972.2800 872.2800 1972.7600 ;
        RECT 870.6800 1977.7200 872.2800 1978.2000 ;
        RECT 825.6800 2010.3600 827.2800 2010.8400 ;
        RECT 825.6800 2015.8000 827.2800 2016.2800 ;
        RECT 825.6800 1994.0400 827.2800 1994.5200 ;
        RECT 825.6800 1999.4800 827.2800 1999.9600 ;
        RECT 825.6800 2004.9200 827.2800 2005.4000 ;
        RECT 825.6800 1983.1600 827.2800 1983.6400 ;
        RECT 825.6800 1988.6000 827.2800 1989.0800 ;
        RECT 825.6800 1966.8400 827.2800 1967.3200 ;
        RECT 825.6800 1972.2800 827.2800 1972.7600 ;
        RECT 825.6800 1977.7200 827.2800 1978.2000 ;
        RECT 882.2200 1955.9600 885.2200 1956.4400 ;
        RECT 882.2200 1961.4000 885.2200 1961.8800 ;
        RECT 870.6800 1955.9600 872.2800 1956.4400 ;
        RECT 870.6800 1961.4000 872.2800 1961.8800 ;
        RECT 882.2200 1939.6400 885.2200 1940.1200 ;
        RECT 882.2200 1945.0800 885.2200 1945.5600 ;
        RECT 882.2200 1950.5200 885.2200 1951.0000 ;
        RECT 870.6800 1939.6400 872.2800 1940.1200 ;
        RECT 870.6800 1945.0800 872.2800 1945.5600 ;
        RECT 870.6800 1950.5200 872.2800 1951.0000 ;
        RECT 882.2200 1928.7600 885.2200 1929.2400 ;
        RECT 882.2200 1934.2000 885.2200 1934.6800 ;
        RECT 870.6800 1928.7600 872.2800 1929.2400 ;
        RECT 870.6800 1934.2000 872.2800 1934.6800 ;
        RECT 882.2200 1923.3200 885.2200 1923.8000 ;
        RECT 870.6800 1923.3200 872.2800 1923.8000 ;
        RECT 825.6800 1955.9600 827.2800 1956.4400 ;
        RECT 825.6800 1961.4000 827.2800 1961.8800 ;
        RECT 825.6800 1939.6400 827.2800 1940.1200 ;
        RECT 825.6800 1945.0800 827.2800 1945.5600 ;
        RECT 825.6800 1950.5200 827.2800 1951.0000 ;
        RECT 825.6800 1928.7600 827.2800 1929.2400 ;
        RECT 825.6800 1934.2000 827.2800 1934.6800 ;
        RECT 825.6800 1923.3200 827.2800 1923.8000 ;
        RECT 780.6800 2010.3600 782.2800 2010.8400 ;
        RECT 780.6800 2015.8000 782.2800 2016.2800 ;
        RECT 780.6800 1994.0400 782.2800 1994.5200 ;
        RECT 780.6800 1999.4800 782.2800 1999.9600 ;
        RECT 780.6800 2004.9200 782.2800 2005.4000 ;
        RECT 735.6800 2010.3600 737.2800 2010.8400 ;
        RECT 735.6800 2015.8000 737.2800 2016.2800 ;
        RECT 735.6800 1994.0400 737.2800 1994.5200 ;
        RECT 735.6800 1999.4800 737.2800 1999.9600 ;
        RECT 735.6800 2004.9200 737.2800 2005.4000 ;
        RECT 780.6800 1983.1600 782.2800 1983.6400 ;
        RECT 780.6800 1988.6000 782.2800 1989.0800 ;
        RECT 780.6800 1966.8400 782.2800 1967.3200 ;
        RECT 780.6800 1972.2800 782.2800 1972.7600 ;
        RECT 780.6800 1977.7200 782.2800 1978.2000 ;
        RECT 735.6800 1983.1600 737.2800 1983.6400 ;
        RECT 735.6800 1988.6000 737.2800 1989.0800 ;
        RECT 735.6800 1966.8400 737.2800 1967.3200 ;
        RECT 735.6800 1972.2800 737.2800 1972.7600 ;
        RECT 735.6800 1977.7200 737.2800 1978.2000 ;
        RECT 686.1200 2010.3600 689.1200 2010.8400 ;
        RECT 686.1200 2015.8000 689.1200 2016.2800 ;
        RECT 686.1200 1999.4800 689.1200 1999.9600 ;
        RECT 686.1200 1994.0400 689.1200 1994.5200 ;
        RECT 686.1200 2004.9200 689.1200 2005.4000 ;
        RECT 686.1200 1983.1600 689.1200 1983.6400 ;
        RECT 686.1200 1988.6000 689.1200 1989.0800 ;
        RECT 686.1200 1972.2800 689.1200 1972.7600 ;
        RECT 686.1200 1966.8400 689.1200 1967.3200 ;
        RECT 686.1200 1977.7200 689.1200 1978.2000 ;
        RECT 780.6800 1955.9600 782.2800 1956.4400 ;
        RECT 780.6800 1961.4000 782.2800 1961.8800 ;
        RECT 780.6800 1939.6400 782.2800 1940.1200 ;
        RECT 780.6800 1945.0800 782.2800 1945.5600 ;
        RECT 780.6800 1950.5200 782.2800 1951.0000 ;
        RECT 735.6800 1955.9600 737.2800 1956.4400 ;
        RECT 735.6800 1961.4000 737.2800 1961.8800 ;
        RECT 735.6800 1939.6400 737.2800 1940.1200 ;
        RECT 735.6800 1945.0800 737.2800 1945.5600 ;
        RECT 735.6800 1950.5200 737.2800 1951.0000 ;
        RECT 780.6800 1934.2000 782.2800 1934.6800 ;
        RECT 780.6800 1928.7600 782.2800 1929.2400 ;
        RECT 780.6800 1923.3200 782.2800 1923.8000 ;
        RECT 735.6800 1934.2000 737.2800 1934.6800 ;
        RECT 735.6800 1928.7600 737.2800 1929.2400 ;
        RECT 735.6800 1923.3200 737.2800 1923.8000 ;
        RECT 686.1200 1955.9600 689.1200 1956.4400 ;
        RECT 686.1200 1961.4000 689.1200 1961.8800 ;
        RECT 686.1200 1945.0800 689.1200 1945.5600 ;
        RECT 686.1200 1939.6400 689.1200 1940.1200 ;
        RECT 686.1200 1950.5200 689.1200 1951.0000 ;
        RECT 686.1200 1928.7600 689.1200 1929.2400 ;
        RECT 686.1200 1934.2000 689.1200 1934.6800 ;
        RECT 686.1200 1923.3200 689.1200 1923.8000 ;
        RECT 686.1200 2121.5100 885.2200 2124.5100 ;
        RECT 686.1200 1916.4100 885.2200 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 1686.7700 872.2800 1894.8700 ;
        RECT 825.6800 1686.7700 827.2800 1894.8700 ;
        RECT 780.6800 1686.7700 782.2800 1894.8700 ;
        RECT 735.6800 1686.7700 737.2800 1894.8700 ;
        RECT 882.2200 1686.7700 885.2200 1894.8700 ;
        RECT 686.1200 1686.7700 689.1200 1894.8700 ;
      LAYER met3 ;
        RECT 882.2200 1889.5200 885.2200 1890.0000 ;
        RECT 870.6800 1889.5200 872.2800 1890.0000 ;
        RECT 882.2200 1878.6400 885.2200 1879.1200 ;
        RECT 882.2200 1884.0800 885.2200 1884.5600 ;
        RECT 870.6800 1878.6400 872.2800 1879.1200 ;
        RECT 870.6800 1884.0800 872.2800 1884.5600 ;
        RECT 882.2200 1862.3200 885.2200 1862.8000 ;
        RECT 882.2200 1867.7600 885.2200 1868.2400 ;
        RECT 870.6800 1862.3200 872.2800 1862.8000 ;
        RECT 870.6800 1867.7600 872.2800 1868.2400 ;
        RECT 882.2200 1851.4400 885.2200 1851.9200 ;
        RECT 882.2200 1856.8800 885.2200 1857.3600 ;
        RECT 870.6800 1851.4400 872.2800 1851.9200 ;
        RECT 870.6800 1856.8800 872.2800 1857.3600 ;
        RECT 882.2200 1873.2000 885.2200 1873.6800 ;
        RECT 870.6800 1873.2000 872.2800 1873.6800 ;
        RECT 825.6800 1878.6400 827.2800 1879.1200 ;
        RECT 825.6800 1884.0800 827.2800 1884.5600 ;
        RECT 825.6800 1889.5200 827.2800 1890.0000 ;
        RECT 825.6800 1862.3200 827.2800 1862.8000 ;
        RECT 825.6800 1867.7600 827.2800 1868.2400 ;
        RECT 825.6800 1856.8800 827.2800 1857.3600 ;
        RECT 825.6800 1851.4400 827.2800 1851.9200 ;
        RECT 825.6800 1873.2000 827.2800 1873.6800 ;
        RECT 882.2200 1835.1200 885.2200 1835.6000 ;
        RECT 882.2200 1840.5600 885.2200 1841.0400 ;
        RECT 870.6800 1835.1200 872.2800 1835.6000 ;
        RECT 870.6800 1840.5600 872.2800 1841.0400 ;
        RECT 882.2200 1818.8000 885.2200 1819.2800 ;
        RECT 882.2200 1824.2400 885.2200 1824.7200 ;
        RECT 882.2200 1829.6800 885.2200 1830.1600 ;
        RECT 870.6800 1818.8000 872.2800 1819.2800 ;
        RECT 870.6800 1824.2400 872.2800 1824.7200 ;
        RECT 870.6800 1829.6800 872.2800 1830.1600 ;
        RECT 882.2200 1807.9200 885.2200 1808.4000 ;
        RECT 882.2200 1813.3600 885.2200 1813.8400 ;
        RECT 870.6800 1807.9200 872.2800 1808.4000 ;
        RECT 870.6800 1813.3600 872.2800 1813.8400 ;
        RECT 882.2200 1791.6000 885.2200 1792.0800 ;
        RECT 882.2200 1797.0400 885.2200 1797.5200 ;
        RECT 882.2200 1802.4800 885.2200 1802.9600 ;
        RECT 870.6800 1791.6000 872.2800 1792.0800 ;
        RECT 870.6800 1797.0400 872.2800 1797.5200 ;
        RECT 870.6800 1802.4800 872.2800 1802.9600 ;
        RECT 825.6800 1835.1200 827.2800 1835.6000 ;
        RECT 825.6800 1840.5600 827.2800 1841.0400 ;
        RECT 825.6800 1818.8000 827.2800 1819.2800 ;
        RECT 825.6800 1824.2400 827.2800 1824.7200 ;
        RECT 825.6800 1829.6800 827.2800 1830.1600 ;
        RECT 825.6800 1807.9200 827.2800 1808.4000 ;
        RECT 825.6800 1813.3600 827.2800 1813.8400 ;
        RECT 825.6800 1791.6000 827.2800 1792.0800 ;
        RECT 825.6800 1797.0400 827.2800 1797.5200 ;
        RECT 825.6800 1802.4800 827.2800 1802.9600 ;
        RECT 882.2200 1846.0000 885.2200 1846.4800 ;
        RECT 825.6800 1846.0000 827.2800 1846.4800 ;
        RECT 870.6800 1846.0000 872.2800 1846.4800 ;
        RECT 780.6800 1878.6400 782.2800 1879.1200 ;
        RECT 780.6800 1884.0800 782.2800 1884.5600 ;
        RECT 780.6800 1889.5200 782.2800 1890.0000 ;
        RECT 735.6800 1878.6400 737.2800 1879.1200 ;
        RECT 735.6800 1884.0800 737.2800 1884.5600 ;
        RECT 735.6800 1889.5200 737.2800 1890.0000 ;
        RECT 780.6800 1862.3200 782.2800 1862.8000 ;
        RECT 780.6800 1867.7600 782.2800 1868.2400 ;
        RECT 780.6800 1851.4400 782.2800 1851.9200 ;
        RECT 780.6800 1856.8800 782.2800 1857.3600 ;
        RECT 735.6800 1862.3200 737.2800 1862.8000 ;
        RECT 735.6800 1867.7600 737.2800 1868.2400 ;
        RECT 735.6800 1851.4400 737.2800 1851.9200 ;
        RECT 735.6800 1856.8800 737.2800 1857.3600 ;
        RECT 735.6800 1873.2000 737.2800 1873.6800 ;
        RECT 780.6800 1873.2000 782.2800 1873.6800 ;
        RECT 686.1200 1889.5200 689.1200 1890.0000 ;
        RECT 686.1200 1884.0800 689.1200 1884.5600 ;
        RECT 686.1200 1878.6400 689.1200 1879.1200 ;
        RECT 686.1200 1867.7600 689.1200 1868.2400 ;
        RECT 686.1200 1862.3200 689.1200 1862.8000 ;
        RECT 686.1200 1856.8800 689.1200 1857.3600 ;
        RECT 686.1200 1851.4400 689.1200 1851.9200 ;
        RECT 686.1200 1873.2000 689.1200 1873.6800 ;
        RECT 780.6800 1835.1200 782.2800 1835.6000 ;
        RECT 780.6800 1840.5600 782.2800 1841.0400 ;
        RECT 780.6800 1818.8000 782.2800 1819.2800 ;
        RECT 780.6800 1824.2400 782.2800 1824.7200 ;
        RECT 780.6800 1829.6800 782.2800 1830.1600 ;
        RECT 735.6800 1835.1200 737.2800 1835.6000 ;
        RECT 735.6800 1840.5600 737.2800 1841.0400 ;
        RECT 735.6800 1818.8000 737.2800 1819.2800 ;
        RECT 735.6800 1824.2400 737.2800 1824.7200 ;
        RECT 735.6800 1829.6800 737.2800 1830.1600 ;
        RECT 780.6800 1807.9200 782.2800 1808.4000 ;
        RECT 780.6800 1813.3600 782.2800 1813.8400 ;
        RECT 780.6800 1791.6000 782.2800 1792.0800 ;
        RECT 780.6800 1797.0400 782.2800 1797.5200 ;
        RECT 780.6800 1802.4800 782.2800 1802.9600 ;
        RECT 735.6800 1807.9200 737.2800 1808.4000 ;
        RECT 735.6800 1813.3600 737.2800 1813.8400 ;
        RECT 735.6800 1791.6000 737.2800 1792.0800 ;
        RECT 735.6800 1797.0400 737.2800 1797.5200 ;
        RECT 735.6800 1802.4800 737.2800 1802.9600 ;
        RECT 686.1200 1835.1200 689.1200 1835.6000 ;
        RECT 686.1200 1840.5600 689.1200 1841.0400 ;
        RECT 686.1200 1824.2400 689.1200 1824.7200 ;
        RECT 686.1200 1818.8000 689.1200 1819.2800 ;
        RECT 686.1200 1829.6800 689.1200 1830.1600 ;
        RECT 686.1200 1807.9200 689.1200 1808.4000 ;
        RECT 686.1200 1813.3600 689.1200 1813.8400 ;
        RECT 686.1200 1797.0400 689.1200 1797.5200 ;
        RECT 686.1200 1791.6000 689.1200 1792.0800 ;
        RECT 686.1200 1802.4800 689.1200 1802.9600 ;
        RECT 686.1200 1846.0000 689.1200 1846.4800 ;
        RECT 735.6800 1846.0000 737.2800 1846.4800 ;
        RECT 780.6800 1846.0000 782.2800 1846.4800 ;
        RECT 882.2200 1780.7200 885.2200 1781.2000 ;
        RECT 882.2200 1786.1600 885.2200 1786.6400 ;
        RECT 870.6800 1780.7200 872.2800 1781.2000 ;
        RECT 870.6800 1786.1600 872.2800 1786.6400 ;
        RECT 882.2200 1764.4000 885.2200 1764.8800 ;
        RECT 882.2200 1769.8400 885.2200 1770.3200 ;
        RECT 882.2200 1775.2800 885.2200 1775.7600 ;
        RECT 870.6800 1764.4000 872.2800 1764.8800 ;
        RECT 870.6800 1769.8400 872.2800 1770.3200 ;
        RECT 870.6800 1775.2800 872.2800 1775.7600 ;
        RECT 882.2200 1753.5200 885.2200 1754.0000 ;
        RECT 882.2200 1758.9600 885.2200 1759.4400 ;
        RECT 870.6800 1753.5200 872.2800 1754.0000 ;
        RECT 870.6800 1758.9600 872.2800 1759.4400 ;
        RECT 882.2200 1737.2000 885.2200 1737.6800 ;
        RECT 882.2200 1742.6400 885.2200 1743.1200 ;
        RECT 882.2200 1748.0800 885.2200 1748.5600 ;
        RECT 870.6800 1737.2000 872.2800 1737.6800 ;
        RECT 870.6800 1742.6400 872.2800 1743.1200 ;
        RECT 870.6800 1748.0800 872.2800 1748.5600 ;
        RECT 825.6800 1780.7200 827.2800 1781.2000 ;
        RECT 825.6800 1786.1600 827.2800 1786.6400 ;
        RECT 825.6800 1764.4000 827.2800 1764.8800 ;
        RECT 825.6800 1769.8400 827.2800 1770.3200 ;
        RECT 825.6800 1775.2800 827.2800 1775.7600 ;
        RECT 825.6800 1753.5200 827.2800 1754.0000 ;
        RECT 825.6800 1758.9600 827.2800 1759.4400 ;
        RECT 825.6800 1737.2000 827.2800 1737.6800 ;
        RECT 825.6800 1742.6400 827.2800 1743.1200 ;
        RECT 825.6800 1748.0800 827.2800 1748.5600 ;
        RECT 882.2200 1726.3200 885.2200 1726.8000 ;
        RECT 882.2200 1731.7600 885.2200 1732.2400 ;
        RECT 870.6800 1726.3200 872.2800 1726.8000 ;
        RECT 870.6800 1731.7600 872.2800 1732.2400 ;
        RECT 882.2200 1710.0000 885.2200 1710.4800 ;
        RECT 882.2200 1715.4400 885.2200 1715.9200 ;
        RECT 882.2200 1720.8800 885.2200 1721.3600 ;
        RECT 870.6800 1710.0000 872.2800 1710.4800 ;
        RECT 870.6800 1715.4400 872.2800 1715.9200 ;
        RECT 870.6800 1720.8800 872.2800 1721.3600 ;
        RECT 882.2200 1699.1200 885.2200 1699.6000 ;
        RECT 882.2200 1704.5600 885.2200 1705.0400 ;
        RECT 870.6800 1699.1200 872.2800 1699.6000 ;
        RECT 870.6800 1704.5600 872.2800 1705.0400 ;
        RECT 882.2200 1693.6800 885.2200 1694.1600 ;
        RECT 870.6800 1693.6800 872.2800 1694.1600 ;
        RECT 825.6800 1726.3200 827.2800 1726.8000 ;
        RECT 825.6800 1731.7600 827.2800 1732.2400 ;
        RECT 825.6800 1710.0000 827.2800 1710.4800 ;
        RECT 825.6800 1715.4400 827.2800 1715.9200 ;
        RECT 825.6800 1720.8800 827.2800 1721.3600 ;
        RECT 825.6800 1699.1200 827.2800 1699.6000 ;
        RECT 825.6800 1704.5600 827.2800 1705.0400 ;
        RECT 825.6800 1693.6800 827.2800 1694.1600 ;
        RECT 780.6800 1780.7200 782.2800 1781.2000 ;
        RECT 780.6800 1786.1600 782.2800 1786.6400 ;
        RECT 780.6800 1764.4000 782.2800 1764.8800 ;
        RECT 780.6800 1769.8400 782.2800 1770.3200 ;
        RECT 780.6800 1775.2800 782.2800 1775.7600 ;
        RECT 735.6800 1780.7200 737.2800 1781.2000 ;
        RECT 735.6800 1786.1600 737.2800 1786.6400 ;
        RECT 735.6800 1764.4000 737.2800 1764.8800 ;
        RECT 735.6800 1769.8400 737.2800 1770.3200 ;
        RECT 735.6800 1775.2800 737.2800 1775.7600 ;
        RECT 780.6800 1753.5200 782.2800 1754.0000 ;
        RECT 780.6800 1758.9600 782.2800 1759.4400 ;
        RECT 780.6800 1737.2000 782.2800 1737.6800 ;
        RECT 780.6800 1742.6400 782.2800 1743.1200 ;
        RECT 780.6800 1748.0800 782.2800 1748.5600 ;
        RECT 735.6800 1753.5200 737.2800 1754.0000 ;
        RECT 735.6800 1758.9600 737.2800 1759.4400 ;
        RECT 735.6800 1737.2000 737.2800 1737.6800 ;
        RECT 735.6800 1742.6400 737.2800 1743.1200 ;
        RECT 735.6800 1748.0800 737.2800 1748.5600 ;
        RECT 686.1200 1780.7200 689.1200 1781.2000 ;
        RECT 686.1200 1786.1600 689.1200 1786.6400 ;
        RECT 686.1200 1769.8400 689.1200 1770.3200 ;
        RECT 686.1200 1764.4000 689.1200 1764.8800 ;
        RECT 686.1200 1775.2800 689.1200 1775.7600 ;
        RECT 686.1200 1753.5200 689.1200 1754.0000 ;
        RECT 686.1200 1758.9600 689.1200 1759.4400 ;
        RECT 686.1200 1742.6400 689.1200 1743.1200 ;
        RECT 686.1200 1737.2000 689.1200 1737.6800 ;
        RECT 686.1200 1748.0800 689.1200 1748.5600 ;
        RECT 780.6800 1726.3200 782.2800 1726.8000 ;
        RECT 780.6800 1731.7600 782.2800 1732.2400 ;
        RECT 780.6800 1710.0000 782.2800 1710.4800 ;
        RECT 780.6800 1715.4400 782.2800 1715.9200 ;
        RECT 780.6800 1720.8800 782.2800 1721.3600 ;
        RECT 735.6800 1726.3200 737.2800 1726.8000 ;
        RECT 735.6800 1731.7600 737.2800 1732.2400 ;
        RECT 735.6800 1710.0000 737.2800 1710.4800 ;
        RECT 735.6800 1715.4400 737.2800 1715.9200 ;
        RECT 735.6800 1720.8800 737.2800 1721.3600 ;
        RECT 780.6800 1704.5600 782.2800 1705.0400 ;
        RECT 780.6800 1699.1200 782.2800 1699.6000 ;
        RECT 780.6800 1693.6800 782.2800 1694.1600 ;
        RECT 735.6800 1704.5600 737.2800 1705.0400 ;
        RECT 735.6800 1699.1200 737.2800 1699.6000 ;
        RECT 735.6800 1693.6800 737.2800 1694.1600 ;
        RECT 686.1200 1726.3200 689.1200 1726.8000 ;
        RECT 686.1200 1731.7600 689.1200 1732.2400 ;
        RECT 686.1200 1715.4400 689.1200 1715.9200 ;
        RECT 686.1200 1710.0000 689.1200 1710.4800 ;
        RECT 686.1200 1720.8800 689.1200 1721.3600 ;
        RECT 686.1200 1699.1200 689.1200 1699.6000 ;
        RECT 686.1200 1704.5600 689.1200 1705.0400 ;
        RECT 686.1200 1693.6800 689.1200 1694.1600 ;
        RECT 686.1200 1891.8700 885.2200 1894.8700 ;
        RECT 686.1200 1686.7700 885.2200 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 1457.1300 872.2800 1665.2300 ;
        RECT 825.6800 1457.1300 827.2800 1665.2300 ;
        RECT 780.6800 1457.1300 782.2800 1665.2300 ;
        RECT 735.6800 1457.1300 737.2800 1665.2300 ;
        RECT 882.2200 1457.1300 885.2200 1665.2300 ;
        RECT 686.1200 1457.1300 689.1200 1665.2300 ;
      LAYER met3 ;
        RECT 882.2200 1659.8800 885.2200 1660.3600 ;
        RECT 870.6800 1659.8800 872.2800 1660.3600 ;
        RECT 882.2200 1649.0000 885.2200 1649.4800 ;
        RECT 882.2200 1654.4400 885.2200 1654.9200 ;
        RECT 870.6800 1649.0000 872.2800 1649.4800 ;
        RECT 870.6800 1654.4400 872.2800 1654.9200 ;
        RECT 882.2200 1632.6800 885.2200 1633.1600 ;
        RECT 882.2200 1638.1200 885.2200 1638.6000 ;
        RECT 870.6800 1632.6800 872.2800 1633.1600 ;
        RECT 870.6800 1638.1200 872.2800 1638.6000 ;
        RECT 882.2200 1621.8000 885.2200 1622.2800 ;
        RECT 882.2200 1627.2400 885.2200 1627.7200 ;
        RECT 870.6800 1621.8000 872.2800 1622.2800 ;
        RECT 870.6800 1627.2400 872.2800 1627.7200 ;
        RECT 882.2200 1643.5600 885.2200 1644.0400 ;
        RECT 870.6800 1643.5600 872.2800 1644.0400 ;
        RECT 825.6800 1649.0000 827.2800 1649.4800 ;
        RECT 825.6800 1654.4400 827.2800 1654.9200 ;
        RECT 825.6800 1659.8800 827.2800 1660.3600 ;
        RECT 825.6800 1632.6800 827.2800 1633.1600 ;
        RECT 825.6800 1638.1200 827.2800 1638.6000 ;
        RECT 825.6800 1627.2400 827.2800 1627.7200 ;
        RECT 825.6800 1621.8000 827.2800 1622.2800 ;
        RECT 825.6800 1643.5600 827.2800 1644.0400 ;
        RECT 882.2200 1605.4800 885.2200 1605.9600 ;
        RECT 882.2200 1610.9200 885.2200 1611.4000 ;
        RECT 870.6800 1605.4800 872.2800 1605.9600 ;
        RECT 870.6800 1610.9200 872.2800 1611.4000 ;
        RECT 882.2200 1589.1600 885.2200 1589.6400 ;
        RECT 882.2200 1594.6000 885.2200 1595.0800 ;
        RECT 882.2200 1600.0400 885.2200 1600.5200 ;
        RECT 870.6800 1589.1600 872.2800 1589.6400 ;
        RECT 870.6800 1594.6000 872.2800 1595.0800 ;
        RECT 870.6800 1600.0400 872.2800 1600.5200 ;
        RECT 882.2200 1578.2800 885.2200 1578.7600 ;
        RECT 882.2200 1583.7200 885.2200 1584.2000 ;
        RECT 870.6800 1578.2800 872.2800 1578.7600 ;
        RECT 870.6800 1583.7200 872.2800 1584.2000 ;
        RECT 882.2200 1561.9600 885.2200 1562.4400 ;
        RECT 882.2200 1567.4000 885.2200 1567.8800 ;
        RECT 882.2200 1572.8400 885.2200 1573.3200 ;
        RECT 870.6800 1561.9600 872.2800 1562.4400 ;
        RECT 870.6800 1567.4000 872.2800 1567.8800 ;
        RECT 870.6800 1572.8400 872.2800 1573.3200 ;
        RECT 825.6800 1605.4800 827.2800 1605.9600 ;
        RECT 825.6800 1610.9200 827.2800 1611.4000 ;
        RECT 825.6800 1589.1600 827.2800 1589.6400 ;
        RECT 825.6800 1594.6000 827.2800 1595.0800 ;
        RECT 825.6800 1600.0400 827.2800 1600.5200 ;
        RECT 825.6800 1578.2800 827.2800 1578.7600 ;
        RECT 825.6800 1583.7200 827.2800 1584.2000 ;
        RECT 825.6800 1561.9600 827.2800 1562.4400 ;
        RECT 825.6800 1567.4000 827.2800 1567.8800 ;
        RECT 825.6800 1572.8400 827.2800 1573.3200 ;
        RECT 882.2200 1616.3600 885.2200 1616.8400 ;
        RECT 825.6800 1616.3600 827.2800 1616.8400 ;
        RECT 870.6800 1616.3600 872.2800 1616.8400 ;
        RECT 780.6800 1649.0000 782.2800 1649.4800 ;
        RECT 780.6800 1654.4400 782.2800 1654.9200 ;
        RECT 780.6800 1659.8800 782.2800 1660.3600 ;
        RECT 735.6800 1649.0000 737.2800 1649.4800 ;
        RECT 735.6800 1654.4400 737.2800 1654.9200 ;
        RECT 735.6800 1659.8800 737.2800 1660.3600 ;
        RECT 780.6800 1632.6800 782.2800 1633.1600 ;
        RECT 780.6800 1638.1200 782.2800 1638.6000 ;
        RECT 780.6800 1621.8000 782.2800 1622.2800 ;
        RECT 780.6800 1627.2400 782.2800 1627.7200 ;
        RECT 735.6800 1632.6800 737.2800 1633.1600 ;
        RECT 735.6800 1638.1200 737.2800 1638.6000 ;
        RECT 735.6800 1621.8000 737.2800 1622.2800 ;
        RECT 735.6800 1627.2400 737.2800 1627.7200 ;
        RECT 735.6800 1643.5600 737.2800 1644.0400 ;
        RECT 780.6800 1643.5600 782.2800 1644.0400 ;
        RECT 686.1200 1659.8800 689.1200 1660.3600 ;
        RECT 686.1200 1654.4400 689.1200 1654.9200 ;
        RECT 686.1200 1649.0000 689.1200 1649.4800 ;
        RECT 686.1200 1638.1200 689.1200 1638.6000 ;
        RECT 686.1200 1632.6800 689.1200 1633.1600 ;
        RECT 686.1200 1627.2400 689.1200 1627.7200 ;
        RECT 686.1200 1621.8000 689.1200 1622.2800 ;
        RECT 686.1200 1643.5600 689.1200 1644.0400 ;
        RECT 780.6800 1605.4800 782.2800 1605.9600 ;
        RECT 780.6800 1610.9200 782.2800 1611.4000 ;
        RECT 780.6800 1589.1600 782.2800 1589.6400 ;
        RECT 780.6800 1594.6000 782.2800 1595.0800 ;
        RECT 780.6800 1600.0400 782.2800 1600.5200 ;
        RECT 735.6800 1605.4800 737.2800 1605.9600 ;
        RECT 735.6800 1610.9200 737.2800 1611.4000 ;
        RECT 735.6800 1589.1600 737.2800 1589.6400 ;
        RECT 735.6800 1594.6000 737.2800 1595.0800 ;
        RECT 735.6800 1600.0400 737.2800 1600.5200 ;
        RECT 780.6800 1578.2800 782.2800 1578.7600 ;
        RECT 780.6800 1583.7200 782.2800 1584.2000 ;
        RECT 780.6800 1561.9600 782.2800 1562.4400 ;
        RECT 780.6800 1567.4000 782.2800 1567.8800 ;
        RECT 780.6800 1572.8400 782.2800 1573.3200 ;
        RECT 735.6800 1578.2800 737.2800 1578.7600 ;
        RECT 735.6800 1583.7200 737.2800 1584.2000 ;
        RECT 735.6800 1561.9600 737.2800 1562.4400 ;
        RECT 735.6800 1567.4000 737.2800 1567.8800 ;
        RECT 735.6800 1572.8400 737.2800 1573.3200 ;
        RECT 686.1200 1605.4800 689.1200 1605.9600 ;
        RECT 686.1200 1610.9200 689.1200 1611.4000 ;
        RECT 686.1200 1594.6000 689.1200 1595.0800 ;
        RECT 686.1200 1589.1600 689.1200 1589.6400 ;
        RECT 686.1200 1600.0400 689.1200 1600.5200 ;
        RECT 686.1200 1578.2800 689.1200 1578.7600 ;
        RECT 686.1200 1583.7200 689.1200 1584.2000 ;
        RECT 686.1200 1567.4000 689.1200 1567.8800 ;
        RECT 686.1200 1561.9600 689.1200 1562.4400 ;
        RECT 686.1200 1572.8400 689.1200 1573.3200 ;
        RECT 686.1200 1616.3600 689.1200 1616.8400 ;
        RECT 735.6800 1616.3600 737.2800 1616.8400 ;
        RECT 780.6800 1616.3600 782.2800 1616.8400 ;
        RECT 882.2200 1551.0800 885.2200 1551.5600 ;
        RECT 882.2200 1556.5200 885.2200 1557.0000 ;
        RECT 870.6800 1551.0800 872.2800 1551.5600 ;
        RECT 870.6800 1556.5200 872.2800 1557.0000 ;
        RECT 882.2200 1534.7600 885.2200 1535.2400 ;
        RECT 882.2200 1540.2000 885.2200 1540.6800 ;
        RECT 882.2200 1545.6400 885.2200 1546.1200 ;
        RECT 870.6800 1534.7600 872.2800 1535.2400 ;
        RECT 870.6800 1540.2000 872.2800 1540.6800 ;
        RECT 870.6800 1545.6400 872.2800 1546.1200 ;
        RECT 882.2200 1523.8800 885.2200 1524.3600 ;
        RECT 882.2200 1529.3200 885.2200 1529.8000 ;
        RECT 870.6800 1523.8800 872.2800 1524.3600 ;
        RECT 870.6800 1529.3200 872.2800 1529.8000 ;
        RECT 882.2200 1507.5600 885.2200 1508.0400 ;
        RECT 882.2200 1513.0000 885.2200 1513.4800 ;
        RECT 882.2200 1518.4400 885.2200 1518.9200 ;
        RECT 870.6800 1507.5600 872.2800 1508.0400 ;
        RECT 870.6800 1513.0000 872.2800 1513.4800 ;
        RECT 870.6800 1518.4400 872.2800 1518.9200 ;
        RECT 825.6800 1551.0800 827.2800 1551.5600 ;
        RECT 825.6800 1556.5200 827.2800 1557.0000 ;
        RECT 825.6800 1534.7600 827.2800 1535.2400 ;
        RECT 825.6800 1540.2000 827.2800 1540.6800 ;
        RECT 825.6800 1545.6400 827.2800 1546.1200 ;
        RECT 825.6800 1523.8800 827.2800 1524.3600 ;
        RECT 825.6800 1529.3200 827.2800 1529.8000 ;
        RECT 825.6800 1507.5600 827.2800 1508.0400 ;
        RECT 825.6800 1513.0000 827.2800 1513.4800 ;
        RECT 825.6800 1518.4400 827.2800 1518.9200 ;
        RECT 882.2200 1496.6800 885.2200 1497.1600 ;
        RECT 882.2200 1502.1200 885.2200 1502.6000 ;
        RECT 870.6800 1496.6800 872.2800 1497.1600 ;
        RECT 870.6800 1502.1200 872.2800 1502.6000 ;
        RECT 882.2200 1480.3600 885.2200 1480.8400 ;
        RECT 882.2200 1485.8000 885.2200 1486.2800 ;
        RECT 882.2200 1491.2400 885.2200 1491.7200 ;
        RECT 870.6800 1480.3600 872.2800 1480.8400 ;
        RECT 870.6800 1485.8000 872.2800 1486.2800 ;
        RECT 870.6800 1491.2400 872.2800 1491.7200 ;
        RECT 882.2200 1469.4800 885.2200 1469.9600 ;
        RECT 882.2200 1474.9200 885.2200 1475.4000 ;
        RECT 870.6800 1469.4800 872.2800 1469.9600 ;
        RECT 870.6800 1474.9200 872.2800 1475.4000 ;
        RECT 882.2200 1464.0400 885.2200 1464.5200 ;
        RECT 870.6800 1464.0400 872.2800 1464.5200 ;
        RECT 825.6800 1496.6800 827.2800 1497.1600 ;
        RECT 825.6800 1502.1200 827.2800 1502.6000 ;
        RECT 825.6800 1480.3600 827.2800 1480.8400 ;
        RECT 825.6800 1485.8000 827.2800 1486.2800 ;
        RECT 825.6800 1491.2400 827.2800 1491.7200 ;
        RECT 825.6800 1469.4800 827.2800 1469.9600 ;
        RECT 825.6800 1474.9200 827.2800 1475.4000 ;
        RECT 825.6800 1464.0400 827.2800 1464.5200 ;
        RECT 780.6800 1551.0800 782.2800 1551.5600 ;
        RECT 780.6800 1556.5200 782.2800 1557.0000 ;
        RECT 780.6800 1534.7600 782.2800 1535.2400 ;
        RECT 780.6800 1540.2000 782.2800 1540.6800 ;
        RECT 780.6800 1545.6400 782.2800 1546.1200 ;
        RECT 735.6800 1551.0800 737.2800 1551.5600 ;
        RECT 735.6800 1556.5200 737.2800 1557.0000 ;
        RECT 735.6800 1534.7600 737.2800 1535.2400 ;
        RECT 735.6800 1540.2000 737.2800 1540.6800 ;
        RECT 735.6800 1545.6400 737.2800 1546.1200 ;
        RECT 780.6800 1523.8800 782.2800 1524.3600 ;
        RECT 780.6800 1529.3200 782.2800 1529.8000 ;
        RECT 780.6800 1507.5600 782.2800 1508.0400 ;
        RECT 780.6800 1513.0000 782.2800 1513.4800 ;
        RECT 780.6800 1518.4400 782.2800 1518.9200 ;
        RECT 735.6800 1523.8800 737.2800 1524.3600 ;
        RECT 735.6800 1529.3200 737.2800 1529.8000 ;
        RECT 735.6800 1507.5600 737.2800 1508.0400 ;
        RECT 735.6800 1513.0000 737.2800 1513.4800 ;
        RECT 735.6800 1518.4400 737.2800 1518.9200 ;
        RECT 686.1200 1551.0800 689.1200 1551.5600 ;
        RECT 686.1200 1556.5200 689.1200 1557.0000 ;
        RECT 686.1200 1540.2000 689.1200 1540.6800 ;
        RECT 686.1200 1534.7600 689.1200 1535.2400 ;
        RECT 686.1200 1545.6400 689.1200 1546.1200 ;
        RECT 686.1200 1523.8800 689.1200 1524.3600 ;
        RECT 686.1200 1529.3200 689.1200 1529.8000 ;
        RECT 686.1200 1513.0000 689.1200 1513.4800 ;
        RECT 686.1200 1507.5600 689.1200 1508.0400 ;
        RECT 686.1200 1518.4400 689.1200 1518.9200 ;
        RECT 780.6800 1496.6800 782.2800 1497.1600 ;
        RECT 780.6800 1502.1200 782.2800 1502.6000 ;
        RECT 780.6800 1480.3600 782.2800 1480.8400 ;
        RECT 780.6800 1485.8000 782.2800 1486.2800 ;
        RECT 780.6800 1491.2400 782.2800 1491.7200 ;
        RECT 735.6800 1496.6800 737.2800 1497.1600 ;
        RECT 735.6800 1502.1200 737.2800 1502.6000 ;
        RECT 735.6800 1480.3600 737.2800 1480.8400 ;
        RECT 735.6800 1485.8000 737.2800 1486.2800 ;
        RECT 735.6800 1491.2400 737.2800 1491.7200 ;
        RECT 780.6800 1474.9200 782.2800 1475.4000 ;
        RECT 780.6800 1469.4800 782.2800 1469.9600 ;
        RECT 780.6800 1464.0400 782.2800 1464.5200 ;
        RECT 735.6800 1474.9200 737.2800 1475.4000 ;
        RECT 735.6800 1469.4800 737.2800 1469.9600 ;
        RECT 735.6800 1464.0400 737.2800 1464.5200 ;
        RECT 686.1200 1496.6800 689.1200 1497.1600 ;
        RECT 686.1200 1502.1200 689.1200 1502.6000 ;
        RECT 686.1200 1485.8000 689.1200 1486.2800 ;
        RECT 686.1200 1480.3600 689.1200 1480.8400 ;
        RECT 686.1200 1491.2400 689.1200 1491.7200 ;
        RECT 686.1200 1469.4800 689.1200 1469.9600 ;
        RECT 686.1200 1474.9200 689.1200 1475.4000 ;
        RECT 686.1200 1464.0400 689.1200 1464.5200 ;
        RECT 686.1200 1662.2300 885.2200 1665.2300 ;
        RECT 686.1200 1457.1300 885.2200 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 1227.4900 872.2800 1435.5900 ;
        RECT 825.6800 1227.4900 827.2800 1435.5900 ;
        RECT 780.6800 1227.4900 782.2800 1435.5900 ;
        RECT 735.6800 1227.4900 737.2800 1435.5900 ;
        RECT 882.2200 1227.4900 885.2200 1435.5900 ;
        RECT 686.1200 1227.4900 689.1200 1435.5900 ;
      LAYER met3 ;
        RECT 882.2200 1430.2400 885.2200 1430.7200 ;
        RECT 870.6800 1430.2400 872.2800 1430.7200 ;
        RECT 882.2200 1419.3600 885.2200 1419.8400 ;
        RECT 882.2200 1424.8000 885.2200 1425.2800 ;
        RECT 870.6800 1419.3600 872.2800 1419.8400 ;
        RECT 870.6800 1424.8000 872.2800 1425.2800 ;
        RECT 882.2200 1403.0400 885.2200 1403.5200 ;
        RECT 882.2200 1408.4800 885.2200 1408.9600 ;
        RECT 870.6800 1403.0400 872.2800 1403.5200 ;
        RECT 870.6800 1408.4800 872.2800 1408.9600 ;
        RECT 882.2200 1392.1600 885.2200 1392.6400 ;
        RECT 882.2200 1397.6000 885.2200 1398.0800 ;
        RECT 870.6800 1392.1600 872.2800 1392.6400 ;
        RECT 870.6800 1397.6000 872.2800 1398.0800 ;
        RECT 882.2200 1413.9200 885.2200 1414.4000 ;
        RECT 870.6800 1413.9200 872.2800 1414.4000 ;
        RECT 825.6800 1419.3600 827.2800 1419.8400 ;
        RECT 825.6800 1424.8000 827.2800 1425.2800 ;
        RECT 825.6800 1430.2400 827.2800 1430.7200 ;
        RECT 825.6800 1403.0400 827.2800 1403.5200 ;
        RECT 825.6800 1408.4800 827.2800 1408.9600 ;
        RECT 825.6800 1397.6000 827.2800 1398.0800 ;
        RECT 825.6800 1392.1600 827.2800 1392.6400 ;
        RECT 825.6800 1413.9200 827.2800 1414.4000 ;
        RECT 882.2200 1375.8400 885.2200 1376.3200 ;
        RECT 882.2200 1381.2800 885.2200 1381.7600 ;
        RECT 870.6800 1375.8400 872.2800 1376.3200 ;
        RECT 870.6800 1381.2800 872.2800 1381.7600 ;
        RECT 882.2200 1359.5200 885.2200 1360.0000 ;
        RECT 882.2200 1364.9600 885.2200 1365.4400 ;
        RECT 882.2200 1370.4000 885.2200 1370.8800 ;
        RECT 870.6800 1359.5200 872.2800 1360.0000 ;
        RECT 870.6800 1364.9600 872.2800 1365.4400 ;
        RECT 870.6800 1370.4000 872.2800 1370.8800 ;
        RECT 882.2200 1348.6400 885.2200 1349.1200 ;
        RECT 882.2200 1354.0800 885.2200 1354.5600 ;
        RECT 870.6800 1348.6400 872.2800 1349.1200 ;
        RECT 870.6800 1354.0800 872.2800 1354.5600 ;
        RECT 882.2200 1332.3200 885.2200 1332.8000 ;
        RECT 882.2200 1337.7600 885.2200 1338.2400 ;
        RECT 882.2200 1343.2000 885.2200 1343.6800 ;
        RECT 870.6800 1332.3200 872.2800 1332.8000 ;
        RECT 870.6800 1337.7600 872.2800 1338.2400 ;
        RECT 870.6800 1343.2000 872.2800 1343.6800 ;
        RECT 825.6800 1375.8400 827.2800 1376.3200 ;
        RECT 825.6800 1381.2800 827.2800 1381.7600 ;
        RECT 825.6800 1359.5200 827.2800 1360.0000 ;
        RECT 825.6800 1364.9600 827.2800 1365.4400 ;
        RECT 825.6800 1370.4000 827.2800 1370.8800 ;
        RECT 825.6800 1348.6400 827.2800 1349.1200 ;
        RECT 825.6800 1354.0800 827.2800 1354.5600 ;
        RECT 825.6800 1332.3200 827.2800 1332.8000 ;
        RECT 825.6800 1337.7600 827.2800 1338.2400 ;
        RECT 825.6800 1343.2000 827.2800 1343.6800 ;
        RECT 882.2200 1386.7200 885.2200 1387.2000 ;
        RECT 825.6800 1386.7200 827.2800 1387.2000 ;
        RECT 870.6800 1386.7200 872.2800 1387.2000 ;
        RECT 780.6800 1419.3600 782.2800 1419.8400 ;
        RECT 780.6800 1424.8000 782.2800 1425.2800 ;
        RECT 780.6800 1430.2400 782.2800 1430.7200 ;
        RECT 735.6800 1419.3600 737.2800 1419.8400 ;
        RECT 735.6800 1424.8000 737.2800 1425.2800 ;
        RECT 735.6800 1430.2400 737.2800 1430.7200 ;
        RECT 780.6800 1403.0400 782.2800 1403.5200 ;
        RECT 780.6800 1408.4800 782.2800 1408.9600 ;
        RECT 780.6800 1392.1600 782.2800 1392.6400 ;
        RECT 780.6800 1397.6000 782.2800 1398.0800 ;
        RECT 735.6800 1403.0400 737.2800 1403.5200 ;
        RECT 735.6800 1408.4800 737.2800 1408.9600 ;
        RECT 735.6800 1392.1600 737.2800 1392.6400 ;
        RECT 735.6800 1397.6000 737.2800 1398.0800 ;
        RECT 735.6800 1413.9200 737.2800 1414.4000 ;
        RECT 780.6800 1413.9200 782.2800 1414.4000 ;
        RECT 686.1200 1430.2400 689.1200 1430.7200 ;
        RECT 686.1200 1424.8000 689.1200 1425.2800 ;
        RECT 686.1200 1419.3600 689.1200 1419.8400 ;
        RECT 686.1200 1408.4800 689.1200 1408.9600 ;
        RECT 686.1200 1403.0400 689.1200 1403.5200 ;
        RECT 686.1200 1397.6000 689.1200 1398.0800 ;
        RECT 686.1200 1392.1600 689.1200 1392.6400 ;
        RECT 686.1200 1413.9200 689.1200 1414.4000 ;
        RECT 780.6800 1375.8400 782.2800 1376.3200 ;
        RECT 780.6800 1381.2800 782.2800 1381.7600 ;
        RECT 780.6800 1359.5200 782.2800 1360.0000 ;
        RECT 780.6800 1364.9600 782.2800 1365.4400 ;
        RECT 780.6800 1370.4000 782.2800 1370.8800 ;
        RECT 735.6800 1375.8400 737.2800 1376.3200 ;
        RECT 735.6800 1381.2800 737.2800 1381.7600 ;
        RECT 735.6800 1359.5200 737.2800 1360.0000 ;
        RECT 735.6800 1364.9600 737.2800 1365.4400 ;
        RECT 735.6800 1370.4000 737.2800 1370.8800 ;
        RECT 780.6800 1348.6400 782.2800 1349.1200 ;
        RECT 780.6800 1354.0800 782.2800 1354.5600 ;
        RECT 780.6800 1332.3200 782.2800 1332.8000 ;
        RECT 780.6800 1337.7600 782.2800 1338.2400 ;
        RECT 780.6800 1343.2000 782.2800 1343.6800 ;
        RECT 735.6800 1348.6400 737.2800 1349.1200 ;
        RECT 735.6800 1354.0800 737.2800 1354.5600 ;
        RECT 735.6800 1332.3200 737.2800 1332.8000 ;
        RECT 735.6800 1337.7600 737.2800 1338.2400 ;
        RECT 735.6800 1343.2000 737.2800 1343.6800 ;
        RECT 686.1200 1375.8400 689.1200 1376.3200 ;
        RECT 686.1200 1381.2800 689.1200 1381.7600 ;
        RECT 686.1200 1364.9600 689.1200 1365.4400 ;
        RECT 686.1200 1359.5200 689.1200 1360.0000 ;
        RECT 686.1200 1370.4000 689.1200 1370.8800 ;
        RECT 686.1200 1348.6400 689.1200 1349.1200 ;
        RECT 686.1200 1354.0800 689.1200 1354.5600 ;
        RECT 686.1200 1337.7600 689.1200 1338.2400 ;
        RECT 686.1200 1332.3200 689.1200 1332.8000 ;
        RECT 686.1200 1343.2000 689.1200 1343.6800 ;
        RECT 686.1200 1386.7200 689.1200 1387.2000 ;
        RECT 735.6800 1386.7200 737.2800 1387.2000 ;
        RECT 780.6800 1386.7200 782.2800 1387.2000 ;
        RECT 882.2200 1321.4400 885.2200 1321.9200 ;
        RECT 882.2200 1326.8800 885.2200 1327.3600 ;
        RECT 870.6800 1321.4400 872.2800 1321.9200 ;
        RECT 870.6800 1326.8800 872.2800 1327.3600 ;
        RECT 882.2200 1305.1200 885.2200 1305.6000 ;
        RECT 882.2200 1310.5600 885.2200 1311.0400 ;
        RECT 882.2200 1316.0000 885.2200 1316.4800 ;
        RECT 870.6800 1305.1200 872.2800 1305.6000 ;
        RECT 870.6800 1310.5600 872.2800 1311.0400 ;
        RECT 870.6800 1316.0000 872.2800 1316.4800 ;
        RECT 882.2200 1294.2400 885.2200 1294.7200 ;
        RECT 882.2200 1299.6800 885.2200 1300.1600 ;
        RECT 870.6800 1294.2400 872.2800 1294.7200 ;
        RECT 870.6800 1299.6800 872.2800 1300.1600 ;
        RECT 882.2200 1277.9200 885.2200 1278.4000 ;
        RECT 882.2200 1283.3600 885.2200 1283.8400 ;
        RECT 882.2200 1288.8000 885.2200 1289.2800 ;
        RECT 870.6800 1277.9200 872.2800 1278.4000 ;
        RECT 870.6800 1283.3600 872.2800 1283.8400 ;
        RECT 870.6800 1288.8000 872.2800 1289.2800 ;
        RECT 825.6800 1321.4400 827.2800 1321.9200 ;
        RECT 825.6800 1326.8800 827.2800 1327.3600 ;
        RECT 825.6800 1305.1200 827.2800 1305.6000 ;
        RECT 825.6800 1310.5600 827.2800 1311.0400 ;
        RECT 825.6800 1316.0000 827.2800 1316.4800 ;
        RECT 825.6800 1294.2400 827.2800 1294.7200 ;
        RECT 825.6800 1299.6800 827.2800 1300.1600 ;
        RECT 825.6800 1277.9200 827.2800 1278.4000 ;
        RECT 825.6800 1283.3600 827.2800 1283.8400 ;
        RECT 825.6800 1288.8000 827.2800 1289.2800 ;
        RECT 882.2200 1267.0400 885.2200 1267.5200 ;
        RECT 882.2200 1272.4800 885.2200 1272.9600 ;
        RECT 870.6800 1267.0400 872.2800 1267.5200 ;
        RECT 870.6800 1272.4800 872.2800 1272.9600 ;
        RECT 882.2200 1250.7200 885.2200 1251.2000 ;
        RECT 882.2200 1256.1600 885.2200 1256.6400 ;
        RECT 882.2200 1261.6000 885.2200 1262.0800 ;
        RECT 870.6800 1250.7200 872.2800 1251.2000 ;
        RECT 870.6800 1256.1600 872.2800 1256.6400 ;
        RECT 870.6800 1261.6000 872.2800 1262.0800 ;
        RECT 882.2200 1239.8400 885.2200 1240.3200 ;
        RECT 882.2200 1245.2800 885.2200 1245.7600 ;
        RECT 870.6800 1239.8400 872.2800 1240.3200 ;
        RECT 870.6800 1245.2800 872.2800 1245.7600 ;
        RECT 882.2200 1234.4000 885.2200 1234.8800 ;
        RECT 870.6800 1234.4000 872.2800 1234.8800 ;
        RECT 825.6800 1267.0400 827.2800 1267.5200 ;
        RECT 825.6800 1272.4800 827.2800 1272.9600 ;
        RECT 825.6800 1250.7200 827.2800 1251.2000 ;
        RECT 825.6800 1256.1600 827.2800 1256.6400 ;
        RECT 825.6800 1261.6000 827.2800 1262.0800 ;
        RECT 825.6800 1239.8400 827.2800 1240.3200 ;
        RECT 825.6800 1245.2800 827.2800 1245.7600 ;
        RECT 825.6800 1234.4000 827.2800 1234.8800 ;
        RECT 780.6800 1321.4400 782.2800 1321.9200 ;
        RECT 780.6800 1326.8800 782.2800 1327.3600 ;
        RECT 780.6800 1305.1200 782.2800 1305.6000 ;
        RECT 780.6800 1310.5600 782.2800 1311.0400 ;
        RECT 780.6800 1316.0000 782.2800 1316.4800 ;
        RECT 735.6800 1321.4400 737.2800 1321.9200 ;
        RECT 735.6800 1326.8800 737.2800 1327.3600 ;
        RECT 735.6800 1305.1200 737.2800 1305.6000 ;
        RECT 735.6800 1310.5600 737.2800 1311.0400 ;
        RECT 735.6800 1316.0000 737.2800 1316.4800 ;
        RECT 780.6800 1294.2400 782.2800 1294.7200 ;
        RECT 780.6800 1299.6800 782.2800 1300.1600 ;
        RECT 780.6800 1277.9200 782.2800 1278.4000 ;
        RECT 780.6800 1283.3600 782.2800 1283.8400 ;
        RECT 780.6800 1288.8000 782.2800 1289.2800 ;
        RECT 735.6800 1294.2400 737.2800 1294.7200 ;
        RECT 735.6800 1299.6800 737.2800 1300.1600 ;
        RECT 735.6800 1277.9200 737.2800 1278.4000 ;
        RECT 735.6800 1283.3600 737.2800 1283.8400 ;
        RECT 735.6800 1288.8000 737.2800 1289.2800 ;
        RECT 686.1200 1321.4400 689.1200 1321.9200 ;
        RECT 686.1200 1326.8800 689.1200 1327.3600 ;
        RECT 686.1200 1310.5600 689.1200 1311.0400 ;
        RECT 686.1200 1305.1200 689.1200 1305.6000 ;
        RECT 686.1200 1316.0000 689.1200 1316.4800 ;
        RECT 686.1200 1294.2400 689.1200 1294.7200 ;
        RECT 686.1200 1299.6800 689.1200 1300.1600 ;
        RECT 686.1200 1283.3600 689.1200 1283.8400 ;
        RECT 686.1200 1277.9200 689.1200 1278.4000 ;
        RECT 686.1200 1288.8000 689.1200 1289.2800 ;
        RECT 780.6800 1267.0400 782.2800 1267.5200 ;
        RECT 780.6800 1272.4800 782.2800 1272.9600 ;
        RECT 780.6800 1250.7200 782.2800 1251.2000 ;
        RECT 780.6800 1256.1600 782.2800 1256.6400 ;
        RECT 780.6800 1261.6000 782.2800 1262.0800 ;
        RECT 735.6800 1267.0400 737.2800 1267.5200 ;
        RECT 735.6800 1272.4800 737.2800 1272.9600 ;
        RECT 735.6800 1250.7200 737.2800 1251.2000 ;
        RECT 735.6800 1256.1600 737.2800 1256.6400 ;
        RECT 735.6800 1261.6000 737.2800 1262.0800 ;
        RECT 780.6800 1245.2800 782.2800 1245.7600 ;
        RECT 780.6800 1239.8400 782.2800 1240.3200 ;
        RECT 780.6800 1234.4000 782.2800 1234.8800 ;
        RECT 735.6800 1245.2800 737.2800 1245.7600 ;
        RECT 735.6800 1239.8400 737.2800 1240.3200 ;
        RECT 735.6800 1234.4000 737.2800 1234.8800 ;
        RECT 686.1200 1267.0400 689.1200 1267.5200 ;
        RECT 686.1200 1272.4800 689.1200 1272.9600 ;
        RECT 686.1200 1256.1600 689.1200 1256.6400 ;
        RECT 686.1200 1250.7200 689.1200 1251.2000 ;
        RECT 686.1200 1261.6000 689.1200 1262.0800 ;
        RECT 686.1200 1239.8400 689.1200 1240.3200 ;
        RECT 686.1200 1245.2800 689.1200 1245.7600 ;
        RECT 686.1200 1234.4000 689.1200 1234.8800 ;
        RECT 686.1200 1432.5900 885.2200 1435.5900 ;
        RECT 686.1200 1227.4900 885.2200 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 997.8500 872.2800 1205.9500 ;
        RECT 825.6800 997.8500 827.2800 1205.9500 ;
        RECT 780.6800 997.8500 782.2800 1205.9500 ;
        RECT 735.6800 997.8500 737.2800 1205.9500 ;
        RECT 882.2200 997.8500 885.2200 1205.9500 ;
        RECT 686.1200 997.8500 689.1200 1205.9500 ;
      LAYER met3 ;
        RECT 882.2200 1200.6000 885.2200 1201.0800 ;
        RECT 870.6800 1200.6000 872.2800 1201.0800 ;
        RECT 882.2200 1189.7200 885.2200 1190.2000 ;
        RECT 882.2200 1195.1600 885.2200 1195.6400 ;
        RECT 870.6800 1189.7200 872.2800 1190.2000 ;
        RECT 870.6800 1195.1600 872.2800 1195.6400 ;
        RECT 882.2200 1173.4000 885.2200 1173.8800 ;
        RECT 882.2200 1178.8400 885.2200 1179.3200 ;
        RECT 870.6800 1173.4000 872.2800 1173.8800 ;
        RECT 870.6800 1178.8400 872.2800 1179.3200 ;
        RECT 882.2200 1162.5200 885.2200 1163.0000 ;
        RECT 882.2200 1167.9600 885.2200 1168.4400 ;
        RECT 870.6800 1162.5200 872.2800 1163.0000 ;
        RECT 870.6800 1167.9600 872.2800 1168.4400 ;
        RECT 882.2200 1184.2800 885.2200 1184.7600 ;
        RECT 870.6800 1184.2800 872.2800 1184.7600 ;
        RECT 825.6800 1189.7200 827.2800 1190.2000 ;
        RECT 825.6800 1195.1600 827.2800 1195.6400 ;
        RECT 825.6800 1200.6000 827.2800 1201.0800 ;
        RECT 825.6800 1173.4000 827.2800 1173.8800 ;
        RECT 825.6800 1178.8400 827.2800 1179.3200 ;
        RECT 825.6800 1167.9600 827.2800 1168.4400 ;
        RECT 825.6800 1162.5200 827.2800 1163.0000 ;
        RECT 825.6800 1184.2800 827.2800 1184.7600 ;
        RECT 882.2200 1146.2000 885.2200 1146.6800 ;
        RECT 882.2200 1151.6400 885.2200 1152.1200 ;
        RECT 870.6800 1146.2000 872.2800 1146.6800 ;
        RECT 870.6800 1151.6400 872.2800 1152.1200 ;
        RECT 882.2200 1129.8800 885.2200 1130.3600 ;
        RECT 882.2200 1135.3200 885.2200 1135.8000 ;
        RECT 882.2200 1140.7600 885.2200 1141.2400 ;
        RECT 870.6800 1129.8800 872.2800 1130.3600 ;
        RECT 870.6800 1135.3200 872.2800 1135.8000 ;
        RECT 870.6800 1140.7600 872.2800 1141.2400 ;
        RECT 882.2200 1119.0000 885.2200 1119.4800 ;
        RECT 882.2200 1124.4400 885.2200 1124.9200 ;
        RECT 870.6800 1119.0000 872.2800 1119.4800 ;
        RECT 870.6800 1124.4400 872.2800 1124.9200 ;
        RECT 882.2200 1102.6800 885.2200 1103.1600 ;
        RECT 882.2200 1108.1200 885.2200 1108.6000 ;
        RECT 882.2200 1113.5600 885.2200 1114.0400 ;
        RECT 870.6800 1102.6800 872.2800 1103.1600 ;
        RECT 870.6800 1108.1200 872.2800 1108.6000 ;
        RECT 870.6800 1113.5600 872.2800 1114.0400 ;
        RECT 825.6800 1146.2000 827.2800 1146.6800 ;
        RECT 825.6800 1151.6400 827.2800 1152.1200 ;
        RECT 825.6800 1129.8800 827.2800 1130.3600 ;
        RECT 825.6800 1135.3200 827.2800 1135.8000 ;
        RECT 825.6800 1140.7600 827.2800 1141.2400 ;
        RECT 825.6800 1119.0000 827.2800 1119.4800 ;
        RECT 825.6800 1124.4400 827.2800 1124.9200 ;
        RECT 825.6800 1102.6800 827.2800 1103.1600 ;
        RECT 825.6800 1108.1200 827.2800 1108.6000 ;
        RECT 825.6800 1113.5600 827.2800 1114.0400 ;
        RECT 882.2200 1157.0800 885.2200 1157.5600 ;
        RECT 825.6800 1157.0800 827.2800 1157.5600 ;
        RECT 870.6800 1157.0800 872.2800 1157.5600 ;
        RECT 780.6800 1189.7200 782.2800 1190.2000 ;
        RECT 780.6800 1195.1600 782.2800 1195.6400 ;
        RECT 780.6800 1200.6000 782.2800 1201.0800 ;
        RECT 735.6800 1189.7200 737.2800 1190.2000 ;
        RECT 735.6800 1195.1600 737.2800 1195.6400 ;
        RECT 735.6800 1200.6000 737.2800 1201.0800 ;
        RECT 780.6800 1173.4000 782.2800 1173.8800 ;
        RECT 780.6800 1178.8400 782.2800 1179.3200 ;
        RECT 780.6800 1162.5200 782.2800 1163.0000 ;
        RECT 780.6800 1167.9600 782.2800 1168.4400 ;
        RECT 735.6800 1173.4000 737.2800 1173.8800 ;
        RECT 735.6800 1178.8400 737.2800 1179.3200 ;
        RECT 735.6800 1162.5200 737.2800 1163.0000 ;
        RECT 735.6800 1167.9600 737.2800 1168.4400 ;
        RECT 735.6800 1184.2800 737.2800 1184.7600 ;
        RECT 780.6800 1184.2800 782.2800 1184.7600 ;
        RECT 686.1200 1200.6000 689.1200 1201.0800 ;
        RECT 686.1200 1195.1600 689.1200 1195.6400 ;
        RECT 686.1200 1189.7200 689.1200 1190.2000 ;
        RECT 686.1200 1178.8400 689.1200 1179.3200 ;
        RECT 686.1200 1173.4000 689.1200 1173.8800 ;
        RECT 686.1200 1167.9600 689.1200 1168.4400 ;
        RECT 686.1200 1162.5200 689.1200 1163.0000 ;
        RECT 686.1200 1184.2800 689.1200 1184.7600 ;
        RECT 780.6800 1146.2000 782.2800 1146.6800 ;
        RECT 780.6800 1151.6400 782.2800 1152.1200 ;
        RECT 780.6800 1129.8800 782.2800 1130.3600 ;
        RECT 780.6800 1135.3200 782.2800 1135.8000 ;
        RECT 780.6800 1140.7600 782.2800 1141.2400 ;
        RECT 735.6800 1146.2000 737.2800 1146.6800 ;
        RECT 735.6800 1151.6400 737.2800 1152.1200 ;
        RECT 735.6800 1129.8800 737.2800 1130.3600 ;
        RECT 735.6800 1135.3200 737.2800 1135.8000 ;
        RECT 735.6800 1140.7600 737.2800 1141.2400 ;
        RECT 780.6800 1119.0000 782.2800 1119.4800 ;
        RECT 780.6800 1124.4400 782.2800 1124.9200 ;
        RECT 780.6800 1102.6800 782.2800 1103.1600 ;
        RECT 780.6800 1108.1200 782.2800 1108.6000 ;
        RECT 780.6800 1113.5600 782.2800 1114.0400 ;
        RECT 735.6800 1119.0000 737.2800 1119.4800 ;
        RECT 735.6800 1124.4400 737.2800 1124.9200 ;
        RECT 735.6800 1102.6800 737.2800 1103.1600 ;
        RECT 735.6800 1108.1200 737.2800 1108.6000 ;
        RECT 735.6800 1113.5600 737.2800 1114.0400 ;
        RECT 686.1200 1146.2000 689.1200 1146.6800 ;
        RECT 686.1200 1151.6400 689.1200 1152.1200 ;
        RECT 686.1200 1135.3200 689.1200 1135.8000 ;
        RECT 686.1200 1129.8800 689.1200 1130.3600 ;
        RECT 686.1200 1140.7600 689.1200 1141.2400 ;
        RECT 686.1200 1119.0000 689.1200 1119.4800 ;
        RECT 686.1200 1124.4400 689.1200 1124.9200 ;
        RECT 686.1200 1108.1200 689.1200 1108.6000 ;
        RECT 686.1200 1102.6800 689.1200 1103.1600 ;
        RECT 686.1200 1113.5600 689.1200 1114.0400 ;
        RECT 686.1200 1157.0800 689.1200 1157.5600 ;
        RECT 735.6800 1157.0800 737.2800 1157.5600 ;
        RECT 780.6800 1157.0800 782.2800 1157.5600 ;
        RECT 882.2200 1091.8000 885.2200 1092.2800 ;
        RECT 882.2200 1097.2400 885.2200 1097.7200 ;
        RECT 870.6800 1091.8000 872.2800 1092.2800 ;
        RECT 870.6800 1097.2400 872.2800 1097.7200 ;
        RECT 882.2200 1075.4800 885.2200 1075.9600 ;
        RECT 882.2200 1080.9200 885.2200 1081.4000 ;
        RECT 882.2200 1086.3600 885.2200 1086.8400 ;
        RECT 870.6800 1075.4800 872.2800 1075.9600 ;
        RECT 870.6800 1080.9200 872.2800 1081.4000 ;
        RECT 870.6800 1086.3600 872.2800 1086.8400 ;
        RECT 882.2200 1064.6000 885.2200 1065.0800 ;
        RECT 882.2200 1070.0400 885.2200 1070.5200 ;
        RECT 870.6800 1064.6000 872.2800 1065.0800 ;
        RECT 870.6800 1070.0400 872.2800 1070.5200 ;
        RECT 882.2200 1048.2800 885.2200 1048.7600 ;
        RECT 882.2200 1053.7200 885.2200 1054.2000 ;
        RECT 882.2200 1059.1600 885.2200 1059.6400 ;
        RECT 870.6800 1048.2800 872.2800 1048.7600 ;
        RECT 870.6800 1053.7200 872.2800 1054.2000 ;
        RECT 870.6800 1059.1600 872.2800 1059.6400 ;
        RECT 825.6800 1091.8000 827.2800 1092.2800 ;
        RECT 825.6800 1097.2400 827.2800 1097.7200 ;
        RECT 825.6800 1075.4800 827.2800 1075.9600 ;
        RECT 825.6800 1080.9200 827.2800 1081.4000 ;
        RECT 825.6800 1086.3600 827.2800 1086.8400 ;
        RECT 825.6800 1064.6000 827.2800 1065.0800 ;
        RECT 825.6800 1070.0400 827.2800 1070.5200 ;
        RECT 825.6800 1048.2800 827.2800 1048.7600 ;
        RECT 825.6800 1053.7200 827.2800 1054.2000 ;
        RECT 825.6800 1059.1600 827.2800 1059.6400 ;
        RECT 882.2200 1037.4000 885.2200 1037.8800 ;
        RECT 882.2200 1042.8400 885.2200 1043.3200 ;
        RECT 870.6800 1037.4000 872.2800 1037.8800 ;
        RECT 870.6800 1042.8400 872.2800 1043.3200 ;
        RECT 882.2200 1021.0800 885.2200 1021.5600 ;
        RECT 882.2200 1026.5200 885.2200 1027.0000 ;
        RECT 882.2200 1031.9600 885.2200 1032.4400 ;
        RECT 870.6800 1021.0800 872.2800 1021.5600 ;
        RECT 870.6800 1026.5200 872.2800 1027.0000 ;
        RECT 870.6800 1031.9600 872.2800 1032.4400 ;
        RECT 882.2200 1010.2000 885.2200 1010.6800 ;
        RECT 882.2200 1015.6400 885.2200 1016.1200 ;
        RECT 870.6800 1010.2000 872.2800 1010.6800 ;
        RECT 870.6800 1015.6400 872.2800 1016.1200 ;
        RECT 882.2200 1004.7600 885.2200 1005.2400 ;
        RECT 870.6800 1004.7600 872.2800 1005.2400 ;
        RECT 825.6800 1037.4000 827.2800 1037.8800 ;
        RECT 825.6800 1042.8400 827.2800 1043.3200 ;
        RECT 825.6800 1021.0800 827.2800 1021.5600 ;
        RECT 825.6800 1026.5200 827.2800 1027.0000 ;
        RECT 825.6800 1031.9600 827.2800 1032.4400 ;
        RECT 825.6800 1010.2000 827.2800 1010.6800 ;
        RECT 825.6800 1015.6400 827.2800 1016.1200 ;
        RECT 825.6800 1004.7600 827.2800 1005.2400 ;
        RECT 780.6800 1091.8000 782.2800 1092.2800 ;
        RECT 780.6800 1097.2400 782.2800 1097.7200 ;
        RECT 780.6800 1075.4800 782.2800 1075.9600 ;
        RECT 780.6800 1080.9200 782.2800 1081.4000 ;
        RECT 780.6800 1086.3600 782.2800 1086.8400 ;
        RECT 735.6800 1091.8000 737.2800 1092.2800 ;
        RECT 735.6800 1097.2400 737.2800 1097.7200 ;
        RECT 735.6800 1075.4800 737.2800 1075.9600 ;
        RECT 735.6800 1080.9200 737.2800 1081.4000 ;
        RECT 735.6800 1086.3600 737.2800 1086.8400 ;
        RECT 780.6800 1064.6000 782.2800 1065.0800 ;
        RECT 780.6800 1070.0400 782.2800 1070.5200 ;
        RECT 780.6800 1048.2800 782.2800 1048.7600 ;
        RECT 780.6800 1053.7200 782.2800 1054.2000 ;
        RECT 780.6800 1059.1600 782.2800 1059.6400 ;
        RECT 735.6800 1064.6000 737.2800 1065.0800 ;
        RECT 735.6800 1070.0400 737.2800 1070.5200 ;
        RECT 735.6800 1048.2800 737.2800 1048.7600 ;
        RECT 735.6800 1053.7200 737.2800 1054.2000 ;
        RECT 735.6800 1059.1600 737.2800 1059.6400 ;
        RECT 686.1200 1091.8000 689.1200 1092.2800 ;
        RECT 686.1200 1097.2400 689.1200 1097.7200 ;
        RECT 686.1200 1080.9200 689.1200 1081.4000 ;
        RECT 686.1200 1075.4800 689.1200 1075.9600 ;
        RECT 686.1200 1086.3600 689.1200 1086.8400 ;
        RECT 686.1200 1064.6000 689.1200 1065.0800 ;
        RECT 686.1200 1070.0400 689.1200 1070.5200 ;
        RECT 686.1200 1053.7200 689.1200 1054.2000 ;
        RECT 686.1200 1048.2800 689.1200 1048.7600 ;
        RECT 686.1200 1059.1600 689.1200 1059.6400 ;
        RECT 780.6800 1037.4000 782.2800 1037.8800 ;
        RECT 780.6800 1042.8400 782.2800 1043.3200 ;
        RECT 780.6800 1021.0800 782.2800 1021.5600 ;
        RECT 780.6800 1026.5200 782.2800 1027.0000 ;
        RECT 780.6800 1031.9600 782.2800 1032.4400 ;
        RECT 735.6800 1037.4000 737.2800 1037.8800 ;
        RECT 735.6800 1042.8400 737.2800 1043.3200 ;
        RECT 735.6800 1021.0800 737.2800 1021.5600 ;
        RECT 735.6800 1026.5200 737.2800 1027.0000 ;
        RECT 735.6800 1031.9600 737.2800 1032.4400 ;
        RECT 780.6800 1015.6400 782.2800 1016.1200 ;
        RECT 780.6800 1010.2000 782.2800 1010.6800 ;
        RECT 780.6800 1004.7600 782.2800 1005.2400 ;
        RECT 735.6800 1015.6400 737.2800 1016.1200 ;
        RECT 735.6800 1010.2000 737.2800 1010.6800 ;
        RECT 735.6800 1004.7600 737.2800 1005.2400 ;
        RECT 686.1200 1037.4000 689.1200 1037.8800 ;
        RECT 686.1200 1042.8400 689.1200 1043.3200 ;
        RECT 686.1200 1026.5200 689.1200 1027.0000 ;
        RECT 686.1200 1021.0800 689.1200 1021.5600 ;
        RECT 686.1200 1031.9600 689.1200 1032.4400 ;
        RECT 686.1200 1010.2000 689.1200 1010.6800 ;
        RECT 686.1200 1015.6400 689.1200 1016.1200 ;
        RECT 686.1200 1004.7600 689.1200 1005.2400 ;
        RECT 686.1200 1202.9500 885.2200 1205.9500 ;
        RECT 686.1200 997.8500 885.2200 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 870.6800 768.2100 872.2800 976.3100 ;
        RECT 825.6800 768.2100 827.2800 976.3100 ;
        RECT 780.6800 768.2100 782.2800 976.3100 ;
        RECT 735.6800 768.2100 737.2800 976.3100 ;
        RECT 882.2200 768.2100 885.2200 976.3100 ;
        RECT 686.1200 768.2100 689.1200 976.3100 ;
      LAYER met3 ;
        RECT 882.2200 970.9600 885.2200 971.4400 ;
        RECT 870.6800 970.9600 872.2800 971.4400 ;
        RECT 882.2200 960.0800 885.2200 960.5600 ;
        RECT 882.2200 965.5200 885.2200 966.0000 ;
        RECT 870.6800 960.0800 872.2800 960.5600 ;
        RECT 870.6800 965.5200 872.2800 966.0000 ;
        RECT 882.2200 943.7600 885.2200 944.2400 ;
        RECT 882.2200 949.2000 885.2200 949.6800 ;
        RECT 870.6800 943.7600 872.2800 944.2400 ;
        RECT 870.6800 949.2000 872.2800 949.6800 ;
        RECT 882.2200 932.8800 885.2200 933.3600 ;
        RECT 882.2200 938.3200 885.2200 938.8000 ;
        RECT 870.6800 932.8800 872.2800 933.3600 ;
        RECT 870.6800 938.3200 872.2800 938.8000 ;
        RECT 882.2200 954.6400 885.2200 955.1200 ;
        RECT 870.6800 954.6400 872.2800 955.1200 ;
        RECT 825.6800 960.0800 827.2800 960.5600 ;
        RECT 825.6800 965.5200 827.2800 966.0000 ;
        RECT 825.6800 970.9600 827.2800 971.4400 ;
        RECT 825.6800 943.7600 827.2800 944.2400 ;
        RECT 825.6800 949.2000 827.2800 949.6800 ;
        RECT 825.6800 938.3200 827.2800 938.8000 ;
        RECT 825.6800 932.8800 827.2800 933.3600 ;
        RECT 825.6800 954.6400 827.2800 955.1200 ;
        RECT 882.2200 916.5600 885.2200 917.0400 ;
        RECT 882.2200 922.0000 885.2200 922.4800 ;
        RECT 870.6800 916.5600 872.2800 917.0400 ;
        RECT 870.6800 922.0000 872.2800 922.4800 ;
        RECT 882.2200 900.2400 885.2200 900.7200 ;
        RECT 882.2200 905.6800 885.2200 906.1600 ;
        RECT 882.2200 911.1200 885.2200 911.6000 ;
        RECT 870.6800 900.2400 872.2800 900.7200 ;
        RECT 870.6800 905.6800 872.2800 906.1600 ;
        RECT 870.6800 911.1200 872.2800 911.6000 ;
        RECT 882.2200 889.3600 885.2200 889.8400 ;
        RECT 882.2200 894.8000 885.2200 895.2800 ;
        RECT 870.6800 889.3600 872.2800 889.8400 ;
        RECT 870.6800 894.8000 872.2800 895.2800 ;
        RECT 882.2200 873.0400 885.2200 873.5200 ;
        RECT 882.2200 878.4800 885.2200 878.9600 ;
        RECT 882.2200 883.9200 885.2200 884.4000 ;
        RECT 870.6800 873.0400 872.2800 873.5200 ;
        RECT 870.6800 878.4800 872.2800 878.9600 ;
        RECT 870.6800 883.9200 872.2800 884.4000 ;
        RECT 825.6800 916.5600 827.2800 917.0400 ;
        RECT 825.6800 922.0000 827.2800 922.4800 ;
        RECT 825.6800 900.2400 827.2800 900.7200 ;
        RECT 825.6800 905.6800 827.2800 906.1600 ;
        RECT 825.6800 911.1200 827.2800 911.6000 ;
        RECT 825.6800 889.3600 827.2800 889.8400 ;
        RECT 825.6800 894.8000 827.2800 895.2800 ;
        RECT 825.6800 873.0400 827.2800 873.5200 ;
        RECT 825.6800 878.4800 827.2800 878.9600 ;
        RECT 825.6800 883.9200 827.2800 884.4000 ;
        RECT 882.2200 927.4400 885.2200 927.9200 ;
        RECT 825.6800 927.4400 827.2800 927.9200 ;
        RECT 870.6800 927.4400 872.2800 927.9200 ;
        RECT 780.6800 960.0800 782.2800 960.5600 ;
        RECT 780.6800 965.5200 782.2800 966.0000 ;
        RECT 780.6800 970.9600 782.2800 971.4400 ;
        RECT 735.6800 960.0800 737.2800 960.5600 ;
        RECT 735.6800 965.5200 737.2800 966.0000 ;
        RECT 735.6800 970.9600 737.2800 971.4400 ;
        RECT 780.6800 943.7600 782.2800 944.2400 ;
        RECT 780.6800 949.2000 782.2800 949.6800 ;
        RECT 780.6800 932.8800 782.2800 933.3600 ;
        RECT 780.6800 938.3200 782.2800 938.8000 ;
        RECT 735.6800 943.7600 737.2800 944.2400 ;
        RECT 735.6800 949.2000 737.2800 949.6800 ;
        RECT 735.6800 932.8800 737.2800 933.3600 ;
        RECT 735.6800 938.3200 737.2800 938.8000 ;
        RECT 735.6800 954.6400 737.2800 955.1200 ;
        RECT 780.6800 954.6400 782.2800 955.1200 ;
        RECT 686.1200 970.9600 689.1200 971.4400 ;
        RECT 686.1200 965.5200 689.1200 966.0000 ;
        RECT 686.1200 960.0800 689.1200 960.5600 ;
        RECT 686.1200 949.2000 689.1200 949.6800 ;
        RECT 686.1200 943.7600 689.1200 944.2400 ;
        RECT 686.1200 938.3200 689.1200 938.8000 ;
        RECT 686.1200 932.8800 689.1200 933.3600 ;
        RECT 686.1200 954.6400 689.1200 955.1200 ;
        RECT 780.6800 916.5600 782.2800 917.0400 ;
        RECT 780.6800 922.0000 782.2800 922.4800 ;
        RECT 780.6800 900.2400 782.2800 900.7200 ;
        RECT 780.6800 905.6800 782.2800 906.1600 ;
        RECT 780.6800 911.1200 782.2800 911.6000 ;
        RECT 735.6800 916.5600 737.2800 917.0400 ;
        RECT 735.6800 922.0000 737.2800 922.4800 ;
        RECT 735.6800 900.2400 737.2800 900.7200 ;
        RECT 735.6800 905.6800 737.2800 906.1600 ;
        RECT 735.6800 911.1200 737.2800 911.6000 ;
        RECT 780.6800 889.3600 782.2800 889.8400 ;
        RECT 780.6800 894.8000 782.2800 895.2800 ;
        RECT 780.6800 873.0400 782.2800 873.5200 ;
        RECT 780.6800 878.4800 782.2800 878.9600 ;
        RECT 780.6800 883.9200 782.2800 884.4000 ;
        RECT 735.6800 889.3600 737.2800 889.8400 ;
        RECT 735.6800 894.8000 737.2800 895.2800 ;
        RECT 735.6800 873.0400 737.2800 873.5200 ;
        RECT 735.6800 878.4800 737.2800 878.9600 ;
        RECT 735.6800 883.9200 737.2800 884.4000 ;
        RECT 686.1200 916.5600 689.1200 917.0400 ;
        RECT 686.1200 922.0000 689.1200 922.4800 ;
        RECT 686.1200 905.6800 689.1200 906.1600 ;
        RECT 686.1200 900.2400 689.1200 900.7200 ;
        RECT 686.1200 911.1200 689.1200 911.6000 ;
        RECT 686.1200 889.3600 689.1200 889.8400 ;
        RECT 686.1200 894.8000 689.1200 895.2800 ;
        RECT 686.1200 878.4800 689.1200 878.9600 ;
        RECT 686.1200 873.0400 689.1200 873.5200 ;
        RECT 686.1200 883.9200 689.1200 884.4000 ;
        RECT 686.1200 927.4400 689.1200 927.9200 ;
        RECT 735.6800 927.4400 737.2800 927.9200 ;
        RECT 780.6800 927.4400 782.2800 927.9200 ;
        RECT 882.2200 862.1600 885.2200 862.6400 ;
        RECT 882.2200 867.6000 885.2200 868.0800 ;
        RECT 870.6800 862.1600 872.2800 862.6400 ;
        RECT 870.6800 867.6000 872.2800 868.0800 ;
        RECT 882.2200 845.8400 885.2200 846.3200 ;
        RECT 882.2200 851.2800 885.2200 851.7600 ;
        RECT 882.2200 856.7200 885.2200 857.2000 ;
        RECT 870.6800 845.8400 872.2800 846.3200 ;
        RECT 870.6800 851.2800 872.2800 851.7600 ;
        RECT 870.6800 856.7200 872.2800 857.2000 ;
        RECT 882.2200 834.9600 885.2200 835.4400 ;
        RECT 882.2200 840.4000 885.2200 840.8800 ;
        RECT 870.6800 834.9600 872.2800 835.4400 ;
        RECT 870.6800 840.4000 872.2800 840.8800 ;
        RECT 882.2200 818.6400 885.2200 819.1200 ;
        RECT 882.2200 824.0800 885.2200 824.5600 ;
        RECT 882.2200 829.5200 885.2200 830.0000 ;
        RECT 870.6800 818.6400 872.2800 819.1200 ;
        RECT 870.6800 824.0800 872.2800 824.5600 ;
        RECT 870.6800 829.5200 872.2800 830.0000 ;
        RECT 825.6800 862.1600 827.2800 862.6400 ;
        RECT 825.6800 867.6000 827.2800 868.0800 ;
        RECT 825.6800 845.8400 827.2800 846.3200 ;
        RECT 825.6800 851.2800 827.2800 851.7600 ;
        RECT 825.6800 856.7200 827.2800 857.2000 ;
        RECT 825.6800 834.9600 827.2800 835.4400 ;
        RECT 825.6800 840.4000 827.2800 840.8800 ;
        RECT 825.6800 818.6400 827.2800 819.1200 ;
        RECT 825.6800 824.0800 827.2800 824.5600 ;
        RECT 825.6800 829.5200 827.2800 830.0000 ;
        RECT 882.2200 807.7600 885.2200 808.2400 ;
        RECT 882.2200 813.2000 885.2200 813.6800 ;
        RECT 870.6800 807.7600 872.2800 808.2400 ;
        RECT 870.6800 813.2000 872.2800 813.6800 ;
        RECT 882.2200 791.4400 885.2200 791.9200 ;
        RECT 882.2200 796.8800 885.2200 797.3600 ;
        RECT 882.2200 802.3200 885.2200 802.8000 ;
        RECT 870.6800 791.4400 872.2800 791.9200 ;
        RECT 870.6800 796.8800 872.2800 797.3600 ;
        RECT 870.6800 802.3200 872.2800 802.8000 ;
        RECT 882.2200 780.5600 885.2200 781.0400 ;
        RECT 882.2200 786.0000 885.2200 786.4800 ;
        RECT 870.6800 780.5600 872.2800 781.0400 ;
        RECT 870.6800 786.0000 872.2800 786.4800 ;
        RECT 882.2200 775.1200 885.2200 775.6000 ;
        RECT 870.6800 775.1200 872.2800 775.6000 ;
        RECT 825.6800 807.7600 827.2800 808.2400 ;
        RECT 825.6800 813.2000 827.2800 813.6800 ;
        RECT 825.6800 791.4400 827.2800 791.9200 ;
        RECT 825.6800 796.8800 827.2800 797.3600 ;
        RECT 825.6800 802.3200 827.2800 802.8000 ;
        RECT 825.6800 780.5600 827.2800 781.0400 ;
        RECT 825.6800 786.0000 827.2800 786.4800 ;
        RECT 825.6800 775.1200 827.2800 775.6000 ;
        RECT 780.6800 862.1600 782.2800 862.6400 ;
        RECT 780.6800 867.6000 782.2800 868.0800 ;
        RECT 780.6800 845.8400 782.2800 846.3200 ;
        RECT 780.6800 851.2800 782.2800 851.7600 ;
        RECT 780.6800 856.7200 782.2800 857.2000 ;
        RECT 735.6800 862.1600 737.2800 862.6400 ;
        RECT 735.6800 867.6000 737.2800 868.0800 ;
        RECT 735.6800 845.8400 737.2800 846.3200 ;
        RECT 735.6800 851.2800 737.2800 851.7600 ;
        RECT 735.6800 856.7200 737.2800 857.2000 ;
        RECT 780.6800 834.9600 782.2800 835.4400 ;
        RECT 780.6800 840.4000 782.2800 840.8800 ;
        RECT 780.6800 818.6400 782.2800 819.1200 ;
        RECT 780.6800 824.0800 782.2800 824.5600 ;
        RECT 780.6800 829.5200 782.2800 830.0000 ;
        RECT 735.6800 834.9600 737.2800 835.4400 ;
        RECT 735.6800 840.4000 737.2800 840.8800 ;
        RECT 735.6800 818.6400 737.2800 819.1200 ;
        RECT 735.6800 824.0800 737.2800 824.5600 ;
        RECT 735.6800 829.5200 737.2800 830.0000 ;
        RECT 686.1200 862.1600 689.1200 862.6400 ;
        RECT 686.1200 867.6000 689.1200 868.0800 ;
        RECT 686.1200 851.2800 689.1200 851.7600 ;
        RECT 686.1200 845.8400 689.1200 846.3200 ;
        RECT 686.1200 856.7200 689.1200 857.2000 ;
        RECT 686.1200 834.9600 689.1200 835.4400 ;
        RECT 686.1200 840.4000 689.1200 840.8800 ;
        RECT 686.1200 824.0800 689.1200 824.5600 ;
        RECT 686.1200 818.6400 689.1200 819.1200 ;
        RECT 686.1200 829.5200 689.1200 830.0000 ;
        RECT 780.6800 807.7600 782.2800 808.2400 ;
        RECT 780.6800 813.2000 782.2800 813.6800 ;
        RECT 780.6800 791.4400 782.2800 791.9200 ;
        RECT 780.6800 796.8800 782.2800 797.3600 ;
        RECT 780.6800 802.3200 782.2800 802.8000 ;
        RECT 735.6800 807.7600 737.2800 808.2400 ;
        RECT 735.6800 813.2000 737.2800 813.6800 ;
        RECT 735.6800 791.4400 737.2800 791.9200 ;
        RECT 735.6800 796.8800 737.2800 797.3600 ;
        RECT 735.6800 802.3200 737.2800 802.8000 ;
        RECT 780.6800 786.0000 782.2800 786.4800 ;
        RECT 780.6800 780.5600 782.2800 781.0400 ;
        RECT 780.6800 775.1200 782.2800 775.6000 ;
        RECT 735.6800 786.0000 737.2800 786.4800 ;
        RECT 735.6800 780.5600 737.2800 781.0400 ;
        RECT 735.6800 775.1200 737.2800 775.6000 ;
        RECT 686.1200 807.7600 689.1200 808.2400 ;
        RECT 686.1200 813.2000 689.1200 813.6800 ;
        RECT 686.1200 796.8800 689.1200 797.3600 ;
        RECT 686.1200 791.4400 689.1200 791.9200 ;
        RECT 686.1200 802.3200 689.1200 802.8000 ;
        RECT 686.1200 780.5600 689.1200 781.0400 ;
        RECT 686.1200 786.0000 689.1200 786.4800 ;
        RECT 686.1200 775.1200 689.1200 775.6000 ;
        RECT 686.1200 973.3100 885.2200 976.3100 ;
        RECT 686.1200 768.2100 885.2200 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single2'
    PORT
      LAYER met4 ;
        RECT 1133.3400 2833.6100 1135.3400 2854.5400 ;
        RECT 906.3400 2833.6100 908.3400 2854.5400 ;
      LAYER met3 ;
        RECT 1133.3400 2850.0400 1135.3400 2850.5200 ;
        RECT 906.3400 2850.0400 908.3400 2850.5200 ;
        RECT 1133.3400 2839.1600 1135.3400 2839.6400 ;
        RECT 906.3400 2839.1600 908.3400 2839.6400 ;
        RECT 906.3400 2844.6000 908.3400 2845.0800 ;
        RECT 1133.3400 2844.6000 1135.3400 2845.0800 ;
        RECT 906.3400 2852.5400 1135.3400 2854.5400 ;
        RECT 906.3400 2833.6100 1135.3400 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single2'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 538.5700 1091.9000 746.6700 ;
        RECT 1045.9000 538.5700 1046.9000 746.6700 ;
        RECT 1000.9000 538.5700 1001.9000 746.6700 ;
        RECT 955.9000 538.5700 956.9000 746.6700 ;
        RECT 1132.3400 538.5700 1135.3400 746.6700 ;
        RECT 906.3400 538.5700 909.3400 746.6700 ;
      LAYER met3 ;
        RECT 1132.3400 735.8800 1135.3400 736.3600 ;
        RECT 1132.3400 741.3200 1135.3400 741.8000 ;
        RECT 1090.9000 735.8800 1091.9000 736.3600 ;
        RECT 1090.9000 741.3200 1091.9000 741.8000 ;
        RECT 1132.3400 719.5600 1135.3400 720.0400 ;
        RECT 1132.3400 725.0000 1135.3400 725.4800 ;
        RECT 1132.3400 730.4400 1135.3400 730.9200 ;
        RECT 1132.3400 714.1200 1135.3400 714.6000 ;
        RECT 1132.3400 703.2400 1135.3400 703.7200 ;
        RECT 1132.3400 708.6800 1135.3400 709.1600 ;
        RECT 1090.9000 719.5600 1091.9000 720.0400 ;
        RECT 1090.9000 725.0000 1091.9000 725.4800 ;
        RECT 1090.9000 730.4400 1091.9000 730.9200 ;
        RECT 1090.9000 703.2400 1091.9000 703.7200 ;
        RECT 1090.9000 708.6800 1091.9000 709.1600 ;
        RECT 1090.9000 714.1200 1091.9000 714.6000 ;
        RECT 1045.9000 735.8800 1046.9000 736.3600 ;
        RECT 1045.9000 741.3200 1046.9000 741.8000 ;
        RECT 1045.9000 719.5600 1046.9000 720.0400 ;
        RECT 1045.9000 725.0000 1046.9000 725.4800 ;
        RECT 1045.9000 730.4400 1046.9000 730.9200 ;
        RECT 1045.9000 703.2400 1046.9000 703.7200 ;
        RECT 1045.9000 708.6800 1046.9000 709.1600 ;
        RECT 1045.9000 714.1200 1046.9000 714.6000 ;
        RECT 1132.3400 692.3600 1135.3400 692.8400 ;
        RECT 1132.3400 697.8000 1135.3400 698.2800 ;
        RECT 1132.3400 686.9200 1135.3400 687.4000 ;
        RECT 1132.3400 681.4800 1135.3400 681.9600 ;
        RECT 1132.3400 676.0400 1135.3400 676.5200 ;
        RECT 1090.9000 692.3600 1091.9000 692.8400 ;
        RECT 1090.9000 697.8000 1091.9000 698.2800 ;
        RECT 1090.9000 676.0400 1091.9000 676.5200 ;
        RECT 1090.9000 681.4800 1091.9000 681.9600 ;
        RECT 1090.9000 686.9200 1091.9000 687.4000 ;
        RECT 1132.3400 659.7200 1135.3400 660.2000 ;
        RECT 1132.3400 665.1600 1135.3400 665.6400 ;
        RECT 1132.3400 670.6000 1135.3400 671.0800 ;
        RECT 1132.3400 654.2800 1135.3400 654.7600 ;
        RECT 1132.3400 643.4000 1135.3400 643.8800 ;
        RECT 1132.3400 648.8400 1135.3400 649.3200 ;
        RECT 1090.9000 659.7200 1091.9000 660.2000 ;
        RECT 1090.9000 665.1600 1091.9000 665.6400 ;
        RECT 1090.9000 670.6000 1091.9000 671.0800 ;
        RECT 1090.9000 643.4000 1091.9000 643.8800 ;
        RECT 1090.9000 648.8400 1091.9000 649.3200 ;
        RECT 1090.9000 654.2800 1091.9000 654.7600 ;
        RECT 1045.9000 692.3600 1046.9000 692.8400 ;
        RECT 1045.9000 697.8000 1046.9000 698.2800 ;
        RECT 1045.9000 676.0400 1046.9000 676.5200 ;
        RECT 1045.9000 681.4800 1046.9000 681.9600 ;
        RECT 1045.9000 686.9200 1046.9000 687.4000 ;
        RECT 1045.9000 659.7200 1046.9000 660.2000 ;
        RECT 1045.9000 665.1600 1046.9000 665.6400 ;
        RECT 1045.9000 670.6000 1046.9000 671.0800 ;
        RECT 1045.9000 643.4000 1046.9000 643.8800 ;
        RECT 1045.9000 648.8400 1046.9000 649.3200 ;
        RECT 1045.9000 654.2800 1046.9000 654.7600 ;
        RECT 1000.9000 735.8800 1001.9000 736.3600 ;
        RECT 1000.9000 741.3200 1001.9000 741.8000 ;
        RECT 1000.9000 719.5600 1001.9000 720.0400 ;
        RECT 1000.9000 725.0000 1001.9000 725.4800 ;
        RECT 1000.9000 730.4400 1001.9000 730.9200 ;
        RECT 1000.9000 703.2400 1001.9000 703.7200 ;
        RECT 1000.9000 708.6800 1001.9000 709.1600 ;
        RECT 1000.9000 714.1200 1001.9000 714.6000 ;
        RECT 955.9000 735.8800 956.9000 736.3600 ;
        RECT 955.9000 741.3200 956.9000 741.8000 ;
        RECT 906.3400 741.3200 909.3400 741.8000 ;
        RECT 906.3400 735.8800 909.3400 736.3600 ;
        RECT 955.9000 719.5600 956.9000 720.0400 ;
        RECT 955.9000 725.0000 956.9000 725.4800 ;
        RECT 955.9000 730.4400 956.9000 730.9200 ;
        RECT 955.9000 703.2400 956.9000 703.7200 ;
        RECT 955.9000 708.6800 956.9000 709.1600 ;
        RECT 955.9000 714.1200 956.9000 714.6000 ;
        RECT 906.3400 730.4400 909.3400 730.9200 ;
        RECT 906.3400 719.5600 909.3400 720.0400 ;
        RECT 906.3400 725.0000 909.3400 725.4800 ;
        RECT 906.3400 714.1200 909.3400 714.6000 ;
        RECT 906.3400 703.2400 909.3400 703.7200 ;
        RECT 906.3400 708.6800 909.3400 709.1600 ;
        RECT 1000.9000 692.3600 1001.9000 692.8400 ;
        RECT 1000.9000 697.8000 1001.9000 698.2800 ;
        RECT 1000.9000 676.0400 1001.9000 676.5200 ;
        RECT 1000.9000 681.4800 1001.9000 681.9600 ;
        RECT 1000.9000 686.9200 1001.9000 687.4000 ;
        RECT 1000.9000 659.7200 1001.9000 660.2000 ;
        RECT 1000.9000 665.1600 1001.9000 665.6400 ;
        RECT 1000.9000 670.6000 1001.9000 671.0800 ;
        RECT 1000.9000 643.4000 1001.9000 643.8800 ;
        RECT 1000.9000 648.8400 1001.9000 649.3200 ;
        RECT 1000.9000 654.2800 1001.9000 654.7600 ;
        RECT 955.9000 692.3600 956.9000 692.8400 ;
        RECT 955.9000 697.8000 956.9000 698.2800 ;
        RECT 955.9000 676.0400 956.9000 676.5200 ;
        RECT 955.9000 681.4800 956.9000 681.9600 ;
        RECT 955.9000 686.9200 956.9000 687.4000 ;
        RECT 906.3400 697.8000 909.3400 698.2800 ;
        RECT 906.3400 692.3600 909.3400 692.8400 ;
        RECT 906.3400 681.4800 909.3400 681.9600 ;
        RECT 906.3400 686.9200 909.3400 687.4000 ;
        RECT 906.3400 676.0400 909.3400 676.5200 ;
        RECT 955.9000 659.7200 956.9000 660.2000 ;
        RECT 955.9000 665.1600 956.9000 665.6400 ;
        RECT 955.9000 670.6000 956.9000 671.0800 ;
        RECT 955.9000 643.4000 956.9000 643.8800 ;
        RECT 955.9000 648.8400 956.9000 649.3200 ;
        RECT 955.9000 654.2800 956.9000 654.7600 ;
        RECT 906.3400 670.6000 909.3400 671.0800 ;
        RECT 906.3400 659.7200 909.3400 660.2000 ;
        RECT 906.3400 665.1600 909.3400 665.6400 ;
        RECT 906.3400 654.2800 909.3400 654.7600 ;
        RECT 906.3400 643.4000 909.3400 643.8800 ;
        RECT 906.3400 648.8400 909.3400 649.3200 ;
        RECT 1132.3400 632.5200 1135.3400 633.0000 ;
        RECT 1132.3400 637.9600 1135.3400 638.4400 ;
        RECT 1132.3400 627.0800 1135.3400 627.5600 ;
        RECT 1132.3400 621.6400 1135.3400 622.1200 ;
        RECT 1132.3400 616.2000 1135.3400 616.6800 ;
        RECT 1090.9000 632.5200 1091.9000 633.0000 ;
        RECT 1090.9000 637.9600 1091.9000 638.4400 ;
        RECT 1090.9000 616.2000 1091.9000 616.6800 ;
        RECT 1090.9000 621.6400 1091.9000 622.1200 ;
        RECT 1090.9000 627.0800 1091.9000 627.5600 ;
        RECT 1132.3400 599.8800 1135.3400 600.3600 ;
        RECT 1132.3400 605.3200 1135.3400 605.8000 ;
        RECT 1132.3400 610.7600 1135.3400 611.2400 ;
        RECT 1132.3400 594.4400 1135.3400 594.9200 ;
        RECT 1132.3400 583.5600 1135.3400 584.0400 ;
        RECT 1132.3400 589.0000 1135.3400 589.4800 ;
        RECT 1090.9000 599.8800 1091.9000 600.3600 ;
        RECT 1090.9000 605.3200 1091.9000 605.8000 ;
        RECT 1090.9000 610.7600 1091.9000 611.2400 ;
        RECT 1090.9000 583.5600 1091.9000 584.0400 ;
        RECT 1090.9000 589.0000 1091.9000 589.4800 ;
        RECT 1090.9000 594.4400 1091.9000 594.9200 ;
        RECT 1045.9000 632.5200 1046.9000 633.0000 ;
        RECT 1045.9000 637.9600 1046.9000 638.4400 ;
        RECT 1045.9000 616.2000 1046.9000 616.6800 ;
        RECT 1045.9000 621.6400 1046.9000 622.1200 ;
        RECT 1045.9000 627.0800 1046.9000 627.5600 ;
        RECT 1045.9000 599.8800 1046.9000 600.3600 ;
        RECT 1045.9000 605.3200 1046.9000 605.8000 ;
        RECT 1045.9000 610.7600 1046.9000 611.2400 ;
        RECT 1045.9000 583.5600 1046.9000 584.0400 ;
        RECT 1045.9000 589.0000 1046.9000 589.4800 ;
        RECT 1045.9000 594.4400 1046.9000 594.9200 ;
        RECT 1132.3400 572.6800 1135.3400 573.1600 ;
        RECT 1132.3400 578.1200 1135.3400 578.6000 ;
        RECT 1132.3400 567.2400 1135.3400 567.7200 ;
        RECT 1132.3400 561.8000 1135.3400 562.2800 ;
        RECT 1132.3400 556.3600 1135.3400 556.8400 ;
        RECT 1090.9000 572.6800 1091.9000 573.1600 ;
        RECT 1090.9000 578.1200 1091.9000 578.6000 ;
        RECT 1090.9000 556.3600 1091.9000 556.8400 ;
        RECT 1090.9000 561.8000 1091.9000 562.2800 ;
        RECT 1090.9000 567.2400 1091.9000 567.7200 ;
        RECT 1132.3400 545.4800 1135.3400 545.9600 ;
        RECT 1132.3400 550.9200 1135.3400 551.4000 ;
        RECT 1090.9000 545.4800 1091.9000 545.9600 ;
        RECT 1090.9000 550.9200 1091.9000 551.4000 ;
        RECT 1045.9000 572.6800 1046.9000 573.1600 ;
        RECT 1045.9000 578.1200 1046.9000 578.6000 ;
        RECT 1045.9000 556.3600 1046.9000 556.8400 ;
        RECT 1045.9000 561.8000 1046.9000 562.2800 ;
        RECT 1045.9000 567.2400 1046.9000 567.7200 ;
        RECT 1045.9000 545.4800 1046.9000 545.9600 ;
        RECT 1045.9000 550.9200 1046.9000 551.4000 ;
        RECT 1000.9000 632.5200 1001.9000 633.0000 ;
        RECT 1000.9000 637.9600 1001.9000 638.4400 ;
        RECT 1000.9000 616.2000 1001.9000 616.6800 ;
        RECT 1000.9000 621.6400 1001.9000 622.1200 ;
        RECT 1000.9000 627.0800 1001.9000 627.5600 ;
        RECT 1000.9000 599.8800 1001.9000 600.3600 ;
        RECT 1000.9000 605.3200 1001.9000 605.8000 ;
        RECT 1000.9000 610.7600 1001.9000 611.2400 ;
        RECT 1000.9000 583.5600 1001.9000 584.0400 ;
        RECT 1000.9000 589.0000 1001.9000 589.4800 ;
        RECT 1000.9000 594.4400 1001.9000 594.9200 ;
        RECT 955.9000 632.5200 956.9000 633.0000 ;
        RECT 955.9000 637.9600 956.9000 638.4400 ;
        RECT 955.9000 616.2000 956.9000 616.6800 ;
        RECT 955.9000 621.6400 956.9000 622.1200 ;
        RECT 955.9000 627.0800 956.9000 627.5600 ;
        RECT 906.3400 637.9600 909.3400 638.4400 ;
        RECT 906.3400 632.5200 909.3400 633.0000 ;
        RECT 906.3400 621.6400 909.3400 622.1200 ;
        RECT 906.3400 627.0800 909.3400 627.5600 ;
        RECT 906.3400 616.2000 909.3400 616.6800 ;
        RECT 955.9000 599.8800 956.9000 600.3600 ;
        RECT 955.9000 605.3200 956.9000 605.8000 ;
        RECT 955.9000 610.7600 956.9000 611.2400 ;
        RECT 955.9000 583.5600 956.9000 584.0400 ;
        RECT 955.9000 589.0000 956.9000 589.4800 ;
        RECT 955.9000 594.4400 956.9000 594.9200 ;
        RECT 906.3400 610.7600 909.3400 611.2400 ;
        RECT 906.3400 599.8800 909.3400 600.3600 ;
        RECT 906.3400 605.3200 909.3400 605.8000 ;
        RECT 906.3400 594.4400 909.3400 594.9200 ;
        RECT 906.3400 583.5600 909.3400 584.0400 ;
        RECT 906.3400 589.0000 909.3400 589.4800 ;
        RECT 1000.9000 572.6800 1001.9000 573.1600 ;
        RECT 1000.9000 578.1200 1001.9000 578.6000 ;
        RECT 1000.9000 556.3600 1001.9000 556.8400 ;
        RECT 1000.9000 561.8000 1001.9000 562.2800 ;
        RECT 1000.9000 567.2400 1001.9000 567.7200 ;
        RECT 1000.9000 545.4800 1001.9000 545.9600 ;
        RECT 1000.9000 550.9200 1001.9000 551.4000 ;
        RECT 955.9000 572.6800 956.9000 573.1600 ;
        RECT 955.9000 578.1200 956.9000 578.6000 ;
        RECT 955.9000 556.3600 956.9000 556.8400 ;
        RECT 955.9000 561.8000 956.9000 562.2800 ;
        RECT 955.9000 567.2400 956.9000 567.7200 ;
        RECT 906.3400 578.1200 909.3400 578.6000 ;
        RECT 906.3400 572.6800 909.3400 573.1600 ;
        RECT 906.3400 561.8000 909.3400 562.2800 ;
        RECT 906.3400 567.2400 909.3400 567.7200 ;
        RECT 906.3400 556.3600 909.3400 556.8400 ;
        RECT 955.9000 545.4800 956.9000 545.9600 ;
        RECT 955.9000 550.9200 956.9000 551.4000 ;
        RECT 906.3400 550.9200 909.3400 551.4000 ;
        RECT 906.3400 545.4800 909.3400 545.9600 ;
        RECT 906.3400 743.6700 1135.3400 746.6700 ;
        RECT 906.3400 538.5700 1135.3400 541.5700 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 308.9300 1091.9000 517.0300 ;
        RECT 1045.9000 308.9300 1046.9000 517.0300 ;
        RECT 1000.9000 308.9300 1001.9000 517.0300 ;
        RECT 955.9000 308.9300 956.9000 517.0300 ;
        RECT 1132.3400 308.9300 1135.3400 517.0300 ;
        RECT 906.3400 308.9300 909.3400 517.0300 ;
      LAYER met3 ;
        RECT 1132.3400 506.2400 1135.3400 506.7200 ;
        RECT 1132.3400 511.6800 1135.3400 512.1600 ;
        RECT 1090.9000 506.2400 1091.9000 506.7200 ;
        RECT 1090.9000 511.6800 1091.9000 512.1600 ;
        RECT 1132.3400 489.9200 1135.3400 490.4000 ;
        RECT 1132.3400 495.3600 1135.3400 495.8400 ;
        RECT 1132.3400 500.8000 1135.3400 501.2800 ;
        RECT 1132.3400 484.4800 1135.3400 484.9600 ;
        RECT 1132.3400 473.6000 1135.3400 474.0800 ;
        RECT 1132.3400 479.0400 1135.3400 479.5200 ;
        RECT 1090.9000 489.9200 1091.9000 490.4000 ;
        RECT 1090.9000 495.3600 1091.9000 495.8400 ;
        RECT 1090.9000 500.8000 1091.9000 501.2800 ;
        RECT 1090.9000 473.6000 1091.9000 474.0800 ;
        RECT 1090.9000 479.0400 1091.9000 479.5200 ;
        RECT 1090.9000 484.4800 1091.9000 484.9600 ;
        RECT 1045.9000 506.2400 1046.9000 506.7200 ;
        RECT 1045.9000 511.6800 1046.9000 512.1600 ;
        RECT 1045.9000 489.9200 1046.9000 490.4000 ;
        RECT 1045.9000 495.3600 1046.9000 495.8400 ;
        RECT 1045.9000 500.8000 1046.9000 501.2800 ;
        RECT 1045.9000 473.6000 1046.9000 474.0800 ;
        RECT 1045.9000 479.0400 1046.9000 479.5200 ;
        RECT 1045.9000 484.4800 1046.9000 484.9600 ;
        RECT 1132.3400 462.7200 1135.3400 463.2000 ;
        RECT 1132.3400 468.1600 1135.3400 468.6400 ;
        RECT 1132.3400 457.2800 1135.3400 457.7600 ;
        RECT 1132.3400 451.8400 1135.3400 452.3200 ;
        RECT 1132.3400 446.4000 1135.3400 446.8800 ;
        RECT 1090.9000 462.7200 1091.9000 463.2000 ;
        RECT 1090.9000 468.1600 1091.9000 468.6400 ;
        RECT 1090.9000 446.4000 1091.9000 446.8800 ;
        RECT 1090.9000 451.8400 1091.9000 452.3200 ;
        RECT 1090.9000 457.2800 1091.9000 457.7600 ;
        RECT 1132.3400 430.0800 1135.3400 430.5600 ;
        RECT 1132.3400 435.5200 1135.3400 436.0000 ;
        RECT 1132.3400 440.9600 1135.3400 441.4400 ;
        RECT 1132.3400 424.6400 1135.3400 425.1200 ;
        RECT 1132.3400 413.7600 1135.3400 414.2400 ;
        RECT 1132.3400 419.2000 1135.3400 419.6800 ;
        RECT 1090.9000 430.0800 1091.9000 430.5600 ;
        RECT 1090.9000 435.5200 1091.9000 436.0000 ;
        RECT 1090.9000 440.9600 1091.9000 441.4400 ;
        RECT 1090.9000 413.7600 1091.9000 414.2400 ;
        RECT 1090.9000 419.2000 1091.9000 419.6800 ;
        RECT 1090.9000 424.6400 1091.9000 425.1200 ;
        RECT 1045.9000 462.7200 1046.9000 463.2000 ;
        RECT 1045.9000 468.1600 1046.9000 468.6400 ;
        RECT 1045.9000 446.4000 1046.9000 446.8800 ;
        RECT 1045.9000 451.8400 1046.9000 452.3200 ;
        RECT 1045.9000 457.2800 1046.9000 457.7600 ;
        RECT 1045.9000 430.0800 1046.9000 430.5600 ;
        RECT 1045.9000 435.5200 1046.9000 436.0000 ;
        RECT 1045.9000 440.9600 1046.9000 441.4400 ;
        RECT 1045.9000 413.7600 1046.9000 414.2400 ;
        RECT 1045.9000 419.2000 1046.9000 419.6800 ;
        RECT 1045.9000 424.6400 1046.9000 425.1200 ;
        RECT 1000.9000 506.2400 1001.9000 506.7200 ;
        RECT 1000.9000 511.6800 1001.9000 512.1600 ;
        RECT 1000.9000 489.9200 1001.9000 490.4000 ;
        RECT 1000.9000 495.3600 1001.9000 495.8400 ;
        RECT 1000.9000 500.8000 1001.9000 501.2800 ;
        RECT 1000.9000 473.6000 1001.9000 474.0800 ;
        RECT 1000.9000 479.0400 1001.9000 479.5200 ;
        RECT 1000.9000 484.4800 1001.9000 484.9600 ;
        RECT 955.9000 506.2400 956.9000 506.7200 ;
        RECT 955.9000 511.6800 956.9000 512.1600 ;
        RECT 906.3400 511.6800 909.3400 512.1600 ;
        RECT 906.3400 506.2400 909.3400 506.7200 ;
        RECT 955.9000 489.9200 956.9000 490.4000 ;
        RECT 955.9000 495.3600 956.9000 495.8400 ;
        RECT 955.9000 500.8000 956.9000 501.2800 ;
        RECT 955.9000 473.6000 956.9000 474.0800 ;
        RECT 955.9000 479.0400 956.9000 479.5200 ;
        RECT 955.9000 484.4800 956.9000 484.9600 ;
        RECT 906.3400 500.8000 909.3400 501.2800 ;
        RECT 906.3400 489.9200 909.3400 490.4000 ;
        RECT 906.3400 495.3600 909.3400 495.8400 ;
        RECT 906.3400 484.4800 909.3400 484.9600 ;
        RECT 906.3400 473.6000 909.3400 474.0800 ;
        RECT 906.3400 479.0400 909.3400 479.5200 ;
        RECT 1000.9000 462.7200 1001.9000 463.2000 ;
        RECT 1000.9000 468.1600 1001.9000 468.6400 ;
        RECT 1000.9000 446.4000 1001.9000 446.8800 ;
        RECT 1000.9000 451.8400 1001.9000 452.3200 ;
        RECT 1000.9000 457.2800 1001.9000 457.7600 ;
        RECT 1000.9000 430.0800 1001.9000 430.5600 ;
        RECT 1000.9000 435.5200 1001.9000 436.0000 ;
        RECT 1000.9000 440.9600 1001.9000 441.4400 ;
        RECT 1000.9000 413.7600 1001.9000 414.2400 ;
        RECT 1000.9000 419.2000 1001.9000 419.6800 ;
        RECT 1000.9000 424.6400 1001.9000 425.1200 ;
        RECT 955.9000 462.7200 956.9000 463.2000 ;
        RECT 955.9000 468.1600 956.9000 468.6400 ;
        RECT 955.9000 446.4000 956.9000 446.8800 ;
        RECT 955.9000 451.8400 956.9000 452.3200 ;
        RECT 955.9000 457.2800 956.9000 457.7600 ;
        RECT 906.3400 468.1600 909.3400 468.6400 ;
        RECT 906.3400 462.7200 909.3400 463.2000 ;
        RECT 906.3400 451.8400 909.3400 452.3200 ;
        RECT 906.3400 457.2800 909.3400 457.7600 ;
        RECT 906.3400 446.4000 909.3400 446.8800 ;
        RECT 955.9000 430.0800 956.9000 430.5600 ;
        RECT 955.9000 435.5200 956.9000 436.0000 ;
        RECT 955.9000 440.9600 956.9000 441.4400 ;
        RECT 955.9000 413.7600 956.9000 414.2400 ;
        RECT 955.9000 419.2000 956.9000 419.6800 ;
        RECT 955.9000 424.6400 956.9000 425.1200 ;
        RECT 906.3400 440.9600 909.3400 441.4400 ;
        RECT 906.3400 430.0800 909.3400 430.5600 ;
        RECT 906.3400 435.5200 909.3400 436.0000 ;
        RECT 906.3400 424.6400 909.3400 425.1200 ;
        RECT 906.3400 413.7600 909.3400 414.2400 ;
        RECT 906.3400 419.2000 909.3400 419.6800 ;
        RECT 1132.3400 402.8800 1135.3400 403.3600 ;
        RECT 1132.3400 408.3200 1135.3400 408.8000 ;
        RECT 1132.3400 397.4400 1135.3400 397.9200 ;
        RECT 1132.3400 392.0000 1135.3400 392.4800 ;
        RECT 1132.3400 386.5600 1135.3400 387.0400 ;
        RECT 1090.9000 402.8800 1091.9000 403.3600 ;
        RECT 1090.9000 408.3200 1091.9000 408.8000 ;
        RECT 1090.9000 386.5600 1091.9000 387.0400 ;
        RECT 1090.9000 392.0000 1091.9000 392.4800 ;
        RECT 1090.9000 397.4400 1091.9000 397.9200 ;
        RECT 1132.3400 370.2400 1135.3400 370.7200 ;
        RECT 1132.3400 375.6800 1135.3400 376.1600 ;
        RECT 1132.3400 381.1200 1135.3400 381.6000 ;
        RECT 1132.3400 364.8000 1135.3400 365.2800 ;
        RECT 1132.3400 353.9200 1135.3400 354.4000 ;
        RECT 1132.3400 359.3600 1135.3400 359.8400 ;
        RECT 1090.9000 370.2400 1091.9000 370.7200 ;
        RECT 1090.9000 375.6800 1091.9000 376.1600 ;
        RECT 1090.9000 381.1200 1091.9000 381.6000 ;
        RECT 1090.9000 353.9200 1091.9000 354.4000 ;
        RECT 1090.9000 359.3600 1091.9000 359.8400 ;
        RECT 1090.9000 364.8000 1091.9000 365.2800 ;
        RECT 1045.9000 402.8800 1046.9000 403.3600 ;
        RECT 1045.9000 408.3200 1046.9000 408.8000 ;
        RECT 1045.9000 386.5600 1046.9000 387.0400 ;
        RECT 1045.9000 392.0000 1046.9000 392.4800 ;
        RECT 1045.9000 397.4400 1046.9000 397.9200 ;
        RECT 1045.9000 370.2400 1046.9000 370.7200 ;
        RECT 1045.9000 375.6800 1046.9000 376.1600 ;
        RECT 1045.9000 381.1200 1046.9000 381.6000 ;
        RECT 1045.9000 353.9200 1046.9000 354.4000 ;
        RECT 1045.9000 359.3600 1046.9000 359.8400 ;
        RECT 1045.9000 364.8000 1046.9000 365.2800 ;
        RECT 1132.3400 343.0400 1135.3400 343.5200 ;
        RECT 1132.3400 348.4800 1135.3400 348.9600 ;
        RECT 1132.3400 337.6000 1135.3400 338.0800 ;
        RECT 1132.3400 332.1600 1135.3400 332.6400 ;
        RECT 1132.3400 326.7200 1135.3400 327.2000 ;
        RECT 1090.9000 343.0400 1091.9000 343.5200 ;
        RECT 1090.9000 348.4800 1091.9000 348.9600 ;
        RECT 1090.9000 326.7200 1091.9000 327.2000 ;
        RECT 1090.9000 332.1600 1091.9000 332.6400 ;
        RECT 1090.9000 337.6000 1091.9000 338.0800 ;
        RECT 1132.3400 315.8400 1135.3400 316.3200 ;
        RECT 1132.3400 321.2800 1135.3400 321.7600 ;
        RECT 1090.9000 315.8400 1091.9000 316.3200 ;
        RECT 1090.9000 321.2800 1091.9000 321.7600 ;
        RECT 1045.9000 343.0400 1046.9000 343.5200 ;
        RECT 1045.9000 348.4800 1046.9000 348.9600 ;
        RECT 1045.9000 326.7200 1046.9000 327.2000 ;
        RECT 1045.9000 332.1600 1046.9000 332.6400 ;
        RECT 1045.9000 337.6000 1046.9000 338.0800 ;
        RECT 1045.9000 315.8400 1046.9000 316.3200 ;
        RECT 1045.9000 321.2800 1046.9000 321.7600 ;
        RECT 1000.9000 402.8800 1001.9000 403.3600 ;
        RECT 1000.9000 408.3200 1001.9000 408.8000 ;
        RECT 1000.9000 386.5600 1001.9000 387.0400 ;
        RECT 1000.9000 392.0000 1001.9000 392.4800 ;
        RECT 1000.9000 397.4400 1001.9000 397.9200 ;
        RECT 1000.9000 370.2400 1001.9000 370.7200 ;
        RECT 1000.9000 375.6800 1001.9000 376.1600 ;
        RECT 1000.9000 381.1200 1001.9000 381.6000 ;
        RECT 1000.9000 353.9200 1001.9000 354.4000 ;
        RECT 1000.9000 359.3600 1001.9000 359.8400 ;
        RECT 1000.9000 364.8000 1001.9000 365.2800 ;
        RECT 955.9000 402.8800 956.9000 403.3600 ;
        RECT 955.9000 408.3200 956.9000 408.8000 ;
        RECT 955.9000 386.5600 956.9000 387.0400 ;
        RECT 955.9000 392.0000 956.9000 392.4800 ;
        RECT 955.9000 397.4400 956.9000 397.9200 ;
        RECT 906.3400 408.3200 909.3400 408.8000 ;
        RECT 906.3400 402.8800 909.3400 403.3600 ;
        RECT 906.3400 392.0000 909.3400 392.4800 ;
        RECT 906.3400 397.4400 909.3400 397.9200 ;
        RECT 906.3400 386.5600 909.3400 387.0400 ;
        RECT 955.9000 370.2400 956.9000 370.7200 ;
        RECT 955.9000 375.6800 956.9000 376.1600 ;
        RECT 955.9000 381.1200 956.9000 381.6000 ;
        RECT 955.9000 353.9200 956.9000 354.4000 ;
        RECT 955.9000 359.3600 956.9000 359.8400 ;
        RECT 955.9000 364.8000 956.9000 365.2800 ;
        RECT 906.3400 381.1200 909.3400 381.6000 ;
        RECT 906.3400 370.2400 909.3400 370.7200 ;
        RECT 906.3400 375.6800 909.3400 376.1600 ;
        RECT 906.3400 364.8000 909.3400 365.2800 ;
        RECT 906.3400 353.9200 909.3400 354.4000 ;
        RECT 906.3400 359.3600 909.3400 359.8400 ;
        RECT 1000.9000 343.0400 1001.9000 343.5200 ;
        RECT 1000.9000 348.4800 1001.9000 348.9600 ;
        RECT 1000.9000 326.7200 1001.9000 327.2000 ;
        RECT 1000.9000 332.1600 1001.9000 332.6400 ;
        RECT 1000.9000 337.6000 1001.9000 338.0800 ;
        RECT 1000.9000 315.8400 1001.9000 316.3200 ;
        RECT 1000.9000 321.2800 1001.9000 321.7600 ;
        RECT 955.9000 343.0400 956.9000 343.5200 ;
        RECT 955.9000 348.4800 956.9000 348.9600 ;
        RECT 955.9000 326.7200 956.9000 327.2000 ;
        RECT 955.9000 332.1600 956.9000 332.6400 ;
        RECT 955.9000 337.6000 956.9000 338.0800 ;
        RECT 906.3400 348.4800 909.3400 348.9600 ;
        RECT 906.3400 343.0400 909.3400 343.5200 ;
        RECT 906.3400 332.1600 909.3400 332.6400 ;
        RECT 906.3400 337.6000 909.3400 338.0800 ;
        RECT 906.3400 326.7200 909.3400 327.2000 ;
        RECT 955.9000 315.8400 956.9000 316.3200 ;
        RECT 955.9000 321.2800 956.9000 321.7600 ;
        RECT 906.3400 321.2800 909.3400 321.7600 ;
        RECT 906.3400 315.8400 909.3400 316.3200 ;
        RECT 906.3400 514.0300 1135.3400 517.0300 ;
        RECT 906.3400 308.9300 1135.3400 311.9300 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 79.2900 1091.9000 287.3900 ;
        RECT 1045.9000 79.2900 1046.9000 287.3900 ;
        RECT 1000.9000 79.2900 1001.9000 287.3900 ;
        RECT 955.9000 79.2900 956.9000 287.3900 ;
        RECT 1132.3400 79.2900 1135.3400 287.3900 ;
        RECT 906.3400 79.2900 909.3400 287.3900 ;
      LAYER met3 ;
        RECT 1132.3400 276.6000 1135.3400 277.0800 ;
        RECT 1132.3400 282.0400 1135.3400 282.5200 ;
        RECT 1090.9000 276.6000 1091.9000 277.0800 ;
        RECT 1090.9000 282.0400 1091.9000 282.5200 ;
        RECT 1132.3400 260.2800 1135.3400 260.7600 ;
        RECT 1132.3400 265.7200 1135.3400 266.2000 ;
        RECT 1132.3400 271.1600 1135.3400 271.6400 ;
        RECT 1132.3400 254.8400 1135.3400 255.3200 ;
        RECT 1132.3400 243.9600 1135.3400 244.4400 ;
        RECT 1132.3400 249.4000 1135.3400 249.8800 ;
        RECT 1090.9000 260.2800 1091.9000 260.7600 ;
        RECT 1090.9000 265.7200 1091.9000 266.2000 ;
        RECT 1090.9000 271.1600 1091.9000 271.6400 ;
        RECT 1090.9000 243.9600 1091.9000 244.4400 ;
        RECT 1090.9000 249.4000 1091.9000 249.8800 ;
        RECT 1090.9000 254.8400 1091.9000 255.3200 ;
        RECT 1045.9000 276.6000 1046.9000 277.0800 ;
        RECT 1045.9000 282.0400 1046.9000 282.5200 ;
        RECT 1045.9000 260.2800 1046.9000 260.7600 ;
        RECT 1045.9000 265.7200 1046.9000 266.2000 ;
        RECT 1045.9000 271.1600 1046.9000 271.6400 ;
        RECT 1045.9000 243.9600 1046.9000 244.4400 ;
        RECT 1045.9000 249.4000 1046.9000 249.8800 ;
        RECT 1045.9000 254.8400 1046.9000 255.3200 ;
        RECT 1132.3400 233.0800 1135.3400 233.5600 ;
        RECT 1132.3400 238.5200 1135.3400 239.0000 ;
        RECT 1132.3400 227.6400 1135.3400 228.1200 ;
        RECT 1132.3400 222.2000 1135.3400 222.6800 ;
        RECT 1132.3400 216.7600 1135.3400 217.2400 ;
        RECT 1090.9000 233.0800 1091.9000 233.5600 ;
        RECT 1090.9000 238.5200 1091.9000 239.0000 ;
        RECT 1090.9000 216.7600 1091.9000 217.2400 ;
        RECT 1090.9000 222.2000 1091.9000 222.6800 ;
        RECT 1090.9000 227.6400 1091.9000 228.1200 ;
        RECT 1132.3400 200.4400 1135.3400 200.9200 ;
        RECT 1132.3400 205.8800 1135.3400 206.3600 ;
        RECT 1132.3400 211.3200 1135.3400 211.8000 ;
        RECT 1132.3400 195.0000 1135.3400 195.4800 ;
        RECT 1132.3400 184.1200 1135.3400 184.6000 ;
        RECT 1132.3400 189.5600 1135.3400 190.0400 ;
        RECT 1090.9000 200.4400 1091.9000 200.9200 ;
        RECT 1090.9000 205.8800 1091.9000 206.3600 ;
        RECT 1090.9000 211.3200 1091.9000 211.8000 ;
        RECT 1090.9000 184.1200 1091.9000 184.6000 ;
        RECT 1090.9000 189.5600 1091.9000 190.0400 ;
        RECT 1090.9000 195.0000 1091.9000 195.4800 ;
        RECT 1045.9000 233.0800 1046.9000 233.5600 ;
        RECT 1045.9000 238.5200 1046.9000 239.0000 ;
        RECT 1045.9000 216.7600 1046.9000 217.2400 ;
        RECT 1045.9000 222.2000 1046.9000 222.6800 ;
        RECT 1045.9000 227.6400 1046.9000 228.1200 ;
        RECT 1045.9000 200.4400 1046.9000 200.9200 ;
        RECT 1045.9000 205.8800 1046.9000 206.3600 ;
        RECT 1045.9000 211.3200 1046.9000 211.8000 ;
        RECT 1045.9000 184.1200 1046.9000 184.6000 ;
        RECT 1045.9000 189.5600 1046.9000 190.0400 ;
        RECT 1045.9000 195.0000 1046.9000 195.4800 ;
        RECT 1000.9000 276.6000 1001.9000 277.0800 ;
        RECT 1000.9000 282.0400 1001.9000 282.5200 ;
        RECT 1000.9000 260.2800 1001.9000 260.7600 ;
        RECT 1000.9000 265.7200 1001.9000 266.2000 ;
        RECT 1000.9000 271.1600 1001.9000 271.6400 ;
        RECT 1000.9000 243.9600 1001.9000 244.4400 ;
        RECT 1000.9000 249.4000 1001.9000 249.8800 ;
        RECT 1000.9000 254.8400 1001.9000 255.3200 ;
        RECT 955.9000 276.6000 956.9000 277.0800 ;
        RECT 955.9000 282.0400 956.9000 282.5200 ;
        RECT 906.3400 282.0400 909.3400 282.5200 ;
        RECT 906.3400 276.6000 909.3400 277.0800 ;
        RECT 955.9000 260.2800 956.9000 260.7600 ;
        RECT 955.9000 265.7200 956.9000 266.2000 ;
        RECT 955.9000 271.1600 956.9000 271.6400 ;
        RECT 955.9000 243.9600 956.9000 244.4400 ;
        RECT 955.9000 249.4000 956.9000 249.8800 ;
        RECT 955.9000 254.8400 956.9000 255.3200 ;
        RECT 906.3400 271.1600 909.3400 271.6400 ;
        RECT 906.3400 260.2800 909.3400 260.7600 ;
        RECT 906.3400 265.7200 909.3400 266.2000 ;
        RECT 906.3400 254.8400 909.3400 255.3200 ;
        RECT 906.3400 243.9600 909.3400 244.4400 ;
        RECT 906.3400 249.4000 909.3400 249.8800 ;
        RECT 1000.9000 233.0800 1001.9000 233.5600 ;
        RECT 1000.9000 238.5200 1001.9000 239.0000 ;
        RECT 1000.9000 216.7600 1001.9000 217.2400 ;
        RECT 1000.9000 222.2000 1001.9000 222.6800 ;
        RECT 1000.9000 227.6400 1001.9000 228.1200 ;
        RECT 1000.9000 200.4400 1001.9000 200.9200 ;
        RECT 1000.9000 205.8800 1001.9000 206.3600 ;
        RECT 1000.9000 211.3200 1001.9000 211.8000 ;
        RECT 1000.9000 184.1200 1001.9000 184.6000 ;
        RECT 1000.9000 189.5600 1001.9000 190.0400 ;
        RECT 1000.9000 195.0000 1001.9000 195.4800 ;
        RECT 955.9000 233.0800 956.9000 233.5600 ;
        RECT 955.9000 238.5200 956.9000 239.0000 ;
        RECT 955.9000 216.7600 956.9000 217.2400 ;
        RECT 955.9000 222.2000 956.9000 222.6800 ;
        RECT 955.9000 227.6400 956.9000 228.1200 ;
        RECT 906.3400 238.5200 909.3400 239.0000 ;
        RECT 906.3400 233.0800 909.3400 233.5600 ;
        RECT 906.3400 222.2000 909.3400 222.6800 ;
        RECT 906.3400 227.6400 909.3400 228.1200 ;
        RECT 906.3400 216.7600 909.3400 217.2400 ;
        RECT 955.9000 200.4400 956.9000 200.9200 ;
        RECT 955.9000 205.8800 956.9000 206.3600 ;
        RECT 955.9000 211.3200 956.9000 211.8000 ;
        RECT 955.9000 184.1200 956.9000 184.6000 ;
        RECT 955.9000 189.5600 956.9000 190.0400 ;
        RECT 955.9000 195.0000 956.9000 195.4800 ;
        RECT 906.3400 211.3200 909.3400 211.8000 ;
        RECT 906.3400 200.4400 909.3400 200.9200 ;
        RECT 906.3400 205.8800 909.3400 206.3600 ;
        RECT 906.3400 195.0000 909.3400 195.4800 ;
        RECT 906.3400 184.1200 909.3400 184.6000 ;
        RECT 906.3400 189.5600 909.3400 190.0400 ;
        RECT 1132.3400 173.2400 1135.3400 173.7200 ;
        RECT 1132.3400 178.6800 1135.3400 179.1600 ;
        RECT 1132.3400 167.8000 1135.3400 168.2800 ;
        RECT 1132.3400 162.3600 1135.3400 162.8400 ;
        RECT 1132.3400 156.9200 1135.3400 157.4000 ;
        RECT 1090.9000 173.2400 1091.9000 173.7200 ;
        RECT 1090.9000 178.6800 1091.9000 179.1600 ;
        RECT 1090.9000 156.9200 1091.9000 157.4000 ;
        RECT 1090.9000 162.3600 1091.9000 162.8400 ;
        RECT 1090.9000 167.8000 1091.9000 168.2800 ;
        RECT 1132.3400 140.6000 1135.3400 141.0800 ;
        RECT 1132.3400 146.0400 1135.3400 146.5200 ;
        RECT 1132.3400 151.4800 1135.3400 151.9600 ;
        RECT 1132.3400 135.1600 1135.3400 135.6400 ;
        RECT 1132.3400 124.2800 1135.3400 124.7600 ;
        RECT 1132.3400 129.7200 1135.3400 130.2000 ;
        RECT 1090.9000 140.6000 1091.9000 141.0800 ;
        RECT 1090.9000 146.0400 1091.9000 146.5200 ;
        RECT 1090.9000 151.4800 1091.9000 151.9600 ;
        RECT 1090.9000 124.2800 1091.9000 124.7600 ;
        RECT 1090.9000 129.7200 1091.9000 130.2000 ;
        RECT 1090.9000 135.1600 1091.9000 135.6400 ;
        RECT 1045.9000 173.2400 1046.9000 173.7200 ;
        RECT 1045.9000 178.6800 1046.9000 179.1600 ;
        RECT 1045.9000 156.9200 1046.9000 157.4000 ;
        RECT 1045.9000 162.3600 1046.9000 162.8400 ;
        RECT 1045.9000 167.8000 1046.9000 168.2800 ;
        RECT 1045.9000 140.6000 1046.9000 141.0800 ;
        RECT 1045.9000 146.0400 1046.9000 146.5200 ;
        RECT 1045.9000 151.4800 1046.9000 151.9600 ;
        RECT 1045.9000 124.2800 1046.9000 124.7600 ;
        RECT 1045.9000 129.7200 1046.9000 130.2000 ;
        RECT 1045.9000 135.1600 1046.9000 135.6400 ;
        RECT 1132.3400 113.4000 1135.3400 113.8800 ;
        RECT 1132.3400 118.8400 1135.3400 119.3200 ;
        RECT 1132.3400 107.9600 1135.3400 108.4400 ;
        RECT 1132.3400 102.5200 1135.3400 103.0000 ;
        RECT 1132.3400 97.0800 1135.3400 97.5600 ;
        RECT 1090.9000 113.4000 1091.9000 113.8800 ;
        RECT 1090.9000 118.8400 1091.9000 119.3200 ;
        RECT 1090.9000 97.0800 1091.9000 97.5600 ;
        RECT 1090.9000 102.5200 1091.9000 103.0000 ;
        RECT 1090.9000 107.9600 1091.9000 108.4400 ;
        RECT 1132.3400 86.2000 1135.3400 86.6800 ;
        RECT 1132.3400 91.6400 1135.3400 92.1200 ;
        RECT 1090.9000 86.2000 1091.9000 86.6800 ;
        RECT 1090.9000 91.6400 1091.9000 92.1200 ;
        RECT 1045.9000 113.4000 1046.9000 113.8800 ;
        RECT 1045.9000 118.8400 1046.9000 119.3200 ;
        RECT 1045.9000 97.0800 1046.9000 97.5600 ;
        RECT 1045.9000 102.5200 1046.9000 103.0000 ;
        RECT 1045.9000 107.9600 1046.9000 108.4400 ;
        RECT 1045.9000 86.2000 1046.9000 86.6800 ;
        RECT 1045.9000 91.6400 1046.9000 92.1200 ;
        RECT 1000.9000 173.2400 1001.9000 173.7200 ;
        RECT 1000.9000 178.6800 1001.9000 179.1600 ;
        RECT 1000.9000 156.9200 1001.9000 157.4000 ;
        RECT 1000.9000 162.3600 1001.9000 162.8400 ;
        RECT 1000.9000 167.8000 1001.9000 168.2800 ;
        RECT 1000.9000 140.6000 1001.9000 141.0800 ;
        RECT 1000.9000 146.0400 1001.9000 146.5200 ;
        RECT 1000.9000 151.4800 1001.9000 151.9600 ;
        RECT 1000.9000 124.2800 1001.9000 124.7600 ;
        RECT 1000.9000 129.7200 1001.9000 130.2000 ;
        RECT 1000.9000 135.1600 1001.9000 135.6400 ;
        RECT 955.9000 173.2400 956.9000 173.7200 ;
        RECT 955.9000 178.6800 956.9000 179.1600 ;
        RECT 955.9000 156.9200 956.9000 157.4000 ;
        RECT 955.9000 162.3600 956.9000 162.8400 ;
        RECT 955.9000 167.8000 956.9000 168.2800 ;
        RECT 906.3400 178.6800 909.3400 179.1600 ;
        RECT 906.3400 173.2400 909.3400 173.7200 ;
        RECT 906.3400 162.3600 909.3400 162.8400 ;
        RECT 906.3400 167.8000 909.3400 168.2800 ;
        RECT 906.3400 156.9200 909.3400 157.4000 ;
        RECT 955.9000 140.6000 956.9000 141.0800 ;
        RECT 955.9000 146.0400 956.9000 146.5200 ;
        RECT 955.9000 151.4800 956.9000 151.9600 ;
        RECT 955.9000 124.2800 956.9000 124.7600 ;
        RECT 955.9000 129.7200 956.9000 130.2000 ;
        RECT 955.9000 135.1600 956.9000 135.6400 ;
        RECT 906.3400 151.4800 909.3400 151.9600 ;
        RECT 906.3400 140.6000 909.3400 141.0800 ;
        RECT 906.3400 146.0400 909.3400 146.5200 ;
        RECT 906.3400 135.1600 909.3400 135.6400 ;
        RECT 906.3400 124.2800 909.3400 124.7600 ;
        RECT 906.3400 129.7200 909.3400 130.2000 ;
        RECT 1000.9000 113.4000 1001.9000 113.8800 ;
        RECT 1000.9000 118.8400 1001.9000 119.3200 ;
        RECT 1000.9000 97.0800 1001.9000 97.5600 ;
        RECT 1000.9000 102.5200 1001.9000 103.0000 ;
        RECT 1000.9000 107.9600 1001.9000 108.4400 ;
        RECT 1000.9000 86.2000 1001.9000 86.6800 ;
        RECT 1000.9000 91.6400 1001.9000 92.1200 ;
        RECT 955.9000 113.4000 956.9000 113.8800 ;
        RECT 955.9000 118.8400 956.9000 119.3200 ;
        RECT 955.9000 97.0800 956.9000 97.5600 ;
        RECT 955.9000 102.5200 956.9000 103.0000 ;
        RECT 955.9000 107.9600 956.9000 108.4400 ;
        RECT 906.3400 118.8400 909.3400 119.3200 ;
        RECT 906.3400 113.4000 909.3400 113.8800 ;
        RECT 906.3400 102.5200 909.3400 103.0000 ;
        RECT 906.3400 107.9600 909.3400 108.4400 ;
        RECT 906.3400 97.0800 909.3400 97.5600 ;
        RECT 955.9000 86.2000 956.9000 86.6800 ;
        RECT 955.9000 91.6400 956.9000 92.1200 ;
        RECT 906.3400 91.6400 909.3400 92.1200 ;
        RECT 906.3400 86.2000 909.3400 86.6800 ;
        RECT 906.3400 284.3900 1135.3400 287.3900 ;
        RECT 906.3400 79.2900 1135.3400 82.2900 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'S_term_single2'
    PORT
      LAYER met4 ;
        RECT 906.3400 37.6700 908.3400 58.6000 ;
        RECT 1133.3400 37.6700 1135.3400 58.6000 ;
      LAYER met3 ;
        RECT 1133.3400 54.1000 1135.3400 54.5800 ;
        RECT 906.3400 54.1000 908.3400 54.5800 ;
        RECT 1133.3400 43.2200 1135.3400 43.7000 ;
        RECT 906.3400 43.2200 908.3400 43.7000 ;
        RECT 1133.3400 48.6600 1135.3400 49.1400 ;
        RECT 906.3400 48.6600 908.3400 49.1400 ;
        RECT 906.3400 56.6000 1135.3400 58.6000 ;
        RECT 906.3400 37.6700 1135.3400 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single2'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 2605.3300 1091.9000 2813.4300 ;
        RECT 1045.9000 2605.3300 1046.9000 2813.4300 ;
        RECT 1000.9000 2605.3300 1001.9000 2813.4300 ;
        RECT 955.9000 2605.3300 956.9000 2813.4300 ;
        RECT 1132.3400 2605.3300 1135.3400 2813.4300 ;
        RECT 906.3400 2605.3300 909.3400 2813.4300 ;
      LAYER met3 ;
        RECT 1132.3400 2802.6400 1135.3400 2803.1200 ;
        RECT 1132.3400 2808.0800 1135.3400 2808.5600 ;
        RECT 1090.9000 2802.6400 1091.9000 2803.1200 ;
        RECT 1090.9000 2808.0800 1091.9000 2808.5600 ;
        RECT 1132.3400 2786.3200 1135.3400 2786.8000 ;
        RECT 1132.3400 2791.7600 1135.3400 2792.2400 ;
        RECT 1132.3400 2797.2000 1135.3400 2797.6800 ;
        RECT 1132.3400 2780.8800 1135.3400 2781.3600 ;
        RECT 1132.3400 2770.0000 1135.3400 2770.4800 ;
        RECT 1132.3400 2775.4400 1135.3400 2775.9200 ;
        RECT 1090.9000 2786.3200 1091.9000 2786.8000 ;
        RECT 1090.9000 2791.7600 1091.9000 2792.2400 ;
        RECT 1090.9000 2797.2000 1091.9000 2797.6800 ;
        RECT 1090.9000 2770.0000 1091.9000 2770.4800 ;
        RECT 1090.9000 2775.4400 1091.9000 2775.9200 ;
        RECT 1090.9000 2780.8800 1091.9000 2781.3600 ;
        RECT 1045.9000 2802.6400 1046.9000 2803.1200 ;
        RECT 1045.9000 2808.0800 1046.9000 2808.5600 ;
        RECT 1045.9000 2786.3200 1046.9000 2786.8000 ;
        RECT 1045.9000 2791.7600 1046.9000 2792.2400 ;
        RECT 1045.9000 2797.2000 1046.9000 2797.6800 ;
        RECT 1045.9000 2770.0000 1046.9000 2770.4800 ;
        RECT 1045.9000 2775.4400 1046.9000 2775.9200 ;
        RECT 1045.9000 2780.8800 1046.9000 2781.3600 ;
        RECT 1132.3400 2759.1200 1135.3400 2759.6000 ;
        RECT 1132.3400 2764.5600 1135.3400 2765.0400 ;
        RECT 1132.3400 2753.6800 1135.3400 2754.1600 ;
        RECT 1132.3400 2748.2400 1135.3400 2748.7200 ;
        RECT 1132.3400 2742.8000 1135.3400 2743.2800 ;
        RECT 1090.9000 2759.1200 1091.9000 2759.6000 ;
        RECT 1090.9000 2764.5600 1091.9000 2765.0400 ;
        RECT 1090.9000 2742.8000 1091.9000 2743.2800 ;
        RECT 1090.9000 2748.2400 1091.9000 2748.7200 ;
        RECT 1090.9000 2753.6800 1091.9000 2754.1600 ;
        RECT 1132.3400 2726.4800 1135.3400 2726.9600 ;
        RECT 1132.3400 2731.9200 1135.3400 2732.4000 ;
        RECT 1132.3400 2737.3600 1135.3400 2737.8400 ;
        RECT 1132.3400 2721.0400 1135.3400 2721.5200 ;
        RECT 1132.3400 2710.1600 1135.3400 2710.6400 ;
        RECT 1132.3400 2715.6000 1135.3400 2716.0800 ;
        RECT 1090.9000 2726.4800 1091.9000 2726.9600 ;
        RECT 1090.9000 2731.9200 1091.9000 2732.4000 ;
        RECT 1090.9000 2737.3600 1091.9000 2737.8400 ;
        RECT 1090.9000 2710.1600 1091.9000 2710.6400 ;
        RECT 1090.9000 2715.6000 1091.9000 2716.0800 ;
        RECT 1090.9000 2721.0400 1091.9000 2721.5200 ;
        RECT 1045.9000 2759.1200 1046.9000 2759.6000 ;
        RECT 1045.9000 2764.5600 1046.9000 2765.0400 ;
        RECT 1045.9000 2742.8000 1046.9000 2743.2800 ;
        RECT 1045.9000 2748.2400 1046.9000 2748.7200 ;
        RECT 1045.9000 2753.6800 1046.9000 2754.1600 ;
        RECT 1045.9000 2726.4800 1046.9000 2726.9600 ;
        RECT 1045.9000 2731.9200 1046.9000 2732.4000 ;
        RECT 1045.9000 2737.3600 1046.9000 2737.8400 ;
        RECT 1045.9000 2710.1600 1046.9000 2710.6400 ;
        RECT 1045.9000 2715.6000 1046.9000 2716.0800 ;
        RECT 1045.9000 2721.0400 1046.9000 2721.5200 ;
        RECT 1000.9000 2802.6400 1001.9000 2803.1200 ;
        RECT 1000.9000 2808.0800 1001.9000 2808.5600 ;
        RECT 1000.9000 2786.3200 1001.9000 2786.8000 ;
        RECT 1000.9000 2791.7600 1001.9000 2792.2400 ;
        RECT 1000.9000 2797.2000 1001.9000 2797.6800 ;
        RECT 1000.9000 2770.0000 1001.9000 2770.4800 ;
        RECT 1000.9000 2775.4400 1001.9000 2775.9200 ;
        RECT 1000.9000 2780.8800 1001.9000 2781.3600 ;
        RECT 955.9000 2802.6400 956.9000 2803.1200 ;
        RECT 955.9000 2808.0800 956.9000 2808.5600 ;
        RECT 906.3400 2808.0800 909.3400 2808.5600 ;
        RECT 906.3400 2802.6400 909.3400 2803.1200 ;
        RECT 955.9000 2786.3200 956.9000 2786.8000 ;
        RECT 955.9000 2791.7600 956.9000 2792.2400 ;
        RECT 955.9000 2797.2000 956.9000 2797.6800 ;
        RECT 955.9000 2770.0000 956.9000 2770.4800 ;
        RECT 955.9000 2775.4400 956.9000 2775.9200 ;
        RECT 955.9000 2780.8800 956.9000 2781.3600 ;
        RECT 906.3400 2797.2000 909.3400 2797.6800 ;
        RECT 906.3400 2786.3200 909.3400 2786.8000 ;
        RECT 906.3400 2791.7600 909.3400 2792.2400 ;
        RECT 906.3400 2780.8800 909.3400 2781.3600 ;
        RECT 906.3400 2770.0000 909.3400 2770.4800 ;
        RECT 906.3400 2775.4400 909.3400 2775.9200 ;
        RECT 1000.9000 2759.1200 1001.9000 2759.6000 ;
        RECT 1000.9000 2764.5600 1001.9000 2765.0400 ;
        RECT 1000.9000 2742.8000 1001.9000 2743.2800 ;
        RECT 1000.9000 2748.2400 1001.9000 2748.7200 ;
        RECT 1000.9000 2753.6800 1001.9000 2754.1600 ;
        RECT 1000.9000 2726.4800 1001.9000 2726.9600 ;
        RECT 1000.9000 2731.9200 1001.9000 2732.4000 ;
        RECT 1000.9000 2737.3600 1001.9000 2737.8400 ;
        RECT 1000.9000 2710.1600 1001.9000 2710.6400 ;
        RECT 1000.9000 2715.6000 1001.9000 2716.0800 ;
        RECT 1000.9000 2721.0400 1001.9000 2721.5200 ;
        RECT 955.9000 2759.1200 956.9000 2759.6000 ;
        RECT 955.9000 2764.5600 956.9000 2765.0400 ;
        RECT 955.9000 2742.8000 956.9000 2743.2800 ;
        RECT 955.9000 2748.2400 956.9000 2748.7200 ;
        RECT 955.9000 2753.6800 956.9000 2754.1600 ;
        RECT 906.3400 2764.5600 909.3400 2765.0400 ;
        RECT 906.3400 2759.1200 909.3400 2759.6000 ;
        RECT 906.3400 2748.2400 909.3400 2748.7200 ;
        RECT 906.3400 2753.6800 909.3400 2754.1600 ;
        RECT 906.3400 2742.8000 909.3400 2743.2800 ;
        RECT 955.9000 2726.4800 956.9000 2726.9600 ;
        RECT 955.9000 2731.9200 956.9000 2732.4000 ;
        RECT 955.9000 2737.3600 956.9000 2737.8400 ;
        RECT 955.9000 2710.1600 956.9000 2710.6400 ;
        RECT 955.9000 2715.6000 956.9000 2716.0800 ;
        RECT 955.9000 2721.0400 956.9000 2721.5200 ;
        RECT 906.3400 2737.3600 909.3400 2737.8400 ;
        RECT 906.3400 2726.4800 909.3400 2726.9600 ;
        RECT 906.3400 2731.9200 909.3400 2732.4000 ;
        RECT 906.3400 2721.0400 909.3400 2721.5200 ;
        RECT 906.3400 2710.1600 909.3400 2710.6400 ;
        RECT 906.3400 2715.6000 909.3400 2716.0800 ;
        RECT 1132.3400 2699.2800 1135.3400 2699.7600 ;
        RECT 1132.3400 2704.7200 1135.3400 2705.2000 ;
        RECT 1132.3400 2693.8400 1135.3400 2694.3200 ;
        RECT 1132.3400 2688.4000 1135.3400 2688.8800 ;
        RECT 1132.3400 2682.9600 1135.3400 2683.4400 ;
        RECT 1090.9000 2699.2800 1091.9000 2699.7600 ;
        RECT 1090.9000 2704.7200 1091.9000 2705.2000 ;
        RECT 1090.9000 2682.9600 1091.9000 2683.4400 ;
        RECT 1090.9000 2688.4000 1091.9000 2688.8800 ;
        RECT 1090.9000 2693.8400 1091.9000 2694.3200 ;
        RECT 1132.3400 2666.6400 1135.3400 2667.1200 ;
        RECT 1132.3400 2672.0800 1135.3400 2672.5600 ;
        RECT 1132.3400 2677.5200 1135.3400 2678.0000 ;
        RECT 1132.3400 2661.2000 1135.3400 2661.6800 ;
        RECT 1132.3400 2650.3200 1135.3400 2650.8000 ;
        RECT 1132.3400 2655.7600 1135.3400 2656.2400 ;
        RECT 1090.9000 2666.6400 1091.9000 2667.1200 ;
        RECT 1090.9000 2672.0800 1091.9000 2672.5600 ;
        RECT 1090.9000 2677.5200 1091.9000 2678.0000 ;
        RECT 1090.9000 2650.3200 1091.9000 2650.8000 ;
        RECT 1090.9000 2655.7600 1091.9000 2656.2400 ;
        RECT 1090.9000 2661.2000 1091.9000 2661.6800 ;
        RECT 1045.9000 2699.2800 1046.9000 2699.7600 ;
        RECT 1045.9000 2704.7200 1046.9000 2705.2000 ;
        RECT 1045.9000 2682.9600 1046.9000 2683.4400 ;
        RECT 1045.9000 2688.4000 1046.9000 2688.8800 ;
        RECT 1045.9000 2693.8400 1046.9000 2694.3200 ;
        RECT 1045.9000 2666.6400 1046.9000 2667.1200 ;
        RECT 1045.9000 2672.0800 1046.9000 2672.5600 ;
        RECT 1045.9000 2677.5200 1046.9000 2678.0000 ;
        RECT 1045.9000 2650.3200 1046.9000 2650.8000 ;
        RECT 1045.9000 2655.7600 1046.9000 2656.2400 ;
        RECT 1045.9000 2661.2000 1046.9000 2661.6800 ;
        RECT 1132.3400 2639.4400 1135.3400 2639.9200 ;
        RECT 1132.3400 2644.8800 1135.3400 2645.3600 ;
        RECT 1132.3400 2634.0000 1135.3400 2634.4800 ;
        RECT 1132.3400 2628.5600 1135.3400 2629.0400 ;
        RECT 1132.3400 2623.1200 1135.3400 2623.6000 ;
        RECT 1090.9000 2639.4400 1091.9000 2639.9200 ;
        RECT 1090.9000 2644.8800 1091.9000 2645.3600 ;
        RECT 1090.9000 2623.1200 1091.9000 2623.6000 ;
        RECT 1090.9000 2628.5600 1091.9000 2629.0400 ;
        RECT 1090.9000 2634.0000 1091.9000 2634.4800 ;
        RECT 1132.3400 2612.2400 1135.3400 2612.7200 ;
        RECT 1132.3400 2617.6800 1135.3400 2618.1600 ;
        RECT 1090.9000 2612.2400 1091.9000 2612.7200 ;
        RECT 1090.9000 2617.6800 1091.9000 2618.1600 ;
        RECT 1045.9000 2639.4400 1046.9000 2639.9200 ;
        RECT 1045.9000 2644.8800 1046.9000 2645.3600 ;
        RECT 1045.9000 2623.1200 1046.9000 2623.6000 ;
        RECT 1045.9000 2628.5600 1046.9000 2629.0400 ;
        RECT 1045.9000 2634.0000 1046.9000 2634.4800 ;
        RECT 1045.9000 2612.2400 1046.9000 2612.7200 ;
        RECT 1045.9000 2617.6800 1046.9000 2618.1600 ;
        RECT 1000.9000 2699.2800 1001.9000 2699.7600 ;
        RECT 1000.9000 2704.7200 1001.9000 2705.2000 ;
        RECT 1000.9000 2682.9600 1001.9000 2683.4400 ;
        RECT 1000.9000 2688.4000 1001.9000 2688.8800 ;
        RECT 1000.9000 2693.8400 1001.9000 2694.3200 ;
        RECT 1000.9000 2666.6400 1001.9000 2667.1200 ;
        RECT 1000.9000 2672.0800 1001.9000 2672.5600 ;
        RECT 1000.9000 2677.5200 1001.9000 2678.0000 ;
        RECT 1000.9000 2650.3200 1001.9000 2650.8000 ;
        RECT 1000.9000 2655.7600 1001.9000 2656.2400 ;
        RECT 1000.9000 2661.2000 1001.9000 2661.6800 ;
        RECT 955.9000 2699.2800 956.9000 2699.7600 ;
        RECT 955.9000 2704.7200 956.9000 2705.2000 ;
        RECT 955.9000 2682.9600 956.9000 2683.4400 ;
        RECT 955.9000 2688.4000 956.9000 2688.8800 ;
        RECT 955.9000 2693.8400 956.9000 2694.3200 ;
        RECT 906.3400 2704.7200 909.3400 2705.2000 ;
        RECT 906.3400 2699.2800 909.3400 2699.7600 ;
        RECT 906.3400 2688.4000 909.3400 2688.8800 ;
        RECT 906.3400 2693.8400 909.3400 2694.3200 ;
        RECT 906.3400 2682.9600 909.3400 2683.4400 ;
        RECT 955.9000 2666.6400 956.9000 2667.1200 ;
        RECT 955.9000 2672.0800 956.9000 2672.5600 ;
        RECT 955.9000 2677.5200 956.9000 2678.0000 ;
        RECT 955.9000 2650.3200 956.9000 2650.8000 ;
        RECT 955.9000 2655.7600 956.9000 2656.2400 ;
        RECT 955.9000 2661.2000 956.9000 2661.6800 ;
        RECT 906.3400 2677.5200 909.3400 2678.0000 ;
        RECT 906.3400 2666.6400 909.3400 2667.1200 ;
        RECT 906.3400 2672.0800 909.3400 2672.5600 ;
        RECT 906.3400 2661.2000 909.3400 2661.6800 ;
        RECT 906.3400 2650.3200 909.3400 2650.8000 ;
        RECT 906.3400 2655.7600 909.3400 2656.2400 ;
        RECT 1000.9000 2639.4400 1001.9000 2639.9200 ;
        RECT 1000.9000 2644.8800 1001.9000 2645.3600 ;
        RECT 1000.9000 2623.1200 1001.9000 2623.6000 ;
        RECT 1000.9000 2628.5600 1001.9000 2629.0400 ;
        RECT 1000.9000 2634.0000 1001.9000 2634.4800 ;
        RECT 1000.9000 2612.2400 1001.9000 2612.7200 ;
        RECT 1000.9000 2617.6800 1001.9000 2618.1600 ;
        RECT 955.9000 2639.4400 956.9000 2639.9200 ;
        RECT 955.9000 2644.8800 956.9000 2645.3600 ;
        RECT 955.9000 2623.1200 956.9000 2623.6000 ;
        RECT 955.9000 2628.5600 956.9000 2629.0400 ;
        RECT 955.9000 2634.0000 956.9000 2634.4800 ;
        RECT 906.3400 2644.8800 909.3400 2645.3600 ;
        RECT 906.3400 2639.4400 909.3400 2639.9200 ;
        RECT 906.3400 2628.5600 909.3400 2629.0400 ;
        RECT 906.3400 2634.0000 909.3400 2634.4800 ;
        RECT 906.3400 2623.1200 909.3400 2623.6000 ;
        RECT 955.9000 2612.2400 956.9000 2612.7200 ;
        RECT 955.9000 2617.6800 956.9000 2618.1600 ;
        RECT 906.3400 2617.6800 909.3400 2618.1600 ;
        RECT 906.3400 2612.2400 909.3400 2612.7200 ;
        RECT 906.3400 2810.4300 1135.3400 2813.4300 ;
        RECT 906.3400 2605.3300 1135.3400 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 2375.6900 1091.9000 2583.7900 ;
        RECT 1045.9000 2375.6900 1046.9000 2583.7900 ;
        RECT 1000.9000 2375.6900 1001.9000 2583.7900 ;
        RECT 955.9000 2375.6900 956.9000 2583.7900 ;
        RECT 1132.3400 2375.6900 1135.3400 2583.7900 ;
        RECT 906.3400 2375.6900 909.3400 2583.7900 ;
      LAYER met3 ;
        RECT 1132.3400 2573.0000 1135.3400 2573.4800 ;
        RECT 1132.3400 2578.4400 1135.3400 2578.9200 ;
        RECT 1090.9000 2573.0000 1091.9000 2573.4800 ;
        RECT 1090.9000 2578.4400 1091.9000 2578.9200 ;
        RECT 1132.3400 2556.6800 1135.3400 2557.1600 ;
        RECT 1132.3400 2562.1200 1135.3400 2562.6000 ;
        RECT 1132.3400 2567.5600 1135.3400 2568.0400 ;
        RECT 1132.3400 2551.2400 1135.3400 2551.7200 ;
        RECT 1132.3400 2540.3600 1135.3400 2540.8400 ;
        RECT 1132.3400 2545.8000 1135.3400 2546.2800 ;
        RECT 1090.9000 2556.6800 1091.9000 2557.1600 ;
        RECT 1090.9000 2562.1200 1091.9000 2562.6000 ;
        RECT 1090.9000 2567.5600 1091.9000 2568.0400 ;
        RECT 1090.9000 2540.3600 1091.9000 2540.8400 ;
        RECT 1090.9000 2545.8000 1091.9000 2546.2800 ;
        RECT 1090.9000 2551.2400 1091.9000 2551.7200 ;
        RECT 1045.9000 2573.0000 1046.9000 2573.4800 ;
        RECT 1045.9000 2578.4400 1046.9000 2578.9200 ;
        RECT 1045.9000 2556.6800 1046.9000 2557.1600 ;
        RECT 1045.9000 2562.1200 1046.9000 2562.6000 ;
        RECT 1045.9000 2567.5600 1046.9000 2568.0400 ;
        RECT 1045.9000 2540.3600 1046.9000 2540.8400 ;
        RECT 1045.9000 2545.8000 1046.9000 2546.2800 ;
        RECT 1045.9000 2551.2400 1046.9000 2551.7200 ;
        RECT 1132.3400 2529.4800 1135.3400 2529.9600 ;
        RECT 1132.3400 2534.9200 1135.3400 2535.4000 ;
        RECT 1132.3400 2524.0400 1135.3400 2524.5200 ;
        RECT 1132.3400 2518.6000 1135.3400 2519.0800 ;
        RECT 1132.3400 2513.1600 1135.3400 2513.6400 ;
        RECT 1090.9000 2529.4800 1091.9000 2529.9600 ;
        RECT 1090.9000 2534.9200 1091.9000 2535.4000 ;
        RECT 1090.9000 2513.1600 1091.9000 2513.6400 ;
        RECT 1090.9000 2518.6000 1091.9000 2519.0800 ;
        RECT 1090.9000 2524.0400 1091.9000 2524.5200 ;
        RECT 1132.3400 2496.8400 1135.3400 2497.3200 ;
        RECT 1132.3400 2502.2800 1135.3400 2502.7600 ;
        RECT 1132.3400 2507.7200 1135.3400 2508.2000 ;
        RECT 1132.3400 2491.4000 1135.3400 2491.8800 ;
        RECT 1132.3400 2480.5200 1135.3400 2481.0000 ;
        RECT 1132.3400 2485.9600 1135.3400 2486.4400 ;
        RECT 1090.9000 2496.8400 1091.9000 2497.3200 ;
        RECT 1090.9000 2502.2800 1091.9000 2502.7600 ;
        RECT 1090.9000 2507.7200 1091.9000 2508.2000 ;
        RECT 1090.9000 2480.5200 1091.9000 2481.0000 ;
        RECT 1090.9000 2485.9600 1091.9000 2486.4400 ;
        RECT 1090.9000 2491.4000 1091.9000 2491.8800 ;
        RECT 1045.9000 2529.4800 1046.9000 2529.9600 ;
        RECT 1045.9000 2534.9200 1046.9000 2535.4000 ;
        RECT 1045.9000 2513.1600 1046.9000 2513.6400 ;
        RECT 1045.9000 2518.6000 1046.9000 2519.0800 ;
        RECT 1045.9000 2524.0400 1046.9000 2524.5200 ;
        RECT 1045.9000 2496.8400 1046.9000 2497.3200 ;
        RECT 1045.9000 2502.2800 1046.9000 2502.7600 ;
        RECT 1045.9000 2507.7200 1046.9000 2508.2000 ;
        RECT 1045.9000 2480.5200 1046.9000 2481.0000 ;
        RECT 1045.9000 2485.9600 1046.9000 2486.4400 ;
        RECT 1045.9000 2491.4000 1046.9000 2491.8800 ;
        RECT 1000.9000 2573.0000 1001.9000 2573.4800 ;
        RECT 1000.9000 2578.4400 1001.9000 2578.9200 ;
        RECT 1000.9000 2556.6800 1001.9000 2557.1600 ;
        RECT 1000.9000 2562.1200 1001.9000 2562.6000 ;
        RECT 1000.9000 2567.5600 1001.9000 2568.0400 ;
        RECT 1000.9000 2540.3600 1001.9000 2540.8400 ;
        RECT 1000.9000 2545.8000 1001.9000 2546.2800 ;
        RECT 1000.9000 2551.2400 1001.9000 2551.7200 ;
        RECT 955.9000 2573.0000 956.9000 2573.4800 ;
        RECT 955.9000 2578.4400 956.9000 2578.9200 ;
        RECT 906.3400 2578.4400 909.3400 2578.9200 ;
        RECT 906.3400 2573.0000 909.3400 2573.4800 ;
        RECT 955.9000 2556.6800 956.9000 2557.1600 ;
        RECT 955.9000 2562.1200 956.9000 2562.6000 ;
        RECT 955.9000 2567.5600 956.9000 2568.0400 ;
        RECT 955.9000 2540.3600 956.9000 2540.8400 ;
        RECT 955.9000 2545.8000 956.9000 2546.2800 ;
        RECT 955.9000 2551.2400 956.9000 2551.7200 ;
        RECT 906.3400 2567.5600 909.3400 2568.0400 ;
        RECT 906.3400 2556.6800 909.3400 2557.1600 ;
        RECT 906.3400 2562.1200 909.3400 2562.6000 ;
        RECT 906.3400 2551.2400 909.3400 2551.7200 ;
        RECT 906.3400 2540.3600 909.3400 2540.8400 ;
        RECT 906.3400 2545.8000 909.3400 2546.2800 ;
        RECT 1000.9000 2529.4800 1001.9000 2529.9600 ;
        RECT 1000.9000 2534.9200 1001.9000 2535.4000 ;
        RECT 1000.9000 2513.1600 1001.9000 2513.6400 ;
        RECT 1000.9000 2518.6000 1001.9000 2519.0800 ;
        RECT 1000.9000 2524.0400 1001.9000 2524.5200 ;
        RECT 1000.9000 2496.8400 1001.9000 2497.3200 ;
        RECT 1000.9000 2502.2800 1001.9000 2502.7600 ;
        RECT 1000.9000 2507.7200 1001.9000 2508.2000 ;
        RECT 1000.9000 2480.5200 1001.9000 2481.0000 ;
        RECT 1000.9000 2485.9600 1001.9000 2486.4400 ;
        RECT 1000.9000 2491.4000 1001.9000 2491.8800 ;
        RECT 955.9000 2529.4800 956.9000 2529.9600 ;
        RECT 955.9000 2534.9200 956.9000 2535.4000 ;
        RECT 955.9000 2513.1600 956.9000 2513.6400 ;
        RECT 955.9000 2518.6000 956.9000 2519.0800 ;
        RECT 955.9000 2524.0400 956.9000 2524.5200 ;
        RECT 906.3400 2534.9200 909.3400 2535.4000 ;
        RECT 906.3400 2529.4800 909.3400 2529.9600 ;
        RECT 906.3400 2518.6000 909.3400 2519.0800 ;
        RECT 906.3400 2524.0400 909.3400 2524.5200 ;
        RECT 906.3400 2513.1600 909.3400 2513.6400 ;
        RECT 955.9000 2496.8400 956.9000 2497.3200 ;
        RECT 955.9000 2502.2800 956.9000 2502.7600 ;
        RECT 955.9000 2507.7200 956.9000 2508.2000 ;
        RECT 955.9000 2480.5200 956.9000 2481.0000 ;
        RECT 955.9000 2485.9600 956.9000 2486.4400 ;
        RECT 955.9000 2491.4000 956.9000 2491.8800 ;
        RECT 906.3400 2507.7200 909.3400 2508.2000 ;
        RECT 906.3400 2496.8400 909.3400 2497.3200 ;
        RECT 906.3400 2502.2800 909.3400 2502.7600 ;
        RECT 906.3400 2491.4000 909.3400 2491.8800 ;
        RECT 906.3400 2480.5200 909.3400 2481.0000 ;
        RECT 906.3400 2485.9600 909.3400 2486.4400 ;
        RECT 1132.3400 2469.6400 1135.3400 2470.1200 ;
        RECT 1132.3400 2475.0800 1135.3400 2475.5600 ;
        RECT 1132.3400 2464.2000 1135.3400 2464.6800 ;
        RECT 1132.3400 2458.7600 1135.3400 2459.2400 ;
        RECT 1132.3400 2453.3200 1135.3400 2453.8000 ;
        RECT 1090.9000 2469.6400 1091.9000 2470.1200 ;
        RECT 1090.9000 2475.0800 1091.9000 2475.5600 ;
        RECT 1090.9000 2453.3200 1091.9000 2453.8000 ;
        RECT 1090.9000 2458.7600 1091.9000 2459.2400 ;
        RECT 1090.9000 2464.2000 1091.9000 2464.6800 ;
        RECT 1132.3400 2437.0000 1135.3400 2437.4800 ;
        RECT 1132.3400 2442.4400 1135.3400 2442.9200 ;
        RECT 1132.3400 2447.8800 1135.3400 2448.3600 ;
        RECT 1132.3400 2431.5600 1135.3400 2432.0400 ;
        RECT 1132.3400 2420.6800 1135.3400 2421.1600 ;
        RECT 1132.3400 2426.1200 1135.3400 2426.6000 ;
        RECT 1090.9000 2437.0000 1091.9000 2437.4800 ;
        RECT 1090.9000 2442.4400 1091.9000 2442.9200 ;
        RECT 1090.9000 2447.8800 1091.9000 2448.3600 ;
        RECT 1090.9000 2420.6800 1091.9000 2421.1600 ;
        RECT 1090.9000 2426.1200 1091.9000 2426.6000 ;
        RECT 1090.9000 2431.5600 1091.9000 2432.0400 ;
        RECT 1045.9000 2469.6400 1046.9000 2470.1200 ;
        RECT 1045.9000 2475.0800 1046.9000 2475.5600 ;
        RECT 1045.9000 2453.3200 1046.9000 2453.8000 ;
        RECT 1045.9000 2458.7600 1046.9000 2459.2400 ;
        RECT 1045.9000 2464.2000 1046.9000 2464.6800 ;
        RECT 1045.9000 2437.0000 1046.9000 2437.4800 ;
        RECT 1045.9000 2442.4400 1046.9000 2442.9200 ;
        RECT 1045.9000 2447.8800 1046.9000 2448.3600 ;
        RECT 1045.9000 2420.6800 1046.9000 2421.1600 ;
        RECT 1045.9000 2426.1200 1046.9000 2426.6000 ;
        RECT 1045.9000 2431.5600 1046.9000 2432.0400 ;
        RECT 1132.3400 2409.8000 1135.3400 2410.2800 ;
        RECT 1132.3400 2415.2400 1135.3400 2415.7200 ;
        RECT 1132.3400 2404.3600 1135.3400 2404.8400 ;
        RECT 1132.3400 2398.9200 1135.3400 2399.4000 ;
        RECT 1132.3400 2393.4800 1135.3400 2393.9600 ;
        RECT 1090.9000 2409.8000 1091.9000 2410.2800 ;
        RECT 1090.9000 2415.2400 1091.9000 2415.7200 ;
        RECT 1090.9000 2393.4800 1091.9000 2393.9600 ;
        RECT 1090.9000 2398.9200 1091.9000 2399.4000 ;
        RECT 1090.9000 2404.3600 1091.9000 2404.8400 ;
        RECT 1132.3400 2382.6000 1135.3400 2383.0800 ;
        RECT 1132.3400 2388.0400 1135.3400 2388.5200 ;
        RECT 1090.9000 2382.6000 1091.9000 2383.0800 ;
        RECT 1090.9000 2388.0400 1091.9000 2388.5200 ;
        RECT 1045.9000 2409.8000 1046.9000 2410.2800 ;
        RECT 1045.9000 2415.2400 1046.9000 2415.7200 ;
        RECT 1045.9000 2393.4800 1046.9000 2393.9600 ;
        RECT 1045.9000 2398.9200 1046.9000 2399.4000 ;
        RECT 1045.9000 2404.3600 1046.9000 2404.8400 ;
        RECT 1045.9000 2382.6000 1046.9000 2383.0800 ;
        RECT 1045.9000 2388.0400 1046.9000 2388.5200 ;
        RECT 1000.9000 2469.6400 1001.9000 2470.1200 ;
        RECT 1000.9000 2475.0800 1001.9000 2475.5600 ;
        RECT 1000.9000 2453.3200 1001.9000 2453.8000 ;
        RECT 1000.9000 2458.7600 1001.9000 2459.2400 ;
        RECT 1000.9000 2464.2000 1001.9000 2464.6800 ;
        RECT 1000.9000 2437.0000 1001.9000 2437.4800 ;
        RECT 1000.9000 2442.4400 1001.9000 2442.9200 ;
        RECT 1000.9000 2447.8800 1001.9000 2448.3600 ;
        RECT 1000.9000 2420.6800 1001.9000 2421.1600 ;
        RECT 1000.9000 2426.1200 1001.9000 2426.6000 ;
        RECT 1000.9000 2431.5600 1001.9000 2432.0400 ;
        RECT 955.9000 2469.6400 956.9000 2470.1200 ;
        RECT 955.9000 2475.0800 956.9000 2475.5600 ;
        RECT 955.9000 2453.3200 956.9000 2453.8000 ;
        RECT 955.9000 2458.7600 956.9000 2459.2400 ;
        RECT 955.9000 2464.2000 956.9000 2464.6800 ;
        RECT 906.3400 2475.0800 909.3400 2475.5600 ;
        RECT 906.3400 2469.6400 909.3400 2470.1200 ;
        RECT 906.3400 2458.7600 909.3400 2459.2400 ;
        RECT 906.3400 2464.2000 909.3400 2464.6800 ;
        RECT 906.3400 2453.3200 909.3400 2453.8000 ;
        RECT 955.9000 2437.0000 956.9000 2437.4800 ;
        RECT 955.9000 2442.4400 956.9000 2442.9200 ;
        RECT 955.9000 2447.8800 956.9000 2448.3600 ;
        RECT 955.9000 2420.6800 956.9000 2421.1600 ;
        RECT 955.9000 2426.1200 956.9000 2426.6000 ;
        RECT 955.9000 2431.5600 956.9000 2432.0400 ;
        RECT 906.3400 2447.8800 909.3400 2448.3600 ;
        RECT 906.3400 2437.0000 909.3400 2437.4800 ;
        RECT 906.3400 2442.4400 909.3400 2442.9200 ;
        RECT 906.3400 2431.5600 909.3400 2432.0400 ;
        RECT 906.3400 2420.6800 909.3400 2421.1600 ;
        RECT 906.3400 2426.1200 909.3400 2426.6000 ;
        RECT 1000.9000 2409.8000 1001.9000 2410.2800 ;
        RECT 1000.9000 2415.2400 1001.9000 2415.7200 ;
        RECT 1000.9000 2393.4800 1001.9000 2393.9600 ;
        RECT 1000.9000 2398.9200 1001.9000 2399.4000 ;
        RECT 1000.9000 2404.3600 1001.9000 2404.8400 ;
        RECT 1000.9000 2382.6000 1001.9000 2383.0800 ;
        RECT 1000.9000 2388.0400 1001.9000 2388.5200 ;
        RECT 955.9000 2409.8000 956.9000 2410.2800 ;
        RECT 955.9000 2415.2400 956.9000 2415.7200 ;
        RECT 955.9000 2393.4800 956.9000 2393.9600 ;
        RECT 955.9000 2398.9200 956.9000 2399.4000 ;
        RECT 955.9000 2404.3600 956.9000 2404.8400 ;
        RECT 906.3400 2415.2400 909.3400 2415.7200 ;
        RECT 906.3400 2409.8000 909.3400 2410.2800 ;
        RECT 906.3400 2398.9200 909.3400 2399.4000 ;
        RECT 906.3400 2404.3600 909.3400 2404.8400 ;
        RECT 906.3400 2393.4800 909.3400 2393.9600 ;
        RECT 955.9000 2382.6000 956.9000 2383.0800 ;
        RECT 955.9000 2388.0400 956.9000 2388.5200 ;
        RECT 906.3400 2388.0400 909.3400 2388.5200 ;
        RECT 906.3400 2382.6000 909.3400 2383.0800 ;
        RECT 906.3400 2580.7900 1135.3400 2583.7900 ;
        RECT 906.3400 2375.6900 1135.3400 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 2146.0500 1091.9000 2354.1500 ;
        RECT 1045.9000 2146.0500 1046.9000 2354.1500 ;
        RECT 1000.9000 2146.0500 1001.9000 2354.1500 ;
        RECT 955.9000 2146.0500 956.9000 2354.1500 ;
        RECT 1132.3400 2146.0500 1135.3400 2354.1500 ;
        RECT 906.3400 2146.0500 909.3400 2354.1500 ;
      LAYER met3 ;
        RECT 1132.3400 2343.3600 1135.3400 2343.8400 ;
        RECT 1132.3400 2348.8000 1135.3400 2349.2800 ;
        RECT 1090.9000 2343.3600 1091.9000 2343.8400 ;
        RECT 1090.9000 2348.8000 1091.9000 2349.2800 ;
        RECT 1132.3400 2327.0400 1135.3400 2327.5200 ;
        RECT 1132.3400 2332.4800 1135.3400 2332.9600 ;
        RECT 1132.3400 2337.9200 1135.3400 2338.4000 ;
        RECT 1132.3400 2321.6000 1135.3400 2322.0800 ;
        RECT 1132.3400 2310.7200 1135.3400 2311.2000 ;
        RECT 1132.3400 2316.1600 1135.3400 2316.6400 ;
        RECT 1090.9000 2327.0400 1091.9000 2327.5200 ;
        RECT 1090.9000 2332.4800 1091.9000 2332.9600 ;
        RECT 1090.9000 2337.9200 1091.9000 2338.4000 ;
        RECT 1090.9000 2310.7200 1091.9000 2311.2000 ;
        RECT 1090.9000 2316.1600 1091.9000 2316.6400 ;
        RECT 1090.9000 2321.6000 1091.9000 2322.0800 ;
        RECT 1045.9000 2343.3600 1046.9000 2343.8400 ;
        RECT 1045.9000 2348.8000 1046.9000 2349.2800 ;
        RECT 1045.9000 2327.0400 1046.9000 2327.5200 ;
        RECT 1045.9000 2332.4800 1046.9000 2332.9600 ;
        RECT 1045.9000 2337.9200 1046.9000 2338.4000 ;
        RECT 1045.9000 2310.7200 1046.9000 2311.2000 ;
        RECT 1045.9000 2316.1600 1046.9000 2316.6400 ;
        RECT 1045.9000 2321.6000 1046.9000 2322.0800 ;
        RECT 1132.3400 2299.8400 1135.3400 2300.3200 ;
        RECT 1132.3400 2305.2800 1135.3400 2305.7600 ;
        RECT 1132.3400 2294.4000 1135.3400 2294.8800 ;
        RECT 1132.3400 2288.9600 1135.3400 2289.4400 ;
        RECT 1132.3400 2283.5200 1135.3400 2284.0000 ;
        RECT 1090.9000 2299.8400 1091.9000 2300.3200 ;
        RECT 1090.9000 2305.2800 1091.9000 2305.7600 ;
        RECT 1090.9000 2283.5200 1091.9000 2284.0000 ;
        RECT 1090.9000 2288.9600 1091.9000 2289.4400 ;
        RECT 1090.9000 2294.4000 1091.9000 2294.8800 ;
        RECT 1132.3400 2267.2000 1135.3400 2267.6800 ;
        RECT 1132.3400 2272.6400 1135.3400 2273.1200 ;
        RECT 1132.3400 2278.0800 1135.3400 2278.5600 ;
        RECT 1132.3400 2261.7600 1135.3400 2262.2400 ;
        RECT 1132.3400 2250.8800 1135.3400 2251.3600 ;
        RECT 1132.3400 2256.3200 1135.3400 2256.8000 ;
        RECT 1090.9000 2267.2000 1091.9000 2267.6800 ;
        RECT 1090.9000 2272.6400 1091.9000 2273.1200 ;
        RECT 1090.9000 2278.0800 1091.9000 2278.5600 ;
        RECT 1090.9000 2250.8800 1091.9000 2251.3600 ;
        RECT 1090.9000 2256.3200 1091.9000 2256.8000 ;
        RECT 1090.9000 2261.7600 1091.9000 2262.2400 ;
        RECT 1045.9000 2299.8400 1046.9000 2300.3200 ;
        RECT 1045.9000 2305.2800 1046.9000 2305.7600 ;
        RECT 1045.9000 2283.5200 1046.9000 2284.0000 ;
        RECT 1045.9000 2288.9600 1046.9000 2289.4400 ;
        RECT 1045.9000 2294.4000 1046.9000 2294.8800 ;
        RECT 1045.9000 2267.2000 1046.9000 2267.6800 ;
        RECT 1045.9000 2272.6400 1046.9000 2273.1200 ;
        RECT 1045.9000 2278.0800 1046.9000 2278.5600 ;
        RECT 1045.9000 2250.8800 1046.9000 2251.3600 ;
        RECT 1045.9000 2256.3200 1046.9000 2256.8000 ;
        RECT 1045.9000 2261.7600 1046.9000 2262.2400 ;
        RECT 1000.9000 2343.3600 1001.9000 2343.8400 ;
        RECT 1000.9000 2348.8000 1001.9000 2349.2800 ;
        RECT 1000.9000 2327.0400 1001.9000 2327.5200 ;
        RECT 1000.9000 2332.4800 1001.9000 2332.9600 ;
        RECT 1000.9000 2337.9200 1001.9000 2338.4000 ;
        RECT 1000.9000 2310.7200 1001.9000 2311.2000 ;
        RECT 1000.9000 2316.1600 1001.9000 2316.6400 ;
        RECT 1000.9000 2321.6000 1001.9000 2322.0800 ;
        RECT 955.9000 2343.3600 956.9000 2343.8400 ;
        RECT 955.9000 2348.8000 956.9000 2349.2800 ;
        RECT 906.3400 2348.8000 909.3400 2349.2800 ;
        RECT 906.3400 2343.3600 909.3400 2343.8400 ;
        RECT 955.9000 2327.0400 956.9000 2327.5200 ;
        RECT 955.9000 2332.4800 956.9000 2332.9600 ;
        RECT 955.9000 2337.9200 956.9000 2338.4000 ;
        RECT 955.9000 2310.7200 956.9000 2311.2000 ;
        RECT 955.9000 2316.1600 956.9000 2316.6400 ;
        RECT 955.9000 2321.6000 956.9000 2322.0800 ;
        RECT 906.3400 2337.9200 909.3400 2338.4000 ;
        RECT 906.3400 2327.0400 909.3400 2327.5200 ;
        RECT 906.3400 2332.4800 909.3400 2332.9600 ;
        RECT 906.3400 2321.6000 909.3400 2322.0800 ;
        RECT 906.3400 2310.7200 909.3400 2311.2000 ;
        RECT 906.3400 2316.1600 909.3400 2316.6400 ;
        RECT 1000.9000 2299.8400 1001.9000 2300.3200 ;
        RECT 1000.9000 2305.2800 1001.9000 2305.7600 ;
        RECT 1000.9000 2283.5200 1001.9000 2284.0000 ;
        RECT 1000.9000 2288.9600 1001.9000 2289.4400 ;
        RECT 1000.9000 2294.4000 1001.9000 2294.8800 ;
        RECT 1000.9000 2267.2000 1001.9000 2267.6800 ;
        RECT 1000.9000 2272.6400 1001.9000 2273.1200 ;
        RECT 1000.9000 2278.0800 1001.9000 2278.5600 ;
        RECT 1000.9000 2250.8800 1001.9000 2251.3600 ;
        RECT 1000.9000 2256.3200 1001.9000 2256.8000 ;
        RECT 1000.9000 2261.7600 1001.9000 2262.2400 ;
        RECT 955.9000 2299.8400 956.9000 2300.3200 ;
        RECT 955.9000 2305.2800 956.9000 2305.7600 ;
        RECT 955.9000 2283.5200 956.9000 2284.0000 ;
        RECT 955.9000 2288.9600 956.9000 2289.4400 ;
        RECT 955.9000 2294.4000 956.9000 2294.8800 ;
        RECT 906.3400 2305.2800 909.3400 2305.7600 ;
        RECT 906.3400 2299.8400 909.3400 2300.3200 ;
        RECT 906.3400 2288.9600 909.3400 2289.4400 ;
        RECT 906.3400 2294.4000 909.3400 2294.8800 ;
        RECT 906.3400 2283.5200 909.3400 2284.0000 ;
        RECT 955.9000 2267.2000 956.9000 2267.6800 ;
        RECT 955.9000 2272.6400 956.9000 2273.1200 ;
        RECT 955.9000 2278.0800 956.9000 2278.5600 ;
        RECT 955.9000 2250.8800 956.9000 2251.3600 ;
        RECT 955.9000 2256.3200 956.9000 2256.8000 ;
        RECT 955.9000 2261.7600 956.9000 2262.2400 ;
        RECT 906.3400 2278.0800 909.3400 2278.5600 ;
        RECT 906.3400 2267.2000 909.3400 2267.6800 ;
        RECT 906.3400 2272.6400 909.3400 2273.1200 ;
        RECT 906.3400 2261.7600 909.3400 2262.2400 ;
        RECT 906.3400 2250.8800 909.3400 2251.3600 ;
        RECT 906.3400 2256.3200 909.3400 2256.8000 ;
        RECT 1132.3400 2240.0000 1135.3400 2240.4800 ;
        RECT 1132.3400 2245.4400 1135.3400 2245.9200 ;
        RECT 1132.3400 2234.5600 1135.3400 2235.0400 ;
        RECT 1132.3400 2229.1200 1135.3400 2229.6000 ;
        RECT 1132.3400 2223.6800 1135.3400 2224.1600 ;
        RECT 1090.9000 2240.0000 1091.9000 2240.4800 ;
        RECT 1090.9000 2245.4400 1091.9000 2245.9200 ;
        RECT 1090.9000 2223.6800 1091.9000 2224.1600 ;
        RECT 1090.9000 2229.1200 1091.9000 2229.6000 ;
        RECT 1090.9000 2234.5600 1091.9000 2235.0400 ;
        RECT 1132.3400 2207.3600 1135.3400 2207.8400 ;
        RECT 1132.3400 2212.8000 1135.3400 2213.2800 ;
        RECT 1132.3400 2218.2400 1135.3400 2218.7200 ;
        RECT 1132.3400 2201.9200 1135.3400 2202.4000 ;
        RECT 1132.3400 2191.0400 1135.3400 2191.5200 ;
        RECT 1132.3400 2196.4800 1135.3400 2196.9600 ;
        RECT 1090.9000 2207.3600 1091.9000 2207.8400 ;
        RECT 1090.9000 2212.8000 1091.9000 2213.2800 ;
        RECT 1090.9000 2218.2400 1091.9000 2218.7200 ;
        RECT 1090.9000 2191.0400 1091.9000 2191.5200 ;
        RECT 1090.9000 2196.4800 1091.9000 2196.9600 ;
        RECT 1090.9000 2201.9200 1091.9000 2202.4000 ;
        RECT 1045.9000 2240.0000 1046.9000 2240.4800 ;
        RECT 1045.9000 2245.4400 1046.9000 2245.9200 ;
        RECT 1045.9000 2223.6800 1046.9000 2224.1600 ;
        RECT 1045.9000 2229.1200 1046.9000 2229.6000 ;
        RECT 1045.9000 2234.5600 1046.9000 2235.0400 ;
        RECT 1045.9000 2207.3600 1046.9000 2207.8400 ;
        RECT 1045.9000 2212.8000 1046.9000 2213.2800 ;
        RECT 1045.9000 2218.2400 1046.9000 2218.7200 ;
        RECT 1045.9000 2191.0400 1046.9000 2191.5200 ;
        RECT 1045.9000 2196.4800 1046.9000 2196.9600 ;
        RECT 1045.9000 2201.9200 1046.9000 2202.4000 ;
        RECT 1132.3400 2180.1600 1135.3400 2180.6400 ;
        RECT 1132.3400 2185.6000 1135.3400 2186.0800 ;
        RECT 1132.3400 2174.7200 1135.3400 2175.2000 ;
        RECT 1132.3400 2169.2800 1135.3400 2169.7600 ;
        RECT 1132.3400 2163.8400 1135.3400 2164.3200 ;
        RECT 1090.9000 2180.1600 1091.9000 2180.6400 ;
        RECT 1090.9000 2185.6000 1091.9000 2186.0800 ;
        RECT 1090.9000 2163.8400 1091.9000 2164.3200 ;
        RECT 1090.9000 2169.2800 1091.9000 2169.7600 ;
        RECT 1090.9000 2174.7200 1091.9000 2175.2000 ;
        RECT 1132.3400 2152.9600 1135.3400 2153.4400 ;
        RECT 1132.3400 2158.4000 1135.3400 2158.8800 ;
        RECT 1090.9000 2152.9600 1091.9000 2153.4400 ;
        RECT 1090.9000 2158.4000 1091.9000 2158.8800 ;
        RECT 1045.9000 2180.1600 1046.9000 2180.6400 ;
        RECT 1045.9000 2185.6000 1046.9000 2186.0800 ;
        RECT 1045.9000 2163.8400 1046.9000 2164.3200 ;
        RECT 1045.9000 2169.2800 1046.9000 2169.7600 ;
        RECT 1045.9000 2174.7200 1046.9000 2175.2000 ;
        RECT 1045.9000 2152.9600 1046.9000 2153.4400 ;
        RECT 1045.9000 2158.4000 1046.9000 2158.8800 ;
        RECT 1000.9000 2240.0000 1001.9000 2240.4800 ;
        RECT 1000.9000 2245.4400 1001.9000 2245.9200 ;
        RECT 1000.9000 2223.6800 1001.9000 2224.1600 ;
        RECT 1000.9000 2229.1200 1001.9000 2229.6000 ;
        RECT 1000.9000 2234.5600 1001.9000 2235.0400 ;
        RECT 1000.9000 2207.3600 1001.9000 2207.8400 ;
        RECT 1000.9000 2212.8000 1001.9000 2213.2800 ;
        RECT 1000.9000 2218.2400 1001.9000 2218.7200 ;
        RECT 1000.9000 2191.0400 1001.9000 2191.5200 ;
        RECT 1000.9000 2196.4800 1001.9000 2196.9600 ;
        RECT 1000.9000 2201.9200 1001.9000 2202.4000 ;
        RECT 955.9000 2240.0000 956.9000 2240.4800 ;
        RECT 955.9000 2245.4400 956.9000 2245.9200 ;
        RECT 955.9000 2223.6800 956.9000 2224.1600 ;
        RECT 955.9000 2229.1200 956.9000 2229.6000 ;
        RECT 955.9000 2234.5600 956.9000 2235.0400 ;
        RECT 906.3400 2245.4400 909.3400 2245.9200 ;
        RECT 906.3400 2240.0000 909.3400 2240.4800 ;
        RECT 906.3400 2229.1200 909.3400 2229.6000 ;
        RECT 906.3400 2234.5600 909.3400 2235.0400 ;
        RECT 906.3400 2223.6800 909.3400 2224.1600 ;
        RECT 955.9000 2207.3600 956.9000 2207.8400 ;
        RECT 955.9000 2212.8000 956.9000 2213.2800 ;
        RECT 955.9000 2218.2400 956.9000 2218.7200 ;
        RECT 955.9000 2191.0400 956.9000 2191.5200 ;
        RECT 955.9000 2196.4800 956.9000 2196.9600 ;
        RECT 955.9000 2201.9200 956.9000 2202.4000 ;
        RECT 906.3400 2218.2400 909.3400 2218.7200 ;
        RECT 906.3400 2207.3600 909.3400 2207.8400 ;
        RECT 906.3400 2212.8000 909.3400 2213.2800 ;
        RECT 906.3400 2201.9200 909.3400 2202.4000 ;
        RECT 906.3400 2191.0400 909.3400 2191.5200 ;
        RECT 906.3400 2196.4800 909.3400 2196.9600 ;
        RECT 1000.9000 2180.1600 1001.9000 2180.6400 ;
        RECT 1000.9000 2185.6000 1001.9000 2186.0800 ;
        RECT 1000.9000 2163.8400 1001.9000 2164.3200 ;
        RECT 1000.9000 2169.2800 1001.9000 2169.7600 ;
        RECT 1000.9000 2174.7200 1001.9000 2175.2000 ;
        RECT 1000.9000 2152.9600 1001.9000 2153.4400 ;
        RECT 1000.9000 2158.4000 1001.9000 2158.8800 ;
        RECT 955.9000 2180.1600 956.9000 2180.6400 ;
        RECT 955.9000 2185.6000 956.9000 2186.0800 ;
        RECT 955.9000 2163.8400 956.9000 2164.3200 ;
        RECT 955.9000 2169.2800 956.9000 2169.7600 ;
        RECT 955.9000 2174.7200 956.9000 2175.2000 ;
        RECT 906.3400 2185.6000 909.3400 2186.0800 ;
        RECT 906.3400 2180.1600 909.3400 2180.6400 ;
        RECT 906.3400 2169.2800 909.3400 2169.7600 ;
        RECT 906.3400 2174.7200 909.3400 2175.2000 ;
        RECT 906.3400 2163.8400 909.3400 2164.3200 ;
        RECT 955.9000 2152.9600 956.9000 2153.4400 ;
        RECT 955.9000 2158.4000 956.9000 2158.8800 ;
        RECT 906.3400 2158.4000 909.3400 2158.8800 ;
        RECT 906.3400 2152.9600 909.3400 2153.4400 ;
        RECT 906.3400 2351.1500 1135.3400 2354.1500 ;
        RECT 906.3400 2146.0500 1135.3400 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 1916.4100 1091.9000 2124.5100 ;
        RECT 1045.9000 1916.4100 1046.9000 2124.5100 ;
        RECT 1000.9000 1916.4100 1001.9000 2124.5100 ;
        RECT 955.9000 1916.4100 956.9000 2124.5100 ;
        RECT 1132.3400 1916.4100 1135.3400 2124.5100 ;
        RECT 906.3400 1916.4100 909.3400 2124.5100 ;
      LAYER met3 ;
        RECT 1132.3400 2113.7200 1135.3400 2114.2000 ;
        RECT 1132.3400 2119.1600 1135.3400 2119.6400 ;
        RECT 1090.9000 2113.7200 1091.9000 2114.2000 ;
        RECT 1090.9000 2119.1600 1091.9000 2119.6400 ;
        RECT 1132.3400 2097.4000 1135.3400 2097.8800 ;
        RECT 1132.3400 2102.8400 1135.3400 2103.3200 ;
        RECT 1132.3400 2108.2800 1135.3400 2108.7600 ;
        RECT 1132.3400 2091.9600 1135.3400 2092.4400 ;
        RECT 1132.3400 2081.0800 1135.3400 2081.5600 ;
        RECT 1132.3400 2086.5200 1135.3400 2087.0000 ;
        RECT 1090.9000 2097.4000 1091.9000 2097.8800 ;
        RECT 1090.9000 2102.8400 1091.9000 2103.3200 ;
        RECT 1090.9000 2108.2800 1091.9000 2108.7600 ;
        RECT 1090.9000 2081.0800 1091.9000 2081.5600 ;
        RECT 1090.9000 2086.5200 1091.9000 2087.0000 ;
        RECT 1090.9000 2091.9600 1091.9000 2092.4400 ;
        RECT 1045.9000 2113.7200 1046.9000 2114.2000 ;
        RECT 1045.9000 2119.1600 1046.9000 2119.6400 ;
        RECT 1045.9000 2097.4000 1046.9000 2097.8800 ;
        RECT 1045.9000 2102.8400 1046.9000 2103.3200 ;
        RECT 1045.9000 2108.2800 1046.9000 2108.7600 ;
        RECT 1045.9000 2081.0800 1046.9000 2081.5600 ;
        RECT 1045.9000 2086.5200 1046.9000 2087.0000 ;
        RECT 1045.9000 2091.9600 1046.9000 2092.4400 ;
        RECT 1132.3400 2070.2000 1135.3400 2070.6800 ;
        RECT 1132.3400 2075.6400 1135.3400 2076.1200 ;
        RECT 1132.3400 2064.7600 1135.3400 2065.2400 ;
        RECT 1132.3400 2059.3200 1135.3400 2059.8000 ;
        RECT 1132.3400 2053.8800 1135.3400 2054.3600 ;
        RECT 1090.9000 2070.2000 1091.9000 2070.6800 ;
        RECT 1090.9000 2075.6400 1091.9000 2076.1200 ;
        RECT 1090.9000 2053.8800 1091.9000 2054.3600 ;
        RECT 1090.9000 2059.3200 1091.9000 2059.8000 ;
        RECT 1090.9000 2064.7600 1091.9000 2065.2400 ;
        RECT 1132.3400 2037.5600 1135.3400 2038.0400 ;
        RECT 1132.3400 2043.0000 1135.3400 2043.4800 ;
        RECT 1132.3400 2048.4400 1135.3400 2048.9200 ;
        RECT 1132.3400 2032.1200 1135.3400 2032.6000 ;
        RECT 1132.3400 2021.2400 1135.3400 2021.7200 ;
        RECT 1132.3400 2026.6800 1135.3400 2027.1600 ;
        RECT 1090.9000 2037.5600 1091.9000 2038.0400 ;
        RECT 1090.9000 2043.0000 1091.9000 2043.4800 ;
        RECT 1090.9000 2048.4400 1091.9000 2048.9200 ;
        RECT 1090.9000 2021.2400 1091.9000 2021.7200 ;
        RECT 1090.9000 2026.6800 1091.9000 2027.1600 ;
        RECT 1090.9000 2032.1200 1091.9000 2032.6000 ;
        RECT 1045.9000 2070.2000 1046.9000 2070.6800 ;
        RECT 1045.9000 2075.6400 1046.9000 2076.1200 ;
        RECT 1045.9000 2053.8800 1046.9000 2054.3600 ;
        RECT 1045.9000 2059.3200 1046.9000 2059.8000 ;
        RECT 1045.9000 2064.7600 1046.9000 2065.2400 ;
        RECT 1045.9000 2037.5600 1046.9000 2038.0400 ;
        RECT 1045.9000 2043.0000 1046.9000 2043.4800 ;
        RECT 1045.9000 2048.4400 1046.9000 2048.9200 ;
        RECT 1045.9000 2021.2400 1046.9000 2021.7200 ;
        RECT 1045.9000 2026.6800 1046.9000 2027.1600 ;
        RECT 1045.9000 2032.1200 1046.9000 2032.6000 ;
        RECT 1000.9000 2113.7200 1001.9000 2114.2000 ;
        RECT 1000.9000 2119.1600 1001.9000 2119.6400 ;
        RECT 1000.9000 2097.4000 1001.9000 2097.8800 ;
        RECT 1000.9000 2102.8400 1001.9000 2103.3200 ;
        RECT 1000.9000 2108.2800 1001.9000 2108.7600 ;
        RECT 1000.9000 2081.0800 1001.9000 2081.5600 ;
        RECT 1000.9000 2086.5200 1001.9000 2087.0000 ;
        RECT 1000.9000 2091.9600 1001.9000 2092.4400 ;
        RECT 955.9000 2113.7200 956.9000 2114.2000 ;
        RECT 955.9000 2119.1600 956.9000 2119.6400 ;
        RECT 906.3400 2119.1600 909.3400 2119.6400 ;
        RECT 906.3400 2113.7200 909.3400 2114.2000 ;
        RECT 955.9000 2097.4000 956.9000 2097.8800 ;
        RECT 955.9000 2102.8400 956.9000 2103.3200 ;
        RECT 955.9000 2108.2800 956.9000 2108.7600 ;
        RECT 955.9000 2081.0800 956.9000 2081.5600 ;
        RECT 955.9000 2086.5200 956.9000 2087.0000 ;
        RECT 955.9000 2091.9600 956.9000 2092.4400 ;
        RECT 906.3400 2108.2800 909.3400 2108.7600 ;
        RECT 906.3400 2097.4000 909.3400 2097.8800 ;
        RECT 906.3400 2102.8400 909.3400 2103.3200 ;
        RECT 906.3400 2091.9600 909.3400 2092.4400 ;
        RECT 906.3400 2081.0800 909.3400 2081.5600 ;
        RECT 906.3400 2086.5200 909.3400 2087.0000 ;
        RECT 1000.9000 2070.2000 1001.9000 2070.6800 ;
        RECT 1000.9000 2075.6400 1001.9000 2076.1200 ;
        RECT 1000.9000 2053.8800 1001.9000 2054.3600 ;
        RECT 1000.9000 2059.3200 1001.9000 2059.8000 ;
        RECT 1000.9000 2064.7600 1001.9000 2065.2400 ;
        RECT 1000.9000 2037.5600 1001.9000 2038.0400 ;
        RECT 1000.9000 2043.0000 1001.9000 2043.4800 ;
        RECT 1000.9000 2048.4400 1001.9000 2048.9200 ;
        RECT 1000.9000 2021.2400 1001.9000 2021.7200 ;
        RECT 1000.9000 2026.6800 1001.9000 2027.1600 ;
        RECT 1000.9000 2032.1200 1001.9000 2032.6000 ;
        RECT 955.9000 2070.2000 956.9000 2070.6800 ;
        RECT 955.9000 2075.6400 956.9000 2076.1200 ;
        RECT 955.9000 2053.8800 956.9000 2054.3600 ;
        RECT 955.9000 2059.3200 956.9000 2059.8000 ;
        RECT 955.9000 2064.7600 956.9000 2065.2400 ;
        RECT 906.3400 2075.6400 909.3400 2076.1200 ;
        RECT 906.3400 2070.2000 909.3400 2070.6800 ;
        RECT 906.3400 2059.3200 909.3400 2059.8000 ;
        RECT 906.3400 2064.7600 909.3400 2065.2400 ;
        RECT 906.3400 2053.8800 909.3400 2054.3600 ;
        RECT 955.9000 2037.5600 956.9000 2038.0400 ;
        RECT 955.9000 2043.0000 956.9000 2043.4800 ;
        RECT 955.9000 2048.4400 956.9000 2048.9200 ;
        RECT 955.9000 2021.2400 956.9000 2021.7200 ;
        RECT 955.9000 2026.6800 956.9000 2027.1600 ;
        RECT 955.9000 2032.1200 956.9000 2032.6000 ;
        RECT 906.3400 2048.4400 909.3400 2048.9200 ;
        RECT 906.3400 2037.5600 909.3400 2038.0400 ;
        RECT 906.3400 2043.0000 909.3400 2043.4800 ;
        RECT 906.3400 2032.1200 909.3400 2032.6000 ;
        RECT 906.3400 2021.2400 909.3400 2021.7200 ;
        RECT 906.3400 2026.6800 909.3400 2027.1600 ;
        RECT 1132.3400 2010.3600 1135.3400 2010.8400 ;
        RECT 1132.3400 2015.8000 1135.3400 2016.2800 ;
        RECT 1132.3400 2004.9200 1135.3400 2005.4000 ;
        RECT 1132.3400 1999.4800 1135.3400 1999.9600 ;
        RECT 1132.3400 1994.0400 1135.3400 1994.5200 ;
        RECT 1090.9000 2010.3600 1091.9000 2010.8400 ;
        RECT 1090.9000 2015.8000 1091.9000 2016.2800 ;
        RECT 1090.9000 1994.0400 1091.9000 1994.5200 ;
        RECT 1090.9000 1999.4800 1091.9000 1999.9600 ;
        RECT 1090.9000 2004.9200 1091.9000 2005.4000 ;
        RECT 1132.3400 1977.7200 1135.3400 1978.2000 ;
        RECT 1132.3400 1983.1600 1135.3400 1983.6400 ;
        RECT 1132.3400 1988.6000 1135.3400 1989.0800 ;
        RECT 1132.3400 1972.2800 1135.3400 1972.7600 ;
        RECT 1132.3400 1961.4000 1135.3400 1961.8800 ;
        RECT 1132.3400 1966.8400 1135.3400 1967.3200 ;
        RECT 1090.9000 1977.7200 1091.9000 1978.2000 ;
        RECT 1090.9000 1983.1600 1091.9000 1983.6400 ;
        RECT 1090.9000 1988.6000 1091.9000 1989.0800 ;
        RECT 1090.9000 1961.4000 1091.9000 1961.8800 ;
        RECT 1090.9000 1966.8400 1091.9000 1967.3200 ;
        RECT 1090.9000 1972.2800 1091.9000 1972.7600 ;
        RECT 1045.9000 2010.3600 1046.9000 2010.8400 ;
        RECT 1045.9000 2015.8000 1046.9000 2016.2800 ;
        RECT 1045.9000 1994.0400 1046.9000 1994.5200 ;
        RECT 1045.9000 1999.4800 1046.9000 1999.9600 ;
        RECT 1045.9000 2004.9200 1046.9000 2005.4000 ;
        RECT 1045.9000 1977.7200 1046.9000 1978.2000 ;
        RECT 1045.9000 1983.1600 1046.9000 1983.6400 ;
        RECT 1045.9000 1988.6000 1046.9000 1989.0800 ;
        RECT 1045.9000 1961.4000 1046.9000 1961.8800 ;
        RECT 1045.9000 1966.8400 1046.9000 1967.3200 ;
        RECT 1045.9000 1972.2800 1046.9000 1972.7600 ;
        RECT 1132.3400 1950.5200 1135.3400 1951.0000 ;
        RECT 1132.3400 1955.9600 1135.3400 1956.4400 ;
        RECT 1132.3400 1945.0800 1135.3400 1945.5600 ;
        RECT 1132.3400 1939.6400 1135.3400 1940.1200 ;
        RECT 1132.3400 1934.2000 1135.3400 1934.6800 ;
        RECT 1090.9000 1950.5200 1091.9000 1951.0000 ;
        RECT 1090.9000 1955.9600 1091.9000 1956.4400 ;
        RECT 1090.9000 1934.2000 1091.9000 1934.6800 ;
        RECT 1090.9000 1939.6400 1091.9000 1940.1200 ;
        RECT 1090.9000 1945.0800 1091.9000 1945.5600 ;
        RECT 1132.3400 1923.3200 1135.3400 1923.8000 ;
        RECT 1132.3400 1928.7600 1135.3400 1929.2400 ;
        RECT 1090.9000 1923.3200 1091.9000 1923.8000 ;
        RECT 1090.9000 1928.7600 1091.9000 1929.2400 ;
        RECT 1045.9000 1950.5200 1046.9000 1951.0000 ;
        RECT 1045.9000 1955.9600 1046.9000 1956.4400 ;
        RECT 1045.9000 1934.2000 1046.9000 1934.6800 ;
        RECT 1045.9000 1939.6400 1046.9000 1940.1200 ;
        RECT 1045.9000 1945.0800 1046.9000 1945.5600 ;
        RECT 1045.9000 1923.3200 1046.9000 1923.8000 ;
        RECT 1045.9000 1928.7600 1046.9000 1929.2400 ;
        RECT 1000.9000 2010.3600 1001.9000 2010.8400 ;
        RECT 1000.9000 2015.8000 1001.9000 2016.2800 ;
        RECT 1000.9000 1994.0400 1001.9000 1994.5200 ;
        RECT 1000.9000 1999.4800 1001.9000 1999.9600 ;
        RECT 1000.9000 2004.9200 1001.9000 2005.4000 ;
        RECT 1000.9000 1977.7200 1001.9000 1978.2000 ;
        RECT 1000.9000 1983.1600 1001.9000 1983.6400 ;
        RECT 1000.9000 1988.6000 1001.9000 1989.0800 ;
        RECT 1000.9000 1961.4000 1001.9000 1961.8800 ;
        RECT 1000.9000 1966.8400 1001.9000 1967.3200 ;
        RECT 1000.9000 1972.2800 1001.9000 1972.7600 ;
        RECT 955.9000 2010.3600 956.9000 2010.8400 ;
        RECT 955.9000 2015.8000 956.9000 2016.2800 ;
        RECT 955.9000 1994.0400 956.9000 1994.5200 ;
        RECT 955.9000 1999.4800 956.9000 1999.9600 ;
        RECT 955.9000 2004.9200 956.9000 2005.4000 ;
        RECT 906.3400 2015.8000 909.3400 2016.2800 ;
        RECT 906.3400 2010.3600 909.3400 2010.8400 ;
        RECT 906.3400 1999.4800 909.3400 1999.9600 ;
        RECT 906.3400 2004.9200 909.3400 2005.4000 ;
        RECT 906.3400 1994.0400 909.3400 1994.5200 ;
        RECT 955.9000 1977.7200 956.9000 1978.2000 ;
        RECT 955.9000 1983.1600 956.9000 1983.6400 ;
        RECT 955.9000 1988.6000 956.9000 1989.0800 ;
        RECT 955.9000 1961.4000 956.9000 1961.8800 ;
        RECT 955.9000 1966.8400 956.9000 1967.3200 ;
        RECT 955.9000 1972.2800 956.9000 1972.7600 ;
        RECT 906.3400 1988.6000 909.3400 1989.0800 ;
        RECT 906.3400 1977.7200 909.3400 1978.2000 ;
        RECT 906.3400 1983.1600 909.3400 1983.6400 ;
        RECT 906.3400 1972.2800 909.3400 1972.7600 ;
        RECT 906.3400 1961.4000 909.3400 1961.8800 ;
        RECT 906.3400 1966.8400 909.3400 1967.3200 ;
        RECT 1000.9000 1950.5200 1001.9000 1951.0000 ;
        RECT 1000.9000 1955.9600 1001.9000 1956.4400 ;
        RECT 1000.9000 1934.2000 1001.9000 1934.6800 ;
        RECT 1000.9000 1939.6400 1001.9000 1940.1200 ;
        RECT 1000.9000 1945.0800 1001.9000 1945.5600 ;
        RECT 1000.9000 1923.3200 1001.9000 1923.8000 ;
        RECT 1000.9000 1928.7600 1001.9000 1929.2400 ;
        RECT 955.9000 1950.5200 956.9000 1951.0000 ;
        RECT 955.9000 1955.9600 956.9000 1956.4400 ;
        RECT 955.9000 1934.2000 956.9000 1934.6800 ;
        RECT 955.9000 1939.6400 956.9000 1940.1200 ;
        RECT 955.9000 1945.0800 956.9000 1945.5600 ;
        RECT 906.3400 1955.9600 909.3400 1956.4400 ;
        RECT 906.3400 1950.5200 909.3400 1951.0000 ;
        RECT 906.3400 1939.6400 909.3400 1940.1200 ;
        RECT 906.3400 1945.0800 909.3400 1945.5600 ;
        RECT 906.3400 1934.2000 909.3400 1934.6800 ;
        RECT 955.9000 1923.3200 956.9000 1923.8000 ;
        RECT 955.9000 1928.7600 956.9000 1929.2400 ;
        RECT 906.3400 1928.7600 909.3400 1929.2400 ;
        RECT 906.3400 1923.3200 909.3400 1923.8000 ;
        RECT 906.3400 2121.5100 1135.3400 2124.5100 ;
        RECT 906.3400 1916.4100 1135.3400 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 1686.7700 1091.9000 1894.8700 ;
        RECT 1045.9000 1686.7700 1046.9000 1894.8700 ;
        RECT 1000.9000 1686.7700 1001.9000 1894.8700 ;
        RECT 955.9000 1686.7700 956.9000 1894.8700 ;
        RECT 1132.3400 1686.7700 1135.3400 1894.8700 ;
        RECT 906.3400 1686.7700 909.3400 1894.8700 ;
      LAYER met3 ;
        RECT 1132.3400 1884.0800 1135.3400 1884.5600 ;
        RECT 1132.3400 1889.5200 1135.3400 1890.0000 ;
        RECT 1090.9000 1884.0800 1091.9000 1884.5600 ;
        RECT 1090.9000 1889.5200 1091.9000 1890.0000 ;
        RECT 1132.3400 1867.7600 1135.3400 1868.2400 ;
        RECT 1132.3400 1873.2000 1135.3400 1873.6800 ;
        RECT 1132.3400 1878.6400 1135.3400 1879.1200 ;
        RECT 1132.3400 1862.3200 1135.3400 1862.8000 ;
        RECT 1132.3400 1851.4400 1135.3400 1851.9200 ;
        RECT 1132.3400 1856.8800 1135.3400 1857.3600 ;
        RECT 1090.9000 1867.7600 1091.9000 1868.2400 ;
        RECT 1090.9000 1873.2000 1091.9000 1873.6800 ;
        RECT 1090.9000 1878.6400 1091.9000 1879.1200 ;
        RECT 1090.9000 1851.4400 1091.9000 1851.9200 ;
        RECT 1090.9000 1856.8800 1091.9000 1857.3600 ;
        RECT 1090.9000 1862.3200 1091.9000 1862.8000 ;
        RECT 1045.9000 1884.0800 1046.9000 1884.5600 ;
        RECT 1045.9000 1889.5200 1046.9000 1890.0000 ;
        RECT 1045.9000 1867.7600 1046.9000 1868.2400 ;
        RECT 1045.9000 1873.2000 1046.9000 1873.6800 ;
        RECT 1045.9000 1878.6400 1046.9000 1879.1200 ;
        RECT 1045.9000 1851.4400 1046.9000 1851.9200 ;
        RECT 1045.9000 1856.8800 1046.9000 1857.3600 ;
        RECT 1045.9000 1862.3200 1046.9000 1862.8000 ;
        RECT 1132.3400 1840.5600 1135.3400 1841.0400 ;
        RECT 1132.3400 1846.0000 1135.3400 1846.4800 ;
        RECT 1132.3400 1835.1200 1135.3400 1835.6000 ;
        RECT 1132.3400 1829.6800 1135.3400 1830.1600 ;
        RECT 1132.3400 1824.2400 1135.3400 1824.7200 ;
        RECT 1090.9000 1840.5600 1091.9000 1841.0400 ;
        RECT 1090.9000 1846.0000 1091.9000 1846.4800 ;
        RECT 1090.9000 1824.2400 1091.9000 1824.7200 ;
        RECT 1090.9000 1829.6800 1091.9000 1830.1600 ;
        RECT 1090.9000 1835.1200 1091.9000 1835.6000 ;
        RECT 1132.3400 1807.9200 1135.3400 1808.4000 ;
        RECT 1132.3400 1813.3600 1135.3400 1813.8400 ;
        RECT 1132.3400 1818.8000 1135.3400 1819.2800 ;
        RECT 1132.3400 1802.4800 1135.3400 1802.9600 ;
        RECT 1132.3400 1791.6000 1135.3400 1792.0800 ;
        RECT 1132.3400 1797.0400 1135.3400 1797.5200 ;
        RECT 1090.9000 1807.9200 1091.9000 1808.4000 ;
        RECT 1090.9000 1813.3600 1091.9000 1813.8400 ;
        RECT 1090.9000 1818.8000 1091.9000 1819.2800 ;
        RECT 1090.9000 1791.6000 1091.9000 1792.0800 ;
        RECT 1090.9000 1797.0400 1091.9000 1797.5200 ;
        RECT 1090.9000 1802.4800 1091.9000 1802.9600 ;
        RECT 1045.9000 1840.5600 1046.9000 1841.0400 ;
        RECT 1045.9000 1846.0000 1046.9000 1846.4800 ;
        RECT 1045.9000 1824.2400 1046.9000 1824.7200 ;
        RECT 1045.9000 1829.6800 1046.9000 1830.1600 ;
        RECT 1045.9000 1835.1200 1046.9000 1835.6000 ;
        RECT 1045.9000 1807.9200 1046.9000 1808.4000 ;
        RECT 1045.9000 1813.3600 1046.9000 1813.8400 ;
        RECT 1045.9000 1818.8000 1046.9000 1819.2800 ;
        RECT 1045.9000 1791.6000 1046.9000 1792.0800 ;
        RECT 1045.9000 1797.0400 1046.9000 1797.5200 ;
        RECT 1045.9000 1802.4800 1046.9000 1802.9600 ;
        RECT 1000.9000 1884.0800 1001.9000 1884.5600 ;
        RECT 1000.9000 1889.5200 1001.9000 1890.0000 ;
        RECT 1000.9000 1867.7600 1001.9000 1868.2400 ;
        RECT 1000.9000 1873.2000 1001.9000 1873.6800 ;
        RECT 1000.9000 1878.6400 1001.9000 1879.1200 ;
        RECT 1000.9000 1851.4400 1001.9000 1851.9200 ;
        RECT 1000.9000 1856.8800 1001.9000 1857.3600 ;
        RECT 1000.9000 1862.3200 1001.9000 1862.8000 ;
        RECT 955.9000 1884.0800 956.9000 1884.5600 ;
        RECT 955.9000 1889.5200 956.9000 1890.0000 ;
        RECT 906.3400 1889.5200 909.3400 1890.0000 ;
        RECT 906.3400 1884.0800 909.3400 1884.5600 ;
        RECT 955.9000 1867.7600 956.9000 1868.2400 ;
        RECT 955.9000 1873.2000 956.9000 1873.6800 ;
        RECT 955.9000 1878.6400 956.9000 1879.1200 ;
        RECT 955.9000 1851.4400 956.9000 1851.9200 ;
        RECT 955.9000 1856.8800 956.9000 1857.3600 ;
        RECT 955.9000 1862.3200 956.9000 1862.8000 ;
        RECT 906.3400 1878.6400 909.3400 1879.1200 ;
        RECT 906.3400 1867.7600 909.3400 1868.2400 ;
        RECT 906.3400 1873.2000 909.3400 1873.6800 ;
        RECT 906.3400 1862.3200 909.3400 1862.8000 ;
        RECT 906.3400 1851.4400 909.3400 1851.9200 ;
        RECT 906.3400 1856.8800 909.3400 1857.3600 ;
        RECT 1000.9000 1840.5600 1001.9000 1841.0400 ;
        RECT 1000.9000 1846.0000 1001.9000 1846.4800 ;
        RECT 1000.9000 1824.2400 1001.9000 1824.7200 ;
        RECT 1000.9000 1829.6800 1001.9000 1830.1600 ;
        RECT 1000.9000 1835.1200 1001.9000 1835.6000 ;
        RECT 1000.9000 1807.9200 1001.9000 1808.4000 ;
        RECT 1000.9000 1813.3600 1001.9000 1813.8400 ;
        RECT 1000.9000 1818.8000 1001.9000 1819.2800 ;
        RECT 1000.9000 1791.6000 1001.9000 1792.0800 ;
        RECT 1000.9000 1797.0400 1001.9000 1797.5200 ;
        RECT 1000.9000 1802.4800 1001.9000 1802.9600 ;
        RECT 955.9000 1840.5600 956.9000 1841.0400 ;
        RECT 955.9000 1846.0000 956.9000 1846.4800 ;
        RECT 955.9000 1824.2400 956.9000 1824.7200 ;
        RECT 955.9000 1829.6800 956.9000 1830.1600 ;
        RECT 955.9000 1835.1200 956.9000 1835.6000 ;
        RECT 906.3400 1846.0000 909.3400 1846.4800 ;
        RECT 906.3400 1840.5600 909.3400 1841.0400 ;
        RECT 906.3400 1829.6800 909.3400 1830.1600 ;
        RECT 906.3400 1835.1200 909.3400 1835.6000 ;
        RECT 906.3400 1824.2400 909.3400 1824.7200 ;
        RECT 955.9000 1807.9200 956.9000 1808.4000 ;
        RECT 955.9000 1813.3600 956.9000 1813.8400 ;
        RECT 955.9000 1818.8000 956.9000 1819.2800 ;
        RECT 955.9000 1791.6000 956.9000 1792.0800 ;
        RECT 955.9000 1797.0400 956.9000 1797.5200 ;
        RECT 955.9000 1802.4800 956.9000 1802.9600 ;
        RECT 906.3400 1818.8000 909.3400 1819.2800 ;
        RECT 906.3400 1807.9200 909.3400 1808.4000 ;
        RECT 906.3400 1813.3600 909.3400 1813.8400 ;
        RECT 906.3400 1802.4800 909.3400 1802.9600 ;
        RECT 906.3400 1791.6000 909.3400 1792.0800 ;
        RECT 906.3400 1797.0400 909.3400 1797.5200 ;
        RECT 1132.3400 1780.7200 1135.3400 1781.2000 ;
        RECT 1132.3400 1786.1600 1135.3400 1786.6400 ;
        RECT 1132.3400 1775.2800 1135.3400 1775.7600 ;
        RECT 1132.3400 1769.8400 1135.3400 1770.3200 ;
        RECT 1132.3400 1764.4000 1135.3400 1764.8800 ;
        RECT 1090.9000 1780.7200 1091.9000 1781.2000 ;
        RECT 1090.9000 1786.1600 1091.9000 1786.6400 ;
        RECT 1090.9000 1764.4000 1091.9000 1764.8800 ;
        RECT 1090.9000 1769.8400 1091.9000 1770.3200 ;
        RECT 1090.9000 1775.2800 1091.9000 1775.7600 ;
        RECT 1132.3400 1748.0800 1135.3400 1748.5600 ;
        RECT 1132.3400 1753.5200 1135.3400 1754.0000 ;
        RECT 1132.3400 1758.9600 1135.3400 1759.4400 ;
        RECT 1132.3400 1742.6400 1135.3400 1743.1200 ;
        RECT 1132.3400 1731.7600 1135.3400 1732.2400 ;
        RECT 1132.3400 1737.2000 1135.3400 1737.6800 ;
        RECT 1090.9000 1748.0800 1091.9000 1748.5600 ;
        RECT 1090.9000 1753.5200 1091.9000 1754.0000 ;
        RECT 1090.9000 1758.9600 1091.9000 1759.4400 ;
        RECT 1090.9000 1731.7600 1091.9000 1732.2400 ;
        RECT 1090.9000 1737.2000 1091.9000 1737.6800 ;
        RECT 1090.9000 1742.6400 1091.9000 1743.1200 ;
        RECT 1045.9000 1780.7200 1046.9000 1781.2000 ;
        RECT 1045.9000 1786.1600 1046.9000 1786.6400 ;
        RECT 1045.9000 1764.4000 1046.9000 1764.8800 ;
        RECT 1045.9000 1769.8400 1046.9000 1770.3200 ;
        RECT 1045.9000 1775.2800 1046.9000 1775.7600 ;
        RECT 1045.9000 1748.0800 1046.9000 1748.5600 ;
        RECT 1045.9000 1753.5200 1046.9000 1754.0000 ;
        RECT 1045.9000 1758.9600 1046.9000 1759.4400 ;
        RECT 1045.9000 1731.7600 1046.9000 1732.2400 ;
        RECT 1045.9000 1737.2000 1046.9000 1737.6800 ;
        RECT 1045.9000 1742.6400 1046.9000 1743.1200 ;
        RECT 1132.3400 1720.8800 1135.3400 1721.3600 ;
        RECT 1132.3400 1726.3200 1135.3400 1726.8000 ;
        RECT 1132.3400 1715.4400 1135.3400 1715.9200 ;
        RECT 1132.3400 1710.0000 1135.3400 1710.4800 ;
        RECT 1132.3400 1704.5600 1135.3400 1705.0400 ;
        RECT 1090.9000 1720.8800 1091.9000 1721.3600 ;
        RECT 1090.9000 1726.3200 1091.9000 1726.8000 ;
        RECT 1090.9000 1704.5600 1091.9000 1705.0400 ;
        RECT 1090.9000 1710.0000 1091.9000 1710.4800 ;
        RECT 1090.9000 1715.4400 1091.9000 1715.9200 ;
        RECT 1132.3400 1693.6800 1135.3400 1694.1600 ;
        RECT 1132.3400 1699.1200 1135.3400 1699.6000 ;
        RECT 1090.9000 1693.6800 1091.9000 1694.1600 ;
        RECT 1090.9000 1699.1200 1091.9000 1699.6000 ;
        RECT 1045.9000 1720.8800 1046.9000 1721.3600 ;
        RECT 1045.9000 1726.3200 1046.9000 1726.8000 ;
        RECT 1045.9000 1704.5600 1046.9000 1705.0400 ;
        RECT 1045.9000 1710.0000 1046.9000 1710.4800 ;
        RECT 1045.9000 1715.4400 1046.9000 1715.9200 ;
        RECT 1045.9000 1693.6800 1046.9000 1694.1600 ;
        RECT 1045.9000 1699.1200 1046.9000 1699.6000 ;
        RECT 1000.9000 1780.7200 1001.9000 1781.2000 ;
        RECT 1000.9000 1786.1600 1001.9000 1786.6400 ;
        RECT 1000.9000 1764.4000 1001.9000 1764.8800 ;
        RECT 1000.9000 1769.8400 1001.9000 1770.3200 ;
        RECT 1000.9000 1775.2800 1001.9000 1775.7600 ;
        RECT 1000.9000 1748.0800 1001.9000 1748.5600 ;
        RECT 1000.9000 1753.5200 1001.9000 1754.0000 ;
        RECT 1000.9000 1758.9600 1001.9000 1759.4400 ;
        RECT 1000.9000 1731.7600 1001.9000 1732.2400 ;
        RECT 1000.9000 1737.2000 1001.9000 1737.6800 ;
        RECT 1000.9000 1742.6400 1001.9000 1743.1200 ;
        RECT 955.9000 1780.7200 956.9000 1781.2000 ;
        RECT 955.9000 1786.1600 956.9000 1786.6400 ;
        RECT 955.9000 1764.4000 956.9000 1764.8800 ;
        RECT 955.9000 1769.8400 956.9000 1770.3200 ;
        RECT 955.9000 1775.2800 956.9000 1775.7600 ;
        RECT 906.3400 1786.1600 909.3400 1786.6400 ;
        RECT 906.3400 1780.7200 909.3400 1781.2000 ;
        RECT 906.3400 1769.8400 909.3400 1770.3200 ;
        RECT 906.3400 1775.2800 909.3400 1775.7600 ;
        RECT 906.3400 1764.4000 909.3400 1764.8800 ;
        RECT 955.9000 1748.0800 956.9000 1748.5600 ;
        RECT 955.9000 1753.5200 956.9000 1754.0000 ;
        RECT 955.9000 1758.9600 956.9000 1759.4400 ;
        RECT 955.9000 1731.7600 956.9000 1732.2400 ;
        RECT 955.9000 1737.2000 956.9000 1737.6800 ;
        RECT 955.9000 1742.6400 956.9000 1743.1200 ;
        RECT 906.3400 1758.9600 909.3400 1759.4400 ;
        RECT 906.3400 1748.0800 909.3400 1748.5600 ;
        RECT 906.3400 1753.5200 909.3400 1754.0000 ;
        RECT 906.3400 1742.6400 909.3400 1743.1200 ;
        RECT 906.3400 1731.7600 909.3400 1732.2400 ;
        RECT 906.3400 1737.2000 909.3400 1737.6800 ;
        RECT 1000.9000 1720.8800 1001.9000 1721.3600 ;
        RECT 1000.9000 1726.3200 1001.9000 1726.8000 ;
        RECT 1000.9000 1704.5600 1001.9000 1705.0400 ;
        RECT 1000.9000 1710.0000 1001.9000 1710.4800 ;
        RECT 1000.9000 1715.4400 1001.9000 1715.9200 ;
        RECT 1000.9000 1693.6800 1001.9000 1694.1600 ;
        RECT 1000.9000 1699.1200 1001.9000 1699.6000 ;
        RECT 955.9000 1720.8800 956.9000 1721.3600 ;
        RECT 955.9000 1726.3200 956.9000 1726.8000 ;
        RECT 955.9000 1704.5600 956.9000 1705.0400 ;
        RECT 955.9000 1710.0000 956.9000 1710.4800 ;
        RECT 955.9000 1715.4400 956.9000 1715.9200 ;
        RECT 906.3400 1726.3200 909.3400 1726.8000 ;
        RECT 906.3400 1720.8800 909.3400 1721.3600 ;
        RECT 906.3400 1710.0000 909.3400 1710.4800 ;
        RECT 906.3400 1715.4400 909.3400 1715.9200 ;
        RECT 906.3400 1704.5600 909.3400 1705.0400 ;
        RECT 955.9000 1693.6800 956.9000 1694.1600 ;
        RECT 955.9000 1699.1200 956.9000 1699.6000 ;
        RECT 906.3400 1699.1200 909.3400 1699.6000 ;
        RECT 906.3400 1693.6800 909.3400 1694.1600 ;
        RECT 906.3400 1891.8700 1135.3400 1894.8700 ;
        RECT 906.3400 1686.7700 1135.3400 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 1457.1300 1091.9000 1665.2300 ;
        RECT 1045.9000 1457.1300 1046.9000 1665.2300 ;
        RECT 1000.9000 1457.1300 1001.9000 1665.2300 ;
        RECT 955.9000 1457.1300 956.9000 1665.2300 ;
        RECT 1132.3400 1457.1300 1135.3400 1665.2300 ;
        RECT 906.3400 1457.1300 909.3400 1665.2300 ;
      LAYER met3 ;
        RECT 1132.3400 1654.4400 1135.3400 1654.9200 ;
        RECT 1132.3400 1659.8800 1135.3400 1660.3600 ;
        RECT 1090.9000 1654.4400 1091.9000 1654.9200 ;
        RECT 1090.9000 1659.8800 1091.9000 1660.3600 ;
        RECT 1132.3400 1638.1200 1135.3400 1638.6000 ;
        RECT 1132.3400 1643.5600 1135.3400 1644.0400 ;
        RECT 1132.3400 1649.0000 1135.3400 1649.4800 ;
        RECT 1132.3400 1632.6800 1135.3400 1633.1600 ;
        RECT 1132.3400 1621.8000 1135.3400 1622.2800 ;
        RECT 1132.3400 1627.2400 1135.3400 1627.7200 ;
        RECT 1090.9000 1638.1200 1091.9000 1638.6000 ;
        RECT 1090.9000 1643.5600 1091.9000 1644.0400 ;
        RECT 1090.9000 1649.0000 1091.9000 1649.4800 ;
        RECT 1090.9000 1621.8000 1091.9000 1622.2800 ;
        RECT 1090.9000 1627.2400 1091.9000 1627.7200 ;
        RECT 1090.9000 1632.6800 1091.9000 1633.1600 ;
        RECT 1045.9000 1654.4400 1046.9000 1654.9200 ;
        RECT 1045.9000 1659.8800 1046.9000 1660.3600 ;
        RECT 1045.9000 1638.1200 1046.9000 1638.6000 ;
        RECT 1045.9000 1643.5600 1046.9000 1644.0400 ;
        RECT 1045.9000 1649.0000 1046.9000 1649.4800 ;
        RECT 1045.9000 1621.8000 1046.9000 1622.2800 ;
        RECT 1045.9000 1627.2400 1046.9000 1627.7200 ;
        RECT 1045.9000 1632.6800 1046.9000 1633.1600 ;
        RECT 1132.3400 1610.9200 1135.3400 1611.4000 ;
        RECT 1132.3400 1616.3600 1135.3400 1616.8400 ;
        RECT 1132.3400 1605.4800 1135.3400 1605.9600 ;
        RECT 1132.3400 1600.0400 1135.3400 1600.5200 ;
        RECT 1132.3400 1594.6000 1135.3400 1595.0800 ;
        RECT 1090.9000 1610.9200 1091.9000 1611.4000 ;
        RECT 1090.9000 1616.3600 1091.9000 1616.8400 ;
        RECT 1090.9000 1594.6000 1091.9000 1595.0800 ;
        RECT 1090.9000 1600.0400 1091.9000 1600.5200 ;
        RECT 1090.9000 1605.4800 1091.9000 1605.9600 ;
        RECT 1132.3400 1578.2800 1135.3400 1578.7600 ;
        RECT 1132.3400 1583.7200 1135.3400 1584.2000 ;
        RECT 1132.3400 1589.1600 1135.3400 1589.6400 ;
        RECT 1132.3400 1572.8400 1135.3400 1573.3200 ;
        RECT 1132.3400 1561.9600 1135.3400 1562.4400 ;
        RECT 1132.3400 1567.4000 1135.3400 1567.8800 ;
        RECT 1090.9000 1578.2800 1091.9000 1578.7600 ;
        RECT 1090.9000 1583.7200 1091.9000 1584.2000 ;
        RECT 1090.9000 1589.1600 1091.9000 1589.6400 ;
        RECT 1090.9000 1561.9600 1091.9000 1562.4400 ;
        RECT 1090.9000 1567.4000 1091.9000 1567.8800 ;
        RECT 1090.9000 1572.8400 1091.9000 1573.3200 ;
        RECT 1045.9000 1610.9200 1046.9000 1611.4000 ;
        RECT 1045.9000 1616.3600 1046.9000 1616.8400 ;
        RECT 1045.9000 1594.6000 1046.9000 1595.0800 ;
        RECT 1045.9000 1600.0400 1046.9000 1600.5200 ;
        RECT 1045.9000 1605.4800 1046.9000 1605.9600 ;
        RECT 1045.9000 1578.2800 1046.9000 1578.7600 ;
        RECT 1045.9000 1583.7200 1046.9000 1584.2000 ;
        RECT 1045.9000 1589.1600 1046.9000 1589.6400 ;
        RECT 1045.9000 1561.9600 1046.9000 1562.4400 ;
        RECT 1045.9000 1567.4000 1046.9000 1567.8800 ;
        RECT 1045.9000 1572.8400 1046.9000 1573.3200 ;
        RECT 1000.9000 1654.4400 1001.9000 1654.9200 ;
        RECT 1000.9000 1659.8800 1001.9000 1660.3600 ;
        RECT 1000.9000 1638.1200 1001.9000 1638.6000 ;
        RECT 1000.9000 1643.5600 1001.9000 1644.0400 ;
        RECT 1000.9000 1649.0000 1001.9000 1649.4800 ;
        RECT 1000.9000 1621.8000 1001.9000 1622.2800 ;
        RECT 1000.9000 1627.2400 1001.9000 1627.7200 ;
        RECT 1000.9000 1632.6800 1001.9000 1633.1600 ;
        RECT 955.9000 1654.4400 956.9000 1654.9200 ;
        RECT 955.9000 1659.8800 956.9000 1660.3600 ;
        RECT 906.3400 1659.8800 909.3400 1660.3600 ;
        RECT 906.3400 1654.4400 909.3400 1654.9200 ;
        RECT 955.9000 1638.1200 956.9000 1638.6000 ;
        RECT 955.9000 1643.5600 956.9000 1644.0400 ;
        RECT 955.9000 1649.0000 956.9000 1649.4800 ;
        RECT 955.9000 1621.8000 956.9000 1622.2800 ;
        RECT 955.9000 1627.2400 956.9000 1627.7200 ;
        RECT 955.9000 1632.6800 956.9000 1633.1600 ;
        RECT 906.3400 1649.0000 909.3400 1649.4800 ;
        RECT 906.3400 1638.1200 909.3400 1638.6000 ;
        RECT 906.3400 1643.5600 909.3400 1644.0400 ;
        RECT 906.3400 1632.6800 909.3400 1633.1600 ;
        RECT 906.3400 1621.8000 909.3400 1622.2800 ;
        RECT 906.3400 1627.2400 909.3400 1627.7200 ;
        RECT 1000.9000 1610.9200 1001.9000 1611.4000 ;
        RECT 1000.9000 1616.3600 1001.9000 1616.8400 ;
        RECT 1000.9000 1594.6000 1001.9000 1595.0800 ;
        RECT 1000.9000 1600.0400 1001.9000 1600.5200 ;
        RECT 1000.9000 1605.4800 1001.9000 1605.9600 ;
        RECT 1000.9000 1578.2800 1001.9000 1578.7600 ;
        RECT 1000.9000 1583.7200 1001.9000 1584.2000 ;
        RECT 1000.9000 1589.1600 1001.9000 1589.6400 ;
        RECT 1000.9000 1561.9600 1001.9000 1562.4400 ;
        RECT 1000.9000 1567.4000 1001.9000 1567.8800 ;
        RECT 1000.9000 1572.8400 1001.9000 1573.3200 ;
        RECT 955.9000 1610.9200 956.9000 1611.4000 ;
        RECT 955.9000 1616.3600 956.9000 1616.8400 ;
        RECT 955.9000 1594.6000 956.9000 1595.0800 ;
        RECT 955.9000 1600.0400 956.9000 1600.5200 ;
        RECT 955.9000 1605.4800 956.9000 1605.9600 ;
        RECT 906.3400 1616.3600 909.3400 1616.8400 ;
        RECT 906.3400 1610.9200 909.3400 1611.4000 ;
        RECT 906.3400 1600.0400 909.3400 1600.5200 ;
        RECT 906.3400 1605.4800 909.3400 1605.9600 ;
        RECT 906.3400 1594.6000 909.3400 1595.0800 ;
        RECT 955.9000 1578.2800 956.9000 1578.7600 ;
        RECT 955.9000 1583.7200 956.9000 1584.2000 ;
        RECT 955.9000 1589.1600 956.9000 1589.6400 ;
        RECT 955.9000 1561.9600 956.9000 1562.4400 ;
        RECT 955.9000 1567.4000 956.9000 1567.8800 ;
        RECT 955.9000 1572.8400 956.9000 1573.3200 ;
        RECT 906.3400 1589.1600 909.3400 1589.6400 ;
        RECT 906.3400 1578.2800 909.3400 1578.7600 ;
        RECT 906.3400 1583.7200 909.3400 1584.2000 ;
        RECT 906.3400 1572.8400 909.3400 1573.3200 ;
        RECT 906.3400 1561.9600 909.3400 1562.4400 ;
        RECT 906.3400 1567.4000 909.3400 1567.8800 ;
        RECT 1132.3400 1551.0800 1135.3400 1551.5600 ;
        RECT 1132.3400 1556.5200 1135.3400 1557.0000 ;
        RECT 1132.3400 1545.6400 1135.3400 1546.1200 ;
        RECT 1132.3400 1540.2000 1135.3400 1540.6800 ;
        RECT 1132.3400 1534.7600 1135.3400 1535.2400 ;
        RECT 1090.9000 1551.0800 1091.9000 1551.5600 ;
        RECT 1090.9000 1556.5200 1091.9000 1557.0000 ;
        RECT 1090.9000 1534.7600 1091.9000 1535.2400 ;
        RECT 1090.9000 1540.2000 1091.9000 1540.6800 ;
        RECT 1090.9000 1545.6400 1091.9000 1546.1200 ;
        RECT 1132.3400 1518.4400 1135.3400 1518.9200 ;
        RECT 1132.3400 1523.8800 1135.3400 1524.3600 ;
        RECT 1132.3400 1529.3200 1135.3400 1529.8000 ;
        RECT 1132.3400 1513.0000 1135.3400 1513.4800 ;
        RECT 1132.3400 1502.1200 1135.3400 1502.6000 ;
        RECT 1132.3400 1507.5600 1135.3400 1508.0400 ;
        RECT 1090.9000 1518.4400 1091.9000 1518.9200 ;
        RECT 1090.9000 1523.8800 1091.9000 1524.3600 ;
        RECT 1090.9000 1529.3200 1091.9000 1529.8000 ;
        RECT 1090.9000 1502.1200 1091.9000 1502.6000 ;
        RECT 1090.9000 1507.5600 1091.9000 1508.0400 ;
        RECT 1090.9000 1513.0000 1091.9000 1513.4800 ;
        RECT 1045.9000 1551.0800 1046.9000 1551.5600 ;
        RECT 1045.9000 1556.5200 1046.9000 1557.0000 ;
        RECT 1045.9000 1534.7600 1046.9000 1535.2400 ;
        RECT 1045.9000 1540.2000 1046.9000 1540.6800 ;
        RECT 1045.9000 1545.6400 1046.9000 1546.1200 ;
        RECT 1045.9000 1518.4400 1046.9000 1518.9200 ;
        RECT 1045.9000 1523.8800 1046.9000 1524.3600 ;
        RECT 1045.9000 1529.3200 1046.9000 1529.8000 ;
        RECT 1045.9000 1502.1200 1046.9000 1502.6000 ;
        RECT 1045.9000 1507.5600 1046.9000 1508.0400 ;
        RECT 1045.9000 1513.0000 1046.9000 1513.4800 ;
        RECT 1132.3400 1491.2400 1135.3400 1491.7200 ;
        RECT 1132.3400 1496.6800 1135.3400 1497.1600 ;
        RECT 1132.3400 1485.8000 1135.3400 1486.2800 ;
        RECT 1132.3400 1480.3600 1135.3400 1480.8400 ;
        RECT 1132.3400 1474.9200 1135.3400 1475.4000 ;
        RECT 1090.9000 1491.2400 1091.9000 1491.7200 ;
        RECT 1090.9000 1496.6800 1091.9000 1497.1600 ;
        RECT 1090.9000 1474.9200 1091.9000 1475.4000 ;
        RECT 1090.9000 1480.3600 1091.9000 1480.8400 ;
        RECT 1090.9000 1485.8000 1091.9000 1486.2800 ;
        RECT 1132.3400 1464.0400 1135.3400 1464.5200 ;
        RECT 1132.3400 1469.4800 1135.3400 1469.9600 ;
        RECT 1090.9000 1464.0400 1091.9000 1464.5200 ;
        RECT 1090.9000 1469.4800 1091.9000 1469.9600 ;
        RECT 1045.9000 1491.2400 1046.9000 1491.7200 ;
        RECT 1045.9000 1496.6800 1046.9000 1497.1600 ;
        RECT 1045.9000 1474.9200 1046.9000 1475.4000 ;
        RECT 1045.9000 1480.3600 1046.9000 1480.8400 ;
        RECT 1045.9000 1485.8000 1046.9000 1486.2800 ;
        RECT 1045.9000 1464.0400 1046.9000 1464.5200 ;
        RECT 1045.9000 1469.4800 1046.9000 1469.9600 ;
        RECT 1000.9000 1551.0800 1001.9000 1551.5600 ;
        RECT 1000.9000 1556.5200 1001.9000 1557.0000 ;
        RECT 1000.9000 1534.7600 1001.9000 1535.2400 ;
        RECT 1000.9000 1540.2000 1001.9000 1540.6800 ;
        RECT 1000.9000 1545.6400 1001.9000 1546.1200 ;
        RECT 1000.9000 1518.4400 1001.9000 1518.9200 ;
        RECT 1000.9000 1523.8800 1001.9000 1524.3600 ;
        RECT 1000.9000 1529.3200 1001.9000 1529.8000 ;
        RECT 1000.9000 1502.1200 1001.9000 1502.6000 ;
        RECT 1000.9000 1507.5600 1001.9000 1508.0400 ;
        RECT 1000.9000 1513.0000 1001.9000 1513.4800 ;
        RECT 955.9000 1551.0800 956.9000 1551.5600 ;
        RECT 955.9000 1556.5200 956.9000 1557.0000 ;
        RECT 955.9000 1534.7600 956.9000 1535.2400 ;
        RECT 955.9000 1540.2000 956.9000 1540.6800 ;
        RECT 955.9000 1545.6400 956.9000 1546.1200 ;
        RECT 906.3400 1556.5200 909.3400 1557.0000 ;
        RECT 906.3400 1551.0800 909.3400 1551.5600 ;
        RECT 906.3400 1540.2000 909.3400 1540.6800 ;
        RECT 906.3400 1545.6400 909.3400 1546.1200 ;
        RECT 906.3400 1534.7600 909.3400 1535.2400 ;
        RECT 955.9000 1518.4400 956.9000 1518.9200 ;
        RECT 955.9000 1523.8800 956.9000 1524.3600 ;
        RECT 955.9000 1529.3200 956.9000 1529.8000 ;
        RECT 955.9000 1502.1200 956.9000 1502.6000 ;
        RECT 955.9000 1507.5600 956.9000 1508.0400 ;
        RECT 955.9000 1513.0000 956.9000 1513.4800 ;
        RECT 906.3400 1529.3200 909.3400 1529.8000 ;
        RECT 906.3400 1518.4400 909.3400 1518.9200 ;
        RECT 906.3400 1523.8800 909.3400 1524.3600 ;
        RECT 906.3400 1513.0000 909.3400 1513.4800 ;
        RECT 906.3400 1502.1200 909.3400 1502.6000 ;
        RECT 906.3400 1507.5600 909.3400 1508.0400 ;
        RECT 1000.9000 1491.2400 1001.9000 1491.7200 ;
        RECT 1000.9000 1496.6800 1001.9000 1497.1600 ;
        RECT 1000.9000 1474.9200 1001.9000 1475.4000 ;
        RECT 1000.9000 1480.3600 1001.9000 1480.8400 ;
        RECT 1000.9000 1485.8000 1001.9000 1486.2800 ;
        RECT 1000.9000 1464.0400 1001.9000 1464.5200 ;
        RECT 1000.9000 1469.4800 1001.9000 1469.9600 ;
        RECT 955.9000 1491.2400 956.9000 1491.7200 ;
        RECT 955.9000 1496.6800 956.9000 1497.1600 ;
        RECT 955.9000 1474.9200 956.9000 1475.4000 ;
        RECT 955.9000 1480.3600 956.9000 1480.8400 ;
        RECT 955.9000 1485.8000 956.9000 1486.2800 ;
        RECT 906.3400 1496.6800 909.3400 1497.1600 ;
        RECT 906.3400 1491.2400 909.3400 1491.7200 ;
        RECT 906.3400 1480.3600 909.3400 1480.8400 ;
        RECT 906.3400 1485.8000 909.3400 1486.2800 ;
        RECT 906.3400 1474.9200 909.3400 1475.4000 ;
        RECT 955.9000 1464.0400 956.9000 1464.5200 ;
        RECT 955.9000 1469.4800 956.9000 1469.9600 ;
        RECT 906.3400 1469.4800 909.3400 1469.9600 ;
        RECT 906.3400 1464.0400 909.3400 1464.5200 ;
        RECT 906.3400 1662.2300 1135.3400 1665.2300 ;
        RECT 906.3400 1457.1300 1135.3400 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 1227.4900 1091.9000 1435.5900 ;
        RECT 1045.9000 1227.4900 1046.9000 1435.5900 ;
        RECT 1000.9000 1227.4900 1001.9000 1435.5900 ;
        RECT 955.9000 1227.4900 956.9000 1435.5900 ;
        RECT 1132.3400 1227.4900 1135.3400 1435.5900 ;
        RECT 906.3400 1227.4900 909.3400 1435.5900 ;
      LAYER met3 ;
        RECT 1132.3400 1424.8000 1135.3400 1425.2800 ;
        RECT 1132.3400 1430.2400 1135.3400 1430.7200 ;
        RECT 1090.9000 1424.8000 1091.9000 1425.2800 ;
        RECT 1090.9000 1430.2400 1091.9000 1430.7200 ;
        RECT 1132.3400 1408.4800 1135.3400 1408.9600 ;
        RECT 1132.3400 1413.9200 1135.3400 1414.4000 ;
        RECT 1132.3400 1419.3600 1135.3400 1419.8400 ;
        RECT 1132.3400 1403.0400 1135.3400 1403.5200 ;
        RECT 1132.3400 1392.1600 1135.3400 1392.6400 ;
        RECT 1132.3400 1397.6000 1135.3400 1398.0800 ;
        RECT 1090.9000 1408.4800 1091.9000 1408.9600 ;
        RECT 1090.9000 1413.9200 1091.9000 1414.4000 ;
        RECT 1090.9000 1419.3600 1091.9000 1419.8400 ;
        RECT 1090.9000 1392.1600 1091.9000 1392.6400 ;
        RECT 1090.9000 1397.6000 1091.9000 1398.0800 ;
        RECT 1090.9000 1403.0400 1091.9000 1403.5200 ;
        RECT 1045.9000 1424.8000 1046.9000 1425.2800 ;
        RECT 1045.9000 1430.2400 1046.9000 1430.7200 ;
        RECT 1045.9000 1408.4800 1046.9000 1408.9600 ;
        RECT 1045.9000 1413.9200 1046.9000 1414.4000 ;
        RECT 1045.9000 1419.3600 1046.9000 1419.8400 ;
        RECT 1045.9000 1392.1600 1046.9000 1392.6400 ;
        RECT 1045.9000 1397.6000 1046.9000 1398.0800 ;
        RECT 1045.9000 1403.0400 1046.9000 1403.5200 ;
        RECT 1132.3400 1381.2800 1135.3400 1381.7600 ;
        RECT 1132.3400 1386.7200 1135.3400 1387.2000 ;
        RECT 1132.3400 1375.8400 1135.3400 1376.3200 ;
        RECT 1132.3400 1370.4000 1135.3400 1370.8800 ;
        RECT 1132.3400 1364.9600 1135.3400 1365.4400 ;
        RECT 1090.9000 1381.2800 1091.9000 1381.7600 ;
        RECT 1090.9000 1386.7200 1091.9000 1387.2000 ;
        RECT 1090.9000 1364.9600 1091.9000 1365.4400 ;
        RECT 1090.9000 1370.4000 1091.9000 1370.8800 ;
        RECT 1090.9000 1375.8400 1091.9000 1376.3200 ;
        RECT 1132.3400 1348.6400 1135.3400 1349.1200 ;
        RECT 1132.3400 1354.0800 1135.3400 1354.5600 ;
        RECT 1132.3400 1359.5200 1135.3400 1360.0000 ;
        RECT 1132.3400 1343.2000 1135.3400 1343.6800 ;
        RECT 1132.3400 1332.3200 1135.3400 1332.8000 ;
        RECT 1132.3400 1337.7600 1135.3400 1338.2400 ;
        RECT 1090.9000 1348.6400 1091.9000 1349.1200 ;
        RECT 1090.9000 1354.0800 1091.9000 1354.5600 ;
        RECT 1090.9000 1359.5200 1091.9000 1360.0000 ;
        RECT 1090.9000 1332.3200 1091.9000 1332.8000 ;
        RECT 1090.9000 1337.7600 1091.9000 1338.2400 ;
        RECT 1090.9000 1343.2000 1091.9000 1343.6800 ;
        RECT 1045.9000 1381.2800 1046.9000 1381.7600 ;
        RECT 1045.9000 1386.7200 1046.9000 1387.2000 ;
        RECT 1045.9000 1364.9600 1046.9000 1365.4400 ;
        RECT 1045.9000 1370.4000 1046.9000 1370.8800 ;
        RECT 1045.9000 1375.8400 1046.9000 1376.3200 ;
        RECT 1045.9000 1348.6400 1046.9000 1349.1200 ;
        RECT 1045.9000 1354.0800 1046.9000 1354.5600 ;
        RECT 1045.9000 1359.5200 1046.9000 1360.0000 ;
        RECT 1045.9000 1332.3200 1046.9000 1332.8000 ;
        RECT 1045.9000 1337.7600 1046.9000 1338.2400 ;
        RECT 1045.9000 1343.2000 1046.9000 1343.6800 ;
        RECT 1000.9000 1424.8000 1001.9000 1425.2800 ;
        RECT 1000.9000 1430.2400 1001.9000 1430.7200 ;
        RECT 1000.9000 1408.4800 1001.9000 1408.9600 ;
        RECT 1000.9000 1413.9200 1001.9000 1414.4000 ;
        RECT 1000.9000 1419.3600 1001.9000 1419.8400 ;
        RECT 1000.9000 1392.1600 1001.9000 1392.6400 ;
        RECT 1000.9000 1397.6000 1001.9000 1398.0800 ;
        RECT 1000.9000 1403.0400 1001.9000 1403.5200 ;
        RECT 955.9000 1424.8000 956.9000 1425.2800 ;
        RECT 955.9000 1430.2400 956.9000 1430.7200 ;
        RECT 906.3400 1430.2400 909.3400 1430.7200 ;
        RECT 906.3400 1424.8000 909.3400 1425.2800 ;
        RECT 955.9000 1408.4800 956.9000 1408.9600 ;
        RECT 955.9000 1413.9200 956.9000 1414.4000 ;
        RECT 955.9000 1419.3600 956.9000 1419.8400 ;
        RECT 955.9000 1392.1600 956.9000 1392.6400 ;
        RECT 955.9000 1397.6000 956.9000 1398.0800 ;
        RECT 955.9000 1403.0400 956.9000 1403.5200 ;
        RECT 906.3400 1419.3600 909.3400 1419.8400 ;
        RECT 906.3400 1408.4800 909.3400 1408.9600 ;
        RECT 906.3400 1413.9200 909.3400 1414.4000 ;
        RECT 906.3400 1403.0400 909.3400 1403.5200 ;
        RECT 906.3400 1392.1600 909.3400 1392.6400 ;
        RECT 906.3400 1397.6000 909.3400 1398.0800 ;
        RECT 1000.9000 1381.2800 1001.9000 1381.7600 ;
        RECT 1000.9000 1386.7200 1001.9000 1387.2000 ;
        RECT 1000.9000 1364.9600 1001.9000 1365.4400 ;
        RECT 1000.9000 1370.4000 1001.9000 1370.8800 ;
        RECT 1000.9000 1375.8400 1001.9000 1376.3200 ;
        RECT 1000.9000 1348.6400 1001.9000 1349.1200 ;
        RECT 1000.9000 1354.0800 1001.9000 1354.5600 ;
        RECT 1000.9000 1359.5200 1001.9000 1360.0000 ;
        RECT 1000.9000 1332.3200 1001.9000 1332.8000 ;
        RECT 1000.9000 1337.7600 1001.9000 1338.2400 ;
        RECT 1000.9000 1343.2000 1001.9000 1343.6800 ;
        RECT 955.9000 1381.2800 956.9000 1381.7600 ;
        RECT 955.9000 1386.7200 956.9000 1387.2000 ;
        RECT 955.9000 1364.9600 956.9000 1365.4400 ;
        RECT 955.9000 1370.4000 956.9000 1370.8800 ;
        RECT 955.9000 1375.8400 956.9000 1376.3200 ;
        RECT 906.3400 1386.7200 909.3400 1387.2000 ;
        RECT 906.3400 1381.2800 909.3400 1381.7600 ;
        RECT 906.3400 1370.4000 909.3400 1370.8800 ;
        RECT 906.3400 1375.8400 909.3400 1376.3200 ;
        RECT 906.3400 1364.9600 909.3400 1365.4400 ;
        RECT 955.9000 1348.6400 956.9000 1349.1200 ;
        RECT 955.9000 1354.0800 956.9000 1354.5600 ;
        RECT 955.9000 1359.5200 956.9000 1360.0000 ;
        RECT 955.9000 1332.3200 956.9000 1332.8000 ;
        RECT 955.9000 1337.7600 956.9000 1338.2400 ;
        RECT 955.9000 1343.2000 956.9000 1343.6800 ;
        RECT 906.3400 1359.5200 909.3400 1360.0000 ;
        RECT 906.3400 1348.6400 909.3400 1349.1200 ;
        RECT 906.3400 1354.0800 909.3400 1354.5600 ;
        RECT 906.3400 1343.2000 909.3400 1343.6800 ;
        RECT 906.3400 1332.3200 909.3400 1332.8000 ;
        RECT 906.3400 1337.7600 909.3400 1338.2400 ;
        RECT 1132.3400 1321.4400 1135.3400 1321.9200 ;
        RECT 1132.3400 1326.8800 1135.3400 1327.3600 ;
        RECT 1132.3400 1316.0000 1135.3400 1316.4800 ;
        RECT 1132.3400 1310.5600 1135.3400 1311.0400 ;
        RECT 1132.3400 1305.1200 1135.3400 1305.6000 ;
        RECT 1090.9000 1321.4400 1091.9000 1321.9200 ;
        RECT 1090.9000 1326.8800 1091.9000 1327.3600 ;
        RECT 1090.9000 1305.1200 1091.9000 1305.6000 ;
        RECT 1090.9000 1310.5600 1091.9000 1311.0400 ;
        RECT 1090.9000 1316.0000 1091.9000 1316.4800 ;
        RECT 1132.3400 1288.8000 1135.3400 1289.2800 ;
        RECT 1132.3400 1294.2400 1135.3400 1294.7200 ;
        RECT 1132.3400 1299.6800 1135.3400 1300.1600 ;
        RECT 1132.3400 1283.3600 1135.3400 1283.8400 ;
        RECT 1132.3400 1272.4800 1135.3400 1272.9600 ;
        RECT 1132.3400 1277.9200 1135.3400 1278.4000 ;
        RECT 1090.9000 1288.8000 1091.9000 1289.2800 ;
        RECT 1090.9000 1294.2400 1091.9000 1294.7200 ;
        RECT 1090.9000 1299.6800 1091.9000 1300.1600 ;
        RECT 1090.9000 1272.4800 1091.9000 1272.9600 ;
        RECT 1090.9000 1277.9200 1091.9000 1278.4000 ;
        RECT 1090.9000 1283.3600 1091.9000 1283.8400 ;
        RECT 1045.9000 1321.4400 1046.9000 1321.9200 ;
        RECT 1045.9000 1326.8800 1046.9000 1327.3600 ;
        RECT 1045.9000 1305.1200 1046.9000 1305.6000 ;
        RECT 1045.9000 1310.5600 1046.9000 1311.0400 ;
        RECT 1045.9000 1316.0000 1046.9000 1316.4800 ;
        RECT 1045.9000 1288.8000 1046.9000 1289.2800 ;
        RECT 1045.9000 1294.2400 1046.9000 1294.7200 ;
        RECT 1045.9000 1299.6800 1046.9000 1300.1600 ;
        RECT 1045.9000 1272.4800 1046.9000 1272.9600 ;
        RECT 1045.9000 1277.9200 1046.9000 1278.4000 ;
        RECT 1045.9000 1283.3600 1046.9000 1283.8400 ;
        RECT 1132.3400 1261.6000 1135.3400 1262.0800 ;
        RECT 1132.3400 1267.0400 1135.3400 1267.5200 ;
        RECT 1132.3400 1256.1600 1135.3400 1256.6400 ;
        RECT 1132.3400 1250.7200 1135.3400 1251.2000 ;
        RECT 1132.3400 1245.2800 1135.3400 1245.7600 ;
        RECT 1090.9000 1261.6000 1091.9000 1262.0800 ;
        RECT 1090.9000 1267.0400 1091.9000 1267.5200 ;
        RECT 1090.9000 1245.2800 1091.9000 1245.7600 ;
        RECT 1090.9000 1250.7200 1091.9000 1251.2000 ;
        RECT 1090.9000 1256.1600 1091.9000 1256.6400 ;
        RECT 1132.3400 1234.4000 1135.3400 1234.8800 ;
        RECT 1132.3400 1239.8400 1135.3400 1240.3200 ;
        RECT 1090.9000 1234.4000 1091.9000 1234.8800 ;
        RECT 1090.9000 1239.8400 1091.9000 1240.3200 ;
        RECT 1045.9000 1261.6000 1046.9000 1262.0800 ;
        RECT 1045.9000 1267.0400 1046.9000 1267.5200 ;
        RECT 1045.9000 1245.2800 1046.9000 1245.7600 ;
        RECT 1045.9000 1250.7200 1046.9000 1251.2000 ;
        RECT 1045.9000 1256.1600 1046.9000 1256.6400 ;
        RECT 1045.9000 1234.4000 1046.9000 1234.8800 ;
        RECT 1045.9000 1239.8400 1046.9000 1240.3200 ;
        RECT 1000.9000 1321.4400 1001.9000 1321.9200 ;
        RECT 1000.9000 1326.8800 1001.9000 1327.3600 ;
        RECT 1000.9000 1305.1200 1001.9000 1305.6000 ;
        RECT 1000.9000 1310.5600 1001.9000 1311.0400 ;
        RECT 1000.9000 1316.0000 1001.9000 1316.4800 ;
        RECT 1000.9000 1288.8000 1001.9000 1289.2800 ;
        RECT 1000.9000 1294.2400 1001.9000 1294.7200 ;
        RECT 1000.9000 1299.6800 1001.9000 1300.1600 ;
        RECT 1000.9000 1272.4800 1001.9000 1272.9600 ;
        RECT 1000.9000 1277.9200 1001.9000 1278.4000 ;
        RECT 1000.9000 1283.3600 1001.9000 1283.8400 ;
        RECT 955.9000 1321.4400 956.9000 1321.9200 ;
        RECT 955.9000 1326.8800 956.9000 1327.3600 ;
        RECT 955.9000 1305.1200 956.9000 1305.6000 ;
        RECT 955.9000 1310.5600 956.9000 1311.0400 ;
        RECT 955.9000 1316.0000 956.9000 1316.4800 ;
        RECT 906.3400 1326.8800 909.3400 1327.3600 ;
        RECT 906.3400 1321.4400 909.3400 1321.9200 ;
        RECT 906.3400 1310.5600 909.3400 1311.0400 ;
        RECT 906.3400 1316.0000 909.3400 1316.4800 ;
        RECT 906.3400 1305.1200 909.3400 1305.6000 ;
        RECT 955.9000 1288.8000 956.9000 1289.2800 ;
        RECT 955.9000 1294.2400 956.9000 1294.7200 ;
        RECT 955.9000 1299.6800 956.9000 1300.1600 ;
        RECT 955.9000 1272.4800 956.9000 1272.9600 ;
        RECT 955.9000 1277.9200 956.9000 1278.4000 ;
        RECT 955.9000 1283.3600 956.9000 1283.8400 ;
        RECT 906.3400 1299.6800 909.3400 1300.1600 ;
        RECT 906.3400 1288.8000 909.3400 1289.2800 ;
        RECT 906.3400 1294.2400 909.3400 1294.7200 ;
        RECT 906.3400 1283.3600 909.3400 1283.8400 ;
        RECT 906.3400 1272.4800 909.3400 1272.9600 ;
        RECT 906.3400 1277.9200 909.3400 1278.4000 ;
        RECT 1000.9000 1261.6000 1001.9000 1262.0800 ;
        RECT 1000.9000 1267.0400 1001.9000 1267.5200 ;
        RECT 1000.9000 1245.2800 1001.9000 1245.7600 ;
        RECT 1000.9000 1250.7200 1001.9000 1251.2000 ;
        RECT 1000.9000 1256.1600 1001.9000 1256.6400 ;
        RECT 1000.9000 1234.4000 1001.9000 1234.8800 ;
        RECT 1000.9000 1239.8400 1001.9000 1240.3200 ;
        RECT 955.9000 1261.6000 956.9000 1262.0800 ;
        RECT 955.9000 1267.0400 956.9000 1267.5200 ;
        RECT 955.9000 1245.2800 956.9000 1245.7600 ;
        RECT 955.9000 1250.7200 956.9000 1251.2000 ;
        RECT 955.9000 1256.1600 956.9000 1256.6400 ;
        RECT 906.3400 1267.0400 909.3400 1267.5200 ;
        RECT 906.3400 1261.6000 909.3400 1262.0800 ;
        RECT 906.3400 1250.7200 909.3400 1251.2000 ;
        RECT 906.3400 1256.1600 909.3400 1256.6400 ;
        RECT 906.3400 1245.2800 909.3400 1245.7600 ;
        RECT 955.9000 1234.4000 956.9000 1234.8800 ;
        RECT 955.9000 1239.8400 956.9000 1240.3200 ;
        RECT 906.3400 1239.8400 909.3400 1240.3200 ;
        RECT 906.3400 1234.4000 909.3400 1234.8800 ;
        RECT 906.3400 1432.5900 1135.3400 1435.5900 ;
        RECT 906.3400 1227.4900 1135.3400 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 997.8500 1091.9000 1205.9500 ;
        RECT 1045.9000 997.8500 1046.9000 1205.9500 ;
        RECT 1000.9000 997.8500 1001.9000 1205.9500 ;
        RECT 955.9000 997.8500 956.9000 1205.9500 ;
        RECT 1132.3400 997.8500 1135.3400 1205.9500 ;
        RECT 906.3400 997.8500 909.3400 1205.9500 ;
      LAYER met3 ;
        RECT 1132.3400 1195.1600 1135.3400 1195.6400 ;
        RECT 1132.3400 1200.6000 1135.3400 1201.0800 ;
        RECT 1090.9000 1195.1600 1091.9000 1195.6400 ;
        RECT 1090.9000 1200.6000 1091.9000 1201.0800 ;
        RECT 1132.3400 1178.8400 1135.3400 1179.3200 ;
        RECT 1132.3400 1184.2800 1135.3400 1184.7600 ;
        RECT 1132.3400 1189.7200 1135.3400 1190.2000 ;
        RECT 1132.3400 1173.4000 1135.3400 1173.8800 ;
        RECT 1132.3400 1162.5200 1135.3400 1163.0000 ;
        RECT 1132.3400 1167.9600 1135.3400 1168.4400 ;
        RECT 1090.9000 1178.8400 1091.9000 1179.3200 ;
        RECT 1090.9000 1184.2800 1091.9000 1184.7600 ;
        RECT 1090.9000 1189.7200 1091.9000 1190.2000 ;
        RECT 1090.9000 1162.5200 1091.9000 1163.0000 ;
        RECT 1090.9000 1167.9600 1091.9000 1168.4400 ;
        RECT 1090.9000 1173.4000 1091.9000 1173.8800 ;
        RECT 1045.9000 1195.1600 1046.9000 1195.6400 ;
        RECT 1045.9000 1200.6000 1046.9000 1201.0800 ;
        RECT 1045.9000 1178.8400 1046.9000 1179.3200 ;
        RECT 1045.9000 1184.2800 1046.9000 1184.7600 ;
        RECT 1045.9000 1189.7200 1046.9000 1190.2000 ;
        RECT 1045.9000 1162.5200 1046.9000 1163.0000 ;
        RECT 1045.9000 1167.9600 1046.9000 1168.4400 ;
        RECT 1045.9000 1173.4000 1046.9000 1173.8800 ;
        RECT 1132.3400 1151.6400 1135.3400 1152.1200 ;
        RECT 1132.3400 1157.0800 1135.3400 1157.5600 ;
        RECT 1132.3400 1146.2000 1135.3400 1146.6800 ;
        RECT 1132.3400 1140.7600 1135.3400 1141.2400 ;
        RECT 1132.3400 1135.3200 1135.3400 1135.8000 ;
        RECT 1090.9000 1151.6400 1091.9000 1152.1200 ;
        RECT 1090.9000 1157.0800 1091.9000 1157.5600 ;
        RECT 1090.9000 1135.3200 1091.9000 1135.8000 ;
        RECT 1090.9000 1140.7600 1091.9000 1141.2400 ;
        RECT 1090.9000 1146.2000 1091.9000 1146.6800 ;
        RECT 1132.3400 1119.0000 1135.3400 1119.4800 ;
        RECT 1132.3400 1124.4400 1135.3400 1124.9200 ;
        RECT 1132.3400 1129.8800 1135.3400 1130.3600 ;
        RECT 1132.3400 1113.5600 1135.3400 1114.0400 ;
        RECT 1132.3400 1102.6800 1135.3400 1103.1600 ;
        RECT 1132.3400 1108.1200 1135.3400 1108.6000 ;
        RECT 1090.9000 1119.0000 1091.9000 1119.4800 ;
        RECT 1090.9000 1124.4400 1091.9000 1124.9200 ;
        RECT 1090.9000 1129.8800 1091.9000 1130.3600 ;
        RECT 1090.9000 1102.6800 1091.9000 1103.1600 ;
        RECT 1090.9000 1108.1200 1091.9000 1108.6000 ;
        RECT 1090.9000 1113.5600 1091.9000 1114.0400 ;
        RECT 1045.9000 1151.6400 1046.9000 1152.1200 ;
        RECT 1045.9000 1157.0800 1046.9000 1157.5600 ;
        RECT 1045.9000 1135.3200 1046.9000 1135.8000 ;
        RECT 1045.9000 1140.7600 1046.9000 1141.2400 ;
        RECT 1045.9000 1146.2000 1046.9000 1146.6800 ;
        RECT 1045.9000 1119.0000 1046.9000 1119.4800 ;
        RECT 1045.9000 1124.4400 1046.9000 1124.9200 ;
        RECT 1045.9000 1129.8800 1046.9000 1130.3600 ;
        RECT 1045.9000 1102.6800 1046.9000 1103.1600 ;
        RECT 1045.9000 1108.1200 1046.9000 1108.6000 ;
        RECT 1045.9000 1113.5600 1046.9000 1114.0400 ;
        RECT 1000.9000 1195.1600 1001.9000 1195.6400 ;
        RECT 1000.9000 1200.6000 1001.9000 1201.0800 ;
        RECT 1000.9000 1178.8400 1001.9000 1179.3200 ;
        RECT 1000.9000 1184.2800 1001.9000 1184.7600 ;
        RECT 1000.9000 1189.7200 1001.9000 1190.2000 ;
        RECT 1000.9000 1162.5200 1001.9000 1163.0000 ;
        RECT 1000.9000 1167.9600 1001.9000 1168.4400 ;
        RECT 1000.9000 1173.4000 1001.9000 1173.8800 ;
        RECT 955.9000 1195.1600 956.9000 1195.6400 ;
        RECT 955.9000 1200.6000 956.9000 1201.0800 ;
        RECT 906.3400 1200.6000 909.3400 1201.0800 ;
        RECT 906.3400 1195.1600 909.3400 1195.6400 ;
        RECT 955.9000 1178.8400 956.9000 1179.3200 ;
        RECT 955.9000 1184.2800 956.9000 1184.7600 ;
        RECT 955.9000 1189.7200 956.9000 1190.2000 ;
        RECT 955.9000 1162.5200 956.9000 1163.0000 ;
        RECT 955.9000 1167.9600 956.9000 1168.4400 ;
        RECT 955.9000 1173.4000 956.9000 1173.8800 ;
        RECT 906.3400 1189.7200 909.3400 1190.2000 ;
        RECT 906.3400 1178.8400 909.3400 1179.3200 ;
        RECT 906.3400 1184.2800 909.3400 1184.7600 ;
        RECT 906.3400 1173.4000 909.3400 1173.8800 ;
        RECT 906.3400 1162.5200 909.3400 1163.0000 ;
        RECT 906.3400 1167.9600 909.3400 1168.4400 ;
        RECT 1000.9000 1151.6400 1001.9000 1152.1200 ;
        RECT 1000.9000 1157.0800 1001.9000 1157.5600 ;
        RECT 1000.9000 1135.3200 1001.9000 1135.8000 ;
        RECT 1000.9000 1140.7600 1001.9000 1141.2400 ;
        RECT 1000.9000 1146.2000 1001.9000 1146.6800 ;
        RECT 1000.9000 1119.0000 1001.9000 1119.4800 ;
        RECT 1000.9000 1124.4400 1001.9000 1124.9200 ;
        RECT 1000.9000 1129.8800 1001.9000 1130.3600 ;
        RECT 1000.9000 1102.6800 1001.9000 1103.1600 ;
        RECT 1000.9000 1108.1200 1001.9000 1108.6000 ;
        RECT 1000.9000 1113.5600 1001.9000 1114.0400 ;
        RECT 955.9000 1151.6400 956.9000 1152.1200 ;
        RECT 955.9000 1157.0800 956.9000 1157.5600 ;
        RECT 955.9000 1135.3200 956.9000 1135.8000 ;
        RECT 955.9000 1140.7600 956.9000 1141.2400 ;
        RECT 955.9000 1146.2000 956.9000 1146.6800 ;
        RECT 906.3400 1157.0800 909.3400 1157.5600 ;
        RECT 906.3400 1151.6400 909.3400 1152.1200 ;
        RECT 906.3400 1140.7600 909.3400 1141.2400 ;
        RECT 906.3400 1146.2000 909.3400 1146.6800 ;
        RECT 906.3400 1135.3200 909.3400 1135.8000 ;
        RECT 955.9000 1119.0000 956.9000 1119.4800 ;
        RECT 955.9000 1124.4400 956.9000 1124.9200 ;
        RECT 955.9000 1129.8800 956.9000 1130.3600 ;
        RECT 955.9000 1102.6800 956.9000 1103.1600 ;
        RECT 955.9000 1108.1200 956.9000 1108.6000 ;
        RECT 955.9000 1113.5600 956.9000 1114.0400 ;
        RECT 906.3400 1129.8800 909.3400 1130.3600 ;
        RECT 906.3400 1119.0000 909.3400 1119.4800 ;
        RECT 906.3400 1124.4400 909.3400 1124.9200 ;
        RECT 906.3400 1113.5600 909.3400 1114.0400 ;
        RECT 906.3400 1102.6800 909.3400 1103.1600 ;
        RECT 906.3400 1108.1200 909.3400 1108.6000 ;
        RECT 1132.3400 1091.8000 1135.3400 1092.2800 ;
        RECT 1132.3400 1097.2400 1135.3400 1097.7200 ;
        RECT 1132.3400 1086.3600 1135.3400 1086.8400 ;
        RECT 1132.3400 1080.9200 1135.3400 1081.4000 ;
        RECT 1132.3400 1075.4800 1135.3400 1075.9600 ;
        RECT 1090.9000 1091.8000 1091.9000 1092.2800 ;
        RECT 1090.9000 1097.2400 1091.9000 1097.7200 ;
        RECT 1090.9000 1075.4800 1091.9000 1075.9600 ;
        RECT 1090.9000 1080.9200 1091.9000 1081.4000 ;
        RECT 1090.9000 1086.3600 1091.9000 1086.8400 ;
        RECT 1132.3400 1059.1600 1135.3400 1059.6400 ;
        RECT 1132.3400 1064.6000 1135.3400 1065.0800 ;
        RECT 1132.3400 1070.0400 1135.3400 1070.5200 ;
        RECT 1132.3400 1053.7200 1135.3400 1054.2000 ;
        RECT 1132.3400 1042.8400 1135.3400 1043.3200 ;
        RECT 1132.3400 1048.2800 1135.3400 1048.7600 ;
        RECT 1090.9000 1059.1600 1091.9000 1059.6400 ;
        RECT 1090.9000 1064.6000 1091.9000 1065.0800 ;
        RECT 1090.9000 1070.0400 1091.9000 1070.5200 ;
        RECT 1090.9000 1042.8400 1091.9000 1043.3200 ;
        RECT 1090.9000 1048.2800 1091.9000 1048.7600 ;
        RECT 1090.9000 1053.7200 1091.9000 1054.2000 ;
        RECT 1045.9000 1091.8000 1046.9000 1092.2800 ;
        RECT 1045.9000 1097.2400 1046.9000 1097.7200 ;
        RECT 1045.9000 1075.4800 1046.9000 1075.9600 ;
        RECT 1045.9000 1080.9200 1046.9000 1081.4000 ;
        RECT 1045.9000 1086.3600 1046.9000 1086.8400 ;
        RECT 1045.9000 1059.1600 1046.9000 1059.6400 ;
        RECT 1045.9000 1064.6000 1046.9000 1065.0800 ;
        RECT 1045.9000 1070.0400 1046.9000 1070.5200 ;
        RECT 1045.9000 1042.8400 1046.9000 1043.3200 ;
        RECT 1045.9000 1048.2800 1046.9000 1048.7600 ;
        RECT 1045.9000 1053.7200 1046.9000 1054.2000 ;
        RECT 1132.3400 1031.9600 1135.3400 1032.4400 ;
        RECT 1132.3400 1037.4000 1135.3400 1037.8800 ;
        RECT 1132.3400 1026.5200 1135.3400 1027.0000 ;
        RECT 1132.3400 1021.0800 1135.3400 1021.5600 ;
        RECT 1132.3400 1015.6400 1135.3400 1016.1200 ;
        RECT 1090.9000 1031.9600 1091.9000 1032.4400 ;
        RECT 1090.9000 1037.4000 1091.9000 1037.8800 ;
        RECT 1090.9000 1015.6400 1091.9000 1016.1200 ;
        RECT 1090.9000 1021.0800 1091.9000 1021.5600 ;
        RECT 1090.9000 1026.5200 1091.9000 1027.0000 ;
        RECT 1132.3400 1004.7600 1135.3400 1005.2400 ;
        RECT 1132.3400 1010.2000 1135.3400 1010.6800 ;
        RECT 1090.9000 1004.7600 1091.9000 1005.2400 ;
        RECT 1090.9000 1010.2000 1091.9000 1010.6800 ;
        RECT 1045.9000 1031.9600 1046.9000 1032.4400 ;
        RECT 1045.9000 1037.4000 1046.9000 1037.8800 ;
        RECT 1045.9000 1015.6400 1046.9000 1016.1200 ;
        RECT 1045.9000 1021.0800 1046.9000 1021.5600 ;
        RECT 1045.9000 1026.5200 1046.9000 1027.0000 ;
        RECT 1045.9000 1004.7600 1046.9000 1005.2400 ;
        RECT 1045.9000 1010.2000 1046.9000 1010.6800 ;
        RECT 1000.9000 1091.8000 1001.9000 1092.2800 ;
        RECT 1000.9000 1097.2400 1001.9000 1097.7200 ;
        RECT 1000.9000 1075.4800 1001.9000 1075.9600 ;
        RECT 1000.9000 1080.9200 1001.9000 1081.4000 ;
        RECT 1000.9000 1086.3600 1001.9000 1086.8400 ;
        RECT 1000.9000 1059.1600 1001.9000 1059.6400 ;
        RECT 1000.9000 1064.6000 1001.9000 1065.0800 ;
        RECT 1000.9000 1070.0400 1001.9000 1070.5200 ;
        RECT 1000.9000 1042.8400 1001.9000 1043.3200 ;
        RECT 1000.9000 1048.2800 1001.9000 1048.7600 ;
        RECT 1000.9000 1053.7200 1001.9000 1054.2000 ;
        RECT 955.9000 1091.8000 956.9000 1092.2800 ;
        RECT 955.9000 1097.2400 956.9000 1097.7200 ;
        RECT 955.9000 1075.4800 956.9000 1075.9600 ;
        RECT 955.9000 1080.9200 956.9000 1081.4000 ;
        RECT 955.9000 1086.3600 956.9000 1086.8400 ;
        RECT 906.3400 1097.2400 909.3400 1097.7200 ;
        RECT 906.3400 1091.8000 909.3400 1092.2800 ;
        RECT 906.3400 1080.9200 909.3400 1081.4000 ;
        RECT 906.3400 1086.3600 909.3400 1086.8400 ;
        RECT 906.3400 1075.4800 909.3400 1075.9600 ;
        RECT 955.9000 1059.1600 956.9000 1059.6400 ;
        RECT 955.9000 1064.6000 956.9000 1065.0800 ;
        RECT 955.9000 1070.0400 956.9000 1070.5200 ;
        RECT 955.9000 1042.8400 956.9000 1043.3200 ;
        RECT 955.9000 1048.2800 956.9000 1048.7600 ;
        RECT 955.9000 1053.7200 956.9000 1054.2000 ;
        RECT 906.3400 1070.0400 909.3400 1070.5200 ;
        RECT 906.3400 1059.1600 909.3400 1059.6400 ;
        RECT 906.3400 1064.6000 909.3400 1065.0800 ;
        RECT 906.3400 1053.7200 909.3400 1054.2000 ;
        RECT 906.3400 1042.8400 909.3400 1043.3200 ;
        RECT 906.3400 1048.2800 909.3400 1048.7600 ;
        RECT 1000.9000 1031.9600 1001.9000 1032.4400 ;
        RECT 1000.9000 1037.4000 1001.9000 1037.8800 ;
        RECT 1000.9000 1015.6400 1001.9000 1016.1200 ;
        RECT 1000.9000 1021.0800 1001.9000 1021.5600 ;
        RECT 1000.9000 1026.5200 1001.9000 1027.0000 ;
        RECT 1000.9000 1004.7600 1001.9000 1005.2400 ;
        RECT 1000.9000 1010.2000 1001.9000 1010.6800 ;
        RECT 955.9000 1031.9600 956.9000 1032.4400 ;
        RECT 955.9000 1037.4000 956.9000 1037.8800 ;
        RECT 955.9000 1015.6400 956.9000 1016.1200 ;
        RECT 955.9000 1021.0800 956.9000 1021.5600 ;
        RECT 955.9000 1026.5200 956.9000 1027.0000 ;
        RECT 906.3400 1037.4000 909.3400 1037.8800 ;
        RECT 906.3400 1031.9600 909.3400 1032.4400 ;
        RECT 906.3400 1021.0800 909.3400 1021.5600 ;
        RECT 906.3400 1026.5200 909.3400 1027.0000 ;
        RECT 906.3400 1015.6400 909.3400 1016.1200 ;
        RECT 955.9000 1004.7600 956.9000 1005.2400 ;
        RECT 955.9000 1010.2000 956.9000 1010.6800 ;
        RECT 906.3400 1010.2000 909.3400 1010.6800 ;
        RECT 906.3400 1004.7600 909.3400 1005.2400 ;
        RECT 906.3400 1202.9500 1135.3400 1205.9500 ;
        RECT 906.3400 997.8500 1135.3400 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1090.9000 768.2100 1091.9000 976.3100 ;
        RECT 1045.9000 768.2100 1046.9000 976.3100 ;
        RECT 1000.9000 768.2100 1001.9000 976.3100 ;
        RECT 955.9000 768.2100 956.9000 976.3100 ;
        RECT 1132.3400 768.2100 1135.3400 976.3100 ;
        RECT 906.3400 768.2100 909.3400 976.3100 ;
      LAYER met3 ;
        RECT 1132.3400 965.5200 1135.3400 966.0000 ;
        RECT 1132.3400 970.9600 1135.3400 971.4400 ;
        RECT 1090.9000 965.5200 1091.9000 966.0000 ;
        RECT 1090.9000 970.9600 1091.9000 971.4400 ;
        RECT 1132.3400 949.2000 1135.3400 949.6800 ;
        RECT 1132.3400 954.6400 1135.3400 955.1200 ;
        RECT 1132.3400 960.0800 1135.3400 960.5600 ;
        RECT 1132.3400 943.7600 1135.3400 944.2400 ;
        RECT 1132.3400 932.8800 1135.3400 933.3600 ;
        RECT 1132.3400 938.3200 1135.3400 938.8000 ;
        RECT 1090.9000 949.2000 1091.9000 949.6800 ;
        RECT 1090.9000 954.6400 1091.9000 955.1200 ;
        RECT 1090.9000 960.0800 1091.9000 960.5600 ;
        RECT 1090.9000 932.8800 1091.9000 933.3600 ;
        RECT 1090.9000 938.3200 1091.9000 938.8000 ;
        RECT 1090.9000 943.7600 1091.9000 944.2400 ;
        RECT 1045.9000 965.5200 1046.9000 966.0000 ;
        RECT 1045.9000 970.9600 1046.9000 971.4400 ;
        RECT 1045.9000 949.2000 1046.9000 949.6800 ;
        RECT 1045.9000 954.6400 1046.9000 955.1200 ;
        RECT 1045.9000 960.0800 1046.9000 960.5600 ;
        RECT 1045.9000 932.8800 1046.9000 933.3600 ;
        RECT 1045.9000 938.3200 1046.9000 938.8000 ;
        RECT 1045.9000 943.7600 1046.9000 944.2400 ;
        RECT 1132.3400 922.0000 1135.3400 922.4800 ;
        RECT 1132.3400 927.4400 1135.3400 927.9200 ;
        RECT 1132.3400 916.5600 1135.3400 917.0400 ;
        RECT 1132.3400 911.1200 1135.3400 911.6000 ;
        RECT 1132.3400 905.6800 1135.3400 906.1600 ;
        RECT 1090.9000 922.0000 1091.9000 922.4800 ;
        RECT 1090.9000 927.4400 1091.9000 927.9200 ;
        RECT 1090.9000 905.6800 1091.9000 906.1600 ;
        RECT 1090.9000 911.1200 1091.9000 911.6000 ;
        RECT 1090.9000 916.5600 1091.9000 917.0400 ;
        RECT 1132.3400 889.3600 1135.3400 889.8400 ;
        RECT 1132.3400 894.8000 1135.3400 895.2800 ;
        RECT 1132.3400 900.2400 1135.3400 900.7200 ;
        RECT 1132.3400 883.9200 1135.3400 884.4000 ;
        RECT 1132.3400 873.0400 1135.3400 873.5200 ;
        RECT 1132.3400 878.4800 1135.3400 878.9600 ;
        RECT 1090.9000 889.3600 1091.9000 889.8400 ;
        RECT 1090.9000 894.8000 1091.9000 895.2800 ;
        RECT 1090.9000 900.2400 1091.9000 900.7200 ;
        RECT 1090.9000 873.0400 1091.9000 873.5200 ;
        RECT 1090.9000 878.4800 1091.9000 878.9600 ;
        RECT 1090.9000 883.9200 1091.9000 884.4000 ;
        RECT 1045.9000 922.0000 1046.9000 922.4800 ;
        RECT 1045.9000 927.4400 1046.9000 927.9200 ;
        RECT 1045.9000 905.6800 1046.9000 906.1600 ;
        RECT 1045.9000 911.1200 1046.9000 911.6000 ;
        RECT 1045.9000 916.5600 1046.9000 917.0400 ;
        RECT 1045.9000 889.3600 1046.9000 889.8400 ;
        RECT 1045.9000 894.8000 1046.9000 895.2800 ;
        RECT 1045.9000 900.2400 1046.9000 900.7200 ;
        RECT 1045.9000 873.0400 1046.9000 873.5200 ;
        RECT 1045.9000 878.4800 1046.9000 878.9600 ;
        RECT 1045.9000 883.9200 1046.9000 884.4000 ;
        RECT 1000.9000 965.5200 1001.9000 966.0000 ;
        RECT 1000.9000 970.9600 1001.9000 971.4400 ;
        RECT 1000.9000 949.2000 1001.9000 949.6800 ;
        RECT 1000.9000 954.6400 1001.9000 955.1200 ;
        RECT 1000.9000 960.0800 1001.9000 960.5600 ;
        RECT 1000.9000 932.8800 1001.9000 933.3600 ;
        RECT 1000.9000 938.3200 1001.9000 938.8000 ;
        RECT 1000.9000 943.7600 1001.9000 944.2400 ;
        RECT 955.9000 965.5200 956.9000 966.0000 ;
        RECT 955.9000 970.9600 956.9000 971.4400 ;
        RECT 906.3400 970.9600 909.3400 971.4400 ;
        RECT 906.3400 965.5200 909.3400 966.0000 ;
        RECT 955.9000 949.2000 956.9000 949.6800 ;
        RECT 955.9000 954.6400 956.9000 955.1200 ;
        RECT 955.9000 960.0800 956.9000 960.5600 ;
        RECT 955.9000 932.8800 956.9000 933.3600 ;
        RECT 955.9000 938.3200 956.9000 938.8000 ;
        RECT 955.9000 943.7600 956.9000 944.2400 ;
        RECT 906.3400 960.0800 909.3400 960.5600 ;
        RECT 906.3400 949.2000 909.3400 949.6800 ;
        RECT 906.3400 954.6400 909.3400 955.1200 ;
        RECT 906.3400 943.7600 909.3400 944.2400 ;
        RECT 906.3400 932.8800 909.3400 933.3600 ;
        RECT 906.3400 938.3200 909.3400 938.8000 ;
        RECT 1000.9000 922.0000 1001.9000 922.4800 ;
        RECT 1000.9000 927.4400 1001.9000 927.9200 ;
        RECT 1000.9000 905.6800 1001.9000 906.1600 ;
        RECT 1000.9000 911.1200 1001.9000 911.6000 ;
        RECT 1000.9000 916.5600 1001.9000 917.0400 ;
        RECT 1000.9000 889.3600 1001.9000 889.8400 ;
        RECT 1000.9000 894.8000 1001.9000 895.2800 ;
        RECT 1000.9000 900.2400 1001.9000 900.7200 ;
        RECT 1000.9000 873.0400 1001.9000 873.5200 ;
        RECT 1000.9000 878.4800 1001.9000 878.9600 ;
        RECT 1000.9000 883.9200 1001.9000 884.4000 ;
        RECT 955.9000 922.0000 956.9000 922.4800 ;
        RECT 955.9000 927.4400 956.9000 927.9200 ;
        RECT 955.9000 905.6800 956.9000 906.1600 ;
        RECT 955.9000 911.1200 956.9000 911.6000 ;
        RECT 955.9000 916.5600 956.9000 917.0400 ;
        RECT 906.3400 927.4400 909.3400 927.9200 ;
        RECT 906.3400 922.0000 909.3400 922.4800 ;
        RECT 906.3400 911.1200 909.3400 911.6000 ;
        RECT 906.3400 916.5600 909.3400 917.0400 ;
        RECT 906.3400 905.6800 909.3400 906.1600 ;
        RECT 955.9000 889.3600 956.9000 889.8400 ;
        RECT 955.9000 894.8000 956.9000 895.2800 ;
        RECT 955.9000 900.2400 956.9000 900.7200 ;
        RECT 955.9000 873.0400 956.9000 873.5200 ;
        RECT 955.9000 878.4800 956.9000 878.9600 ;
        RECT 955.9000 883.9200 956.9000 884.4000 ;
        RECT 906.3400 900.2400 909.3400 900.7200 ;
        RECT 906.3400 889.3600 909.3400 889.8400 ;
        RECT 906.3400 894.8000 909.3400 895.2800 ;
        RECT 906.3400 883.9200 909.3400 884.4000 ;
        RECT 906.3400 873.0400 909.3400 873.5200 ;
        RECT 906.3400 878.4800 909.3400 878.9600 ;
        RECT 1132.3400 862.1600 1135.3400 862.6400 ;
        RECT 1132.3400 867.6000 1135.3400 868.0800 ;
        RECT 1132.3400 856.7200 1135.3400 857.2000 ;
        RECT 1132.3400 851.2800 1135.3400 851.7600 ;
        RECT 1132.3400 845.8400 1135.3400 846.3200 ;
        RECT 1090.9000 862.1600 1091.9000 862.6400 ;
        RECT 1090.9000 867.6000 1091.9000 868.0800 ;
        RECT 1090.9000 845.8400 1091.9000 846.3200 ;
        RECT 1090.9000 851.2800 1091.9000 851.7600 ;
        RECT 1090.9000 856.7200 1091.9000 857.2000 ;
        RECT 1132.3400 829.5200 1135.3400 830.0000 ;
        RECT 1132.3400 834.9600 1135.3400 835.4400 ;
        RECT 1132.3400 840.4000 1135.3400 840.8800 ;
        RECT 1132.3400 824.0800 1135.3400 824.5600 ;
        RECT 1132.3400 813.2000 1135.3400 813.6800 ;
        RECT 1132.3400 818.6400 1135.3400 819.1200 ;
        RECT 1090.9000 829.5200 1091.9000 830.0000 ;
        RECT 1090.9000 834.9600 1091.9000 835.4400 ;
        RECT 1090.9000 840.4000 1091.9000 840.8800 ;
        RECT 1090.9000 813.2000 1091.9000 813.6800 ;
        RECT 1090.9000 818.6400 1091.9000 819.1200 ;
        RECT 1090.9000 824.0800 1091.9000 824.5600 ;
        RECT 1045.9000 862.1600 1046.9000 862.6400 ;
        RECT 1045.9000 867.6000 1046.9000 868.0800 ;
        RECT 1045.9000 845.8400 1046.9000 846.3200 ;
        RECT 1045.9000 851.2800 1046.9000 851.7600 ;
        RECT 1045.9000 856.7200 1046.9000 857.2000 ;
        RECT 1045.9000 829.5200 1046.9000 830.0000 ;
        RECT 1045.9000 834.9600 1046.9000 835.4400 ;
        RECT 1045.9000 840.4000 1046.9000 840.8800 ;
        RECT 1045.9000 813.2000 1046.9000 813.6800 ;
        RECT 1045.9000 818.6400 1046.9000 819.1200 ;
        RECT 1045.9000 824.0800 1046.9000 824.5600 ;
        RECT 1132.3400 802.3200 1135.3400 802.8000 ;
        RECT 1132.3400 807.7600 1135.3400 808.2400 ;
        RECT 1132.3400 796.8800 1135.3400 797.3600 ;
        RECT 1132.3400 791.4400 1135.3400 791.9200 ;
        RECT 1132.3400 786.0000 1135.3400 786.4800 ;
        RECT 1090.9000 802.3200 1091.9000 802.8000 ;
        RECT 1090.9000 807.7600 1091.9000 808.2400 ;
        RECT 1090.9000 786.0000 1091.9000 786.4800 ;
        RECT 1090.9000 791.4400 1091.9000 791.9200 ;
        RECT 1090.9000 796.8800 1091.9000 797.3600 ;
        RECT 1132.3400 775.1200 1135.3400 775.6000 ;
        RECT 1132.3400 780.5600 1135.3400 781.0400 ;
        RECT 1090.9000 775.1200 1091.9000 775.6000 ;
        RECT 1090.9000 780.5600 1091.9000 781.0400 ;
        RECT 1045.9000 802.3200 1046.9000 802.8000 ;
        RECT 1045.9000 807.7600 1046.9000 808.2400 ;
        RECT 1045.9000 786.0000 1046.9000 786.4800 ;
        RECT 1045.9000 791.4400 1046.9000 791.9200 ;
        RECT 1045.9000 796.8800 1046.9000 797.3600 ;
        RECT 1045.9000 775.1200 1046.9000 775.6000 ;
        RECT 1045.9000 780.5600 1046.9000 781.0400 ;
        RECT 1000.9000 862.1600 1001.9000 862.6400 ;
        RECT 1000.9000 867.6000 1001.9000 868.0800 ;
        RECT 1000.9000 845.8400 1001.9000 846.3200 ;
        RECT 1000.9000 851.2800 1001.9000 851.7600 ;
        RECT 1000.9000 856.7200 1001.9000 857.2000 ;
        RECT 1000.9000 829.5200 1001.9000 830.0000 ;
        RECT 1000.9000 834.9600 1001.9000 835.4400 ;
        RECT 1000.9000 840.4000 1001.9000 840.8800 ;
        RECT 1000.9000 813.2000 1001.9000 813.6800 ;
        RECT 1000.9000 818.6400 1001.9000 819.1200 ;
        RECT 1000.9000 824.0800 1001.9000 824.5600 ;
        RECT 955.9000 862.1600 956.9000 862.6400 ;
        RECT 955.9000 867.6000 956.9000 868.0800 ;
        RECT 955.9000 845.8400 956.9000 846.3200 ;
        RECT 955.9000 851.2800 956.9000 851.7600 ;
        RECT 955.9000 856.7200 956.9000 857.2000 ;
        RECT 906.3400 867.6000 909.3400 868.0800 ;
        RECT 906.3400 862.1600 909.3400 862.6400 ;
        RECT 906.3400 851.2800 909.3400 851.7600 ;
        RECT 906.3400 856.7200 909.3400 857.2000 ;
        RECT 906.3400 845.8400 909.3400 846.3200 ;
        RECT 955.9000 829.5200 956.9000 830.0000 ;
        RECT 955.9000 834.9600 956.9000 835.4400 ;
        RECT 955.9000 840.4000 956.9000 840.8800 ;
        RECT 955.9000 813.2000 956.9000 813.6800 ;
        RECT 955.9000 818.6400 956.9000 819.1200 ;
        RECT 955.9000 824.0800 956.9000 824.5600 ;
        RECT 906.3400 840.4000 909.3400 840.8800 ;
        RECT 906.3400 829.5200 909.3400 830.0000 ;
        RECT 906.3400 834.9600 909.3400 835.4400 ;
        RECT 906.3400 824.0800 909.3400 824.5600 ;
        RECT 906.3400 813.2000 909.3400 813.6800 ;
        RECT 906.3400 818.6400 909.3400 819.1200 ;
        RECT 1000.9000 802.3200 1001.9000 802.8000 ;
        RECT 1000.9000 807.7600 1001.9000 808.2400 ;
        RECT 1000.9000 786.0000 1001.9000 786.4800 ;
        RECT 1000.9000 791.4400 1001.9000 791.9200 ;
        RECT 1000.9000 796.8800 1001.9000 797.3600 ;
        RECT 1000.9000 775.1200 1001.9000 775.6000 ;
        RECT 1000.9000 780.5600 1001.9000 781.0400 ;
        RECT 955.9000 802.3200 956.9000 802.8000 ;
        RECT 955.9000 807.7600 956.9000 808.2400 ;
        RECT 955.9000 786.0000 956.9000 786.4800 ;
        RECT 955.9000 791.4400 956.9000 791.9200 ;
        RECT 955.9000 796.8800 956.9000 797.3600 ;
        RECT 906.3400 807.7600 909.3400 808.2400 ;
        RECT 906.3400 802.3200 909.3400 802.8000 ;
        RECT 906.3400 791.4400 909.3400 791.9200 ;
        RECT 906.3400 796.8800 909.3400 797.3600 ;
        RECT 906.3400 786.0000 909.3400 786.4800 ;
        RECT 955.9000 775.1200 956.9000 775.6000 ;
        RECT 955.9000 780.5600 956.9000 781.0400 ;
        RECT 906.3400 780.5600 909.3400 781.0400 ;
        RECT 906.3400 775.1200 909.3400 775.6000 ;
        RECT 906.3400 973.3100 1135.3400 976.3100 ;
        RECT 906.3400 768.2100 1135.3400 771.2100 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1156.4600 2833.6100 1158.4600 2854.5400 ;
        RECT 1353.5600 2833.6100 1355.5600 2854.5400 ;
      LAYER met3 ;
        RECT 1353.5600 2850.0400 1355.5600 2850.5200 ;
        RECT 1156.4600 2850.0400 1158.4600 2850.5200 ;
        RECT 1353.5600 2839.1600 1355.5600 2839.6400 ;
        RECT 1156.4600 2839.1600 1158.4600 2839.6400 ;
        RECT 1353.5600 2844.6000 1355.5600 2845.0800 ;
        RECT 1156.4600 2844.6000 1158.4600 2845.0800 ;
        RECT 1156.4600 2852.5400 1355.5600 2854.5400 ;
        RECT 1156.4600 2833.6100 1355.5600 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 538.5700 1342.6200 746.6700 ;
        RECT 1296.0200 538.5700 1297.6200 746.6700 ;
        RECT 1251.0200 538.5700 1252.6200 746.6700 ;
        RECT 1206.0200 538.5700 1207.6200 746.6700 ;
        RECT 1352.5600 538.5700 1355.5600 746.6700 ;
        RECT 1156.4600 538.5700 1159.4600 746.6700 ;
      LAYER met3 ;
        RECT 1352.5600 741.3200 1355.5600 741.8000 ;
        RECT 1341.0200 741.3200 1342.6200 741.8000 ;
        RECT 1352.5600 730.4400 1355.5600 730.9200 ;
        RECT 1352.5600 735.8800 1355.5600 736.3600 ;
        RECT 1341.0200 730.4400 1342.6200 730.9200 ;
        RECT 1341.0200 735.8800 1342.6200 736.3600 ;
        RECT 1352.5600 714.1200 1355.5600 714.6000 ;
        RECT 1352.5600 719.5600 1355.5600 720.0400 ;
        RECT 1341.0200 714.1200 1342.6200 714.6000 ;
        RECT 1341.0200 719.5600 1342.6200 720.0400 ;
        RECT 1352.5600 703.2400 1355.5600 703.7200 ;
        RECT 1352.5600 708.6800 1355.5600 709.1600 ;
        RECT 1341.0200 703.2400 1342.6200 703.7200 ;
        RECT 1341.0200 708.6800 1342.6200 709.1600 ;
        RECT 1352.5600 725.0000 1355.5600 725.4800 ;
        RECT 1341.0200 725.0000 1342.6200 725.4800 ;
        RECT 1296.0200 730.4400 1297.6200 730.9200 ;
        RECT 1296.0200 735.8800 1297.6200 736.3600 ;
        RECT 1296.0200 741.3200 1297.6200 741.8000 ;
        RECT 1296.0200 714.1200 1297.6200 714.6000 ;
        RECT 1296.0200 719.5600 1297.6200 720.0400 ;
        RECT 1296.0200 708.6800 1297.6200 709.1600 ;
        RECT 1296.0200 703.2400 1297.6200 703.7200 ;
        RECT 1296.0200 725.0000 1297.6200 725.4800 ;
        RECT 1352.5600 686.9200 1355.5600 687.4000 ;
        RECT 1352.5600 692.3600 1355.5600 692.8400 ;
        RECT 1341.0200 686.9200 1342.6200 687.4000 ;
        RECT 1341.0200 692.3600 1342.6200 692.8400 ;
        RECT 1352.5600 670.6000 1355.5600 671.0800 ;
        RECT 1352.5600 676.0400 1355.5600 676.5200 ;
        RECT 1352.5600 681.4800 1355.5600 681.9600 ;
        RECT 1341.0200 670.6000 1342.6200 671.0800 ;
        RECT 1341.0200 676.0400 1342.6200 676.5200 ;
        RECT 1341.0200 681.4800 1342.6200 681.9600 ;
        RECT 1352.5600 659.7200 1355.5600 660.2000 ;
        RECT 1352.5600 665.1600 1355.5600 665.6400 ;
        RECT 1341.0200 659.7200 1342.6200 660.2000 ;
        RECT 1341.0200 665.1600 1342.6200 665.6400 ;
        RECT 1352.5600 643.4000 1355.5600 643.8800 ;
        RECT 1352.5600 648.8400 1355.5600 649.3200 ;
        RECT 1352.5600 654.2800 1355.5600 654.7600 ;
        RECT 1341.0200 643.4000 1342.6200 643.8800 ;
        RECT 1341.0200 648.8400 1342.6200 649.3200 ;
        RECT 1341.0200 654.2800 1342.6200 654.7600 ;
        RECT 1296.0200 686.9200 1297.6200 687.4000 ;
        RECT 1296.0200 692.3600 1297.6200 692.8400 ;
        RECT 1296.0200 670.6000 1297.6200 671.0800 ;
        RECT 1296.0200 676.0400 1297.6200 676.5200 ;
        RECT 1296.0200 681.4800 1297.6200 681.9600 ;
        RECT 1296.0200 659.7200 1297.6200 660.2000 ;
        RECT 1296.0200 665.1600 1297.6200 665.6400 ;
        RECT 1296.0200 643.4000 1297.6200 643.8800 ;
        RECT 1296.0200 648.8400 1297.6200 649.3200 ;
        RECT 1296.0200 654.2800 1297.6200 654.7600 ;
        RECT 1352.5600 697.8000 1355.5600 698.2800 ;
        RECT 1296.0200 697.8000 1297.6200 698.2800 ;
        RECT 1341.0200 697.8000 1342.6200 698.2800 ;
        RECT 1251.0200 730.4400 1252.6200 730.9200 ;
        RECT 1251.0200 735.8800 1252.6200 736.3600 ;
        RECT 1251.0200 741.3200 1252.6200 741.8000 ;
        RECT 1206.0200 730.4400 1207.6200 730.9200 ;
        RECT 1206.0200 735.8800 1207.6200 736.3600 ;
        RECT 1206.0200 741.3200 1207.6200 741.8000 ;
        RECT 1251.0200 714.1200 1252.6200 714.6000 ;
        RECT 1251.0200 719.5600 1252.6200 720.0400 ;
        RECT 1251.0200 703.2400 1252.6200 703.7200 ;
        RECT 1251.0200 708.6800 1252.6200 709.1600 ;
        RECT 1206.0200 714.1200 1207.6200 714.6000 ;
        RECT 1206.0200 719.5600 1207.6200 720.0400 ;
        RECT 1206.0200 703.2400 1207.6200 703.7200 ;
        RECT 1206.0200 708.6800 1207.6200 709.1600 ;
        RECT 1206.0200 725.0000 1207.6200 725.4800 ;
        RECT 1251.0200 725.0000 1252.6200 725.4800 ;
        RECT 1156.4600 741.3200 1159.4600 741.8000 ;
        RECT 1156.4600 735.8800 1159.4600 736.3600 ;
        RECT 1156.4600 730.4400 1159.4600 730.9200 ;
        RECT 1156.4600 719.5600 1159.4600 720.0400 ;
        RECT 1156.4600 714.1200 1159.4600 714.6000 ;
        RECT 1156.4600 708.6800 1159.4600 709.1600 ;
        RECT 1156.4600 703.2400 1159.4600 703.7200 ;
        RECT 1156.4600 725.0000 1159.4600 725.4800 ;
        RECT 1251.0200 686.9200 1252.6200 687.4000 ;
        RECT 1251.0200 692.3600 1252.6200 692.8400 ;
        RECT 1251.0200 670.6000 1252.6200 671.0800 ;
        RECT 1251.0200 676.0400 1252.6200 676.5200 ;
        RECT 1251.0200 681.4800 1252.6200 681.9600 ;
        RECT 1206.0200 686.9200 1207.6200 687.4000 ;
        RECT 1206.0200 692.3600 1207.6200 692.8400 ;
        RECT 1206.0200 670.6000 1207.6200 671.0800 ;
        RECT 1206.0200 676.0400 1207.6200 676.5200 ;
        RECT 1206.0200 681.4800 1207.6200 681.9600 ;
        RECT 1251.0200 659.7200 1252.6200 660.2000 ;
        RECT 1251.0200 665.1600 1252.6200 665.6400 ;
        RECT 1251.0200 643.4000 1252.6200 643.8800 ;
        RECT 1251.0200 648.8400 1252.6200 649.3200 ;
        RECT 1251.0200 654.2800 1252.6200 654.7600 ;
        RECT 1206.0200 659.7200 1207.6200 660.2000 ;
        RECT 1206.0200 665.1600 1207.6200 665.6400 ;
        RECT 1206.0200 643.4000 1207.6200 643.8800 ;
        RECT 1206.0200 648.8400 1207.6200 649.3200 ;
        RECT 1206.0200 654.2800 1207.6200 654.7600 ;
        RECT 1156.4600 686.9200 1159.4600 687.4000 ;
        RECT 1156.4600 692.3600 1159.4600 692.8400 ;
        RECT 1156.4600 676.0400 1159.4600 676.5200 ;
        RECT 1156.4600 670.6000 1159.4600 671.0800 ;
        RECT 1156.4600 681.4800 1159.4600 681.9600 ;
        RECT 1156.4600 659.7200 1159.4600 660.2000 ;
        RECT 1156.4600 665.1600 1159.4600 665.6400 ;
        RECT 1156.4600 648.8400 1159.4600 649.3200 ;
        RECT 1156.4600 643.4000 1159.4600 643.8800 ;
        RECT 1156.4600 654.2800 1159.4600 654.7600 ;
        RECT 1156.4600 697.8000 1159.4600 698.2800 ;
        RECT 1206.0200 697.8000 1207.6200 698.2800 ;
        RECT 1251.0200 697.8000 1252.6200 698.2800 ;
        RECT 1352.5600 632.5200 1355.5600 633.0000 ;
        RECT 1352.5600 637.9600 1355.5600 638.4400 ;
        RECT 1341.0200 632.5200 1342.6200 633.0000 ;
        RECT 1341.0200 637.9600 1342.6200 638.4400 ;
        RECT 1352.5600 616.2000 1355.5600 616.6800 ;
        RECT 1352.5600 621.6400 1355.5600 622.1200 ;
        RECT 1352.5600 627.0800 1355.5600 627.5600 ;
        RECT 1341.0200 616.2000 1342.6200 616.6800 ;
        RECT 1341.0200 621.6400 1342.6200 622.1200 ;
        RECT 1341.0200 627.0800 1342.6200 627.5600 ;
        RECT 1352.5600 605.3200 1355.5600 605.8000 ;
        RECT 1352.5600 610.7600 1355.5600 611.2400 ;
        RECT 1341.0200 605.3200 1342.6200 605.8000 ;
        RECT 1341.0200 610.7600 1342.6200 611.2400 ;
        RECT 1352.5600 589.0000 1355.5600 589.4800 ;
        RECT 1352.5600 594.4400 1355.5600 594.9200 ;
        RECT 1352.5600 599.8800 1355.5600 600.3600 ;
        RECT 1341.0200 589.0000 1342.6200 589.4800 ;
        RECT 1341.0200 594.4400 1342.6200 594.9200 ;
        RECT 1341.0200 599.8800 1342.6200 600.3600 ;
        RECT 1296.0200 632.5200 1297.6200 633.0000 ;
        RECT 1296.0200 637.9600 1297.6200 638.4400 ;
        RECT 1296.0200 616.2000 1297.6200 616.6800 ;
        RECT 1296.0200 621.6400 1297.6200 622.1200 ;
        RECT 1296.0200 627.0800 1297.6200 627.5600 ;
        RECT 1296.0200 605.3200 1297.6200 605.8000 ;
        RECT 1296.0200 610.7600 1297.6200 611.2400 ;
        RECT 1296.0200 589.0000 1297.6200 589.4800 ;
        RECT 1296.0200 594.4400 1297.6200 594.9200 ;
        RECT 1296.0200 599.8800 1297.6200 600.3600 ;
        RECT 1352.5600 578.1200 1355.5600 578.6000 ;
        RECT 1352.5600 583.5600 1355.5600 584.0400 ;
        RECT 1341.0200 578.1200 1342.6200 578.6000 ;
        RECT 1341.0200 583.5600 1342.6200 584.0400 ;
        RECT 1352.5600 561.8000 1355.5600 562.2800 ;
        RECT 1352.5600 567.2400 1355.5600 567.7200 ;
        RECT 1352.5600 572.6800 1355.5600 573.1600 ;
        RECT 1341.0200 561.8000 1342.6200 562.2800 ;
        RECT 1341.0200 567.2400 1342.6200 567.7200 ;
        RECT 1341.0200 572.6800 1342.6200 573.1600 ;
        RECT 1352.5600 550.9200 1355.5600 551.4000 ;
        RECT 1352.5600 556.3600 1355.5600 556.8400 ;
        RECT 1341.0200 550.9200 1342.6200 551.4000 ;
        RECT 1341.0200 556.3600 1342.6200 556.8400 ;
        RECT 1352.5600 545.4800 1355.5600 545.9600 ;
        RECT 1341.0200 545.4800 1342.6200 545.9600 ;
        RECT 1296.0200 578.1200 1297.6200 578.6000 ;
        RECT 1296.0200 583.5600 1297.6200 584.0400 ;
        RECT 1296.0200 561.8000 1297.6200 562.2800 ;
        RECT 1296.0200 567.2400 1297.6200 567.7200 ;
        RECT 1296.0200 572.6800 1297.6200 573.1600 ;
        RECT 1296.0200 550.9200 1297.6200 551.4000 ;
        RECT 1296.0200 556.3600 1297.6200 556.8400 ;
        RECT 1296.0200 545.4800 1297.6200 545.9600 ;
        RECT 1251.0200 632.5200 1252.6200 633.0000 ;
        RECT 1251.0200 637.9600 1252.6200 638.4400 ;
        RECT 1251.0200 616.2000 1252.6200 616.6800 ;
        RECT 1251.0200 621.6400 1252.6200 622.1200 ;
        RECT 1251.0200 627.0800 1252.6200 627.5600 ;
        RECT 1206.0200 632.5200 1207.6200 633.0000 ;
        RECT 1206.0200 637.9600 1207.6200 638.4400 ;
        RECT 1206.0200 616.2000 1207.6200 616.6800 ;
        RECT 1206.0200 621.6400 1207.6200 622.1200 ;
        RECT 1206.0200 627.0800 1207.6200 627.5600 ;
        RECT 1251.0200 605.3200 1252.6200 605.8000 ;
        RECT 1251.0200 610.7600 1252.6200 611.2400 ;
        RECT 1251.0200 589.0000 1252.6200 589.4800 ;
        RECT 1251.0200 594.4400 1252.6200 594.9200 ;
        RECT 1251.0200 599.8800 1252.6200 600.3600 ;
        RECT 1206.0200 605.3200 1207.6200 605.8000 ;
        RECT 1206.0200 610.7600 1207.6200 611.2400 ;
        RECT 1206.0200 589.0000 1207.6200 589.4800 ;
        RECT 1206.0200 594.4400 1207.6200 594.9200 ;
        RECT 1206.0200 599.8800 1207.6200 600.3600 ;
        RECT 1156.4600 632.5200 1159.4600 633.0000 ;
        RECT 1156.4600 637.9600 1159.4600 638.4400 ;
        RECT 1156.4600 621.6400 1159.4600 622.1200 ;
        RECT 1156.4600 616.2000 1159.4600 616.6800 ;
        RECT 1156.4600 627.0800 1159.4600 627.5600 ;
        RECT 1156.4600 605.3200 1159.4600 605.8000 ;
        RECT 1156.4600 610.7600 1159.4600 611.2400 ;
        RECT 1156.4600 594.4400 1159.4600 594.9200 ;
        RECT 1156.4600 589.0000 1159.4600 589.4800 ;
        RECT 1156.4600 599.8800 1159.4600 600.3600 ;
        RECT 1251.0200 578.1200 1252.6200 578.6000 ;
        RECT 1251.0200 583.5600 1252.6200 584.0400 ;
        RECT 1251.0200 561.8000 1252.6200 562.2800 ;
        RECT 1251.0200 567.2400 1252.6200 567.7200 ;
        RECT 1251.0200 572.6800 1252.6200 573.1600 ;
        RECT 1206.0200 578.1200 1207.6200 578.6000 ;
        RECT 1206.0200 583.5600 1207.6200 584.0400 ;
        RECT 1206.0200 561.8000 1207.6200 562.2800 ;
        RECT 1206.0200 567.2400 1207.6200 567.7200 ;
        RECT 1206.0200 572.6800 1207.6200 573.1600 ;
        RECT 1251.0200 556.3600 1252.6200 556.8400 ;
        RECT 1251.0200 550.9200 1252.6200 551.4000 ;
        RECT 1251.0200 545.4800 1252.6200 545.9600 ;
        RECT 1206.0200 556.3600 1207.6200 556.8400 ;
        RECT 1206.0200 550.9200 1207.6200 551.4000 ;
        RECT 1206.0200 545.4800 1207.6200 545.9600 ;
        RECT 1156.4600 578.1200 1159.4600 578.6000 ;
        RECT 1156.4600 583.5600 1159.4600 584.0400 ;
        RECT 1156.4600 567.2400 1159.4600 567.7200 ;
        RECT 1156.4600 561.8000 1159.4600 562.2800 ;
        RECT 1156.4600 572.6800 1159.4600 573.1600 ;
        RECT 1156.4600 550.9200 1159.4600 551.4000 ;
        RECT 1156.4600 556.3600 1159.4600 556.8400 ;
        RECT 1156.4600 545.4800 1159.4600 545.9600 ;
        RECT 1156.4600 743.6700 1355.5600 746.6700 ;
        RECT 1156.4600 538.5700 1355.5600 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 308.9300 1342.6200 517.0300 ;
        RECT 1296.0200 308.9300 1297.6200 517.0300 ;
        RECT 1251.0200 308.9300 1252.6200 517.0300 ;
        RECT 1206.0200 308.9300 1207.6200 517.0300 ;
        RECT 1352.5600 308.9300 1355.5600 517.0300 ;
        RECT 1156.4600 308.9300 1159.4600 517.0300 ;
      LAYER met3 ;
        RECT 1352.5600 511.6800 1355.5600 512.1600 ;
        RECT 1341.0200 511.6800 1342.6200 512.1600 ;
        RECT 1352.5600 500.8000 1355.5600 501.2800 ;
        RECT 1352.5600 506.2400 1355.5600 506.7200 ;
        RECT 1341.0200 500.8000 1342.6200 501.2800 ;
        RECT 1341.0200 506.2400 1342.6200 506.7200 ;
        RECT 1352.5600 484.4800 1355.5600 484.9600 ;
        RECT 1352.5600 489.9200 1355.5600 490.4000 ;
        RECT 1341.0200 484.4800 1342.6200 484.9600 ;
        RECT 1341.0200 489.9200 1342.6200 490.4000 ;
        RECT 1352.5600 473.6000 1355.5600 474.0800 ;
        RECT 1352.5600 479.0400 1355.5600 479.5200 ;
        RECT 1341.0200 473.6000 1342.6200 474.0800 ;
        RECT 1341.0200 479.0400 1342.6200 479.5200 ;
        RECT 1352.5600 495.3600 1355.5600 495.8400 ;
        RECT 1341.0200 495.3600 1342.6200 495.8400 ;
        RECT 1296.0200 500.8000 1297.6200 501.2800 ;
        RECT 1296.0200 506.2400 1297.6200 506.7200 ;
        RECT 1296.0200 511.6800 1297.6200 512.1600 ;
        RECT 1296.0200 484.4800 1297.6200 484.9600 ;
        RECT 1296.0200 489.9200 1297.6200 490.4000 ;
        RECT 1296.0200 479.0400 1297.6200 479.5200 ;
        RECT 1296.0200 473.6000 1297.6200 474.0800 ;
        RECT 1296.0200 495.3600 1297.6200 495.8400 ;
        RECT 1352.5600 457.2800 1355.5600 457.7600 ;
        RECT 1352.5600 462.7200 1355.5600 463.2000 ;
        RECT 1341.0200 457.2800 1342.6200 457.7600 ;
        RECT 1341.0200 462.7200 1342.6200 463.2000 ;
        RECT 1352.5600 440.9600 1355.5600 441.4400 ;
        RECT 1352.5600 446.4000 1355.5600 446.8800 ;
        RECT 1352.5600 451.8400 1355.5600 452.3200 ;
        RECT 1341.0200 440.9600 1342.6200 441.4400 ;
        RECT 1341.0200 446.4000 1342.6200 446.8800 ;
        RECT 1341.0200 451.8400 1342.6200 452.3200 ;
        RECT 1352.5600 430.0800 1355.5600 430.5600 ;
        RECT 1352.5600 435.5200 1355.5600 436.0000 ;
        RECT 1341.0200 430.0800 1342.6200 430.5600 ;
        RECT 1341.0200 435.5200 1342.6200 436.0000 ;
        RECT 1352.5600 413.7600 1355.5600 414.2400 ;
        RECT 1352.5600 419.2000 1355.5600 419.6800 ;
        RECT 1352.5600 424.6400 1355.5600 425.1200 ;
        RECT 1341.0200 413.7600 1342.6200 414.2400 ;
        RECT 1341.0200 419.2000 1342.6200 419.6800 ;
        RECT 1341.0200 424.6400 1342.6200 425.1200 ;
        RECT 1296.0200 457.2800 1297.6200 457.7600 ;
        RECT 1296.0200 462.7200 1297.6200 463.2000 ;
        RECT 1296.0200 440.9600 1297.6200 441.4400 ;
        RECT 1296.0200 446.4000 1297.6200 446.8800 ;
        RECT 1296.0200 451.8400 1297.6200 452.3200 ;
        RECT 1296.0200 430.0800 1297.6200 430.5600 ;
        RECT 1296.0200 435.5200 1297.6200 436.0000 ;
        RECT 1296.0200 413.7600 1297.6200 414.2400 ;
        RECT 1296.0200 419.2000 1297.6200 419.6800 ;
        RECT 1296.0200 424.6400 1297.6200 425.1200 ;
        RECT 1352.5600 468.1600 1355.5600 468.6400 ;
        RECT 1296.0200 468.1600 1297.6200 468.6400 ;
        RECT 1341.0200 468.1600 1342.6200 468.6400 ;
        RECT 1251.0200 500.8000 1252.6200 501.2800 ;
        RECT 1251.0200 506.2400 1252.6200 506.7200 ;
        RECT 1251.0200 511.6800 1252.6200 512.1600 ;
        RECT 1206.0200 500.8000 1207.6200 501.2800 ;
        RECT 1206.0200 506.2400 1207.6200 506.7200 ;
        RECT 1206.0200 511.6800 1207.6200 512.1600 ;
        RECT 1251.0200 484.4800 1252.6200 484.9600 ;
        RECT 1251.0200 489.9200 1252.6200 490.4000 ;
        RECT 1251.0200 473.6000 1252.6200 474.0800 ;
        RECT 1251.0200 479.0400 1252.6200 479.5200 ;
        RECT 1206.0200 484.4800 1207.6200 484.9600 ;
        RECT 1206.0200 489.9200 1207.6200 490.4000 ;
        RECT 1206.0200 473.6000 1207.6200 474.0800 ;
        RECT 1206.0200 479.0400 1207.6200 479.5200 ;
        RECT 1206.0200 495.3600 1207.6200 495.8400 ;
        RECT 1251.0200 495.3600 1252.6200 495.8400 ;
        RECT 1156.4600 511.6800 1159.4600 512.1600 ;
        RECT 1156.4600 506.2400 1159.4600 506.7200 ;
        RECT 1156.4600 500.8000 1159.4600 501.2800 ;
        RECT 1156.4600 489.9200 1159.4600 490.4000 ;
        RECT 1156.4600 484.4800 1159.4600 484.9600 ;
        RECT 1156.4600 479.0400 1159.4600 479.5200 ;
        RECT 1156.4600 473.6000 1159.4600 474.0800 ;
        RECT 1156.4600 495.3600 1159.4600 495.8400 ;
        RECT 1251.0200 457.2800 1252.6200 457.7600 ;
        RECT 1251.0200 462.7200 1252.6200 463.2000 ;
        RECT 1251.0200 440.9600 1252.6200 441.4400 ;
        RECT 1251.0200 446.4000 1252.6200 446.8800 ;
        RECT 1251.0200 451.8400 1252.6200 452.3200 ;
        RECT 1206.0200 457.2800 1207.6200 457.7600 ;
        RECT 1206.0200 462.7200 1207.6200 463.2000 ;
        RECT 1206.0200 440.9600 1207.6200 441.4400 ;
        RECT 1206.0200 446.4000 1207.6200 446.8800 ;
        RECT 1206.0200 451.8400 1207.6200 452.3200 ;
        RECT 1251.0200 430.0800 1252.6200 430.5600 ;
        RECT 1251.0200 435.5200 1252.6200 436.0000 ;
        RECT 1251.0200 413.7600 1252.6200 414.2400 ;
        RECT 1251.0200 419.2000 1252.6200 419.6800 ;
        RECT 1251.0200 424.6400 1252.6200 425.1200 ;
        RECT 1206.0200 430.0800 1207.6200 430.5600 ;
        RECT 1206.0200 435.5200 1207.6200 436.0000 ;
        RECT 1206.0200 413.7600 1207.6200 414.2400 ;
        RECT 1206.0200 419.2000 1207.6200 419.6800 ;
        RECT 1206.0200 424.6400 1207.6200 425.1200 ;
        RECT 1156.4600 457.2800 1159.4600 457.7600 ;
        RECT 1156.4600 462.7200 1159.4600 463.2000 ;
        RECT 1156.4600 446.4000 1159.4600 446.8800 ;
        RECT 1156.4600 440.9600 1159.4600 441.4400 ;
        RECT 1156.4600 451.8400 1159.4600 452.3200 ;
        RECT 1156.4600 430.0800 1159.4600 430.5600 ;
        RECT 1156.4600 435.5200 1159.4600 436.0000 ;
        RECT 1156.4600 419.2000 1159.4600 419.6800 ;
        RECT 1156.4600 413.7600 1159.4600 414.2400 ;
        RECT 1156.4600 424.6400 1159.4600 425.1200 ;
        RECT 1156.4600 468.1600 1159.4600 468.6400 ;
        RECT 1206.0200 468.1600 1207.6200 468.6400 ;
        RECT 1251.0200 468.1600 1252.6200 468.6400 ;
        RECT 1352.5600 402.8800 1355.5600 403.3600 ;
        RECT 1352.5600 408.3200 1355.5600 408.8000 ;
        RECT 1341.0200 402.8800 1342.6200 403.3600 ;
        RECT 1341.0200 408.3200 1342.6200 408.8000 ;
        RECT 1352.5600 386.5600 1355.5600 387.0400 ;
        RECT 1352.5600 392.0000 1355.5600 392.4800 ;
        RECT 1352.5600 397.4400 1355.5600 397.9200 ;
        RECT 1341.0200 386.5600 1342.6200 387.0400 ;
        RECT 1341.0200 392.0000 1342.6200 392.4800 ;
        RECT 1341.0200 397.4400 1342.6200 397.9200 ;
        RECT 1352.5600 375.6800 1355.5600 376.1600 ;
        RECT 1352.5600 381.1200 1355.5600 381.6000 ;
        RECT 1341.0200 375.6800 1342.6200 376.1600 ;
        RECT 1341.0200 381.1200 1342.6200 381.6000 ;
        RECT 1352.5600 359.3600 1355.5600 359.8400 ;
        RECT 1352.5600 364.8000 1355.5600 365.2800 ;
        RECT 1352.5600 370.2400 1355.5600 370.7200 ;
        RECT 1341.0200 359.3600 1342.6200 359.8400 ;
        RECT 1341.0200 364.8000 1342.6200 365.2800 ;
        RECT 1341.0200 370.2400 1342.6200 370.7200 ;
        RECT 1296.0200 402.8800 1297.6200 403.3600 ;
        RECT 1296.0200 408.3200 1297.6200 408.8000 ;
        RECT 1296.0200 386.5600 1297.6200 387.0400 ;
        RECT 1296.0200 392.0000 1297.6200 392.4800 ;
        RECT 1296.0200 397.4400 1297.6200 397.9200 ;
        RECT 1296.0200 375.6800 1297.6200 376.1600 ;
        RECT 1296.0200 381.1200 1297.6200 381.6000 ;
        RECT 1296.0200 359.3600 1297.6200 359.8400 ;
        RECT 1296.0200 364.8000 1297.6200 365.2800 ;
        RECT 1296.0200 370.2400 1297.6200 370.7200 ;
        RECT 1352.5600 348.4800 1355.5600 348.9600 ;
        RECT 1352.5600 353.9200 1355.5600 354.4000 ;
        RECT 1341.0200 348.4800 1342.6200 348.9600 ;
        RECT 1341.0200 353.9200 1342.6200 354.4000 ;
        RECT 1352.5600 332.1600 1355.5600 332.6400 ;
        RECT 1352.5600 337.6000 1355.5600 338.0800 ;
        RECT 1352.5600 343.0400 1355.5600 343.5200 ;
        RECT 1341.0200 332.1600 1342.6200 332.6400 ;
        RECT 1341.0200 337.6000 1342.6200 338.0800 ;
        RECT 1341.0200 343.0400 1342.6200 343.5200 ;
        RECT 1352.5600 321.2800 1355.5600 321.7600 ;
        RECT 1352.5600 326.7200 1355.5600 327.2000 ;
        RECT 1341.0200 321.2800 1342.6200 321.7600 ;
        RECT 1341.0200 326.7200 1342.6200 327.2000 ;
        RECT 1352.5600 315.8400 1355.5600 316.3200 ;
        RECT 1341.0200 315.8400 1342.6200 316.3200 ;
        RECT 1296.0200 348.4800 1297.6200 348.9600 ;
        RECT 1296.0200 353.9200 1297.6200 354.4000 ;
        RECT 1296.0200 332.1600 1297.6200 332.6400 ;
        RECT 1296.0200 337.6000 1297.6200 338.0800 ;
        RECT 1296.0200 343.0400 1297.6200 343.5200 ;
        RECT 1296.0200 321.2800 1297.6200 321.7600 ;
        RECT 1296.0200 326.7200 1297.6200 327.2000 ;
        RECT 1296.0200 315.8400 1297.6200 316.3200 ;
        RECT 1251.0200 402.8800 1252.6200 403.3600 ;
        RECT 1251.0200 408.3200 1252.6200 408.8000 ;
        RECT 1251.0200 386.5600 1252.6200 387.0400 ;
        RECT 1251.0200 392.0000 1252.6200 392.4800 ;
        RECT 1251.0200 397.4400 1252.6200 397.9200 ;
        RECT 1206.0200 402.8800 1207.6200 403.3600 ;
        RECT 1206.0200 408.3200 1207.6200 408.8000 ;
        RECT 1206.0200 386.5600 1207.6200 387.0400 ;
        RECT 1206.0200 392.0000 1207.6200 392.4800 ;
        RECT 1206.0200 397.4400 1207.6200 397.9200 ;
        RECT 1251.0200 375.6800 1252.6200 376.1600 ;
        RECT 1251.0200 381.1200 1252.6200 381.6000 ;
        RECT 1251.0200 359.3600 1252.6200 359.8400 ;
        RECT 1251.0200 364.8000 1252.6200 365.2800 ;
        RECT 1251.0200 370.2400 1252.6200 370.7200 ;
        RECT 1206.0200 375.6800 1207.6200 376.1600 ;
        RECT 1206.0200 381.1200 1207.6200 381.6000 ;
        RECT 1206.0200 359.3600 1207.6200 359.8400 ;
        RECT 1206.0200 364.8000 1207.6200 365.2800 ;
        RECT 1206.0200 370.2400 1207.6200 370.7200 ;
        RECT 1156.4600 402.8800 1159.4600 403.3600 ;
        RECT 1156.4600 408.3200 1159.4600 408.8000 ;
        RECT 1156.4600 392.0000 1159.4600 392.4800 ;
        RECT 1156.4600 386.5600 1159.4600 387.0400 ;
        RECT 1156.4600 397.4400 1159.4600 397.9200 ;
        RECT 1156.4600 375.6800 1159.4600 376.1600 ;
        RECT 1156.4600 381.1200 1159.4600 381.6000 ;
        RECT 1156.4600 364.8000 1159.4600 365.2800 ;
        RECT 1156.4600 359.3600 1159.4600 359.8400 ;
        RECT 1156.4600 370.2400 1159.4600 370.7200 ;
        RECT 1251.0200 348.4800 1252.6200 348.9600 ;
        RECT 1251.0200 353.9200 1252.6200 354.4000 ;
        RECT 1251.0200 332.1600 1252.6200 332.6400 ;
        RECT 1251.0200 337.6000 1252.6200 338.0800 ;
        RECT 1251.0200 343.0400 1252.6200 343.5200 ;
        RECT 1206.0200 348.4800 1207.6200 348.9600 ;
        RECT 1206.0200 353.9200 1207.6200 354.4000 ;
        RECT 1206.0200 332.1600 1207.6200 332.6400 ;
        RECT 1206.0200 337.6000 1207.6200 338.0800 ;
        RECT 1206.0200 343.0400 1207.6200 343.5200 ;
        RECT 1251.0200 326.7200 1252.6200 327.2000 ;
        RECT 1251.0200 321.2800 1252.6200 321.7600 ;
        RECT 1251.0200 315.8400 1252.6200 316.3200 ;
        RECT 1206.0200 326.7200 1207.6200 327.2000 ;
        RECT 1206.0200 321.2800 1207.6200 321.7600 ;
        RECT 1206.0200 315.8400 1207.6200 316.3200 ;
        RECT 1156.4600 348.4800 1159.4600 348.9600 ;
        RECT 1156.4600 353.9200 1159.4600 354.4000 ;
        RECT 1156.4600 337.6000 1159.4600 338.0800 ;
        RECT 1156.4600 332.1600 1159.4600 332.6400 ;
        RECT 1156.4600 343.0400 1159.4600 343.5200 ;
        RECT 1156.4600 321.2800 1159.4600 321.7600 ;
        RECT 1156.4600 326.7200 1159.4600 327.2000 ;
        RECT 1156.4600 315.8400 1159.4600 316.3200 ;
        RECT 1156.4600 514.0300 1355.5600 517.0300 ;
        RECT 1156.4600 308.9300 1355.5600 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 79.2900 1342.6200 287.3900 ;
        RECT 1296.0200 79.2900 1297.6200 287.3900 ;
        RECT 1251.0200 79.2900 1252.6200 287.3900 ;
        RECT 1206.0200 79.2900 1207.6200 287.3900 ;
        RECT 1352.5600 79.2900 1355.5600 287.3900 ;
        RECT 1156.4600 79.2900 1159.4600 287.3900 ;
      LAYER met3 ;
        RECT 1352.5600 282.0400 1355.5600 282.5200 ;
        RECT 1341.0200 282.0400 1342.6200 282.5200 ;
        RECT 1352.5600 271.1600 1355.5600 271.6400 ;
        RECT 1352.5600 276.6000 1355.5600 277.0800 ;
        RECT 1341.0200 271.1600 1342.6200 271.6400 ;
        RECT 1341.0200 276.6000 1342.6200 277.0800 ;
        RECT 1352.5600 254.8400 1355.5600 255.3200 ;
        RECT 1352.5600 260.2800 1355.5600 260.7600 ;
        RECT 1341.0200 254.8400 1342.6200 255.3200 ;
        RECT 1341.0200 260.2800 1342.6200 260.7600 ;
        RECT 1352.5600 243.9600 1355.5600 244.4400 ;
        RECT 1352.5600 249.4000 1355.5600 249.8800 ;
        RECT 1341.0200 243.9600 1342.6200 244.4400 ;
        RECT 1341.0200 249.4000 1342.6200 249.8800 ;
        RECT 1352.5600 265.7200 1355.5600 266.2000 ;
        RECT 1341.0200 265.7200 1342.6200 266.2000 ;
        RECT 1296.0200 271.1600 1297.6200 271.6400 ;
        RECT 1296.0200 276.6000 1297.6200 277.0800 ;
        RECT 1296.0200 282.0400 1297.6200 282.5200 ;
        RECT 1296.0200 254.8400 1297.6200 255.3200 ;
        RECT 1296.0200 260.2800 1297.6200 260.7600 ;
        RECT 1296.0200 249.4000 1297.6200 249.8800 ;
        RECT 1296.0200 243.9600 1297.6200 244.4400 ;
        RECT 1296.0200 265.7200 1297.6200 266.2000 ;
        RECT 1352.5600 227.6400 1355.5600 228.1200 ;
        RECT 1352.5600 233.0800 1355.5600 233.5600 ;
        RECT 1341.0200 227.6400 1342.6200 228.1200 ;
        RECT 1341.0200 233.0800 1342.6200 233.5600 ;
        RECT 1352.5600 211.3200 1355.5600 211.8000 ;
        RECT 1352.5600 216.7600 1355.5600 217.2400 ;
        RECT 1352.5600 222.2000 1355.5600 222.6800 ;
        RECT 1341.0200 211.3200 1342.6200 211.8000 ;
        RECT 1341.0200 216.7600 1342.6200 217.2400 ;
        RECT 1341.0200 222.2000 1342.6200 222.6800 ;
        RECT 1352.5600 200.4400 1355.5600 200.9200 ;
        RECT 1352.5600 205.8800 1355.5600 206.3600 ;
        RECT 1341.0200 200.4400 1342.6200 200.9200 ;
        RECT 1341.0200 205.8800 1342.6200 206.3600 ;
        RECT 1352.5600 184.1200 1355.5600 184.6000 ;
        RECT 1352.5600 189.5600 1355.5600 190.0400 ;
        RECT 1352.5600 195.0000 1355.5600 195.4800 ;
        RECT 1341.0200 184.1200 1342.6200 184.6000 ;
        RECT 1341.0200 189.5600 1342.6200 190.0400 ;
        RECT 1341.0200 195.0000 1342.6200 195.4800 ;
        RECT 1296.0200 227.6400 1297.6200 228.1200 ;
        RECT 1296.0200 233.0800 1297.6200 233.5600 ;
        RECT 1296.0200 211.3200 1297.6200 211.8000 ;
        RECT 1296.0200 216.7600 1297.6200 217.2400 ;
        RECT 1296.0200 222.2000 1297.6200 222.6800 ;
        RECT 1296.0200 200.4400 1297.6200 200.9200 ;
        RECT 1296.0200 205.8800 1297.6200 206.3600 ;
        RECT 1296.0200 184.1200 1297.6200 184.6000 ;
        RECT 1296.0200 189.5600 1297.6200 190.0400 ;
        RECT 1296.0200 195.0000 1297.6200 195.4800 ;
        RECT 1352.5600 238.5200 1355.5600 239.0000 ;
        RECT 1296.0200 238.5200 1297.6200 239.0000 ;
        RECT 1341.0200 238.5200 1342.6200 239.0000 ;
        RECT 1251.0200 271.1600 1252.6200 271.6400 ;
        RECT 1251.0200 276.6000 1252.6200 277.0800 ;
        RECT 1251.0200 282.0400 1252.6200 282.5200 ;
        RECT 1206.0200 271.1600 1207.6200 271.6400 ;
        RECT 1206.0200 276.6000 1207.6200 277.0800 ;
        RECT 1206.0200 282.0400 1207.6200 282.5200 ;
        RECT 1251.0200 254.8400 1252.6200 255.3200 ;
        RECT 1251.0200 260.2800 1252.6200 260.7600 ;
        RECT 1251.0200 243.9600 1252.6200 244.4400 ;
        RECT 1251.0200 249.4000 1252.6200 249.8800 ;
        RECT 1206.0200 254.8400 1207.6200 255.3200 ;
        RECT 1206.0200 260.2800 1207.6200 260.7600 ;
        RECT 1206.0200 243.9600 1207.6200 244.4400 ;
        RECT 1206.0200 249.4000 1207.6200 249.8800 ;
        RECT 1206.0200 265.7200 1207.6200 266.2000 ;
        RECT 1251.0200 265.7200 1252.6200 266.2000 ;
        RECT 1156.4600 282.0400 1159.4600 282.5200 ;
        RECT 1156.4600 276.6000 1159.4600 277.0800 ;
        RECT 1156.4600 271.1600 1159.4600 271.6400 ;
        RECT 1156.4600 260.2800 1159.4600 260.7600 ;
        RECT 1156.4600 254.8400 1159.4600 255.3200 ;
        RECT 1156.4600 249.4000 1159.4600 249.8800 ;
        RECT 1156.4600 243.9600 1159.4600 244.4400 ;
        RECT 1156.4600 265.7200 1159.4600 266.2000 ;
        RECT 1251.0200 227.6400 1252.6200 228.1200 ;
        RECT 1251.0200 233.0800 1252.6200 233.5600 ;
        RECT 1251.0200 211.3200 1252.6200 211.8000 ;
        RECT 1251.0200 216.7600 1252.6200 217.2400 ;
        RECT 1251.0200 222.2000 1252.6200 222.6800 ;
        RECT 1206.0200 227.6400 1207.6200 228.1200 ;
        RECT 1206.0200 233.0800 1207.6200 233.5600 ;
        RECT 1206.0200 211.3200 1207.6200 211.8000 ;
        RECT 1206.0200 216.7600 1207.6200 217.2400 ;
        RECT 1206.0200 222.2000 1207.6200 222.6800 ;
        RECT 1251.0200 200.4400 1252.6200 200.9200 ;
        RECT 1251.0200 205.8800 1252.6200 206.3600 ;
        RECT 1251.0200 184.1200 1252.6200 184.6000 ;
        RECT 1251.0200 189.5600 1252.6200 190.0400 ;
        RECT 1251.0200 195.0000 1252.6200 195.4800 ;
        RECT 1206.0200 200.4400 1207.6200 200.9200 ;
        RECT 1206.0200 205.8800 1207.6200 206.3600 ;
        RECT 1206.0200 184.1200 1207.6200 184.6000 ;
        RECT 1206.0200 189.5600 1207.6200 190.0400 ;
        RECT 1206.0200 195.0000 1207.6200 195.4800 ;
        RECT 1156.4600 227.6400 1159.4600 228.1200 ;
        RECT 1156.4600 233.0800 1159.4600 233.5600 ;
        RECT 1156.4600 216.7600 1159.4600 217.2400 ;
        RECT 1156.4600 211.3200 1159.4600 211.8000 ;
        RECT 1156.4600 222.2000 1159.4600 222.6800 ;
        RECT 1156.4600 200.4400 1159.4600 200.9200 ;
        RECT 1156.4600 205.8800 1159.4600 206.3600 ;
        RECT 1156.4600 189.5600 1159.4600 190.0400 ;
        RECT 1156.4600 184.1200 1159.4600 184.6000 ;
        RECT 1156.4600 195.0000 1159.4600 195.4800 ;
        RECT 1156.4600 238.5200 1159.4600 239.0000 ;
        RECT 1206.0200 238.5200 1207.6200 239.0000 ;
        RECT 1251.0200 238.5200 1252.6200 239.0000 ;
        RECT 1352.5600 173.2400 1355.5600 173.7200 ;
        RECT 1352.5600 178.6800 1355.5600 179.1600 ;
        RECT 1341.0200 173.2400 1342.6200 173.7200 ;
        RECT 1341.0200 178.6800 1342.6200 179.1600 ;
        RECT 1352.5600 156.9200 1355.5600 157.4000 ;
        RECT 1352.5600 162.3600 1355.5600 162.8400 ;
        RECT 1352.5600 167.8000 1355.5600 168.2800 ;
        RECT 1341.0200 156.9200 1342.6200 157.4000 ;
        RECT 1341.0200 162.3600 1342.6200 162.8400 ;
        RECT 1341.0200 167.8000 1342.6200 168.2800 ;
        RECT 1352.5600 146.0400 1355.5600 146.5200 ;
        RECT 1352.5600 151.4800 1355.5600 151.9600 ;
        RECT 1341.0200 146.0400 1342.6200 146.5200 ;
        RECT 1341.0200 151.4800 1342.6200 151.9600 ;
        RECT 1352.5600 129.7200 1355.5600 130.2000 ;
        RECT 1352.5600 135.1600 1355.5600 135.6400 ;
        RECT 1352.5600 140.6000 1355.5600 141.0800 ;
        RECT 1341.0200 129.7200 1342.6200 130.2000 ;
        RECT 1341.0200 135.1600 1342.6200 135.6400 ;
        RECT 1341.0200 140.6000 1342.6200 141.0800 ;
        RECT 1296.0200 173.2400 1297.6200 173.7200 ;
        RECT 1296.0200 178.6800 1297.6200 179.1600 ;
        RECT 1296.0200 156.9200 1297.6200 157.4000 ;
        RECT 1296.0200 162.3600 1297.6200 162.8400 ;
        RECT 1296.0200 167.8000 1297.6200 168.2800 ;
        RECT 1296.0200 146.0400 1297.6200 146.5200 ;
        RECT 1296.0200 151.4800 1297.6200 151.9600 ;
        RECT 1296.0200 129.7200 1297.6200 130.2000 ;
        RECT 1296.0200 135.1600 1297.6200 135.6400 ;
        RECT 1296.0200 140.6000 1297.6200 141.0800 ;
        RECT 1352.5600 118.8400 1355.5600 119.3200 ;
        RECT 1352.5600 124.2800 1355.5600 124.7600 ;
        RECT 1341.0200 118.8400 1342.6200 119.3200 ;
        RECT 1341.0200 124.2800 1342.6200 124.7600 ;
        RECT 1352.5600 102.5200 1355.5600 103.0000 ;
        RECT 1352.5600 107.9600 1355.5600 108.4400 ;
        RECT 1352.5600 113.4000 1355.5600 113.8800 ;
        RECT 1341.0200 102.5200 1342.6200 103.0000 ;
        RECT 1341.0200 107.9600 1342.6200 108.4400 ;
        RECT 1341.0200 113.4000 1342.6200 113.8800 ;
        RECT 1352.5600 91.6400 1355.5600 92.1200 ;
        RECT 1352.5600 97.0800 1355.5600 97.5600 ;
        RECT 1341.0200 91.6400 1342.6200 92.1200 ;
        RECT 1341.0200 97.0800 1342.6200 97.5600 ;
        RECT 1352.5600 86.2000 1355.5600 86.6800 ;
        RECT 1341.0200 86.2000 1342.6200 86.6800 ;
        RECT 1296.0200 118.8400 1297.6200 119.3200 ;
        RECT 1296.0200 124.2800 1297.6200 124.7600 ;
        RECT 1296.0200 102.5200 1297.6200 103.0000 ;
        RECT 1296.0200 107.9600 1297.6200 108.4400 ;
        RECT 1296.0200 113.4000 1297.6200 113.8800 ;
        RECT 1296.0200 91.6400 1297.6200 92.1200 ;
        RECT 1296.0200 97.0800 1297.6200 97.5600 ;
        RECT 1296.0200 86.2000 1297.6200 86.6800 ;
        RECT 1251.0200 173.2400 1252.6200 173.7200 ;
        RECT 1251.0200 178.6800 1252.6200 179.1600 ;
        RECT 1251.0200 156.9200 1252.6200 157.4000 ;
        RECT 1251.0200 162.3600 1252.6200 162.8400 ;
        RECT 1251.0200 167.8000 1252.6200 168.2800 ;
        RECT 1206.0200 173.2400 1207.6200 173.7200 ;
        RECT 1206.0200 178.6800 1207.6200 179.1600 ;
        RECT 1206.0200 156.9200 1207.6200 157.4000 ;
        RECT 1206.0200 162.3600 1207.6200 162.8400 ;
        RECT 1206.0200 167.8000 1207.6200 168.2800 ;
        RECT 1251.0200 146.0400 1252.6200 146.5200 ;
        RECT 1251.0200 151.4800 1252.6200 151.9600 ;
        RECT 1251.0200 129.7200 1252.6200 130.2000 ;
        RECT 1251.0200 135.1600 1252.6200 135.6400 ;
        RECT 1251.0200 140.6000 1252.6200 141.0800 ;
        RECT 1206.0200 146.0400 1207.6200 146.5200 ;
        RECT 1206.0200 151.4800 1207.6200 151.9600 ;
        RECT 1206.0200 129.7200 1207.6200 130.2000 ;
        RECT 1206.0200 135.1600 1207.6200 135.6400 ;
        RECT 1206.0200 140.6000 1207.6200 141.0800 ;
        RECT 1156.4600 173.2400 1159.4600 173.7200 ;
        RECT 1156.4600 178.6800 1159.4600 179.1600 ;
        RECT 1156.4600 162.3600 1159.4600 162.8400 ;
        RECT 1156.4600 156.9200 1159.4600 157.4000 ;
        RECT 1156.4600 167.8000 1159.4600 168.2800 ;
        RECT 1156.4600 146.0400 1159.4600 146.5200 ;
        RECT 1156.4600 151.4800 1159.4600 151.9600 ;
        RECT 1156.4600 135.1600 1159.4600 135.6400 ;
        RECT 1156.4600 129.7200 1159.4600 130.2000 ;
        RECT 1156.4600 140.6000 1159.4600 141.0800 ;
        RECT 1251.0200 118.8400 1252.6200 119.3200 ;
        RECT 1251.0200 124.2800 1252.6200 124.7600 ;
        RECT 1251.0200 102.5200 1252.6200 103.0000 ;
        RECT 1251.0200 107.9600 1252.6200 108.4400 ;
        RECT 1251.0200 113.4000 1252.6200 113.8800 ;
        RECT 1206.0200 118.8400 1207.6200 119.3200 ;
        RECT 1206.0200 124.2800 1207.6200 124.7600 ;
        RECT 1206.0200 102.5200 1207.6200 103.0000 ;
        RECT 1206.0200 107.9600 1207.6200 108.4400 ;
        RECT 1206.0200 113.4000 1207.6200 113.8800 ;
        RECT 1251.0200 97.0800 1252.6200 97.5600 ;
        RECT 1251.0200 91.6400 1252.6200 92.1200 ;
        RECT 1251.0200 86.2000 1252.6200 86.6800 ;
        RECT 1206.0200 97.0800 1207.6200 97.5600 ;
        RECT 1206.0200 91.6400 1207.6200 92.1200 ;
        RECT 1206.0200 86.2000 1207.6200 86.6800 ;
        RECT 1156.4600 118.8400 1159.4600 119.3200 ;
        RECT 1156.4600 124.2800 1159.4600 124.7600 ;
        RECT 1156.4600 107.9600 1159.4600 108.4400 ;
        RECT 1156.4600 102.5200 1159.4600 103.0000 ;
        RECT 1156.4600 113.4000 1159.4600 113.8800 ;
        RECT 1156.4600 91.6400 1159.4600 92.1200 ;
        RECT 1156.4600 97.0800 1159.4600 97.5600 ;
        RECT 1156.4600 86.2000 1159.4600 86.6800 ;
        RECT 1156.4600 284.3900 1355.5600 287.3900 ;
        RECT 1156.4600 79.2900 1355.5600 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1156.4600 37.6700 1158.4600 58.6000 ;
        RECT 1353.5600 37.6700 1355.5600 58.6000 ;
      LAYER met3 ;
        RECT 1353.5600 54.1000 1355.5600 54.5800 ;
        RECT 1156.4600 54.1000 1158.4600 54.5800 ;
        RECT 1353.5600 43.2200 1355.5600 43.7000 ;
        RECT 1156.4600 43.2200 1158.4600 43.7000 ;
        RECT 1353.5600 48.6600 1355.5600 49.1400 ;
        RECT 1156.4600 48.6600 1158.4600 49.1400 ;
        RECT 1156.4600 56.6000 1355.5600 58.6000 ;
        RECT 1156.4600 37.6700 1355.5600 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 2605.3300 1342.6200 2813.4300 ;
        RECT 1296.0200 2605.3300 1297.6200 2813.4300 ;
        RECT 1251.0200 2605.3300 1252.6200 2813.4300 ;
        RECT 1206.0200 2605.3300 1207.6200 2813.4300 ;
        RECT 1352.5600 2605.3300 1355.5600 2813.4300 ;
        RECT 1156.4600 2605.3300 1159.4600 2813.4300 ;
      LAYER met3 ;
        RECT 1352.5600 2808.0800 1355.5600 2808.5600 ;
        RECT 1341.0200 2808.0800 1342.6200 2808.5600 ;
        RECT 1352.5600 2797.2000 1355.5600 2797.6800 ;
        RECT 1352.5600 2802.6400 1355.5600 2803.1200 ;
        RECT 1341.0200 2797.2000 1342.6200 2797.6800 ;
        RECT 1341.0200 2802.6400 1342.6200 2803.1200 ;
        RECT 1352.5600 2780.8800 1355.5600 2781.3600 ;
        RECT 1352.5600 2786.3200 1355.5600 2786.8000 ;
        RECT 1341.0200 2780.8800 1342.6200 2781.3600 ;
        RECT 1341.0200 2786.3200 1342.6200 2786.8000 ;
        RECT 1352.5600 2770.0000 1355.5600 2770.4800 ;
        RECT 1352.5600 2775.4400 1355.5600 2775.9200 ;
        RECT 1341.0200 2770.0000 1342.6200 2770.4800 ;
        RECT 1341.0200 2775.4400 1342.6200 2775.9200 ;
        RECT 1352.5600 2791.7600 1355.5600 2792.2400 ;
        RECT 1341.0200 2791.7600 1342.6200 2792.2400 ;
        RECT 1296.0200 2797.2000 1297.6200 2797.6800 ;
        RECT 1296.0200 2802.6400 1297.6200 2803.1200 ;
        RECT 1296.0200 2808.0800 1297.6200 2808.5600 ;
        RECT 1296.0200 2780.8800 1297.6200 2781.3600 ;
        RECT 1296.0200 2786.3200 1297.6200 2786.8000 ;
        RECT 1296.0200 2775.4400 1297.6200 2775.9200 ;
        RECT 1296.0200 2770.0000 1297.6200 2770.4800 ;
        RECT 1296.0200 2791.7600 1297.6200 2792.2400 ;
        RECT 1352.5600 2753.6800 1355.5600 2754.1600 ;
        RECT 1352.5600 2759.1200 1355.5600 2759.6000 ;
        RECT 1341.0200 2753.6800 1342.6200 2754.1600 ;
        RECT 1341.0200 2759.1200 1342.6200 2759.6000 ;
        RECT 1352.5600 2737.3600 1355.5600 2737.8400 ;
        RECT 1352.5600 2742.8000 1355.5600 2743.2800 ;
        RECT 1352.5600 2748.2400 1355.5600 2748.7200 ;
        RECT 1341.0200 2737.3600 1342.6200 2737.8400 ;
        RECT 1341.0200 2742.8000 1342.6200 2743.2800 ;
        RECT 1341.0200 2748.2400 1342.6200 2748.7200 ;
        RECT 1352.5600 2726.4800 1355.5600 2726.9600 ;
        RECT 1352.5600 2731.9200 1355.5600 2732.4000 ;
        RECT 1341.0200 2726.4800 1342.6200 2726.9600 ;
        RECT 1341.0200 2731.9200 1342.6200 2732.4000 ;
        RECT 1352.5600 2710.1600 1355.5600 2710.6400 ;
        RECT 1352.5600 2715.6000 1355.5600 2716.0800 ;
        RECT 1352.5600 2721.0400 1355.5600 2721.5200 ;
        RECT 1341.0200 2710.1600 1342.6200 2710.6400 ;
        RECT 1341.0200 2715.6000 1342.6200 2716.0800 ;
        RECT 1341.0200 2721.0400 1342.6200 2721.5200 ;
        RECT 1296.0200 2753.6800 1297.6200 2754.1600 ;
        RECT 1296.0200 2759.1200 1297.6200 2759.6000 ;
        RECT 1296.0200 2737.3600 1297.6200 2737.8400 ;
        RECT 1296.0200 2742.8000 1297.6200 2743.2800 ;
        RECT 1296.0200 2748.2400 1297.6200 2748.7200 ;
        RECT 1296.0200 2726.4800 1297.6200 2726.9600 ;
        RECT 1296.0200 2731.9200 1297.6200 2732.4000 ;
        RECT 1296.0200 2710.1600 1297.6200 2710.6400 ;
        RECT 1296.0200 2715.6000 1297.6200 2716.0800 ;
        RECT 1296.0200 2721.0400 1297.6200 2721.5200 ;
        RECT 1352.5600 2764.5600 1355.5600 2765.0400 ;
        RECT 1296.0200 2764.5600 1297.6200 2765.0400 ;
        RECT 1341.0200 2764.5600 1342.6200 2765.0400 ;
        RECT 1251.0200 2797.2000 1252.6200 2797.6800 ;
        RECT 1251.0200 2802.6400 1252.6200 2803.1200 ;
        RECT 1251.0200 2808.0800 1252.6200 2808.5600 ;
        RECT 1206.0200 2797.2000 1207.6200 2797.6800 ;
        RECT 1206.0200 2802.6400 1207.6200 2803.1200 ;
        RECT 1206.0200 2808.0800 1207.6200 2808.5600 ;
        RECT 1251.0200 2780.8800 1252.6200 2781.3600 ;
        RECT 1251.0200 2786.3200 1252.6200 2786.8000 ;
        RECT 1251.0200 2770.0000 1252.6200 2770.4800 ;
        RECT 1251.0200 2775.4400 1252.6200 2775.9200 ;
        RECT 1206.0200 2780.8800 1207.6200 2781.3600 ;
        RECT 1206.0200 2786.3200 1207.6200 2786.8000 ;
        RECT 1206.0200 2770.0000 1207.6200 2770.4800 ;
        RECT 1206.0200 2775.4400 1207.6200 2775.9200 ;
        RECT 1206.0200 2791.7600 1207.6200 2792.2400 ;
        RECT 1251.0200 2791.7600 1252.6200 2792.2400 ;
        RECT 1156.4600 2808.0800 1159.4600 2808.5600 ;
        RECT 1156.4600 2802.6400 1159.4600 2803.1200 ;
        RECT 1156.4600 2797.2000 1159.4600 2797.6800 ;
        RECT 1156.4600 2786.3200 1159.4600 2786.8000 ;
        RECT 1156.4600 2780.8800 1159.4600 2781.3600 ;
        RECT 1156.4600 2775.4400 1159.4600 2775.9200 ;
        RECT 1156.4600 2770.0000 1159.4600 2770.4800 ;
        RECT 1156.4600 2791.7600 1159.4600 2792.2400 ;
        RECT 1251.0200 2753.6800 1252.6200 2754.1600 ;
        RECT 1251.0200 2759.1200 1252.6200 2759.6000 ;
        RECT 1251.0200 2737.3600 1252.6200 2737.8400 ;
        RECT 1251.0200 2742.8000 1252.6200 2743.2800 ;
        RECT 1251.0200 2748.2400 1252.6200 2748.7200 ;
        RECT 1206.0200 2753.6800 1207.6200 2754.1600 ;
        RECT 1206.0200 2759.1200 1207.6200 2759.6000 ;
        RECT 1206.0200 2737.3600 1207.6200 2737.8400 ;
        RECT 1206.0200 2742.8000 1207.6200 2743.2800 ;
        RECT 1206.0200 2748.2400 1207.6200 2748.7200 ;
        RECT 1251.0200 2726.4800 1252.6200 2726.9600 ;
        RECT 1251.0200 2731.9200 1252.6200 2732.4000 ;
        RECT 1251.0200 2710.1600 1252.6200 2710.6400 ;
        RECT 1251.0200 2715.6000 1252.6200 2716.0800 ;
        RECT 1251.0200 2721.0400 1252.6200 2721.5200 ;
        RECT 1206.0200 2726.4800 1207.6200 2726.9600 ;
        RECT 1206.0200 2731.9200 1207.6200 2732.4000 ;
        RECT 1206.0200 2710.1600 1207.6200 2710.6400 ;
        RECT 1206.0200 2715.6000 1207.6200 2716.0800 ;
        RECT 1206.0200 2721.0400 1207.6200 2721.5200 ;
        RECT 1156.4600 2753.6800 1159.4600 2754.1600 ;
        RECT 1156.4600 2759.1200 1159.4600 2759.6000 ;
        RECT 1156.4600 2742.8000 1159.4600 2743.2800 ;
        RECT 1156.4600 2737.3600 1159.4600 2737.8400 ;
        RECT 1156.4600 2748.2400 1159.4600 2748.7200 ;
        RECT 1156.4600 2726.4800 1159.4600 2726.9600 ;
        RECT 1156.4600 2731.9200 1159.4600 2732.4000 ;
        RECT 1156.4600 2715.6000 1159.4600 2716.0800 ;
        RECT 1156.4600 2710.1600 1159.4600 2710.6400 ;
        RECT 1156.4600 2721.0400 1159.4600 2721.5200 ;
        RECT 1156.4600 2764.5600 1159.4600 2765.0400 ;
        RECT 1206.0200 2764.5600 1207.6200 2765.0400 ;
        RECT 1251.0200 2764.5600 1252.6200 2765.0400 ;
        RECT 1352.5600 2699.2800 1355.5600 2699.7600 ;
        RECT 1352.5600 2704.7200 1355.5600 2705.2000 ;
        RECT 1341.0200 2699.2800 1342.6200 2699.7600 ;
        RECT 1341.0200 2704.7200 1342.6200 2705.2000 ;
        RECT 1352.5600 2682.9600 1355.5600 2683.4400 ;
        RECT 1352.5600 2688.4000 1355.5600 2688.8800 ;
        RECT 1352.5600 2693.8400 1355.5600 2694.3200 ;
        RECT 1341.0200 2682.9600 1342.6200 2683.4400 ;
        RECT 1341.0200 2688.4000 1342.6200 2688.8800 ;
        RECT 1341.0200 2693.8400 1342.6200 2694.3200 ;
        RECT 1352.5600 2672.0800 1355.5600 2672.5600 ;
        RECT 1352.5600 2677.5200 1355.5600 2678.0000 ;
        RECT 1341.0200 2672.0800 1342.6200 2672.5600 ;
        RECT 1341.0200 2677.5200 1342.6200 2678.0000 ;
        RECT 1352.5600 2655.7600 1355.5600 2656.2400 ;
        RECT 1352.5600 2661.2000 1355.5600 2661.6800 ;
        RECT 1352.5600 2666.6400 1355.5600 2667.1200 ;
        RECT 1341.0200 2655.7600 1342.6200 2656.2400 ;
        RECT 1341.0200 2661.2000 1342.6200 2661.6800 ;
        RECT 1341.0200 2666.6400 1342.6200 2667.1200 ;
        RECT 1296.0200 2699.2800 1297.6200 2699.7600 ;
        RECT 1296.0200 2704.7200 1297.6200 2705.2000 ;
        RECT 1296.0200 2682.9600 1297.6200 2683.4400 ;
        RECT 1296.0200 2688.4000 1297.6200 2688.8800 ;
        RECT 1296.0200 2693.8400 1297.6200 2694.3200 ;
        RECT 1296.0200 2672.0800 1297.6200 2672.5600 ;
        RECT 1296.0200 2677.5200 1297.6200 2678.0000 ;
        RECT 1296.0200 2655.7600 1297.6200 2656.2400 ;
        RECT 1296.0200 2661.2000 1297.6200 2661.6800 ;
        RECT 1296.0200 2666.6400 1297.6200 2667.1200 ;
        RECT 1352.5600 2644.8800 1355.5600 2645.3600 ;
        RECT 1352.5600 2650.3200 1355.5600 2650.8000 ;
        RECT 1341.0200 2644.8800 1342.6200 2645.3600 ;
        RECT 1341.0200 2650.3200 1342.6200 2650.8000 ;
        RECT 1352.5600 2628.5600 1355.5600 2629.0400 ;
        RECT 1352.5600 2634.0000 1355.5600 2634.4800 ;
        RECT 1352.5600 2639.4400 1355.5600 2639.9200 ;
        RECT 1341.0200 2628.5600 1342.6200 2629.0400 ;
        RECT 1341.0200 2634.0000 1342.6200 2634.4800 ;
        RECT 1341.0200 2639.4400 1342.6200 2639.9200 ;
        RECT 1352.5600 2617.6800 1355.5600 2618.1600 ;
        RECT 1352.5600 2623.1200 1355.5600 2623.6000 ;
        RECT 1341.0200 2617.6800 1342.6200 2618.1600 ;
        RECT 1341.0200 2623.1200 1342.6200 2623.6000 ;
        RECT 1352.5600 2612.2400 1355.5600 2612.7200 ;
        RECT 1341.0200 2612.2400 1342.6200 2612.7200 ;
        RECT 1296.0200 2644.8800 1297.6200 2645.3600 ;
        RECT 1296.0200 2650.3200 1297.6200 2650.8000 ;
        RECT 1296.0200 2628.5600 1297.6200 2629.0400 ;
        RECT 1296.0200 2634.0000 1297.6200 2634.4800 ;
        RECT 1296.0200 2639.4400 1297.6200 2639.9200 ;
        RECT 1296.0200 2617.6800 1297.6200 2618.1600 ;
        RECT 1296.0200 2623.1200 1297.6200 2623.6000 ;
        RECT 1296.0200 2612.2400 1297.6200 2612.7200 ;
        RECT 1251.0200 2699.2800 1252.6200 2699.7600 ;
        RECT 1251.0200 2704.7200 1252.6200 2705.2000 ;
        RECT 1251.0200 2682.9600 1252.6200 2683.4400 ;
        RECT 1251.0200 2688.4000 1252.6200 2688.8800 ;
        RECT 1251.0200 2693.8400 1252.6200 2694.3200 ;
        RECT 1206.0200 2699.2800 1207.6200 2699.7600 ;
        RECT 1206.0200 2704.7200 1207.6200 2705.2000 ;
        RECT 1206.0200 2682.9600 1207.6200 2683.4400 ;
        RECT 1206.0200 2688.4000 1207.6200 2688.8800 ;
        RECT 1206.0200 2693.8400 1207.6200 2694.3200 ;
        RECT 1251.0200 2672.0800 1252.6200 2672.5600 ;
        RECT 1251.0200 2677.5200 1252.6200 2678.0000 ;
        RECT 1251.0200 2655.7600 1252.6200 2656.2400 ;
        RECT 1251.0200 2661.2000 1252.6200 2661.6800 ;
        RECT 1251.0200 2666.6400 1252.6200 2667.1200 ;
        RECT 1206.0200 2672.0800 1207.6200 2672.5600 ;
        RECT 1206.0200 2677.5200 1207.6200 2678.0000 ;
        RECT 1206.0200 2655.7600 1207.6200 2656.2400 ;
        RECT 1206.0200 2661.2000 1207.6200 2661.6800 ;
        RECT 1206.0200 2666.6400 1207.6200 2667.1200 ;
        RECT 1156.4600 2699.2800 1159.4600 2699.7600 ;
        RECT 1156.4600 2704.7200 1159.4600 2705.2000 ;
        RECT 1156.4600 2688.4000 1159.4600 2688.8800 ;
        RECT 1156.4600 2682.9600 1159.4600 2683.4400 ;
        RECT 1156.4600 2693.8400 1159.4600 2694.3200 ;
        RECT 1156.4600 2672.0800 1159.4600 2672.5600 ;
        RECT 1156.4600 2677.5200 1159.4600 2678.0000 ;
        RECT 1156.4600 2661.2000 1159.4600 2661.6800 ;
        RECT 1156.4600 2655.7600 1159.4600 2656.2400 ;
        RECT 1156.4600 2666.6400 1159.4600 2667.1200 ;
        RECT 1251.0200 2644.8800 1252.6200 2645.3600 ;
        RECT 1251.0200 2650.3200 1252.6200 2650.8000 ;
        RECT 1251.0200 2628.5600 1252.6200 2629.0400 ;
        RECT 1251.0200 2634.0000 1252.6200 2634.4800 ;
        RECT 1251.0200 2639.4400 1252.6200 2639.9200 ;
        RECT 1206.0200 2644.8800 1207.6200 2645.3600 ;
        RECT 1206.0200 2650.3200 1207.6200 2650.8000 ;
        RECT 1206.0200 2628.5600 1207.6200 2629.0400 ;
        RECT 1206.0200 2634.0000 1207.6200 2634.4800 ;
        RECT 1206.0200 2639.4400 1207.6200 2639.9200 ;
        RECT 1251.0200 2623.1200 1252.6200 2623.6000 ;
        RECT 1251.0200 2617.6800 1252.6200 2618.1600 ;
        RECT 1251.0200 2612.2400 1252.6200 2612.7200 ;
        RECT 1206.0200 2623.1200 1207.6200 2623.6000 ;
        RECT 1206.0200 2617.6800 1207.6200 2618.1600 ;
        RECT 1206.0200 2612.2400 1207.6200 2612.7200 ;
        RECT 1156.4600 2644.8800 1159.4600 2645.3600 ;
        RECT 1156.4600 2650.3200 1159.4600 2650.8000 ;
        RECT 1156.4600 2634.0000 1159.4600 2634.4800 ;
        RECT 1156.4600 2628.5600 1159.4600 2629.0400 ;
        RECT 1156.4600 2639.4400 1159.4600 2639.9200 ;
        RECT 1156.4600 2617.6800 1159.4600 2618.1600 ;
        RECT 1156.4600 2623.1200 1159.4600 2623.6000 ;
        RECT 1156.4600 2612.2400 1159.4600 2612.7200 ;
        RECT 1156.4600 2810.4300 1355.5600 2813.4300 ;
        RECT 1156.4600 2605.3300 1355.5600 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 2375.6900 1342.6200 2583.7900 ;
        RECT 1296.0200 2375.6900 1297.6200 2583.7900 ;
        RECT 1251.0200 2375.6900 1252.6200 2583.7900 ;
        RECT 1206.0200 2375.6900 1207.6200 2583.7900 ;
        RECT 1352.5600 2375.6900 1355.5600 2583.7900 ;
        RECT 1156.4600 2375.6900 1159.4600 2583.7900 ;
      LAYER met3 ;
        RECT 1352.5600 2578.4400 1355.5600 2578.9200 ;
        RECT 1341.0200 2578.4400 1342.6200 2578.9200 ;
        RECT 1352.5600 2567.5600 1355.5600 2568.0400 ;
        RECT 1352.5600 2573.0000 1355.5600 2573.4800 ;
        RECT 1341.0200 2567.5600 1342.6200 2568.0400 ;
        RECT 1341.0200 2573.0000 1342.6200 2573.4800 ;
        RECT 1352.5600 2551.2400 1355.5600 2551.7200 ;
        RECT 1352.5600 2556.6800 1355.5600 2557.1600 ;
        RECT 1341.0200 2551.2400 1342.6200 2551.7200 ;
        RECT 1341.0200 2556.6800 1342.6200 2557.1600 ;
        RECT 1352.5600 2540.3600 1355.5600 2540.8400 ;
        RECT 1352.5600 2545.8000 1355.5600 2546.2800 ;
        RECT 1341.0200 2540.3600 1342.6200 2540.8400 ;
        RECT 1341.0200 2545.8000 1342.6200 2546.2800 ;
        RECT 1352.5600 2562.1200 1355.5600 2562.6000 ;
        RECT 1341.0200 2562.1200 1342.6200 2562.6000 ;
        RECT 1296.0200 2567.5600 1297.6200 2568.0400 ;
        RECT 1296.0200 2573.0000 1297.6200 2573.4800 ;
        RECT 1296.0200 2578.4400 1297.6200 2578.9200 ;
        RECT 1296.0200 2551.2400 1297.6200 2551.7200 ;
        RECT 1296.0200 2556.6800 1297.6200 2557.1600 ;
        RECT 1296.0200 2545.8000 1297.6200 2546.2800 ;
        RECT 1296.0200 2540.3600 1297.6200 2540.8400 ;
        RECT 1296.0200 2562.1200 1297.6200 2562.6000 ;
        RECT 1352.5600 2524.0400 1355.5600 2524.5200 ;
        RECT 1352.5600 2529.4800 1355.5600 2529.9600 ;
        RECT 1341.0200 2524.0400 1342.6200 2524.5200 ;
        RECT 1341.0200 2529.4800 1342.6200 2529.9600 ;
        RECT 1352.5600 2507.7200 1355.5600 2508.2000 ;
        RECT 1352.5600 2513.1600 1355.5600 2513.6400 ;
        RECT 1352.5600 2518.6000 1355.5600 2519.0800 ;
        RECT 1341.0200 2507.7200 1342.6200 2508.2000 ;
        RECT 1341.0200 2513.1600 1342.6200 2513.6400 ;
        RECT 1341.0200 2518.6000 1342.6200 2519.0800 ;
        RECT 1352.5600 2496.8400 1355.5600 2497.3200 ;
        RECT 1352.5600 2502.2800 1355.5600 2502.7600 ;
        RECT 1341.0200 2496.8400 1342.6200 2497.3200 ;
        RECT 1341.0200 2502.2800 1342.6200 2502.7600 ;
        RECT 1352.5600 2480.5200 1355.5600 2481.0000 ;
        RECT 1352.5600 2485.9600 1355.5600 2486.4400 ;
        RECT 1352.5600 2491.4000 1355.5600 2491.8800 ;
        RECT 1341.0200 2480.5200 1342.6200 2481.0000 ;
        RECT 1341.0200 2485.9600 1342.6200 2486.4400 ;
        RECT 1341.0200 2491.4000 1342.6200 2491.8800 ;
        RECT 1296.0200 2524.0400 1297.6200 2524.5200 ;
        RECT 1296.0200 2529.4800 1297.6200 2529.9600 ;
        RECT 1296.0200 2507.7200 1297.6200 2508.2000 ;
        RECT 1296.0200 2513.1600 1297.6200 2513.6400 ;
        RECT 1296.0200 2518.6000 1297.6200 2519.0800 ;
        RECT 1296.0200 2496.8400 1297.6200 2497.3200 ;
        RECT 1296.0200 2502.2800 1297.6200 2502.7600 ;
        RECT 1296.0200 2480.5200 1297.6200 2481.0000 ;
        RECT 1296.0200 2485.9600 1297.6200 2486.4400 ;
        RECT 1296.0200 2491.4000 1297.6200 2491.8800 ;
        RECT 1352.5600 2534.9200 1355.5600 2535.4000 ;
        RECT 1296.0200 2534.9200 1297.6200 2535.4000 ;
        RECT 1341.0200 2534.9200 1342.6200 2535.4000 ;
        RECT 1251.0200 2567.5600 1252.6200 2568.0400 ;
        RECT 1251.0200 2573.0000 1252.6200 2573.4800 ;
        RECT 1251.0200 2578.4400 1252.6200 2578.9200 ;
        RECT 1206.0200 2567.5600 1207.6200 2568.0400 ;
        RECT 1206.0200 2573.0000 1207.6200 2573.4800 ;
        RECT 1206.0200 2578.4400 1207.6200 2578.9200 ;
        RECT 1251.0200 2551.2400 1252.6200 2551.7200 ;
        RECT 1251.0200 2556.6800 1252.6200 2557.1600 ;
        RECT 1251.0200 2540.3600 1252.6200 2540.8400 ;
        RECT 1251.0200 2545.8000 1252.6200 2546.2800 ;
        RECT 1206.0200 2551.2400 1207.6200 2551.7200 ;
        RECT 1206.0200 2556.6800 1207.6200 2557.1600 ;
        RECT 1206.0200 2540.3600 1207.6200 2540.8400 ;
        RECT 1206.0200 2545.8000 1207.6200 2546.2800 ;
        RECT 1206.0200 2562.1200 1207.6200 2562.6000 ;
        RECT 1251.0200 2562.1200 1252.6200 2562.6000 ;
        RECT 1156.4600 2578.4400 1159.4600 2578.9200 ;
        RECT 1156.4600 2573.0000 1159.4600 2573.4800 ;
        RECT 1156.4600 2567.5600 1159.4600 2568.0400 ;
        RECT 1156.4600 2556.6800 1159.4600 2557.1600 ;
        RECT 1156.4600 2551.2400 1159.4600 2551.7200 ;
        RECT 1156.4600 2545.8000 1159.4600 2546.2800 ;
        RECT 1156.4600 2540.3600 1159.4600 2540.8400 ;
        RECT 1156.4600 2562.1200 1159.4600 2562.6000 ;
        RECT 1251.0200 2524.0400 1252.6200 2524.5200 ;
        RECT 1251.0200 2529.4800 1252.6200 2529.9600 ;
        RECT 1251.0200 2507.7200 1252.6200 2508.2000 ;
        RECT 1251.0200 2513.1600 1252.6200 2513.6400 ;
        RECT 1251.0200 2518.6000 1252.6200 2519.0800 ;
        RECT 1206.0200 2524.0400 1207.6200 2524.5200 ;
        RECT 1206.0200 2529.4800 1207.6200 2529.9600 ;
        RECT 1206.0200 2507.7200 1207.6200 2508.2000 ;
        RECT 1206.0200 2513.1600 1207.6200 2513.6400 ;
        RECT 1206.0200 2518.6000 1207.6200 2519.0800 ;
        RECT 1251.0200 2496.8400 1252.6200 2497.3200 ;
        RECT 1251.0200 2502.2800 1252.6200 2502.7600 ;
        RECT 1251.0200 2480.5200 1252.6200 2481.0000 ;
        RECT 1251.0200 2485.9600 1252.6200 2486.4400 ;
        RECT 1251.0200 2491.4000 1252.6200 2491.8800 ;
        RECT 1206.0200 2496.8400 1207.6200 2497.3200 ;
        RECT 1206.0200 2502.2800 1207.6200 2502.7600 ;
        RECT 1206.0200 2480.5200 1207.6200 2481.0000 ;
        RECT 1206.0200 2485.9600 1207.6200 2486.4400 ;
        RECT 1206.0200 2491.4000 1207.6200 2491.8800 ;
        RECT 1156.4600 2524.0400 1159.4600 2524.5200 ;
        RECT 1156.4600 2529.4800 1159.4600 2529.9600 ;
        RECT 1156.4600 2513.1600 1159.4600 2513.6400 ;
        RECT 1156.4600 2507.7200 1159.4600 2508.2000 ;
        RECT 1156.4600 2518.6000 1159.4600 2519.0800 ;
        RECT 1156.4600 2496.8400 1159.4600 2497.3200 ;
        RECT 1156.4600 2502.2800 1159.4600 2502.7600 ;
        RECT 1156.4600 2485.9600 1159.4600 2486.4400 ;
        RECT 1156.4600 2480.5200 1159.4600 2481.0000 ;
        RECT 1156.4600 2491.4000 1159.4600 2491.8800 ;
        RECT 1156.4600 2534.9200 1159.4600 2535.4000 ;
        RECT 1206.0200 2534.9200 1207.6200 2535.4000 ;
        RECT 1251.0200 2534.9200 1252.6200 2535.4000 ;
        RECT 1352.5600 2469.6400 1355.5600 2470.1200 ;
        RECT 1352.5600 2475.0800 1355.5600 2475.5600 ;
        RECT 1341.0200 2469.6400 1342.6200 2470.1200 ;
        RECT 1341.0200 2475.0800 1342.6200 2475.5600 ;
        RECT 1352.5600 2453.3200 1355.5600 2453.8000 ;
        RECT 1352.5600 2458.7600 1355.5600 2459.2400 ;
        RECT 1352.5600 2464.2000 1355.5600 2464.6800 ;
        RECT 1341.0200 2453.3200 1342.6200 2453.8000 ;
        RECT 1341.0200 2458.7600 1342.6200 2459.2400 ;
        RECT 1341.0200 2464.2000 1342.6200 2464.6800 ;
        RECT 1352.5600 2442.4400 1355.5600 2442.9200 ;
        RECT 1352.5600 2447.8800 1355.5600 2448.3600 ;
        RECT 1341.0200 2442.4400 1342.6200 2442.9200 ;
        RECT 1341.0200 2447.8800 1342.6200 2448.3600 ;
        RECT 1352.5600 2426.1200 1355.5600 2426.6000 ;
        RECT 1352.5600 2431.5600 1355.5600 2432.0400 ;
        RECT 1352.5600 2437.0000 1355.5600 2437.4800 ;
        RECT 1341.0200 2426.1200 1342.6200 2426.6000 ;
        RECT 1341.0200 2431.5600 1342.6200 2432.0400 ;
        RECT 1341.0200 2437.0000 1342.6200 2437.4800 ;
        RECT 1296.0200 2469.6400 1297.6200 2470.1200 ;
        RECT 1296.0200 2475.0800 1297.6200 2475.5600 ;
        RECT 1296.0200 2453.3200 1297.6200 2453.8000 ;
        RECT 1296.0200 2458.7600 1297.6200 2459.2400 ;
        RECT 1296.0200 2464.2000 1297.6200 2464.6800 ;
        RECT 1296.0200 2442.4400 1297.6200 2442.9200 ;
        RECT 1296.0200 2447.8800 1297.6200 2448.3600 ;
        RECT 1296.0200 2426.1200 1297.6200 2426.6000 ;
        RECT 1296.0200 2431.5600 1297.6200 2432.0400 ;
        RECT 1296.0200 2437.0000 1297.6200 2437.4800 ;
        RECT 1352.5600 2415.2400 1355.5600 2415.7200 ;
        RECT 1352.5600 2420.6800 1355.5600 2421.1600 ;
        RECT 1341.0200 2415.2400 1342.6200 2415.7200 ;
        RECT 1341.0200 2420.6800 1342.6200 2421.1600 ;
        RECT 1352.5600 2398.9200 1355.5600 2399.4000 ;
        RECT 1352.5600 2404.3600 1355.5600 2404.8400 ;
        RECT 1352.5600 2409.8000 1355.5600 2410.2800 ;
        RECT 1341.0200 2398.9200 1342.6200 2399.4000 ;
        RECT 1341.0200 2404.3600 1342.6200 2404.8400 ;
        RECT 1341.0200 2409.8000 1342.6200 2410.2800 ;
        RECT 1352.5600 2388.0400 1355.5600 2388.5200 ;
        RECT 1352.5600 2393.4800 1355.5600 2393.9600 ;
        RECT 1341.0200 2388.0400 1342.6200 2388.5200 ;
        RECT 1341.0200 2393.4800 1342.6200 2393.9600 ;
        RECT 1352.5600 2382.6000 1355.5600 2383.0800 ;
        RECT 1341.0200 2382.6000 1342.6200 2383.0800 ;
        RECT 1296.0200 2415.2400 1297.6200 2415.7200 ;
        RECT 1296.0200 2420.6800 1297.6200 2421.1600 ;
        RECT 1296.0200 2398.9200 1297.6200 2399.4000 ;
        RECT 1296.0200 2404.3600 1297.6200 2404.8400 ;
        RECT 1296.0200 2409.8000 1297.6200 2410.2800 ;
        RECT 1296.0200 2388.0400 1297.6200 2388.5200 ;
        RECT 1296.0200 2393.4800 1297.6200 2393.9600 ;
        RECT 1296.0200 2382.6000 1297.6200 2383.0800 ;
        RECT 1251.0200 2469.6400 1252.6200 2470.1200 ;
        RECT 1251.0200 2475.0800 1252.6200 2475.5600 ;
        RECT 1251.0200 2453.3200 1252.6200 2453.8000 ;
        RECT 1251.0200 2458.7600 1252.6200 2459.2400 ;
        RECT 1251.0200 2464.2000 1252.6200 2464.6800 ;
        RECT 1206.0200 2469.6400 1207.6200 2470.1200 ;
        RECT 1206.0200 2475.0800 1207.6200 2475.5600 ;
        RECT 1206.0200 2453.3200 1207.6200 2453.8000 ;
        RECT 1206.0200 2458.7600 1207.6200 2459.2400 ;
        RECT 1206.0200 2464.2000 1207.6200 2464.6800 ;
        RECT 1251.0200 2442.4400 1252.6200 2442.9200 ;
        RECT 1251.0200 2447.8800 1252.6200 2448.3600 ;
        RECT 1251.0200 2426.1200 1252.6200 2426.6000 ;
        RECT 1251.0200 2431.5600 1252.6200 2432.0400 ;
        RECT 1251.0200 2437.0000 1252.6200 2437.4800 ;
        RECT 1206.0200 2442.4400 1207.6200 2442.9200 ;
        RECT 1206.0200 2447.8800 1207.6200 2448.3600 ;
        RECT 1206.0200 2426.1200 1207.6200 2426.6000 ;
        RECT 1206.0200 2431.5600 1207.6200 2432.0400 ;
        RECT 1206.0200 2437.0000 1207.6200 2437.4800 ;
        RECT 1156.4600 2469.6400 1159.4600 2470.1200 ;
        RECT 1156.4600 2475.0800 1159.4600 2475.5600 ;
        RECT 1156.4600 2458.7600 1159.4600 2459.2400 ;
        RECT 1156.4600 2453.3200 1159.4600 2453.8000 ;
        RECT 1156.4600 2464.2000 1159.4600 2464.6800 ;
        RECT 1156.4600 2442.4400 1159.4600 2442.9200 ;
        RECT 1156.4600 2447.8800 1159.4600 2448.3600 ;
        RECT 1156.4600 2431.5600 1159.4600 2432.0400 ;
        RECT 1156.4600 2426.1200 1159.4600 2426.6000 ;
        RECT 1156.4600 2437.0000 1159.4600 2437.4800 ;
        RECT 1251.0200 2415.2400 1252.6200 2415.7200 ;
        RECT 1251.0200 2420.6800 1252.6200 2421.1600 ;
        RECT 1251.0200 2398.9200 1252.6200 2399.4000 ;
        RECT 1251.0200 2404.3600 1252.6200 2404.8400 ;
        RECT 1251.0200 2409.8000 1252.6200 2410.2800 ;
        RECT 1206.0200 2415.2400 1207.6200 2415.7200 ;
        RECT 1206.0200 2420.6800 1207.6200 2421.1600 ;
        RECT 1206.0200 2398.9200 1207.6200 2399.4000 ;
        RECT 1206.0200 2404.3600 1207.6200 2404.8400 ;
        RECT 1206.0200 2409.8000 1207.6200 2410.2800 ;
        RECT 1251.0200 2393.4800 1252.6200 2393.9600 ;
        RECT 1251.0200 2388.0400 1252.6200 2388.5200 ;
        RECT 1251.0200 2382.6000 1252.6200 2383.0800 ;
        RECT 1206.0200 2393.4800 1207.6200 2393.9600 ;
        RECT 1206.0200 2388.0400 1207.6200 2388.5200 ;
        RECT 1206.0200 2382.6000 1207.6200 2383.0800 ;
        RECT 1156.4600 2415.2400 1159.4600 2415.7200 ;
        RECT 1156.4600 2420.6800 1159.4600 2421.1600 ;
        RECT 1156.4600 2404.3600 1159.4600 2404.8400 ;
        RECT 1156.4600 2398.9200 1159.4600 2399.4000 ;
        RECT 1156.4600 2409.8000 1159.4600 2410.2800 ;
        RECT 1156.4600 2388.0400 1159.4600 2388.5200 ;
        RECT 1156.4600 2393.4800 1159.4600 2393.9600 ;
        RECT 1156.4600 2382.6000 1159.4600 2383.0800 ;
        RECT 1156.4600 2580.7900 1355.5600 2583.7900 ;
        RECT 1156.4600 2375.6900 1355.5600 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 2146.0500 1342.6200 2354.1500 ;
        RECT 1296.0200 2146.0500 1297.6200 2354.1500 ;
        RECT 1251.0200 2146.0500 1252.6200 2354.1500 ;
        RECT 1206.0200 2146.0500 1207.6200 2354.1500 ;
        RECT 1352.5600 2146.0500 1355.5600 2354.1500 ;
        RECT 1156.4600 2146.0500 1159.4600 2354.1500 ;
      LAYER met3 ;
        RECT 1352.5600 2348.8000 1355.5600 2349.2800 ;
        RECT 1341.0200 2348.8000 1342.6200 2349.2800 ;
        RECT 1352.5600 2337.9200 1355.5600 2338.4000 ;
        RECT 1352.5600 2343.3600 1355.5600 2343.8400 ;
        RECT 1341.0200 2337.9200 1342.6200 2338.4000 ;
        RECT 1341.0200 2343.3600 1342.6200 2343.8400 ;
        RECT 1352.5600 2321.6000 1355.5600 2322.0800 ;
        RECT 1352.5600 2327.0400 1355.5600 2327.5200 ;
        RECT 1341.0200 2321.6000 1342.6200 2322.0800 ;
        RECT 1341.0200 2327.0400 1342.6200 2327.5200 ;
        RECT 1352.5600 2310.7200 1355.5600 2311.2000 ;
        RECT 1352.5600 2316.1600 1355.5600 2316.6400 ;
        RECT 1341.0200 2310.7200 1342.6200 2311.2000 ;
        RECT 1341.0200 2316.1600 1342.6200 2316.6400 ;
        RECT 1352.5600 2332.4800 1355.5600 2332.9600 ;
        RECT 1341.0200 2332.4800 1342.6200 2332.9600 ;
        RECT 1296.0200 2337.9200 1297.6200 2338.4000 ;
        RECT 1296.0200 2343.3600 1297.6200 2343.8400 ;
        RECT 1296.0200 2348.8000 1297.6200 2349.2800 ;
        RECT 1296.0200 2321.6000 1297.6200 2322.0800 ;
        RECT 1296.0200 2327.0400 1297.6200 2327.5200 ;
        RECT 1296.0200 2316.1600 1297.6200 2316.6400 ;
        RECT 1296.0200 2310.7200 1297.6200 2311.2000 ;
        RECT 1296.0200 2332.4800 1297.6200 2332.9600 ;
        RECT 1352.5600 2294.4000 1355.5600 2294.8800 ;
        RECT 1352.5600 2299.8400 1355.5600 2300.3200 ;
        RECT 1341.0200 2294.4000 1342.6200 2294.8800 ;
        RECT 1341.0200 2299.8400 1342.6200 2300.3200 ;
        RECT 1352.5600 2278.0800 1355.5600 2278.5600 ;
        RECT 1352.5600 2283.5200 1355.5600 2284.0000 ;
        RECT 1352.5600 2288.9600 1355.5600 2289.4400 ;
        RECT 1341.0200 2278.0800 1342.6200 2278.5600 ;
        RECT 1341.0200 2283.5200 1342.6200 2284.0000 ;
        RECT 1341.0200 2288.9600 1342.6200 2289.4400 ;
        RECT 1352.5600 2267.2000 1355.5600 2267.6800 ;
        RECT 1352.5600 2272.6400 1355.5600 2273.1200 ;
        RECT 1341.0200 2267.2000 1342.6200 2267.6800 ;
        RECT 1341.0200 2272.6400 1342.6200 2273.1200 ;
        RECT 1352.5600 2250.8800 1355.5600 2251.3600 ;
        RECT 1352.5600 2256.3200 1355.5600 2256.8000 ;
        RECT 1352.5600 2261.7600 1355.5600 2262.2400 ;
        RECT 1341.0200 2250.8800 1342.6200 2251.3600 ;
        RECT 1341.0200 2256.3200 1342.6200 2256.8000 ;
        RECT 1341.0200 2261.7600 1342.6200 2262.2400 ;
        RECT 1296.0200 2294.4000 1297.6200 2294.8800 ;
        RECT 1296.0200 2299.8400 1297.6200 2300.3200 ;
        RECT 1296.0200 2278.0800 1297.6200 2278.5600 ;
        RECT 1296.0200 2283.5200 1297.6200 2284.0000 ;
        RECT 1296.0200 2288.9600 1297.6200 2289.4400 ;
        RECT 1296.0200 2267.2000 1297.6200 2267.6800 ;
        RECT 1296.0200 2272.6400 1297.6200 2273.1200 ;
        RECT 1296.0200 2250.8800 1297.6200 2251.3600 ;
        RECT 1296.0200 2256.3200 1297.6200 2256.8000 ;
        RECT 1296.0200 2261.7600 1297.6200 2262.2400 ;
        RECT 1352.5600 2305.2800 1355.5600 2305.7600 ;
        RECT 1296.0200 2305.2800 1297.6200 2305.7600 ;
        RECT 1341.0200 2305.2800 1342.6200 2305.7600 ;
        RECT 1251.0200 2337.9200 1252.6200 2338.4000 ;
        RECT 1251.0200 2343.3600 1252.6200 2343.8400 ;
        RECT 1251.0200 2348.8000 1252.6200 2349.2800 ;
        RECT 1206.0200 2337.9200 1207.6200 2338.4000 ;
        RECT 1206.0200 2343.3600 1207.6200 2343.8400 ;
        RECT 1206.0200 2348.8000 1207.6200 2349.2800 ;
        RECT 1251.0200 2321.6000 1252.6200 2322.0800 ;
        RECT 1251.0200 2327.0400 1252.6200 2327.5200 ;
        RECT 1251.0200 2310.7200 1252.6200 2311.2000 ;
        RECT 1251.0200 2316.1600 1252.6200 2316.6400 ;
        RECT 1206.0200 2321.6000 1207.6200 2322.0800 ;
        RECT 1206.0200 2327.0400 1207.6200 2327.5200 ;
        RECT 1206.0200 2310.7200 1207.6200 2311.2000 ;
        RECT 1206.0200 2316.1600 1207.6200 2316.6400 ;
        RECT 1206.0200 2332.4800 1207.6200 2332.9600 ;
        RECT 1251.0200 2332.4800 1252.6200 2332.9600 ;
        RECT 1156.4600 2348.8000 1159.4600 2349.2800 ;
        RECT 1156.4600 2343.3600 1159.4600 2343.8400 ;
        RECT 1156.4600 2337.9200 1159.4600 2338.4000 ;
        RECT 1156.4600 2327.0400 1159.4600 2327.5200 ;
        RECT 1156.4600 2321.6000 1159.4600 2322.0800 ;
        RECT 1156.4600 2316.1600 1159.4600 2316.6400 ;
        RECT 1156.4600 2310.7200 1159.4600 2311.2000 ;
        RECT 1156.4600 2332.4800 1159.4600 2332.9600 ;
        RECT 1251.0200 2294.4000 1252.6200 2294.8800 ;
        RECT 1251.0200 2299.8400 1252.6200 2300.3200 ;
        RECT 1251.0200 2278.0800 1252.6200 2278.5600 ;
        RECT 1251.0200 2283.5200 1252.6200 2284.0000 ;
        RECT 1251.0200 2288.9600 1252.6200 2289.4400 ;
        RECT 1206.0200 2294.4000 1207.6200 2294.8800 ;
        RECT 1206.0200 2299.8400 1207.6200 2300.3200 ;
        RECT 1206.0200 2278.0800 1207.6200 2278.5600 ;
        RECT 1206.0200 2283.5200 1207.6200 2284.0000 ;
        RECT 1206.0200 2288.9600 1207.6200 2289.4400 ;
        RECT 1251.0200 2267.2000 1252.6200 2267.6800 ;
        RECT 1251.0200 2272.6400 1252.6200 2273.1200 ;
        RECT 1251.0200 2250.8800 1252.6200 2251.3600 ;
        RECT 1251.0200 2256.3200 1252.6200 2256.8000 ;
        RECT 1251.0200 2261.7600 1252.6200 2262.2400 ;
        RECT 1206.0200 2267.2000 1207.6200 2267.6800 ;
        RECT 1206.0200 2272.6400 1207.6200 2273.1200 ;
        RECT 1206.0200 2250.8800 1207.6200 2251.3600 ;
        RECT 1206.0200 2256.3200 1207.6200 2256.8000 ;
        RECT 1206.0200 2261.7600 1207.6200 2262.2400 ;
        RECT 1156.4600 2294.4000 1159.4600 2294.8800 ;
        RECT 1156.4600 2299.8400 1159.4600 2300.3200 ;
        RECT 1156.4600 2283.5200 1159.4600 2284.0000 ;
        RECT 1156.4600 2278.0800 1159.4600 2278.5600 ;
        RECT 1156.4600 2288.9600 1159.4600 2289.4400 ;
        RECT 1156.4600 2267.2000 1159.4600 2267.6800 ;
        RECT 1156.4600 2272.6400 1159.4600 2273.1200 ;
        RECT 1156.4600 2256.3200 1159.4600 2256.8000 ;
        RECT 1156.4600 2250.8800 1159.4600 2251.3600 ;
        RECT 1156.4600 2261.7600 1159.4600 2262.2400 ;
        RECT 1156.4600 2305.2800 1159.4600 2305.7600 ;
        RECT 1206.0200 2305.2800 1207.6200 2305.7600 ;
        RECT 1251.0200 2305.2800 1252.6200 2305.7600 ;
        RECT 1352.5600 2240.0000 1355.5600 2240.4800 ;
        RECT 1352.5600 2245.4400 1355.5600 2245.9200 ;
        RECT 1341.0200 2240.0000 1342.6200 2240.4800 ;
        RECT 1341.0200 2245.4400 1342.6200 2245.9200 ;
        RECT 1352.5600 2223.6800 1355.5600 2224.1600 ;
        RECT 1352.5600 2229.1200 1355.5600 2229.6000 ;
        RECT 1352.5600 2234.5600 1355.5600 2235.0400 ;
        RECT 1341.0200 2223.6800 1342.6200 2224.1600 ;
        RECT 1341.0200 2229.1200 1342.6200 2229.6000 ;
        RECT 1341.0200 2234.5600 1342.6200 2235.0400 ;
        RECT 1352.5600 2212.8000 1355.5600 2213.2800 ;
        RECT 1352.5600 2218.2400 1355.5600 2218.7200 ;
        RECT 1341.0200 2212.8000 1342.6200 2213.2800 ;
        RECT 1341.0200 2218.2400 1342.6200 2218.7200 ;
        RECT 1352.5600 2196.4800 1355.5600 2196.9600 ;
        RECT 1352.5600 2201.9200 1355.5600 2202.4000 ;
        RECT 1352.5600 2207.3600 1355.5600 2207.8400 ;
        RECT 1341.0200 2196.4800 1342.6200 2196.9600 ;
        RECT 1341.0200 2201.9200 1342.6200 2202.4000 ;
        RECT 1341.0200 2207.3600 1342.6200 2207.8400 ;
        RECT 1296.0200 2240.0000 1297.6200 2240.4800 ;
        RECT 1296.0200 2245.4400 1297.6200 2245.9200 ;
        RECT 1296.0200 2223.6800 1297.6200 2224.1600 ;
        RECT 1296.0200 2229.1200 1297.6200 2229.6000 ;
        RECT 1296.0200 2234.5600 1297.6200 2235.0400 ;
        RECT 1296.0200 2212.8000 1297.6200 2213.2800 ;
        RECT 1296.0200 2218.2400 1297.6200 2218.7200 ;
        RECT 1296.0200 2196.4800 1297.6200 2196.9600 ;
        RECT 1296.0200 2201.9200 1297.6200 2202.4000 ;
        RECT 1296.0200 2207.3600 1297.6200 2207.8400 ;
        RECT 1352.5600 2185.6000 1355.5600 2186.0800 ;
        RECT 1352.5600 2191.0400 1355.5600 2191.5200 ;
        RECT 1341.0200 2185.6000 1342.6200 2186.0800 ;
        RECT 1341.0200 2191.0400 1342.6200 2191.5200 ;
        RECT 1352.5600 2169.2800 1355.5600 2169.7600 ;
        RECT 1352.5600 2174.7200 1355.5600 2175.2000 ;
        RECT 1352.5600 2180.1600 1355.5600 2180.6400 ;
        RECT 1341.0200 2169.2800 1342.6200 2169.7600 ;
        RECT 1341.0200 2174.7200 1342.6200 2175.2000 ;
        RECT 1341.0200 2180.1600 1342.6200 2180.6400 ;
        RECT 1352.5600 2158.4000 1355.5600 2158.8800 ;
        RECT 1352.5600 2163.8400 1355.5600 2164.3200 ;
        RECT 1341.0200 2158.4000 1342.6200 2158.8800 ;
        RECT 1341.0200 2163.8400 1342.6200 2164.3200 ;
        RECT 1352.5600 2152.9600 1355.5600 2153.4400 ;
        RECT 1341.0200 2152.9600 1342.6200 2153.4400 ;
        RECT 1296.0200 2185.6000 1297.6200 2186.0800 ;
        RECT 1296.0200 2191.0400 1297.6200 2191.5200 ;
        RECT 1296.0200 2169.2800 1297.6200 2169.7600 ;
        RECT 1296.0200 2174.7200 1297.6200 2175.2000 ;
        RECT 1296.0200 2180.1600 1297.6200 2180.6400 ;
        RECT 1296.0200 2158.4000 1297.6200 2158.8800 ;
        RECT 1296.0200 2163.8400 1297.6200 2164.3200 ;
        RECT 1296.0200 2152.9600 1297.6200 2153.4400 ;
        RECT 1251.0200 2240.0000 1252.6200 2240.4800 ;
        RECT 1251.0200 2245.4400 1252.6200 2245.9200 ;
        RECT 1251.0200 2223.6800 1252.6200 2224.1600 ;
        RECT 1251.0200 2229.1200 1252.6200 2229.6000 ;
        RECT 1251.0200 2234.5600 1252.6200 2235.0400 ;
        RECT 1206.0200 2240.0000 1207.6200 2240.4800 ;
        RECT 1206.0200 2245.4400 1207.6200 2245.9200 ;
        RECT 1206.0200 2223.6800 1207.6200 2224.1600 ;
        RECT 1206.0200 2229.1200 1207.6200 2229.6000 ;
        RECT 1206.0200 2234.5600 1207.6200 2235.0400 ;
        RECT 1251.0200 2212.8000 1252.6200 2213.2800 ;
        RECT 1251.0200 2218.2400 1252.6200 2218.7200 ;
        RECT 1251.0200 2196.4800 1252.6200 2196.9600 ;
        RECT 1251.0200 2201.9200 1252.6200 2202.4000 ;
        RECT 1251.0200 2207.3600 1252.6200 2207.8400 ;
        RECT 1206.0200 2212.8000 1207.6200 2213.2800 ;
        RECT 1206.0200 2218.2400 1207.6200 2218.7200 ;
        RECT 1206.0200 2196.4800 1207.6200 2196.9600 ;
        RECT 1206.0200 2201.9200 1207.6200 2202.4000 ;
        RECT 1206.0200 2207.3600 1207.6200 2207.8400 ;
        RECT 1156.4600 2240.0000 1159.4600 2240.4800 ;
        RECT 1156.4600 2245.4400 1159.4600 2245.9200 ;
        RECT 1156.4600 2229.1200 1159.4600 2229.6000 ;
        RECT 1156.4600 2223.6800 1159.4600 2224.1600 ;
        RECT 1156.4600 2234.5600 1159.4600 2235.0400 ;
        RECT 1156.4600 2212.8000 1159.4600 2213.2800 ;
        RECT 1156.4600 2218.2400 1159.4600 2218.7200 ;
        RECT 1156.4600 2201.9200 1159.4600 2202.4000 ;
        RECT 1156.4600 2196.4800 1159.4600 2196.9600 ;
        RECT 1156.4600 2207.3600 1159.4600 2207.8400 ;
        RECT 1251.0200 2185.6000 1252.6200 2186.0800 ;
        RECT 1251.0200 2191.0400 1252.6200 2191.5200 ;
        RECT 1251.0200 2169.2800 1252.6200 2169.7600 ;
        RECT 1251.0200 2174.7200 1252.6200 2175.2000 ;
        RECT 1251.0200 2180.1600 1252.6200 2180.6400 ;
        RECT 1206.0200 2185.6000 1207.6200 2186.0800 ;
        RECT 1206.0200 2191.0400 1207.6200 2191.5200 ;
        RECT 1206.0200 2169.2800 1207.6200 2169.7600 ;
        RECT 1206.0200 2174.7200 1207.6200 2175.2000 ;
        RECT 1206.0200 2180.1600 1207.6200 2180.6400 ;
        RECT 1251.0200 2163.8400 1252.6200 2164.3200 ;
        RECT 1251.0200 2158.4000 1252.6200 2158.8800 ;
        RECT 1251.0200 2152.9600 1252.6200 2153.4400 ;
        RECT 1206.0200 2163.8400 1207.6200 2164.3200 ;
        RECT 1206.0200 2158.4000 1207.6200 2158.8800 ;
        RECT 1206.0200 2152.9600 1207.6200 2153.4400 ;
        RECT 1156.4600 2185.6000 1159.4600 2186.0800 ;
        RECT 1156.4600 2191.0400 1159.4600 2191.5200 ;
        RECT 1156.4600 2174.7200 1159.4600 2175.2000 ;
        RECT 1156.4600 2169.2800 1159.4600 2169.7600 ;
        RECT 1156.4600 2180.1600 1159.4600 2180.6400 ;
        RECT 1156.4600 2158.4000 1159.4600 2158.8800 ;
        RECT 1156.4600 2163.8400 1159.4600 2164.3200 ;
        RECT 1156.4600 2152.9600 1159.4600 2153.4400 ;
        RECT 1156.4600 2351.1500 1355.5600 2354.1500 ;
        RECT 1156.4600 2146.0500 1355.5600 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 1916.4100 1342.6200 2124.5100 ;
        RECT 1296.0200 1916.4100 1297.6200 2124.5100 ;
        RECT 1251.0200 1916.4100 1252.6200 2124.5100 ;
        RECT 1206.0200 1916.4100 1207.6200 2124.5100 ;
        RECT 1352.5600 1916.4100 1355.5600 2124.5100 ;
        RECT 1156.4600 1916.4100 1159.4600 2124.5100 ;
      LAYER met3 ;
        RECT 1352.5600 2119.1600 1355.5600 2119.6400 ;
        RECT 1341.0200 2119.1600 1342.6200 2119.6400 ;
        RECT 1352.5600 2108.2800 1355.5600 2108.7600 ;
        RECT 1352.5600 2113.7200 1355.5600 2114.2000 ;
        RECT 1341.0200 2108.2800 1342.6200 2108.7600 ;
        RECT 1341.0200 2113.7200 1342.6200 2114.2000 ;
        RECT 1352.5600 2091.9600 1355.5600 2092.4400 ;
        RECT 1352.5600 2097.4000 1355.5600 2097.8800 ;
        RECT 1341.0200 2091.9600 1342.6200 2092.4400 ;
        RECT 1341.0200 2097.4000 1342.6200 2097.8800 ;
        RECT 1352.5600 2081.0800 1355.5600 2081.5600 ;
        RECT 1352.5600 2086.5200 1355.5600 2087.0000 ;
        RECT 1341.0200 2081.0800 1342.6200 2081.5600 ;
        RECT 1341.0200 2086.5200 1342.6200 2087.0000 ;
        RECT 1352.5600 2102.8400 1355.5600 2103.3200 ;
        RECT 1341.0200 2102.8400 1342.6200 2103.3200 ;
        RECT 1296.0200 2108.2800 1297.6200 2108.7600 ;
        RECT 1296.0200 2113.7200 1297.6200 2114.2000 ;
        RECT 1296.0200 2119.1600 1297.6200 2119.6400 ;
        RECT 1296.0200 2091.9600 1297.6200 2092.4400 ;
        RECT 1296.0200 2097.4000 1297.6200 2097.8800 ;
        RECT 1296.0200 2086.5200 1297.6200 2087.0000 ;
        RECT 1296.0200 2081.0800 1297.6200 2081.5600 ;
        RECT 1296.0200 2102.8400 1297.6200 2103.3200 ;
        RECT 1352.5600 2064.7600 1355.5600 2065.2400 ;
        RECT 1352.5600 2070.2000 1355.5600 2070.6800 ;
        RECT 1341.0200 2064.7600 1342.6200 2065.2400 ;
        RECT 1341.0200 2070.2000 1342.6200 2070.6800 ;
        RECT 1352.5600 2048.4400 1355.5600 2048.9200 ;
        RECT 1352.5600 2053.8800 1355.5600 2054.3600 ;
        RECT 1352.5600 2059.3200 1355.5600 2059.8000 ;
        RECT 1341.0200 2048.4400 1342.6200 2048.9200 ;
        RECT 1341.0200 2053.8800 1342.6200 2054.3600 ;
        RECT 1341.0200 2059.3200 1342.6200 2059.8000 ;
        RECT 1352.5600 2037.5600 1355.5600 2038.0400 ;
        RECT 1352.5600 2043.0000 1355.5600 2043.4800 ;
        RECT 1341.0200 2037.5600 1342.6200 2038.0400 ;
        RECT 1341.0200 2043.0000 1342.6200 2043.4800 ;
        RECT 1352.5600 2021.2400 1355.5600 2021.7200 ;
        RECT 1352.5600 2026.6800 1355.5600 2027.1600 ;
        RECT 1352.5600 2032.1200 1355.5600 2032.6000 ;
        RECT 1341.0200 2021.2400 1342.6200 2021.7200 ;
        RECT 1341.0200 2026.6800 1342.6200 2027.1600 ;
        RECT 1341.0200 2032.1200 1342.6200 2032.6000 ;
        RECT 1296.0200 2064.7600 1297.6200 2065.2400 ;
        RECT 1296.0200 2070.2000 1297.6200 2070.6800 ;
        RECT 1296.0200 2048.4400 1297.6200 2048.9200 ;
        RECT 1296.0200 2053.8800 1297.6200 2054.3600 ;
        RECT 1296.0200 2059.3200 1297.6200 2059.8000 ;
        RECT 1296.0200 2037.5600 1297.6200 2038.0400 ;
        RECT 1296.0200 2043.0000 1297.6200 2043.4800 ;
        RECT 1296.0200 2021.2400 1297.6200 2021.7200 ;
        RECT 1296.0200 2026.6800 1297.6200 2027.1600 ;
        RECT 1296.0200 2032.1200 1297.6200 2032.6000 ;
        RECT 1352.5600 2075.6400 1355.5600 2076.1200 ;
        RECT 1296.0200 2075.6400 1297.6200 2076.1200 ;
        RECT 1341.0200 2075.6400 1342.6200 2076.1200 ;
        RECT 1251.0200 2108.2800 1252.6200 2108.7600 ;
        RECT 1251.0200 2113.7200 1252.6200 2114.2000 ;
        RECT 1251.0200 2119.1600 1252.6200 2119.6400 ;
        RECT 1206.0200 2108.2800 1207.6200 2108.7600 ;
        RECT 1206.0200 2113.7200 1207.6200 2114.2000 ;
        RECT 1206.0200 2119.1600 1207.6200 2119.6400 ;
        RECT 1251.0200 2091.9600 1252.6200 2092.4400 ;
        RECT 1251.0200 2097.4000 1252.6200 2097.8800 ;
        RECT 1251.0200 2081.0800 1252.6200 2081.5600 ;
        RECT 1251.0200 2086.5200 1252.6200 2087.0000 ;
        RECT 1206.0200 2091.9600 1207.6200 2092.4400 ;
        RECT 1206.0200 2097.4000 1207.6200 2097.8800 ;
        RECT 1206.0200 2081.0800 1207.6200 2081.5600 ;
        RECT 1206.0200 2086.5200 1207.6200 2087.0000 ;
        RECT 1206.0200 2102.8400 1207.6200 2103.3200 ;
        RECT 1251.0200 2102.8400 1252.6200 2103.3200 ;
        RECT 1156.4600 2119.1600 1159.4600 2119.6400 ;
        RECT 1156.4600 2113.7200 1159.4600 2114.2000 ;
        RECT 1156.4600 2108.2800 1159.4600 2108.7600 ;
        RECT 1156.4600 2097.4000 1159.4600 2097.8800 ;
        RECT 1156.4600 2091.9600 1159.4600 2092.4400 ;
        RECT 1156.4600 2086.5200 1159.4600 2087.0000 ;
        RECT 1156.4600 2081.0800 1159.4600 2081.5600 ;
        RECT 1156.4600 2102.8400 1159.4600 2103.3200 ;
        RECT 1251.0200 2064.7600 1252.6200 2065.2400 ;
        RECT 1251.0200 2070.2000 1252.6200 2070.6800 ;
        RECT 1251.0200 2048.4400 1252.6200 2048.9200 ;
        RECT 1251.0200 2053.8800 1252.6200 2054.3600 ;
        RECT 1251.0200 2059.3200 1252.6200 2059.8000 ;
        RECT 1206.0200 2064.7600 1207.6200 2065.2400 ;
        RECT 1206.0200 2070.2000 1207.6200 2070.6800 ;
        RECT 1206.0200 2048.4400 1207.6200 2048.9200 ;
        RECT 1206.0200 2053.8800 1207.6200 2054.3600 ;
        RECT 1206.0200 2059.3200 1207.6200 2059.8000 ;
        RECT 1251.0200 2037.5600 1252.6200 2038.0400 ;
        RECT 1251.0200 2043.0000 1252.6200 2043.4800 ;
        RECT 1251.0200 2021.2400 1252.6200 2021.7200 ;
        RECT 1251.0200 2026.6800 1252.6200 2027.1600 ;
        RECT 1251.0200 2032.1200 1252.6200 2032.6000 ;
        RECT 1206.0200 2037.5600 1207.6200 2038.0400 ;
        RECT 1206.0200 2043.0000 1207.6200 2043.4800 ;
        RECT 1206.0200 2021.2400 1207.6200 2021.7200 ;
        RECT 1206.0200 2026.6800 1207.6200 2027.1600 ;
        RECT 1206.0200 2032.1200 1207.6200 2032.6000 ;
        RECT 1156.4600 2064.7600 1159.4600 2065.2400 ;
        RECT 1156.4600 2070.2000 1159.4600 2070.6800 ;
        RECT 1156.4600 2053.8800 1159.4600 2054.3600 ;
        RECT 1156.4600 2048.4400 1159.4600 2048.9200 ;
        RECT 1156.4600 2059.3200 1159.4600 2059.8000 ;
        RECT 1156.4600 2037.5600 1159.4600 2038.0400 ;
        RECT 1156.4600 2043.0000 1159.4600 2043.4800 ;
        RECT 1156.4600 2026.6800 1159.4600 2027.1600 ;
        RECT 1156.4600 2021.2400 1159.4600 2021.7200 ;
        RECT 1156.4600 2032.1200 1159.4600 2032.6000 ;
        RECT 1156.4600 2075.6400 1159.4600 2076.1200 ;
        RECT 1206.0200 2075.6400 1207.6200 2076.1200 ;
        RECT 1251.0200 2075.6400 1252.6200 2076.1200 ;
        RECT 1352.5600 2010.3600 1355.5600 2010.8400 ;
        RECT 1352.5600 2015.8000 1355.5600 2016.2800 ;
        RECT 1341.0200 2010.3600 1342.6200 2010.8400 ;
        RECT 1341.0200 2015.8000 1342.6200 2016.2800 ;
        RECT 1352.5600 1994.0400 1355.5600 1994.5200 ;
        RECT 1352.5600 1999.4800 1355.5600 1999.9600 ;
        RECT 1352.5600 2004.9200 1355.5600 2005.4000 ;
        RECT 1341.0200 1994.0400 1342.6200 1994.5200 ;
        RECT 1341.0200 1999.4800 1342.6200 1999.9600 ;
        RECT 1341.0200 2004.9200 1342.6200 2005.4000 ;
        RECT 1352.5600 1983.1600 1355.5600 1983.6400 ;
        RECT 1352.5600 1988.6000 1355.5600 1989.0800 ;
        RECT 1341.0200 1983.1600 1342.6200 1983.6400 ;
        RECT 1341.0200 1988.6000 1342.6200 1989.0800 ;
        RECT 1352.5600 1966.8400 1355.5600 1967.3200 ;
        RECT 1352.5600 1972.2800 1355.5600 1972.7600 ;
        RECT 1352.5600 1977.7200 1355.5600 1978.2000 ;
        RECT 1341.0200 1966.8400 1342.6200 1967.3200 ;
        RECT 1341.0200 1972.2800 1342.6200 1972.7600 ;
        RECT 1341.0200 1977.7200 1342.6200 1978.2000 ;
        RECT 1296.0200 2010.3600 1297.6200 2010.8400 ;
        RECT 1296.0200 2015.8000 1297.6200 2016.2800 ;
        RECT 1296.0200 1994.0400 1297.6200 1994.5200 ;
        RECT 1296.0200 1999.4800 1297.6200 1999.9600 ;
        RECT 1296.0200 2004.9200 1297.6200 2005.4000 ;
        RECT 1296.0200 1983.1600 1297.6200 1983.6400 ;
        RECT 1296.0200 1988.6000 1297.6200 1989.0800 ;
        RECT 1296.0200 1966.8400 1297.6200 1967.3200 ;
        RECT 1296.0200 1972.2800 1297.6200 1972.7600 ;
        RECT 1296.0200 1977.7200 1297.6200 1978.2000 ;
        RECT 1352.5600 1955.9600 1355.5600 1956.4400 ;
        RECT 1352.5600 1961.4000 1355.5600 1961.8800 ;
        RECT 1341.0200 1955.9600 1342.6200 1956.4400 ;
        RECT 1341.0200 1961.4000 1342.6200 1961.8800 ;
        RECT 1352.5600 1939.6400 1355.5600 1940.1200 ;
        RECT 1352.5600 1945.0800 1355.5600 1945.5600 ;
        RECT 1352.5600 1950.5200 1355.5600 1951.0000 ;
        RECT 1341.0200 1939.6400 1342.6200 1940.1200 ;
        RECT 1341.0200 1945.0800 1342.6200 1945.5600 ;
        RECT 1341.0200 1950.5200 1342.6200 1951.0000 ;
        RECT 1352.5600 1928.7600 1355.5600 1929.2400 ;
        RECT 1352.5600 1934.2000 1355.5600 1934.6800 ;
        RECT 1341.0200 1928.7600 1342.6200 1929.2400 ;
        RECT 1341.0200 1934.2000 1342.6200 1934.6800 ;
        RECT 1352.5600 1923.3200 1355.5600 1923.8000 ;
        RECT 1341.0200 1923.3200 1342.6200 1923.8000 ;
        RECT 1296.0200 1955.9600 1297.6200 1956.4400 ;
        RECT 1296.0200 1961.4000 1297.6200 1961.8800 ;
        RECT 1296.0200 1939.6400 1297.6200 1940.1200 ;
        RECT 1296.0200 1945.0800 1297.6200 1945.5600 ;
        RECT 1296.0200 1950.5200 1297.6200 1951.0000 ;
        RECT 1296.0200 1928.7600 1297.6200 1929.2400 ;
        RECT 1296.0200 1934.2000 1297.6200 1934.6800 ;
        RECT 1296.0200 1923.3200 1297.6200 1923.8000 ;
        RECT 1251.0200 2010.3600 1252.6200 2010.8400 ;
        RECT 1251.0200 2015.8000 1252.6200 2016.2800 ;
        RECT 1251.0200 1994.0400 1252.6200 1994.5200 ;
        RECT 1251.0200 1999.4800 1252.6200 1999.9600 ;
        RECT 1251.0200 2004.9200 1252.6200 2005.4000 ;
        RECT 1206.0200 2010.3600 1207.6200 2010.8400 ;
        RECT 1206.0200 2015.8000 1207.6200 2016.2800 ;
        RECT 1206.0200 1994.0400 1207.6200 1994.5200 ;
        RECT 1206.0200 1999.4800 1207.6200 1999.9600 ;
        RECT 1206.0200 2004.9200 1207.6200 2005.4000 ;
        RECT 1251.0200 1983.1600 1252.6200 1983.6400 ;
        RECT 1251.0200 1988.6000 1252.6200 1989.0800 ;
        RECT 1251.0200 1966.8400 1252.6200 1967.3200 ;
        RECT 1251.0200 1972.2800 1252.6200 1972.7600 ;
        RECT 1251.0200 1977.7200 1252.6200 1978.2000 ;
        RECT 1206.0200 1983.1600 1207.6200 1983.6400 ;
        RECT 1206.0200 1988.6000 1207.6200 1989.0800 ;
        RECT 1206.0200 1966.8400 1207.6200 1967.3200 ;
        RECT 1206.0200 1972.2800 1207.6200 1972.7600 ;
        RECT 1206.0200 1977.7200 1207.6200 1978.2000 ;
        RECT 1156.4600 2010.3600 1159.4600 2010.8400 ;
        RECT 1156.4600 2015.8000 1159.4600 2016.2800 ;
        RECT 1156.4600 1999.4800 1159.4600 1999.9600 ;
        RECT 1156.4600 1994.0400 1159.4600 1994.5200 ;
        RECT 1156.4600 2004.9200 1159.4600 2005.4000 ;
        RECT 1156.4600 1983.1600 1159.4600 1983.6400 ;
        RECT 1156.4600 1988.6000 1159.4600 1989.0800 ;
        RECT 1156.4600 1972.2800 1159.4600 1972.7600 ;
        RECT 1156.4600 1966.8400 1159.4600 1967.3200 ;
        RECT 1156.4600 1977.7200 1159.4600 1978.2000 ;
        RECT 1251.0200 1955.9600 1252.6200 1956.4400 ;
        RECT 1251.0200 1961.4000 1252.6200 1961.8800 ;
        RECT 1251.0200 1939.6400 1252.6200 1940.1200 ;
        RECT 1251.0200 1945.0800 1252.6200 1945.5600 ;
        RECT 1251.0200 1950.5200 1252.6200 1951.0000 ;
        RECT 1206.0200 1955.9600 1207.6200 1956.4400 ;
        RECT 1206.0200 1961.4000 1207.6200 1961.8800 ;
        RECT 1206.0200 1939.6400 1207.6200 1940.1200 ;
        RECT 1206.0200 1945.0800 1207.6200 1945.5600 ;
        RECT 1206.0200 1950.5200 1207.6200 1951.0000 ;
        RECT 1251.0200 1934.2000 1252.6200 1934.6800 ;
        RECT 1251.0200 1928.7600 1252.6200 1929.2400 ;
        RECT 1251.0200 1923.3200 1252.6200 1923.8000 ;
        RECT 1206.0200 1934.2000 1207.6200 1934.6800 ;
        RECT 1206.0200 1928.7600 1207.6200 1929.2400 ;
        RECT 1206.0200 1923.3200 1207.6200 1923.8000 ;
        RECT 1156.4600 1955.9600 1159.4600 1956.4400 ;
        RECT 1156.4600 1961.4000 1159.4600 1961.8800 ;
        RECT 1156.4600 1945.0800 1159.4600 1945.5600 ;
        RECT 1156.4600 1939.6400 1159.4600 1940.1200 ;
        RECT 1156.4600 1950.5200 1159.4600 1951.0000 ;
        RECT 1156.4600 1928.7600 1159.4600 1929.2400 ;
        RECT 1156.4600 1934.2000 1159.4600 1934.6800 ;
        RECT 1156.4600 1923.3200 1159.4600 1923.8000 ;
        RECT 1156.4600 2121.5100 1355.5600 2124.5100 ;
        RECT 1156.4600 1916.4100 1355.5600 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 1686.7700 1342.6200 1894.8700 ;
        RECT 1296.0200 1686.7700 1297.6200 1894.8700 ;
        RECT 1251.0200 1686.7700 1252.6200 1894.8700 ;
        RECT 1206.0200 1686.7700 1207.6200 1894.8700 ;
        RECT 1352.5600 1686.7700 1355.5600 1894.8700 ;
        RECT 1156.4600 1686.7700 1159.4600 1894.8700 ;
      LAYER met3 ;
        RECT 1352.5600 1889.5200 1355.5600 1890.0000 ;
        RECT 1341.0200 1889.5200 1342.6200 1890.0000 ;
        RECT 1352.5600 1878.6400 1355.5600 1879.1200 ;
        RECT 1352.5600 1884.0800 1355.5600 1884.5600 ;
        RECT 1341.0200 1878.6400 1342.6200 1879.1200 ;
        RECT 1341.0200 1884.0800 1342.6200 1884.5600 ;
        RECT 1352.5600 1862.3200 1355.5600 1862.8000 ;
        RECT 1352.5600 1867.7600 1355.5600 1868.2400 ;
        RECT 1341.0200 1862.3200 1342.6200 1862.8000 ;
        RECT 1341.0200 1867.7600 1342.6200 1868.2400 ;
        RECT 1352.5600 1851.4400 1355.5600 1851.9200 ;
        RECT 1352.5600 1856.8800 1355.5600 1857.3600 ;
        RECT 1341.0200 1851.4400 1342.6200 1851.9200 ;
        RECT 1341.0200 1856.8800 1342.6200 1857.3600 ;
        RECT 1352.5600 1873.2000 1355.5600 1873.6800 ;
        RECT 1341.0200 1873.2000 1342.6200 1873.6800 ;
        RECT 1296.0200 1878.6400 1297.6200 1879.1200 ;
        RECT 1296.0200 1884.0800 1297.6200 1884.5600 ;
        RECT 1296.0200 1889.5200 1297.6200 1890.0000 ;
        RECT 1296.0200 1862.3200 1297.6200 1862.8000 ;
        RECT 1296.0200 1867.7600 1297.6200 1868.2400 ;
        RECT 1296.0200 1856.8800 1297.6200 1857.3600 ;
        RECT 1296.0200 1851.4400 1297.6200 1851.9200 ;
        RECT 1296.0200 1873.2000 1297.6200 1873.6800 ;
        RECT 1352.5600 1835.1200 1355.5600 1835.6000 ;
        RECT 1352.5600 1840.5600 1355.5600 1841.0400 ;
        RECT 1341.0200 1835.1200 1342.6200 1835.6000 ;
        RECT 1341.0200 1840.5600 1342.6200 1841.0400 ;
        RECT 1352.5600 1818.8000 1355.5600 1819.2800 ;
        RECT 1352.5600 1824.2400 1355.5600 1824.7200 ;
        RECT 1352.5600 1829.6800 1355.5600 1830.1600 ;
        RECT 1341.0200 1818.8000 1342.6200 1819.2800 ;
        RECT 1341.0200 1824.2400 1342.6200 1824.7200 ;
        RECT 1341.0200 1829.6800 1342.6200 1830.1600 ;
        RECT 1352.5600 1807.9200 1355.5600 1808.4000 ;
        RECT 1352.5600 1813.3600 1355.5600 1813.8400 ;
        RECT 1341.0200 1807.9200 1342.6200 1808.4000 ;
        RECT 1341.0200 1813.3600 1342.6200 1813.8400 ;
        RECT 1352.5600 1791.6000 1355.5600 1792.0800 ;
        RECT 1352.5600 1797.0400 1355.5600 1797.5200 ;
        RECT 1352.5600 1802.4800 1355.5600 1802.9600 ;
        RECT 1341.0200 1791.6000 1342.6200 1792.0800 ;
        RECT 1341.0200 1797.0400 1342.6200 1797.5200 ;
        RECT 1341.0200 1802.4800 1342.6200 1802.9600 ;
        RECT 1296.0200 1835.1200 1297.6200 1835.6000 ;
        RECT 1296.0200 1840.5600 1297.6200 1841.0400 ;
        RECT 1296.0200 1818.8000 1297.6200 1819.2800 ;
        RECT 1296.0200 1824.2400 1297.6200 1824.7200 ;
        RECT 1296.0200 1829.6800 1297.6200 1830.1600 ;
        RECT 1296.0200 1807.9200 1297.6200 1808.4000 ;
        RECT 1296.0200 1813.3600 1297.6200 1813.8400 ;
        RECT 1296.0200 1791.6000 1297.6200 1792.0800 ;
        RECT 1296.0200 1797.0400 1297.6200 1797.5200 ;
        RECT 1296.0200 1802.4800 1297.6200 1802.9600 ;
        RECT 1352.5600 1846.0000 1355.5600 1846.4800 ;
        RECT 1296.0200 1846.0000 1297.6200 1846.4800 ;
        RECT 1341.0200 1846.0000 1342.6200 1846.4800 ;
        RECT 1251.0200 1878.6400 1252.6200 1879.1200 ;
        RECT 1251.0200 1884.0800 1252.6200 1884.5600 ;
        RECT 1251.0200 1889.5200 1252.6200 1890.0000 ;
        RECT 1206.0200 1878.6400 1207.6200 1879.1200 ;
        RECT 1206.0200 1884.0800 1207.6200 1884.5600 ;
        RECT 1206.0200 1889.5200 1207.6200 1890.0000 ;
        RECT 1251.0200 1862.3200 1252.6200 1862.8000 ;
        RECT 1251.0200 1867.7600 1252.6200 1868.2400 ;
        RECT 1251.0200 1851.4400 1252.6200 1851.9200 ;
        RECT 1251.0200 1856.8800 1252.6200 1857.3600 ;
        RECT 1206.0200 1862.3200 1207.6200 1862.8000 ;
        RECT 1206.0200 1867.7600 1207.6200 1868.2400 ;
        RECT 1206.0200 1851.4400 1207.6200 1851.9200 ;
        RECT 1206.0200 1856.8800 1207.6200 1857.3600 ;
        RECT 1206.0200 1873.2000 1207.6200 1873.6800 ;
        RECT 1251.0200 1873.2000 1252.6200 1873.6800 ;
        RECT 1156.4600 1889.5200 1159.4600 1890.0000 ;
        RECT 1156.4600 1884.0800 1159.4600 1884.5600 ;
        RECT 1156.4600 1878.6400 1159.4600 1879.1200 ;
        RECT 1156.4600 1867.7600 1159.4600 1868.2400 ;
        RECT 1156.4600 1862.3200 1159.4600 1862.8000 ;
        RECT 1156.4600 1856.8800 1159.4600 1857.3600 ;
        RECT 1156.4600 1851.4400 1159.4600 1851.9200 ;
        RECT 1156.4600 1873.2000 1159.4600 1873.6800 ;
        RECT 1251.0200 1835.1200 1252.6200 1835.6000 ;
        RECT 1251.0200 1840.5600 1252.6200 1841.0400 ;
        RECT 1251.0200 1818.8000 1252.6200 1819.2800 ;
        RECT 1251.0200 1824.2400 1252.6200 1824.7200 ;
        RECT 1251.0200 1829.6800 1252.6200 1830.1600 ;
        RECT 1206.0200 1835.1200 1207.6200 1835.6000 ;
        RECT 1206.0200 1840.5600 1207.6200 1841.0400 ;
        RECT 1206.0200 1818.8000 1207.6200 1819.2800 ;
        RECT 1206.0200 1824.2400 1207.6200 1824.7200 ;
        RECT 1206.0200 1829.6800 1207.6200 1830.1600 ;
        RECT 1251.0200 1807.9200 1252.6200 1808.4000 ;
        RECT 1251.0200 1813.3600 1252.6200 1813.8400 ;
        RECT 1251.0200 1791.6000 1252.6200 1792.0800 ;
        RECT 1251.0200 1797.0400 1252.6200 1797.5200 ;
        RECT 1251.0200 1802.4800 1252.6200 1802.9600 ;
        RECT 1206.0200 1807.9200 1207.6200 1808.4000 ;
        RECT 1206.0200 1813.3600 1207.6200 1813.8400 ;
        RECT 1206.0200 1791.6000 1207.6200 1792.0800 ;
        RECT 1206.0200 1797.0400 1207.6200 1797.5200 ;
        RECT 1206.0200 1802.4800 1207.6200 1802.9600 ;
        RECT 1156.4600 1835.1200 1159.4600 1835.6000 ;
        RECT 1156.4600 1840.5600 1159.4600 1841.0400 ;
        RECT 1156.4600 1824.2400 1159.4600 1824.7200 ;
        RECT 1156.4600 1818.8000 1159.4600 1819.2800 ;
        RECT 1156.4600 1829.6800 1159.4600 1830.1600 ;
        RECT 1156.4600 1807.9200 1159.4600 1808.4000 ;
        RECT 1156.4600 1813.3600 1159.4600 1813.8400 ;
        RECT 1156.4600 1797.0400 1159.4600 1797.5200 ;
        RECT 1156.4600 1791.6000 1159.4600 1792.0800 ;
        RECT 1156.4600 1802.4800 1159.4600 1802.9600 ;
        RECT 1156.4600 1846.0000 1159.4600 1846.4800 ;
        RECT 1206.0200 1846.0000 1207.6200 1846.4800 ;
        RECT 1251.0200 1846.0000 1252.6200 1846.4800 ;
        RECT 1352.5600 1780.7200 1355.5600 1781.2000 ;
        RECT 1352.5600 1786.1600 1355.5600 1786.6400 ;
        RECT 1341.0200 1780.7200 1342.6200 1781.2000 ;
        RECT 1341.0200 1786.1600 1342.6200 1786.6400 ;
        RECT 1352.5600 1764.4000 1355.5600 1764.8800 ;
        RECT 1352.5600 1769.8400 1355.5600 1770.3200 ;
        RECT 1352.5600 1775.2800 1355.5600 1775.7600 ;
        RECT 1341.0200 1764.4000 1342.6200 1764.8800 ;
        RECT 1341.0200 1769.8400 1342.6200 1770.3200 ;
        RECT 1341.0200 1775.2800 1342.6200 1775.7600 ;
        RECT 1352.5600 1753.5200 1355.5600 1754.0000 ;
        RECT 1352.5600 1758.9600 1355.5600 1759.4400 ;
        RECT 1341.0200 1753.5200 1342.6200 1754.0000 ;
        RECT 1341.0200 1758.9600 1342.6200 1759.4400 ;
        RECT 1352.5600 1737.2000 1355.5600 1737.6800 ;
        RECT 1352.5600 1742.6400 1355.5600 1743.1200 ;
        RECT 1352.5600 1748.0800 1355.5600 1748.5600 ;
        RECT 1341.0200 1737.2000 1342.6200 1737.6800 ;
        RECT 1341.0200 1742.6400 1342.6200 1743.1200 ;
        RECT 1341.0200 1748.0800 1342.6200 1748.5600 ;
        RECT 1296.0200 1780.7200 1297.6200 1781.2000 ;
        RECT 1296.0200 1786.1600 1297.6200 1786.6400 ;
        RECT 1296.0200 1764.4000 1297.6200 1764.8800 ;
        RECT 1296.0200 1769.8400 1297.6200 1770.3200 ;
        RECT 1296.0200 1775.2800 1297.6200 1775.7600 ;
        RECT 1296.0200 1753.5200 1297.6200 1754.0000 ;
        RECT 1296.0200 1758.9600 1297.6200 1759.4400 ;
        RECT 1296.0200 1737.2000 1297.6200 1737.6800 ;
        RECT 1296.0200 1742.6400 1297.6200 1743.1200 ;
        RECT 1296.0200 1748.0800 1297.6200 1748.5600 ;
        RECT 1352.5600 1726.3200 1355.5600 1726.8000 ;
        RECT 1352.5600 1731.7600 1355.5600 1732.2400 ;
        RECT 1341.0200 1726.3200 1342.6200 1726.8000 ;
        RECT 1341.0200 1731.7600 1342.6200 1732.2400 ;
        RECT 1352.5600 1710.0000 1355.5600 1710.4800 ;
        RECT 1352.5600 1715.4400 1355.5600 1715.9200 ;
        RECT 1352.5600 1720.8800 1355.5600 1721.3600 ;
        RECT 1341.0200 1710.0000 1342.6200 1710.4800 ;
        RECT 1341.0200 1715.4400 1342.6200 1715.9200 ;
        RECT 1341.0200 1720.8800 1342.6200 1721.3600 ;
        RECT 1352.5600 1699.1200 1355.5600 1699.6000 ;
        RECT 1352.5600 1704.5600 1355.5600 1705.0400 ;
        RECT 1341.0200 1699.1200 1342.6200 1699.6000 ;
        RECT 1341.0200 1704.5600 1342.6200 1705.0400 ;
        RECT 1352.5600 1693.6800 1355.5600 1694.1600 ;
        RECT 1341.0200 1693.6800 1342.6200 1694.1600 ;
        RECT 1296.0200 1726.3200 1297.6200 1726.8000 ;
        RECT 1296.0200 1731.7600 1297.6200 1732.2400 ;
        RECT 1296.0200 1710.0000 1297.6200 1710.4800 ;
        RECT 1296.0200 1715.4400 1297.6200 1715.9200 ;
        RECT 1296.0200 1720.8800 1297.6200 1721.3600 ;
        RECT 1296.0200 1699.1200 1297.6200 1699.6000 ;
        RECT 1296.0200 1704.5600 1297.6200 1705.0400 ;
        RECT 1296.0200 1693.6800 1297.6200 1694.1600 ;
        RECT 1251.0200 1780.7200 1252.6200 1781.2000 ;
        RECT 1251.0200 1786.1600 1252.6200 1786.6400 ;
        RECT 1251.0200 1764.4000 1252.6200 1764.8800 ;
        RECT 1251.0200 1769.8400 1252.6200 1770.3200 ;
        RECT 1251.0200 1775.2800 1252.6200 1775.7600 ;
        RECT 1206.0200 1780.7200 1207.6200 1781.2000 ;
        RECT 1206.0200 1786.1600 1207.6200 1786.6400 ;
        RECT 1206.0200 1764.4000 1207.6200 1764.8800 ;
        RECT 1206.0200 1769.8400 1207.6200 1770.3200 ;
        RECT 1206.0200 1775.2800 1207.6200 1775.7600 ;
        RECT 1251.0200 1753.5200 1252.6200 1754.0000 ;
        RECT 1251.0200 1758.9600 1252.6200 1759.4400 ;
        RECT 1251.0200 1737.2000 1252.6200 1737.6800 ;
        RECT 1251.0200 1742.6400 1252.6200 1743.1200 ;
        RECT 1251.0200 1748.0800 1252.6200 1748.5600 ;
        RECT 1206.0200 1753.5200 1207.6200 1754.0000 ;
        RECT 1206.0200 1758.9600 1207.6200 1759.4400 ;
        RECT 1206.0200 1737.2000 1207.6200 1737.6800 ;
        RECT 1206.0200 1742.6400 1207.6200 1743.1200 ;
        RECT 1206.0200 1748.0800 1207.6200 1748.5600 ;
        RECT 1156.4600 1780.7200 1159.4600 1781.2000 ;
        RECT 1156.4600 1786.1600 1159.4600 1786.6400 ;
        RECT 1156.4600 1769.8400 1159.4600 1770.3200 ;
        RECT 1156.4600 1764.4000 1159.4600 1764.8800 ;
        RECT 1156.4600 1775.2800 1159.4600 1775.7600 ;
        RECT 1156.4600 1753.5200 1159.4600 1754.0000 ;
        RECT 1156.4600 1758.9600 1159.4600 1759.4400 ;
        RECT 1156.4600 1742.6400 1159.4600 1743.1200 ;
        RECT 1156.4600 1737.2000 1159.4600 1737.6800 ;
        RECT 1156.4600 1748.0800 1159.4600 1748.5600 ;
        RECT 1251.0200 1726.3200 1252.6200 1726.8000 ;
        RECT 1251.0200 1731.7600 1252.6200 1732.2400 ;
        RECT 1251.0200 1710.0000 1252.6200 1710.4800 ;
        RECT 1251.0200 1715.4400 1252.6200 1715.9200 ;
        RECT 1251.0200 1720.8800 1252.6200 1721.3600 ;
        RECT 1206.0200 1726.3200 1207.6200 1726.8000 ;
        RECT 1206.0200 1731.7600 1207.6200 1732.2400 ;
        RECT 1206.0200 1710.0000 1207.6200 1710.4800 ;
        RECT 1206.0200 1715.4400 1207.6200 1715.9200 ;
        RECT 1206.0200 1720.8800 1207.6200 1721.3600 ;
        RECT 1251.0200 1704.5600 1252.6200 1705.0400 ;
        RECT 1251.0200 1699.1200 1252.6200 1699.6000 ;
        RECT 1251.0200 1693.6800 1252.6200 1694.1600 ;
        RECT 1206.0200 1704.5600 1207.6200 1705.0400 ;
        RECT 1206.0200 1699.1200 1207.6200 1699.6000 ;
        RECT 1206.0200 1693.6800 1207.6200 1694.1600 ;
        RECT 1156.4600 1726.3200 1159.4600 1726.8000 ;
        RECT 1156.4600 1731.7600 1159.4600 1732.2400 ;
        RECT 1156.4600 1715.4400 1159.4600 1715.9200 ;
        RECT 1156.4600 1710.0000 1159.4600 1710.4800 ;
        RECT 1156.4600 1720.8800 1159.4600 1721.3600 ;
        RECT 1156.4600 1699.1200 1159.4600 1699.6000 ;
        RECT 1156.4600 1704.5600 1159.4600 1705.0400 ;
        RECT 1156.4600 1693.6800 1159.4600 1694.1600 ;
        RECT 1156.4600 1891.8700 1355.5600 1894.8700 ;
        RECT 1156.4600 1686.7700 1355.5600 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 1457.1300 1342.6200 1665.2300 ;
        RECT 1296.0200 1457.1300 1297.6200 1665.2300 ;
        RECT 1251.0200 1457.1300 1252.6200 1665.2300 ;
        RECT 1206.0200 1457.1300 1207.6200 1665.2300 ;
        RECT 1352.5600 1457.1300 1355.5600 1665.2300 ;
        RECT 1156.4600 1457.1300 1159.4600 1665.2300 ;
      LAYER met3 ;
        RECT 1352.5600 1659.8800 1355.5600 1660.3600 ;
        RECT 1341.0200 1659.8800 1342.6200 1660.3600 ;
        RECT 1352.5600 1649.0000 1355.5600 1649.4800 ;
        RECT 1352.5600 1654.4400 1355.5600 1654.9200 ;
        RECT 1341.0200 1649.0000 1342.6200 1649.4800 ;
        RECT 1341.0200 1654.4400 1342.6200 1654.9200 ;
        RECT 1352.5600 1632.6800 1355.5600 1633.1600 ;
        RECT 1352.5600 1638.1200 1355.5600 1638.6000 ;
        RECT 1341.0200 1632.6800 1342.6200 1633.1600 ;
        RECT 1341.0200 1638.1200 1342.6200 1638.6000 ;
        RECT 1352.5600 1621.8000 1355.5600 1622.2800 ;
        RECT 1352.5600 1627.2400 1355.5600 1627.7200 ;
        RECT 1341.0200 1621.8000 1342.6200 1622.2800 ;
        RECT 1341.0200 1627.2400 1342.6200 1627.7200 ;
        RECT 1352.5600 1643.5600 1355.5600 1644.0400 ;
        RECT 1341.0200 1643.5600 1342.6200 1644.0400 ;
        RECT 1296.0200 1649.0000 1297.6200 1649.4800 ;
        RECT 1296.0200 1654.4400 1297.6200 1654.9200 ;
        RECT 1296.0200 1659.8800 1297.6200 1660.3600 ;
        RECT 1296.0200 1632.6800 1297.6200 1633.1600 ;
        RECT 1296.0200 1638.1200 1297.6200 1638.6000 ;
        RECT 1296.0200 1627.2400 1297.6200 1627.7200 ;
        RECT 1296.0200 1621.8000 1297.6200 1622.2800 ;
        RECT 1296.0200 1643.5600 1297.6200 1644.0400 ;
        RECT 1352.5600 1605.4800 1355.5600 1605.9600 ;
        RECT 1352.5600 1610.9200 1355.5600 1611.4000 ;
        RECT 1341.0200 1605.4800 1342.6200 1605.9600 ;
        RECT 1341.0200 1610.9200 1342.6200 1611.4000 ;
        RECT 1352.5600 1589.1600 1355.5600 1589.6400 ;
        RECT 1352.5600 1594.6000 1355.5600 1595.0800 ;
        RECT 1352.5600 1600.0400 1355.5600 1600.5200 ;
        RECT 1341.0200 1589.1600 1342.6200 1589.6400 ;
        RECT 1341.0200 1594.6000 1342.6200 1595.0800 ;
        RECT 1341.0200 1600.0400 1342.6200 1600.5200 ;
        RECT 1352.5600 1578.2800 1355.5600 1578.7600 ;
        RECT 1352.5600 1583.7200 1355.5600 1584.2000 ;
        RECT 1341.0200 1578.2800 1342.6200 1578.7600 ;
        RECT 1341.0200 1583.7200 1342.6200 1584.2000 ;
        RECT 1352.5600 1561.9600 1355.5600 1562.4400 ;
        RECT 1352.5600 1567.4000 1355.5600 1567.8800 ;
        RECT 1352.5600 1572.8400 1355.5600 1573.3200 ;
        RECT 1341.0200 1561.9600 1342.6200 1562.4400 ;
        RECT 1341.0200 1567.4000 1342.6200 1567.8800 ;
        RECT 1341.0200 1572.8400 1342.6200 1573.3200 ;
        RECT 1296.0200 1605.4800 1297.6200 1605.9600 ;
        RECT 1296.0200 1610.9200 1297.6200 1611.4000 ;
        RECT 1296.0200 1589.1600 1297.6200 1589.6400 ;
        RECT 1296.0200 1594.6000 1297.6200 1595.0800 ;
        RECT 1296.0200 1600.0400 1297.6200 1600.5200 ;
        RECT 1296.0200 1578.2800 1297.6200 1578.7600 ;
        RECT 1296.0200 1583.7200 1297.6200 1584.2000 ;
        RECT 1296.0200 1561.9600 1297.6200 1562.4400 ;
        RECT 1296.0200 1567.4000 1297.6200 1567.8800 ;
        RECT 1296.0200 1572.8400 1297.6200 1573.3200 ;
        RECT 1352.5600 1616.3600 1355.5600 1616.8400 ;
        RECT 1296.0200 1616.3600 1297.6200 1616.8400 ;
        RECT 1341.0200 1616.3600 1342.6200 1616.8400 ;
        RECT 1251.0200 1649.0000 1252.6200 1649.4800 ;
        RECT 1251.0200 1654.4400 1252.6200 1654.9200 ;
        RECT 1251.0200 1659.8800 1252.6200 1660.3600 ;
        RECT 1206.0200 1649.0000 1207.6200 1649.4800 ;
        RECT 1206.0200 1654.4400 1207.6200 1654.9200 ;
        RECT 1206.0200 1659.8800 1207.6200 1660.3600 ;
        RECT 1251.0200 1632.6800 1252.6200 1633.1600 ;
        RECT 1251.0200 1638.1200 1252.6200 1638.6000 ;
        RECT 1251.0200 1621.8000 1252.6200 1622.2800 ;
        RECT 1251.0200 1627.2400 1252.6200 1627.7200 ;
        RECT 1206.0200 1632.6800 1207.6200 1633.1600 ;
        RECT 1206.0200 1638.1200 1207.6200 1638.6000 ;
        RECT 1206.0200 1621.8000 1207.6200 1622.2800 ;
        RECT 1206.0200 1627.2400 1207.6200 1627.7200 ;
        RECT 1206.0200 1643.5600 1207.6200 1644.0400 ;
        RECT 1251.0200 1643.5600 1252.6200 1644.0400 ;
        RECT 1156.4600 1659.8800 1159.4600 1660.3600 ;
        RECT 1156.4600 1654.4400 1159.4600 1654.9200 ;
        RECT 1156.4600 1649.0000 1159.4600 1649.4800 ;
        RECT 1156.4600 1638.1200 1159.4600 1638.6000 ;
        RECT 1156.4600 1632.6800 1159.4600 1633.1600 ;
        RECT 1156.4600 1627.2400 1159.4600 1627.7200 ;
        RECT 1156.4600 1621.8000 1159.4600 1622.2800 ;
        RECT 1156.4600 1643.5600 1159.4600 1644.0400 ;
        RECT 1251.0200 1605.4800 1252.6200 1605.9600 ;
        RECT 1251.0200 1610.9200 1252.6200 1611.4000 ;
        RECT 1251.0200 1589.1600 1252.6200 1589.6400 ;
        RECT 1251.0200 1594.6000 1252.6200 1595.0800 ;
        RECT 1251.0200 1600.0400 1252.6200 1600.5200 ;
        RECT 1206.0200 1605.4800 1207.6200 1605.9600 ;
        RECT 1206.0200 1610.9200 1207.6200 1611.4000 ;
        RECT 1206.0200 1589.1600 1207.6200 1589.6400 ;
        RECT 1206.0200 1594.6000 1207.6200 1595.0800 ;
        RECT 1206.0200 1600.0400 1207.6200 1600.5200 ;
        RECT 1251.0200 1578.2800 1252.6200 1578.7600 ;
        RECT 1251.0200 1583.7200 1252.6200 1584.2000 ;
        RECT 1251.0200 1561.9600 1252.6200 1562.4400 ;
        RECT 1251.0200 1567.4000 1252.6200 1567.8800 ;
        RECT 1251.0200 1572.8400 1252.6200 1573.3200 ;
        RECT 1206.0200 1578.2800 1207.6200 1578.7600 ;
        RECT 1206.0200 1583.7200 1207.6200 1584.2000 ;
        RECT 1206.0200 1561.9600 1207.6200 1562.4400 ;
        RECT 1206.0200 1567.4000 1207.6200 1567.8800 ;
        RECT 1206.0200 1572.8400 1207.6200 1573.3200 ;
        RECT 1156.4600 1605.4800 1159.4600 1605.9600 ;
        RECT 1156.4600 1610.9200 1159.4600 1611.4000 ;
        RECT 1156.4600 1594.6000 1159.4600 1595.0800 ;
        RECT 1156.4600 1589.1600 1159.4600 1589.6400 ;
        RECT 1156.4600 1600.0400 1159.4600 1600.5200 ;
        RECT 1156.4600 1578.2800 1159.4600 1578.7600 ;
        RECT 1156.4600 1583.7200 1159.4600 1584.2000 ;
        RECT 1156.4600 1567.4000 1159.4600 1567.8800 ;
        RECT 1156.4600 1561.9600 1159.4600 1562.4400 ;
        RECT 1156.4600 1572.8400 1159.4600 1573.3200 ;
        RECT 1156.4600 1616.3600 1159.4600 1616.8400 ;
        RECT 1206.0200 1616.3600 1207.6200 1616.8400 ;
        RECT 1251.0200 1616.3600 1252.6200 1616.8400 ;
        RECT 1352.5600 1551.0800 1355.5600 1551.5600 ;
        RECT 1352.5600 1556.5200 1355.5600 1557.0000 ;
        RECT 1341.0200 1551.0800 1342.6200 1551.5600 ;
        RECT 1341.0200 1556.5200 1342.6200 1557.0000 ;
        RECT 1352.5600 1534.7600 1355.5600 1535.2400 ;
        RECT 1352.5600 1540.2000 1355.5600 1540.6800 ;
        RECT 1352.5600 1545.6400 1355.5600 1546.1200 ;
        RECT 1341.0200 1534.7600 1342.6200 1535.2400 ;
        RECT 1341.0200 1540.2000 1342.6200 1540.6800 ;
        RECT 1341.0200 1545.6400 1342.6200 1546.1200 ;
        RECT 1352.5600 1523.8800 1355.5600 1524.3600 ;
        RECT 1352.5600 1529.3200 1355.5600 1529.8000 ;
        RECT 1341.0200 1523.8800 1342.6200 1524.3600 ;
        RECT 1341.0200 1529.3200 1342.6200 1529.8000 ;
        RECT 1352.5600 1507.5600 1355.5600 1508.0400 ;
        RECT 1352.5600 1513.0000 1355.5600 1513.4800 ;
        RECT 1352.5600 1518.4400 1355.5600 1518.9200 ;
        RECT 1341.0200 1507.5600 1342.6200 1508.0400 ;
        RECT 1341.0200 1513.0000 1342.6200 1513.4800 ;
        RECT 1341.0200 1518.4400 1342.6200 1518.9200 ;
        RECT 1296.0200 1551.0800 1297.6200 1551.5600 ;
        RECT 1296.0200 1556.5200 1297.6200 1557.0000 ;
        RECT 1296.0200 1534.7600 1297.6200 1535.2400 ;
        RECT 1296.0200 1540.2000 1297.6200 1540.6800 ;
        RECT 1296.0200 1545.6400 1297.6200 1546.1200 ;
        RECT 1296.0200 1523.8800 1297.6200 1524.3600 ;
        RECT 1296.0200 1529.3200 1297.6200 1529.8000 ;
        RECT 1296.0200 1507.5600 1297.6200 1508.0400 ;
        RECT 1296.0200 1513.0000 1297.6200 1513.4800 ;
        RECT 1296.0200 1518.4400 1297.6200 1518.9200 ;
        RECT 1352.5600 1496.6800 1355.5600 1497.1600 ;
        RECT 1352.5600 1502.1200 1355.5600 1502.6000 ;
        RECT 1341.0200 1496.6800 1342.6200 1497.1600 ;
        RECT 1341.0200 1502.1200 1342.6200 1502.6000 ;
        RECT 1352.5600 1480.3600 1355.5600 1480.8400 ;
        RECT 1352.5600 1485.8000 1355.5600 1486.2800 ;
        RECT 1352.5600 1491.2400 1355.5600 1491.7200 ;
        RECT 1341.0200 1480.3600 1342.6200 1480.8400 ;
        RECT 1341.0200 1485.8000 1342.6200 1486.2800 ;
        RECT 1341.0200 1491.2400 1342.6200 1491.7200 ;
        RECT 1352.5600 1469.4800 1355.5600 1469.9600 ;
        RECT 1352.5600 1474.9200 1355.5600 1475.4000 ;
        RECT 1341.0200 1469.4800 1342.6200 1469.9600 ;
        RECT 1341.0200 1474.9200 1342.6200 1475.4000 ;
        RECT 1352.5600 1464.0400 1355.5600 1464.5200 ;
        RECT 1341.0200 1464.0400 1342.6200 1464.5200 ;
        RECT 1296.0200 1496.6800 1297.6200 1497.1600 ;
        RECT 1296.0200 1502.1200 1297.6200 1502.6000 ;
        RECT 1296.0200 1480.3600 1297.6200 1480.8400 ;
        RECT 1296.0200 1485.8000 1297.6200 1486.2800 ;
        RECT 1296.0200 1491.2400 1297.6200 1491.7200 ;
        RECT 1296.0200 1469.4800 1297.6200 1469.9600 ;
        RECT 1296.0200 1474.9200 1297.6200 1475.4000 ;
        RECT 1296.0200 1464.0400 1297.6200 1464.5200 ;
        RECT 1251.0200 1551.0800 1252.6200 1551.5600 ;
        RECT 1251.0200 1556.5200 1252.6200 1557.0000 ;
        RECT 1251.0200 1534.7600 1252.6200 1535.2400 ;
        RECT 1251.0200 1540.2000 1252.6200 1540.6800 ;
        RECT 1251.0200 1545.6400 1252.6200 1546.1200 ;
        RECT 1206.0200 1551.0800 1207.6200 1551.5600 ;
        RECT 1206.0200 1556.5200 1207.6200 1557.0000 ;
        RECT 1206.0200 1534.7600 1207.6200 1535.2400 ;
        RECT 1206.0200 1540.2000 1207.6200 1540.6800 ;
        RECT 1206.0200 1545.6400 1207.6200 1546.1200 ;
        RECT 1251.0200 1523.8800 1252.6200 1524.3600 ;
        RECT 1251.0200 1529.3200 1252.6200 1529.8000 ;
        RECT 1251.0200 1507.5600 1252.6200 1508.0400 ;
        RECT 1251.0200 1513.0000 1252.6200 1513.4800 ;
        RECT 1251.0200 1518.4400 1252.6200 1518.9200 ;
        RECT 1206.0200 1523.8800 1207.6200 1524.3600 ;
        RECT 1206.0200 1529.3200 1207.6200 1529.8000 ;
        RECT 1206.0200 1507.5600 1207.6200 1508.0400 ;
        RECT 1206.0200 1513.0000 1207.6200 1513.4800 ;
        RECT 1206.0200 1518.4400 1207.6200 1518.9200 ;
        RECT 1156.4600 1551.0800 1159.4600 1551.5600 ;
        RECT 1156.4600 1556.5200 1159.4600 1557.0000 ;
        RECT 1156.4600 1540.2000 1159.4600 1540.6800 ;
        RECT 1156.4600 1534.7600 1159.4600 1535.2400 ;
        RECT 1156.4600 1545.6400 1159.4600 1546.1200 ;
        RECT 1156.4600 1523.8800 1159.4600 1524.3600 ;
        RECT 1156.4600 1529.3200 1159.4600 1529.8000 ;
        RECT 1156.4600 1513.0000 1159.4600 1513.4800 ;
        RECT 1156.4600 1507.5600 1159.4600 1508.0400 ;
        RECT 1156.4600 1518.4400 1159.4600 1518.9200 ;
        RECT 1251.0200 1496.6800 1252.6200 1497.1600 ;
        RECT 1251.0200 1502.1200 1252.6200 1502.6000 ;
        RECT 1251.0200 1480.3600 1252.6200 1480.8400 ;
        RECT 1251.0200 1485.8000 1252.6200 1486.2800 ;
        RECT 1251.0200 1491.2400 1252.6200 1491.7200 ;
        RECT 1206.0200 1496.6800 1207.6200 1497.1600 ;
        RECT 1206.0200 1502.1200 1207.6200 1502.6000 ;
        RECT 1206.0200 1480.3600 1207.6200 1480.8400 ;
        RECT 1206.0200 1485.8000 1207.6200 1486.2800 ;
        RECT 1206.0200 1491.2400 1207.6200 1491.7200 ;
        RECT 1251.0200 1474.9200 1252.6200 1475.4000 ;
        RECT 1251.0200 1469.4800 1252.6200 1469.9600 ;
        RECT 1251.0200 1464.0400 1252.6200 1464.5200 ;
        RECT 1206.0200 1474.9200 1207.6200 1475.4000 ;
        RECT 1206.0200 1469.4800 1207.6200 1469.9600 ;
        RECT 1206.0200 1464.0400 1207.6200 1464.5200 ;
        RECT 1156.4600 1496.6800 1159.4600 1497.1600 ;
        RECT 1156.4600 1502.1200 1159.4600 1502.6000 ;
        RECT 1156.4600 1485.8000 1159.4600 1486.2800 ;
        RECT 1156.4600 1480.3600 1159.4600 1480.8400 ;
        RECT 1156.4600 1491.2400 1159.4600 1491.7200 ;
        RECT 1156.4600 1469.4800 1159.4600 1469.9600 ;
        RECT 1156.4600 1474.9200 1159.4600 1475.4000 ;
        RECT 1156.4600 1464.0400 1159.4600 1464.5200 ;
        RECT 1156.4600 1662.2300 1355.5600 1665.2300 ;
        RECT 1156.4600 1457.1300 1355.5600 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 1227.4900 1342.6200 1435.5900 ;
        RECT 1296.0200 1227.4900 1297.6200 1435.5900 ;
        RECT 1251.0200 1227.4900 1252.6200 1435.5900 ;
        RECT 1206.0200 1227.4900 1207.6200 1435.5900 ;
        RECT 1352.5600 1227.4900 1355.5600 1435.5900 ;
        RECT 1156.4600 1227.4900 1159.4600 1435.5900 ;
      LAYER met3 ;
        RECT 1352.5600 1430.2400 1355.5600 1430.7200 ;
        RECT 1341.0200 1430.2400 1342.6200 1430.7200 ;
        RECT 1352.5600 1419.3600 1355.5600 1419.8400 ;
        RECT 1352.5600 1424.8000 1355.5600 1425.2800 ;
        RECT 1341.0200 1419.3600 1342.6200 1419.8400 ;
        RECT 1341.0200 1424.8000 1342.6200 1425.2800 ;
        RECT 1352.5600 1403.0400 1355.5600 1403.5200 ;
        RECT 1352.5600 1408.4800 1355.5600 1408.9600 ;
        RECT 1341.0200 1403.0400 1342.6200 1403.5200 ;
        RECT 1341.0200 1408.4800 1342.6200 1408.9600 ;
        RECT 1352.5600 1392.1600 1355.5600 1392.6400 ;
        RECT 1352.5600 1397.6000 1355.5600 1398.0800 ;
        RECT 1341.0200 1392.1600 1342.6200 1392.6400 ;
        RECT 1341.0200 1397.6000 1342.6200 1398.0800 ;
        RECT 1352.5600 1413.9200 1355.5600 1414.4000 ;
        RECT 1341.0200 1413.9200 1342.6200 1414.4000 ;
        RECT 1296.0200 1419.3600 1297.6200 1419.8400 ;
        RECT 1296.0200 1424.8000 1297.6200 1425.2800 ;
        RECT 1296.0200 1430.2400 1297.6200 1430.7200 ;
        RECT 1296.0200 1403.0400 1297.6200 1403.5200 ;
        RECT 1296.0200 1408.4800 1297.6200 1408.9600 ;
        RECT 1296.0200 1397.6000 1297.6200 1398.0800 ;
        RECT 1296.0200 1392.1600 1297.6200 1392.6400 ;
        RECT 1296.0200 1413.9200 1297.6200 1414.4000 ;
        RECT 1352.5600 1375.8400 1355.5600 1376.3200 ;
        RECT 1352.5600 1381.2800 1355.5600 1381.7600 ;
        RECT 1341.0200 1375.8400 1342.6200 1376.3200 ;
        RECT 1341.0200 1381.2800 1342.6200 1381.7600 ;
        RECT 1352.5600 1359.5200 1355.5600 1360.0000 ;
        RECT 1352.5600 1364.9600 1355.5600 1365.4400 ;
        RECT 1352.5600 1370.4000 1355.5600 1370.8800 ;
        RECT 1341.0200 1359.5200 1342.6200 1360.0000 ;
        RECT 1341.0200 1364.9600 1342.6200 1365.4400 ;
        RECT 1341.0200 1370.4000 1342.6200 1370.8800 ;
        RECT 1352.5600 1348.6400 1355.5600 1349.1200 ;
        RECT 1352.5600 1354.0800 1355.5600 1354.5600 ;
        RECT 1341.0200 1348.6400 1342.6200 1349.1200 ;
        RECT 1341.0200 1354.0800 1342.6200 1354.5600 ;
        RECT 1352.5600 1332.3200 1355.5600 1332.8000 ;
        RECT 1352.5600 1337.7600 1355.5600 1338.2400 ;
        RECT 1352.5600 1343.2000 1355.5600 1343.6800 ;
        RECT 1341.0200 1332.3200 1342.6200 1332.8000 ;
        RECT 1341.0200 1337.7600 1342.6200 1338.2400 ;
        RECT 1341.0200 1343.2000 1342.6200 1343.6800 ;
        RECT 1296.0200 1375.8400 1297.6200 1376.3200 ;
        RECT 1296.0200 1381.2800 1297.6200 1381.7600 ;
        RECT 1296.0200 1359.5200 1297.6200 1360.0000 ;
        RECT 1296.0200 1364.9600 1297.6200 1365.4400 ;
        RECT 1296.0200 1370.4000 1297.6200 1370.8800 ;
        RECT 1296.0200 1348.6400 1297.6200 1349.1200 ;
        RECT 1296.0200 1354.0800 1297.6200 1354.5600 ;
        RECT 1296.0200 1332.3200 1297.6200 1332.8000 ;
        RECT 1296.0200 1337.7600 1297.6200 1338.2400 ;
        RECT 1296.0200 1343.2000 1297.6200 1343.6800 ;
        RECT 1352.5600 1386.7200 1355.5600 1387.2000 ;
        RECT 1296.0200 1386.7200 1297.6200 1387.2000 ;
        RECT 1341.0200 1386.7200 1342.6200 1387.2000 ;
        RECT 1251.0200 1419.3600 1252.6200 1419.8400 ;
        RECT 1251.0200 1424.8000 1252.6200 1425.2800 ;
        RECT 1251.0200 1430.2400 1252.6200 1430.7200 ;
        RECT 1206.0200 1419.3600 1207.6200 1419.8400 ;
        RECT 1206.0200 1424.8000 1207.6200 1425.2800 ;
        RECT 1206.0200 1430.2400 1207.6200 1430.7200 ;
        RECT 1251.0200 1403.0400 1252.6200 1403.5200 ;
        RECT 1251.0200 1408.4800 1252.6200 1408.9600 ;
        RECT 1251.0200 1392.1600 1252.6200 1392.6400 ;
        RECT 1251.0200 1397.6000 1252.6200 1398.0800 ;
        RECT 1206.0200 1403.0400 1207.6200 1403.5200 ;
        RECT 1206.0200 1408.4800 1207.6200 1408.9600 ;
        RECT 1206.0200 1392.1600 1207.6200 1392.6400 ;
        RECT 1206.0200 1397.6000 1207.6200 1398.0800 ;
        RECT 1206.0200 1413.9200 1207.6200 1414.4000 ;
        RECT 1251.0200 1413.9200 1252.6200 1414.4000 ;
        RECT 1156.4600 1430.2400 1159.4600 1430.7200 ;
        RECT 1156.4600 1424.8000 1159.4600 1425.2800 ;
        RECT 1156.4600 1419.3600 1159.4600 1419.8400 ;
        RECT 1156.4600 1408.4800 1159.4600 1408.9600 ;
        RECT 1156.4600 1403.0400 1159.4600 1403.5200 ;
        RECT 1156.4600 1397.6000 1159.4600 1398.0800 ;
        RECT 1156.4600 1392.1600 1159.4600 1392.6400 ;
        RECT 1156.4600 1413.9200 1159.4600 1414.4000 ;
        RECT 1251.0200 1375.8400 1252.6200 1376.3200 ;
        RECT 1251.0200 1381.2800 1252.6200 1381.7600 ;
        RECT 1251.0200 1359.5200 1252.6200 1360.0000 ;
        RECT 1251.0200 1364.9600 1252.6200 1365.4400 ;
        RECT 1251.0200 1370.4000 1252.6200 1370.8800 ;
        RECT 1206.0200 1375.8400 1207.6200 1376.3200 ;
        RECT 1206.0200 1381.2800 1207.6200 1381.7600 ;
        RECT 1206.0200 1359.5200 1207.6200 1360.0000 ;
        RECT 1206.0200 1364.9600 1207.6200 1365.4400 ;
        RECT 1206.0200 1370.4000 1207.6200 1370.8800 ;
        RECT 1251.0200 1348.6400 1252.6200 1349.1200 ;
        RECT 1251.0200 1354.0800 1252.6200 1354.5600 ;
        RECT 1251.0200 1332.3200 1252.6200 1332.8000 ;
        RECT 1251.0200 1337.7600 1252.6200 1338.2400 ;
        RECT 1251.0200 1343.2000 1252.6200 1343.6800 ;
        RECT 1206.0200 1348.6400 1207.6200 1349.1200 ;
        RECT 1206.0200 1354.0800 1207.6200 1354.5600 ;
        RECT 1206.0200 1332.3200 1207.6200 1332.8000 ;
        RECT 1206.0200 1337.7600 1207.6200 1338.2400 ;
        RECT 1206.0200 1343.2000 1207.6200 1343.6800 ;
        RECT 1156.4600 1375.8400 1159.4600 1376.3200 ;
        RECT 1156.4600 1381.2800 1159.4600 1381.7600 ;
        RECT 1156.4600 1364.9600 1159.4600 1365.4400 ;
        RECT 1156.4600 1359.5200 1159.4600 1360.0000 ;
        RECT 1156.4600 1370.4000 1159.4600 1370.8800 ;
        RECT 1156.4600 1348.6400 1159.4600 1349.1200 ;
        RECT 1156.4600 1354.0800 1159.4600 1354.5600 ;
        RECT 1156.4600 1337.7600 1159.4600 1338.2400 ;
        RECT 1156.4600 1332.3200 1159.4600 1332.8000 ;
        RECT 1156.4600 1343.2000 1159.4600 1343.6800 ;
        RECT 1156.4600 1386.7200 1159.4600 1387.2000 ;
        RECT 1206.0200 1386.7200 1207.6200 1387.2000 ;
        RECT 1251.0200 1386.7200 1252.6200 1387.2000 ;
        RECT 1352.5600 1321.4400 1355.5600 1321.9200 ;
        RECT 1352.5600 1326.8800 1355.5600 1327.3600 ;
        RECT 1341.0200 1321.4400 1342.6200 1321.9200 ;
        RECT 1341.0200 1326.8800 1342.6200 1327.3600 ;
        RECT 1352.5600 1305.1200 1355.5600 1305.6000 ;
        RECT 1352.5600 1310.5600 1355.5600 1311.0400 ;
        RECT 1352.5600 1316.0000 1355.5600 1316.4800 ;
        RECT 1341.0200 1305.1200 1342.6200 1305.6000 ;
        RECT 1341.0200 1310.5600 1342.6200 1311.0400 ;
        RECT 1341.0200 1316.0000 1342.6200 1316.4800 ;
        RECT 1352.5600 1294.2400 1355.5600 1294.7200 ;
        RECT 1352.5600 1299.6800 1355.5600 1300.1600 ;
        RECT 1341.0200 1294.2400 1342.6200 1294.7200 ;
        RECT 1341.0200 1299.6800 1342.6200 1300.1600 ;
        RECT 1352.5600 1277.9200 1355.5600 1278.4000 ;
        RECT 1352.5600 1283.3600 1355.5600 1283.8400 ;
        RECT 1352.5600 1288.8000 1355.5600 1289.2800 ;
        RECT 1341.0200 1277.9200 1342.6200 1278.4000 ;
        RECT 1341.0200 1283.3600 1342.6200 1283.8400 ;
        RECT 1341.0200 1288.8000 1342.6200 1289.2800 ;
        RECT 1296.0200 1321.4400 1297.6200 1321.9200 ;
        RECT 1296.0200 1326.8800 1297.6200 1327.3600 ;
        RECT 1296.0200 1305.1200 1297.6200 1305.6000 ;
        RECT 1296.0200 1310.5600 1297.6200 1311.0400 ;
        RECT 1296.0200 1316.0000 1297.6200 1316.4800 ;
        RECT 1296.0200 1294.2400 1297.6200 1294.7200 ;
        RECT 1296.0200 1299.6800 1297.6200 1300.1600 ;
        RECT 1296.0200 1277.9200 1297.6200 1278.4000 ;
        RECT 1296.0200 1283.3600 1297.6200 1283.8400 ;
        RECT 1296.0200 1288.8000 1297.6200 1289.2800 ;
        RECT 1352.5600 1267.0400 1355.5600 1267.5200 ;
        RECT 1352.5600 1272.4800 1355.5600 1272.9600 ;
        RECT 1341.0200 1267.0400 1342.6200 1267.5200 ;
        RECT 1341.0200 1272.4800 1342.6200 1272.9600 ;
        RECT 1352.5600 1250.7200 1355.5600 1251.2000 ;
        RECT 1352.5600 1256.1600 1355.5600 1256.6400 ;
        RECT 1352.5600 1261.6000 1355.5600 1262.0800 ;
        RECT 1341.0200 1250.7200 1342.6200 1251.2000 ;
        RECT 1341.0200 1256.1600 1342.6200 1256.6400 ;
        RECT 1341.0200 1261.6000 1342.6200 1262.0800 ;
        RECT 1352.5600 1239.8400 1355.5600 1240.3200 ;
        RECT 1352.5600 1245.2800 1355.5600 1245.7600 ;
        RECT 1341.0200 1239.8400 1342.6200 1240.3200 ;
        RECT 1341.0200 1245.2800 1342.6200 1245.7600 ;
        RECT 1352.5600 1234.4000 1355.5600 1234.8800 ;
        RECT 1341.0200 1234.4000 1342.6200 1234.8800 ;
        RECT 1296.0200 1267.0400 1297.6200 1267.5200 ;
        RECT 1296.0200 1272.4800 1297.6200 1272.9600 ;
        RECT 1296.0200 1250.7200 1297.6200 1251.2000 ;
        RECT 1296.0200 1256.1600 1297.6200 1256.6400 ;
        RECT 1296.0200 1261.6000 1297.6200 1262.0800 ;
        RECT 1296.0200 1239.8400 1297.6200 1240.3200 ;
        RECT 1296.0200 1245.2800 1297.6200 1245.7600 ;
        RECT 1296.0200 1234.4000 1297.6200 1234.8800 ;
        RECT 1251.0200 1321.4400 1252.6200 1321.9200 ;
        RECT 1251.0200 1326.8800 1252.6200 1327.3600 ;
        RECT 1251.0200 1305.1200 1252.6200 1305.6000 ;
        RECT 1251.0200 1310.5600 1252.6200 1311.0400 ;
        RECT 1251.0200 1316.0000 1252.6200 1316.4800 ;
        RECT 1206.0200 1321.4400 1207.6200 1321.9200 ;
        RECT 1206.0200 1326.8800 1207.6200 1327.3600 ;
        RECT 1206.0200 1305.1200 1207.6200 1305.6000 ;
        RECT 1206.0200 1310.5600 1207.6200 1311.0400 ;
        RECT 1206.0200 1316.0000 1207.6200 1316.4800 ;
        RECT 1251.0200 1294.2400 1252.6200 1294.7200 ;
        RECT 1251.0200 1299.6800 1252.6200 1300.1600 ;
        RECT 1251.0200 1277.9200 1252.6200 1278.4000 ;
        RECT 1251.0200 1283.3600 1252.6200 1283.8400 ;
        RECT 1251.0200 1288.8000 1252.6200 1289.2800 ;
        RECT 1206.0200 1294.2400 1207.6200 1294.7200 ;
        RECT 1206.0200 1299.6800 1207.6200 1300.1600 ;
        RECT 1206.0200 1277.9200 1207.6200 1278.4000 ;
        RECT 1206.0200 1283.3600 1207.6200 1283.8400 ;
        RECT 1206.0200 1288.8000 1207.6200 1289.2800 ;
        RECT 1156.4600 1321.4400 1159.4600 1321.9200 ;
        RECT 1156.4600 1326.8800 1159.4600 1327.3600 ;
        RECT 1156.4600 1310.5600 1159.4600 1311.0400 ;
        RECT 1156.4600 1305.1200 1159.4600 1305.6000 ;
        RECT 1156.4600 1316.0000 1159.4600 1316.4800 ;
        RECT 1156.4600 1294.2400 1159.4600 1294.7200 ;
        RECT 1156.4600 1299.6800 1159.4600 1300.1600 ;
        RECT 1156.4600 1283.3600 1159.4600 1283.8400 ;
        RECT 1156.4600 1277.9200 1159.4600 1278.4000 ;
        RECT 1156.4600 1288.8000 1159.4600 1289.2800 ;
        RECT 1251.0200 1267.0400 1252.6200 1267.5200 ;
        RECT 1251.0200 1272.4800 1252.6200 1272.9600 ;
        RECT 1251.0200 1250.7200 1252.6200 1251.2000 ;
        RECT 1251.0200 1256.1600 1252.6200 1256.6400 ;
        RECT 1251.0200 1261.6000 1252.6200 1262.0800 ;
        RECT 1206.0200 1267.0400 1207.6200 1267.5200 ;
        RECT 1206.0200 1272.4800 1207.6200 1272.9600 ;
        RECT 1206.0200 1250.7200 1207.6200 1251.2000 ;
        RECT 1206.0200 1256.1600 1207.6200 1256.6400 ;
        RECT 1206.0200 1261.6000 1207.6200 1262.0800 ;
        RECT 1251.0200 1245.2800 1252.6200 1245.7600 ;
        RECT 1251.0200 1239.8400 1252.6200 1240.3200 ;
        RECT 1251.0200 1234.4000 1252.6200 1234.8800 ;
        RECT 1206.0200 1245.2800 1207.6200 1245.7600 ;
        RECT 1206.0200 1239.8400 1207.6200 1240.3200 ;
        RECT 1206.0200 1234.4000 1207.6200 1234.8800 ;
        RECT 1156.4600 1267.0400 1159.4600 1267.5200 ;
        RECT 1156.4600 1272.4800 1159.4600 1272.9600 ;
        RECT 1156.4600 1256.1600 1159.4600 1256.6400 ;
        RECT 1156.4600 1250.7200 1159.4600 1251.2000 ;
        RECT 1156.4600 1261.6000 1159.4600 1262.0800 ;
        RECT 1156.4600 1239.8400 1159.4600 1240.3200 ;
        RECT 1156.4600 1245.2800 1159.4600 1245.7600 ;
        RECT 1156.4600 1234.4000 1159.4600 1234.8800 ;
        RECT 1156.4600 1432.5900 1355.5600 1435.5900 ;
        RECT 1156.4600 1227.4900 1355.5600 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 997.8500 1342.6200 1205.9500 ;
        RECT 1296.0200 997.8500 1297.6200 1205.9500 ;
        RECT 1251.0200 997.8500 1252.6200 1205.9500 ;
        RECT 1206.0200 997.8500 1207.6200 1205.9500 ;
        RECT 1352.5600 997.8500 1355.5600 1205.9500 ;
        RECT 1156.4600 997.8500 1159.4600 1205.9500 ;
      LAYER met3 ;
        RECT 1352.5600 1200.6000 1355.5600 1201.0800 ;
        RECT 1341.0200 1200.6000 1342.6200 1201.0800 ;
        RECT 1352.5600 1189.7200 1355.5600 1190.2000 ;
        RECT 1352.5600 1195.1600 1355.5600 1195.6400 ;
        RECT 1341.0200 1189.7200 1342.6200 1190.2000 ;
        RECT 1341.0200 1195.1600 1342.6200 1195.6400 ;
        RECT 1352.5600 1173.4000 1355.5600 1173.8800 ;
        RECT 1352.5600 1178.8400 1355.5600 1179.3200 ;
        RECT 1341.0200 1173.4000 1342.6200 1173.8800 ;
        RECT 1341.0200 1178.8400 1342.6200 1179.3200 ;
        RECT 1352.5600 1162.5200 1355.5600 1163.0000 ;
        RECT 1352.5600 1167.9600 1355.5600 1168.4400 ;
        RECT 1341.0200 1162.5200 1342.6200 1163.0000 ;
        RECT 1341.0200 1167.9600 1342.6200 1168.4400 ;
        RECT 1352.5600 1184.2800 1355.5600 1184.7600 ;
        RECT 1341.0200 1184.2800 1342.6200 1184.7600 ;
        RECT 1296.0200 1189.7200 1297.6200 1190.2000 ;
        RECT 1296.0200 1195.1600 1297.6200 1195.6400 ;
        RECT 1296.0200 1200.6000 1297.6200 1201.0800 ;
        RECT 1296.0200 1173.4000 1297.6200 1173.8800 ;
        RECT 1296.0200 1178.8400 1297.6200 1179.3200 ;
        RECT 1296.0200 1167.9600 1297.6200 1168.4400 ;
        RECT 1296.0200 1162.5200 1297.6200 1163.0000 ;
        RECT 1296.0200 1184.2800 1297.6200 1184.7600 ;
        RECT 1352.5600 1146.2000 1355.5600 1146.6800 ;
        RECT 1352.5600 1151.6400 1355.5600 1152.1200 ;
        RECT 1341.0200 1146.2000 1342.6200 1146.6800 ;
        RECT 1341.0200 1151.6400 1342.6200 1152.1200 ;
        RECT 1352.5600 1129.8800 1355.5600 1130.3600 ;
        RECT 1352.5600 1135.3200 1355.5600 1135.8000 ;
        RECT 1352.5600 1140.7600 1355.5600 1141.2400 ;
        RECT 1341.0200 1129.8800 1342.6200 1130.3600 ;
        RECT 1341.0200 1135.3200 1342.6200 1135.8000 ;
        RECT 1341.0200 1140.7600 1342.6200 1141.2400 ;
        RECT 1352.5600 1119.0000 1355.5600 1119.4800 ;
        RECT 1352.5600 1124.4400 1355.5600 1124.9200 ;
        RECT 1341.0200 1119.0000 1342.6200 1119.4800 ;
        RECT 1341.0200 1124.4400 1342.6200 1124.9200 ;
        RECT 1352.5600 1102.6800 1355.5600 1103.1600 ;
        RECT 1352.5600 1108.1200 1355.5600 1108.6000 ;
        RECT 1352.5600 1113.5600 1355.5600 1114.0400 ;
        RECT 1341.0200 1102.6800 1342.6200 1103.1600 ;
        RECT 1341.0200 1108.1200 1342.6200 1108.6000 ;
        RECT 1341.0200 1113.5600 1342.6200 1114.0400 ;
        RECT 1296.0200 1146.2000 1297.6200 1146.6800 ;
        RECT 1296.0200 1151.6400 1297.6200 1152.1200 ;
        RECT 1296.0200 1129.8800 1297.6200 1130.3600 ;
        RECT 1296.0200 1135.3200 1297.6200 1135.8000 ;
        RECT 1296.0200 1140.7600 1297.6200 1141.2400 ;
        RECT 1296.0200 1119.0000 1297.6200 1119.4800 ;
        RECT 1296.0200 1124.4400 1297.6200 1124.9200 ;
        RECT 1296.0200 1102.6800 1297.6200 1103.1600 ;
        RECT 1296.0200 1108.1200 1297.6200 1108.6000 ;
        RECT 1296.0200 1113.5600 1297.6200 1114.0400 ;
        RECT 1352.5600 1157.0800 1355.5600 1157.5600 ;
        RECT 1296.0200 1157.0800 1297.6200 1157.5600 ;
        RECT 1341.0200 1157.0800 1342.6200 1157.5600 ;
        RECT 1251.0200 1189.7200 1252.6200 1190.2000 ;
        RECT 1251.0200 1195.1600 1252.6200 1195.6400 ;
        RECT 1251.0200 1200.6000 1252.6200 1201.0800 ;
        RECT 1206.0200 1189.7200 1207.6200 1190.2000 ;
        RECT 1206.0200 1195.1600 1207.6200 1195.6400 ;
        RECT 1206.0200 1200.6000 1207.6200 1201.0800 ;
        RECT 1251.0200 1173.4000 1252.6200 1173.8800 ;
        RECT 1251.0200 1178.8400 1252.6200 1179.3200 ;
        RECT 1251.0200 1162.5200 1252.6200 1163.0000 ;
        RECT 1251.0200 1167.9600 1252.6200 1168.4400 ;
        RECT 1206.0200 1173.4000 1207.6200 1173.8800 ;
        RECT 1206.0200 1178.8400 1207.6200 1179.3200 ;
        RECT 1206.0200 1162.5200 1207.6200 1163.0000 ;
        RECT 1206.0200 1167.9600 1207.6200 1168.4400 ;
        RECT 1206.0200 1184.2800 1207.6200 1184.7600 ;
        RECT 1251.0200 1184.2800 1252.6200 1184.7600 ;
        RECT 1156.4600 1200.6000 1159.4600 1201.0800 ;
        RECT 1156.4600 1195.1600 1159.4600 1195.6400 ;
        RECT 1156.4600 1189.7200 1159.4600 1190.2000 ;
        RECT 1156.4600 1178.8400 1159.4600 1179.3200 ;
        RECT 1156.4600 1173.4000 1159.4600 1173.8800 ;
        RECT 1156.4600 1167.9600 1159.4600 1168.4400 ;
        RECT 1156.4600 1162.5200 1159.4600 1163.0000 ;
        RECT 1156.4600 1184.2800 1159.4600 1184.7600 ;
        RECT 1251.0200 1146.2000 1252.6200 1146.6800 ;
        RECT 1251.0200 1151.6400 1252.6200 1152.1200 ;
        RECT 1251.0200 1129.8800 1252.6200 1130.3600 ;
        RECT 1251.0200 1135.3200 1252.6200 1135.8000 ;
        RECT 1251.0200 1140.7600 1252.6200 1141.2400 ;
        RECT 1206.0200 1146.2000 1207.6200 1146.6800 ;
        RECT 1206.0200 1151.6400 1207.6200 1152.1200 ;
        RECT 1206.0200 1129.8800 1207.6200 1130.3600 ;
        RECT 1206.0200 1135.3200 1207.6200 1135.8000 ;
        RECT 1206.0200 1140.7600 1207.6200 1141.2400 ;
        RECT 1251.0200 1119.0000 1252.6200 1119.4800 ;
        RECT 1251.0200 1124.4400 1252.6200 1124.9200 ;
        RECT 1251.0200 1102.6800 1252.6200 1103.1600 ;
        RECT 1251.0200 1108.1200 1252.6200 1108.6000 ;
        RECT 1251.0200 1113.5600 1252.6200 1114.0400 ;
        RECT 1206.0200 1119.0000 1207.6200 1119.4800 ;
        RECT 1206.0200 1124.4400 1207.6200 1124.9200 ;
        RECT 1206.0200 1102.6800 1207.6200 1103.1600 ;
        RECT 1206.0200 1108.1200 1207.6200 1108.6000 ;
        RECT 1206.0200 1113.5600 1207.6200 1114.0400 ;
        RECT 1156.4600 1146.2000 1159.4600 1146.6800 ;
        RECT 1156.4600 1151.6400 1159.4600 1152.1200 ;
        RECT 1156.4600 1135.3200 1159.4600 1135.8000 ;
        RECT 1156.4600 1129.8800 1159.4600 1130.3600 ;
        RECT 1156.4600 1140.7600 1159.4600 1141.2400 ;
        RECT 1156.4600 1119.0000 1159.4600 1119.4800 ;
        RECT 1156.4600 1124.4400 1159.4600 1124.9200 ;
        RECT 1156.4600 1108.1200 1159.4600 1108.6000 ;
        RECT 1156.4600 1102.6800 1159.4600 1103.1600 ;
        RECT 1156.4600 1113.5600 1159.4600 1114.0400 ;
        RECT 1156.4600 1157.0800 1159.4600 1157.5600 ;
        RECT 1206.0200 1157.0800 1207.6200 1157.5600 ;
        RECT 1251.0200 1157.0800 1252.6200 1157.5600 ;
        RECT 1352.5600 1091.8000 1355.5600 1092.2800 ;
        RECT 1352.5600 1097.2400 1355.5600 1097.7200 ;
        RECT 1341.0200 1091.8000 1342.6200 1092.2800 ;
        RECT 1341.0200 1097.2400 1342.6200 1097.7200 ;
        RECT 1352.5600 1075.4800 1355.5600 1075.9600 ;
        RECT 1352.5600 1080.9200 1355.5600 1081.4000 ;
        RECT 1352.5600 1086.3600 1355.5600 1086.8400 ;
        RECT 1341.0200 1075.4800 1342.6200 1075.9600 ;
        RECT 1341.0200 1080.9200 1342.6200 1081.4000 ;
        RECT 1341.0200 1086.3600 1342.6200 1086.8400 ;
        RECT 1352.5600 1064.6000 1355.5600 1065.0800 ;
        RECT 1352.5600 1070.0400 1355.5600 1070.5200 ;
        RECT 1341.0200 1064.6000 1342.6200 1065.0800 ;
        RECT 1341.0200 1070.0400 1342.6200 1070.5200 ;
        RECT 1352.5600 1048.2800 1355.5600 1048.7600 ;
        RECT 1352.5600 1053.7200 1355.5600 1054.2000 ;
        RECT 1352.5600 1059.1600 1355.5600 1059.6400 ;
        RECT 1341.0200 1048.2800 1342.6200 1048.7600 ;
        RECT 1341.0200 1053.7200 1342.6200 1054.2000 ;
        RECT 1341.0200 1059.1600 1342.6200 1059.6400 ;
        RECT 1296.0200 1091.8000 1297.6200 1092.2800 ;
        RECT 1296.0200 1097.2400 1297.6200 1097.7200 ;
        RECT 1296.0200 1075.4800 1297.6200 1075.9600 ;
        RECT 1296.0200 1080.9200 1297.6200 1081.4000 ;
        RECT 1296.0200 1086.3600 1297.6200 1086.8400 ;
        RECT 1296.0200 1064.6000 1297.6200 1065.0800 ;
        RECT 1296.0200 1070.0400 1297.6200 1070.5200 ;
        RECT 1296.0200 1048.2800 1297.6200 1048.7600 ;
        RECT 1296.0200 1053.7200 1297.6200 1054.2000 ;
        RECT 1296.0200 1059.1600 1297.6200 1059.6400 ;
        RECT 1352.5600 1037.4000 1355.5600 1037.8800 ;
        RECT 1352.5600 1042.8400 1355.5600 1043.3200 ;
        RECT 1341.0200 1037.4000 1342.6200 1037.8800 ;
        RECT 1341.0200 1042.8400 1342.6200 1043.3200 ;
        RECT 1352.5600 1021.0800 1355.5600 1021.5600 ;
        RECT 1352.5600 1026.5200 1355.5600 1027.0000 ;
        RECT 1352.5600 1031.9600 1355.5600 1032.4400 ;
        RECT 1341.0200 1021.0800 1342.6200 1021.5600 ;
        RECT 1341.0200 1026.5200 1342.6200 1027.0000 ;
        RECT 1341.0200 1031.9600 1342.6200 1032.4400 ;
        RECT 1352.5600 1010.2000 1355.5600 1010.6800 ;
        RECT 1352.5600 1015.6400 1355.5600 1016.1200 ;
        RECT 1341.0200 1010.2000 1342.6200 1010.6800 ;
        RECT 1341.0200 1015.6400 1342.6200 1016.1200 ;
        RECT 1352.5600 1004.7600 1355.5600 1005.2400 ;
        RECT 1341.0200 1004.7600 1342.6200 1005.2400 ;
        RECT 1296.0200 1037.4000 1297.6200 1037.8800 ;
        RECT 1296.0200 1042.8400 1297.6200 1043.3200 ;
        RECT 1296.0200 1021.0800 1297.6200 1021.5600 ;
        RECT 1296.0200 1026.5200 1297.6200 1027.0000 ;
        RECT 1296.0200 1031.9600 1297.6200 1032.4400 ;
        RECT 1296.0200 1010.2000 1297.6200 1010.6800 ;
        RECT 1296.0200 1015.6400 1297.6200 1016.1200 ;
        RECT 1296.0200 1004.7600 1297.6200 1005.2400 ;
        RECT 1251.0200 1091.8000 1252.6200 1092.2800 ;
        RECT 1251.0200 1097.2400 1252.6200 1097.7200 ;
        RECT 1251.0200 1075.4800 1252.6200 1075.9600 ;
        RECT 1251.0200 1080.9200 1252.6200 1081.4000 ;
        RECT 1251.0200 1086.3600 1252.6200 1086.8400 ;
        RECT 1206.0200 1091.8000 1207.6200 1092.2800 ;
        RECT 1206.0200 1097.2400 1207.6200 1097.7200 ;
        RECT 1206.0200 1075.4800 1207.6200 1075.9600 ;
        RECT 1206.0200 1080.9200 1207.6200 1081.4000 ;
        RECT 1206.0200 1086.3600 1207.6200 1086.8400 ;
        RECT 1251.0200 1064.6000 1252.6200 1065.0800 ;
        RECT 1251.0200 1070.0400 1252.6200 1070.5200 ;
        RECT 1251.0200 1048.2800 1252.6200 1048.7600 ;
        RECT 1251.0200 1053.7200 1252.6200 1054.2000 ;
        RECT 1251.0200 1059.1600 1252.6200 1059.6400 ;
        RECT 1206.0200 1064.6000 1207.6200 1065.0800 ;
        RECT 1206.0200 1070.0400 1207.6200 1070.5200 ;
        RECT 1206.0200 1048.2800 1207.6200 1048.7600 ;
        RECT 1206.0200 1053.7200 1207.6200 1054.2000 ;
        RECT 1206.0200 1059.1600 1207.6200 1059.6400 ;
        RECT 1156.4600 1091.8000 1159.4600 1092.2800 ;
        RECT 1156.4600 1097.2400 1159.4600 1097.7200 ;
        RECT 1156.4600 1080.9200 1159.4600 1081.4000 ;
        RECT 1156.4600 1075.4800 1159.4600 1075.9600 ;
        RECT 1156.4600 1086.3600 1159.4600 1086.8400 ;
        RECT 1156.4600 1064.6000 1159.4600 1065.0800 ;
        RECT 1156.4600 1070.0400 1159.4600 1070.5200 ;
        RECT 1156.4600 1053.7200 1159.4600 1054.2000 ;
        RECT 1156.4600 1048.2800 1159.4600 1048.7600 ;
        RECT 1156.4600 1059.1600 1159.4600 1059.6400 ;
        RECT 1251.0200 1037.4000 1252.6200 1037.8800 ;
        RECT 1251.0200 1042.8400 1252.6200 1043.3200 ;
        RECT 1251.0200 1021.0800 1252.6200 1021.5600 ;
        RECT 1251.0200 1026.5200 1252.6200 1027.0000 ;
        RECT 1251.0200 1031.9600 1252.6200 1032.4400 ;
        RECT 1206.0200 1037.4000 1207.6200 1037.8800 ;
        RECT 1206.0200 1042.8400 1207.6200 1043.3200 ;
        RECT 1206.0200 1021.0800 1207.6200 1021.5600 ;
        RECT 1206.0200 1026.5200 1207.6200 1027.0000 ;
        RECT 1206.0200 1031.9600 1207.6200 1032.4400 ;
        RECT 1251.0200 1015.6400 1252.6200 1016.1200 ;
        RECT 1251.0200 1010.2000 1252.6200 1010.6800 ;
        RECT 1251.0200 1004.7600 1252.6200 1005.2400 ;
        RECT 1206.0200 1015.6400 1207.6200 1016.1200 ;
        RECT 1206.0200 1010.2000 1207.6200 1010.6800 ;
        RECT 1206.0200 1004.7600 1207.6200 1005.2400 ;
        RECT 1156.4600 1037.4000 1159.4600 1037.8800 ;
        RECT 1156.4600 1042.8400 1159.4600 1043.3200 ;
        RECT 1156.4600 1026.5200 1159.4600 1027.0000 ;
        RECT 1156.4600 1021.0800 1159.4600 1021.5600 ;
        RECT 1156.4600 1031.9600 1159.4600 1032.4400 ;
        RECT 1156.4600 1010.2000 1159.4600 1010.6800 ;
        RECT 1156.4600 1015.6400 1159.4600 1016.1200 ;
        RECT 1156.4600 1004.7600 1159.4600 1005.2400 ;
        RECT 1156.4600 1202.9500 1355.5600 1205.9500 ;
        RECT 1156.4600 997.8500 1355.5600 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1341.0200 768.2100 1342.6200 976.3100 ;
        RECT 1296.0200 768.2100 1297.6200 976.3100 ;
        RECT 1251.0200 768.2100 1252.6200 976.3100 ;
        RECT 1206.0200 768.2100 1207.6200 976.3100 ;
        RECT 1352.5600 768.2100 1355.5600 976.3100 ;
        RECT 1156.4600 768.2100 1159.4600 976.3100 ;
      LAYER met3 ;
        RECT 1352.5600 970.9600 1355.5600 971.4400 ;
        RECT 1341.0200 970.9600 1342.6200 971.4400 ;
        RECT 1352.5600 960.0800 1355.5600 960.5600 ;
        RECT 1352.5600 965.5200 1355.5600 966.0000 ;
        RECT 1341.0200 960.0800 1342.6200 960.5600 ;
        RECT 1341.0200 965.5200 1342.6200 966.0000 ;
        RECT 1352.5600 943.7600 1355.5600 944.2400 ;
        RECT 1352.5600 949.2000 1355.5600 949.6800 ;
        RECT 1341.0200 943.7600 1342.6200 944.2400 ;
        RECT 1341.0200 949.2000 1342.6200 949.6800 ;
        RECT 1352.5600 932.8800 1355.5600 933.3600 ;
        RECT 1352.5600 938.3200 1355.5600 938.8000 ;
        RECT 1341.0200 932.8800 1342.6200 933.3600 ;
        RECT 1341.0200 938.3200 1342.6200 938.8000 ;
        RECT 1352.5600 954.6400 1355.5600 955.1200 ;
        RECT 1341.0200 954.6400 1342.6200 955.1200 ;
        RECT 1296.0200 960.0800 1297.6200 960.5600 ;
        RECT 1296.0200 965.5200 1297.6200 966.0000 ;
        RECT 1296.0200 970.9600 1297.6200 971.4400 ;
        RECT 1296.0200 943.7600 1297.6200 944.2400 ;
        RECT 1296.0200 949.2000 1297.6200 949.6800 ;
        RECT 1296.0200 938.3200 1297.6200 938.8000 ;
        RECT 1296.0200 932.8800 1297.6200 933.3600 ;
        RECT 1296.0200 954.6400 1297.6200 955.1200 ;
        RECT 1352.5600 916.5600 1355.5600 917.0400 ;
        RECT 1352.5600 922.0000 1355.5600 922.4800 ;
        RECT 1341.0200 916.5600 1342.6200 917.0400 ;
        RECT 1341.0200 922.0000 1342.6200 922.4800 ;
        RECT 1352.5600 900.2400 1355.5600 900.7200 ;
        RECT 1352.5600 905.6800 1355.5600 906.1600 ;
        RECT 1352.5600 911.1200 1355.5600 911.6000 ;
        RECT 1341.0200 900.2400 1342.6200 900.7200 ;
        RECT 1341.0200 905.6800 1342.6200 906.1600 ;
        RECT 1341.0200 911.1200 1342.6200 911.6000 ;
        RECT 1352.5600 889.3600 1355.5600 889.8400 ;
        RECT 1352.5600 894.8000 1355.5600 895.2800 ;
        RECT 1341.0200 889.3600 1342.6200 889.8400 ;
        RECT 1341.0200 894.8000 1342.6200 895.2800 ;
        RECT 1352.5600 873.0400 1355.5600 873.5200 ;
        RECT 1352.5600 878.4800 1355.5600 878.9600 ;
        RECT 1352.5600 883.9200 1355.5600 884.4000 ;
        RECT 1341.0200 873.0400 1342.6200 873.5200 ;
        RECT 1341.0200 878.4800 1342.6200 878.9600 ;
        RECT 1341.0200 883.9200 1342.6200 884.4000 ;
        RECT 1296.0200 916.5600 1297.6200 917.0400 ;
        RECT 1296.0200 922.0000 1297.6200 922.4800 ;
        RECT 1296.0200 900.2400 1297.6200 900.7200 ;
        RECT 1296.0200 905.6800 1297.6200 906.1600 ;
        RECT 1296.0200 911.1200 1297.6200 911.6000 ;
        RECT 1296.0200 889.3600 1297.6200 889.8400 ;
        RECT 1296.0200 894.8000 1297.6200 895.2800 ;
        RECT 1296.0200 873.0400 1297.6200 873.5200 ;
        RECT 1296.0200 878.4800 1297.6200 878.9600 ;
        RECT 1296.0200 883.9200 1297.6200 884.4000 ;
        RECT 1352.5600 927.4400 1355.5600 927.9200 ;
        RECT 1296.0200 927.4400 1297.6200 927.9200 ;
        RECT 1341.0200 927.4400 1342.6200 927.9200 ;
        RECT 1251.0200 960.0800 1252.6200 960.5600 ;
        RECT 1251.0200 965.5200 1252.6200 966.0000 ;
        RECT 1251.0200 970.9600 1252.6200 971.4400 ;
        RECT 1206.0200 960.0800 1207.6200 960.5600 ;
        RECT 1206.0200 965.5200 1207.6200 966.0000 ;
        RECT 1206.0200 970.9600 1207.6200 971.4400 ;
        RECT 1251.0200 943.7600 1252.6200 944.2400 ;
        RECT 1251.0200 949.2000 1252.6200 949.6800 ;
        RECT 1251.0200 932.8800 1252.6200 933.3600 ;
        RECT 1251.0200 938.3200 1252.6200 938.8000 ;
        RECT 1206.0200 943.7600 1207.6200 944.2400 ;
        RECT 1206.0200 949.2000 1207.6200 949.6800 ;
        RECT 1206.0200 932.8800 1207.6200 933.3600 ;
        RECT 1206.0200 938.3200 1207.6200 938.8000 ;
        RECT 1206.0200 954.6400 1207.6200 955.1200 ;
        RECT 1251.0200 954.6400 1252.6200 955.1200 ;
        RECT 1156.4600 970.9600 1159.4600 971.4400 ;
        RECT 1156.4600 965.5200 1159.4600 966.0000 ;
        RECT 1156.4600 960.0800 1159.4600 960.5600 ;
        RECT 1156.4600 949.2000 1159.4600 949.6800 ;
        RECT 1156.4600 943.7600 1159.4600 944.2400 ;
        RECT 1156.4600 938.3200 1159.4600 938.8000 ;
        RECT 1156.4600 932.8800 1159.4600 933.3600 ;
        RECT 1156.4600 954.6400 1159.4600 955.1200 ;
        RECT 1251.0200 916.5600 1252.6200 917.0400 ;
        RECT 1251.0200 922.0000 1252.6200 922.4800 ;
        RECT 1251.0200 900.2400 1252.6200 900.7200 ;
        RECT 1251.0200 905.6800 1252.6200 906.1600 ;
        RECT 1251.0200 911.1200 1252.6200 911.6000 ;
        RECT 1206.0200 916.5600 1207.6200 917.0400 ;
        RECT 1206.0200 922.0000 1207.6200 922.4800 ;
        RECT 1206.0200 900.2400 1207.6200 900.7200 ;
        RECT 1206.0200 905.6800 1207.6200 906.1600 ;
        RECT 1206.0200 911.1200 1207.6200 911.6000 ;
        RECT 1251.0200 889.3600 1252.6200 889.8400 ;
        RECT 1251.0200 894.8000 1252.6200 895.2800 ;
        RECT 1251.0200 873.0400 1252.6200 873.5200 ;
        RECT 1251.0200 878.4800 1252.6200 878.9600 ;
        RECT 1251.0200 883.9200 1252.6200 884.4000 ;
        RECT 1206.0200 889.3600 1207.6200 889.8400 ;
        RECT 1206.0200 894.8000 1207.6200 895.2800 ;
        RECT 1206.0200 873.0400 1207.6200 873.5200 ;
        RECT 1206.0200 878.4800 1207.6200 878.9600 ;
        RECT 1206.0200 883.9200 1207.6200 884.4000 ;
        RECT 1156.4600 916.5600 1159.4600 917.0400 ;
        RECT 1156.4600 922.0000 1159.4600 922.4800 ;
        RECT 1156.4600 905.6800 1159.4600 906.1600 ;
        RECT 1156.4600 900.2400 1159.4600 900.7200 ;
        RECT 1156.4600 911.1200 1159.4600 911.6000 ;
        RECT 1156.4600 889.3600 1159.4600 889.8400 ;
        RECT 1156.4600 894.8000 1159.4600 895.2800 ;
        RECT 1156.4600 878.4800 1159.4600 878.9600 ;
        RECT 1156.4600 873.0400 1159.4600 873.5200 ;
        RECT 1156.4600 883.9200 1159.4600 884.4000 ;
        RECT 1156.4600 927.4400 1159.4600 927.9200 ;
        RECT 1206.0200 927.4400 1207.6200 927.9200 ;
        RECT 1251.0200 927.4400 1252.6200 927.9200 ;
        RECT 1352.5600 862.1600 1355.5600 862.6400 ;
        RECT 1352.5600 867.6000 1355.5600 868.0800 ;
        RECT 1341.0200 862.1600 1342.6200 862.6400 ;
        RECT 1341.0200 867.6000 1342.6200 868.0800 ;
        RECT 1352.5600 845.8400 1355.5600 846.3200 ;
        RECT 1352.5600 851.2800 1355.5600 851.7600 ;
        RECT 1352.5600 856.7200 1355.5600 857.2000 ;
        RECT 1341.0200 845.8400 1342.6200 846.3200 ;
        RECT 1341.0200 851.2800 1342.6200 851.7600 ;
        RECT 1341.0200 856.7200 1342.6200 857.2000 ;
        RECT 1352.5600 834.9600 1355.5600 835.4400 ;
        RECT 1352.5600 840.4000 1355.5600 840.8800 ;
        RECT 1341.0200 834.9600 1342.6200 835.4400 ;
        RECT 1341.0200 840.4000 1342.6200 840.8800 ;
        RECT 1352.5600 818.6400 1355.5600 819.1200 ;
        RECT 1352.5600 824.0800 1355.5600 824.5600 ;
        RECT 1352.5600 829.5200 1355.5600 830.0000 ;
        RECT 1341.0200 818.6400 1342.6200 819.1200 ;
        RECT 1341.0200 824.0800 1342.6200 824.5600 ;
        RECT 1341.0200 829.5200 1342.6200 830.0000 ;
        RECT 1296.0200 862.1600 1297.6200 862.6400 ;
        RECT 1296.0200 867.6000 1297.6200 868.0800 ;
        RECT 1296.0200 845.8400 1297.6200 846.3200 ;
        RECT 1296.0200 851.2800 1297.6200 851.7600 ;
        RECT 1296.0200 856.7200 1297.6200 857.2000 ;
        RECT 1296.0200 834.9600 1297.6200 835.4400 ;
        RECT 1296.0200 840.4000 1297.6200 840.8800 ;
        RECT 1296.0200 818.6400 1297.6200 819.1200 ;
        RECT 1296.0200 824.0800 1297.6200 824.5600 ;
        RECT 1296.0200 829.5200 1297.6200 830.0000 ;
        RECT 1352.5600 807.7600 1355.5600 808.2400 ;
        RECT 1352.5600 813.2000 1355.5600 813.6800 ;
        RECT 1341.0200 807.7600 1342.6200 808.2400 ;
        RECT 1341.0200 813.2000 1342.6200 813.6800 ;
        RECT 1352.5600 791.4400 1355.5600 791.9200 ;
        RECT 1352.5600 796.8800 1355.5600 797.3600 ;
        RECT 1352.5600 802.3200 1355.5600 802.8000 ;
        RECT 1341.0200 791.4400 1342.6200 791.9200 ;
        RECT 1341.0200 796.8800 1342.6200 797.3600 ;
        RECT 1341.0200 802.3200 1342.6200 802.8000 ;
        RECT 1352.5600 780.5600 1355.5600 781.0400 ;
        RECT 1352.5600 786.0000 1355.5600 786.4800 ;
        RECT 1341.0200 780.5600 1342.6200 781.0400 ;
        RECT 1341.0200 786.0000 1342.6200 786.4800 ;
        RECT 1352.5600 775.1200 1355.5600 775.6000 ;
        RECT 1341.0200 775.1200 1342.6200 775.6000 ;
        RECT 1296.0200 807.7600 1297.6200 808.2400 ;
        RECT 1296.0200 813.2000 1297.6200 813.6800 ;
        RECT 1296.0200 791.4400 1297.6200 791.9200 ;
        RECT 1296.0200 796.8800 1297.6200 797.3600 ;
        RECT 1296.0200 802.3200 1297.6200 802.8000 ;
        RECT 1296.0200 780.5600 1297.6200 781.0400 ;
        RECT 1296.0200 786.0000 1297.6200 786.4800 ;
        RECT 1296.0200 775.1200 1297.6200 775.6000 ;
        RECT 1251.0200 862.1600 1252.6200 862.6400 ;
        RECT 1251.0200 867.6000 1252.6200 868.0800 ;
        RECT 1251.0200 845.8400 1252.6200 846.3200 ;
        RECT 1251.0200 851.2800 1252.6200 851.7600 ;
        RECT 1251.0200 856.7200 1252.6200 857.2000 ;
        RECT 1206.0200 862.1600 1207.6200 862.6400 ;
        RECT 1206.0200 867.6000 1207.6200 868.0800 ;
        RECT 1206.0200 845.8400 1207.6200 846.3200 ;
        RECT 1206.0200 851.2800 1207.6200 851.7600 ;
        RECT 1206.0200 856.7200 1207.6200 857.2000 ;
        RECT 1251.0200 834.9600 1252.6200 835.4400 ;
        RECT 1251.0200 840.4000 1252.6200 840.8800 ;
        RECT 1251.0200 818.6400 1252.6200 819.1200 ;
        RECT 1251.0200 824.0800 1252.6200 824.5600 ;
        RECT 1251.0200 829.5200 1252.6200 830.0000 ;
        RECT 1206.0200 834.9600 1207.6200 835.4400 ;
        RECT 1206.0200 840.4000 1207.6200 840.8800 ;
        RECT 1206.0200 818.6400 1207.6200 819.1200 ;
        RECT 1206.0200 824.0800 1207.6200 824.5600 ;
        RECT 1206.0200 829.5200 1207.6200 830.0000 ;
        RECT 1156.4600 862.1600 1159.4600 862.6400 ;
        RECT 1156.4600 867.6000 1159.4600 868.0800 ;
        RECT 1156.4600 851.2800 1159.4600 851.7600 ;
        RECT 1156.4600 845.8400 1159.4600 846.3200 ;
        RECT 1156.4600 856.7200 1159.4600 857.2000 ;
        RECT 1156.4600 834.9600 1159.4600 835.4400 ;
        RECT 1156.4600 840.4000 1159.4600 840.8800 ;
        RECT 1156.4600 824.0800 1159.4600 824.5600 ;
        RECT 1156.4600 818.6400 1159.4600 819.1200 ;
        RECT 1156.4600 829.5200 1159.4600 830.0000 ;
        RECT 1251.0200 807.7600 1252.6200 808.2400 ;
        RECT 1251.0200 813.2000 1252.6200 813.6800 ;
        RECT 1251.0200 791.4400 1252.6200 791.9200 ;
        RECT 1251.0200 796.8800 1252.6200 797.3600 ;
        RECT 1251.0200 802.3200 1252.6200 802.8000 ;
        RECT 1206.0200 807.7600 1207.6200 808.2400 ;
        RECT 1206.0200 813.2000 1207.6200 813.6800 ;
        RECT 1206.0200 791.4400 1207.6200 791.9200 ;
        RECT 1206.0200 796.8800 1207.6200 797.3600 ;
        RECT 1206.0200 802.3200 1207.6200 802.8000 ;
        RECT 1251.0200 786.0000 1252.6200 786.4800 ;
        RECT 1251.0200 780.5600 1252.6200 781.0400 ;
        RECT 1251.0200 775.1200 1252.6200 775.6000 ;
        RECT 1206.0200 786.0000 1207.6200 786.4800 ;
        RECT 1206.0200 780.5600 1207.6200 781.0400 ;
        RECT 1206.0200 775.1200 1207.6200 775.6000 ;
        RECT 1156.4600 807.7600 1159.4600 808.2400 ;
        RECT 1156.4600 813.2000 1159.4600 813.6800 ;
        RECT 1156.4600 796.8800 1159.4600 797.3600 ;
        RECT 1156.4600 791.4400 1159.4600 791.9200 ;
        RECT 1156.4600 802.3200 1159.4600 802.8000 ;
        RECT 1156.4600 780.5600 1159.4600 781.0400 ;
        RECT 1156.4600 786.0000 1159.4600 786.4800 ;
        RECT 1156.4600 775.1200 1159.4600 775.6000 ;
        RECT 1156.4600 973.3100 1355.5600 976.3100 ;
        RECT 1156.4600 768.2100 1355.5600 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1376.6800 2833.6100 1378.6800 2854.5400 ;
        RECT 1573.7800 2833.6100 1575.7800 2854.5400 ;
      LAYER met3 ;
        RECT 1573.7800 2850.0400 1575.7800 2850.5200 ;
        RECT 1376.6800 2850.0400 1378.6800 2850.5200 ;
        RECT 1573.7800 2839.1600 1575.7800 2839.6400 ;
        RECT 1376.6800 2839.1600 1378.6800 2839.6400 ;
        RECT 1573.7800 2844.6000 1575.7800 2845.0800 ;
        RECT 1376.6800 2844.6000 1378.6800 2845.0800 ;
        RECT 1376.6800 2852.5400 1575.7800 2854.5400 ;
        RECT 1376.6800 2833.6100 1575.7800 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 538.5700 1562.8400 746.6700 ;
        RECT 1516.2400 538.5700 1517.8400 746.6700 ;
        RECT 1471.2400 538.5700 1472.8400 746.6700 ;
        RECT 1426.2400 538.5700 1427.8400 746.6700 ;
        RECT 1572.7800 538.5700 1575.7800 746.6700 ;
        RECT 1376.6800 538.5700 1379.6800 746.6700 ;
      LAYER met3 ;
        RECT 1572.7800 741.3200 1575.7800 741.8000 ;
        RECT 1561.2400 741.3200 1562.8400 741.8000 ;
        RECT 1572.7800 730.4400 1575.7800 730.9200 ;
        RECT 1572.7800 735.8800 1575.7800 736.3600 ;
        RECT 1561.2400 730.4400 1562.8400 730.9200 ;
        RECT 1561.2400 735.8800 1562.8400 736.3600 ;
        RECT 1572.7800 714.1200 1575.7800 714.6000 ;
        RECT 1572.7800 719.5600 1575.7800 720.0400 ;
        RECT 1561.2400 714.1200 1562.8400 714.6000 ;
        RECT 1561.2400 719.5600 1562.8400 720.0400 ;
        RECT 1572.7800 703.2400 1575.7800 703.7200 ;
        RECT 1572.7800 708.6800 1575.7800 709.1600 ;
        RECT 1561.2400 703.2400 1562.8400 703.7200 ;
        RECT 1561.2400 708.6800 1562.8400 709.1600 ;
        RECT 1572.7800 725.0000 1575.7800 725.4800 ;
        RECT 1561.2400 725.0000 1562.8400 725.4800 ;
        RECT 1516.2400 730.4400 1517.8400 730.9200 ;
        RECT 1516.2400 735.8800 1517.8400 736.3600 ;
        RECT 1516.2400 741.3200 1517.8400 741.8000 ;
        RECT 1516.2400 714.1200 1517.8400 714.6000 ;
        RECT 1516.2400 719.5600 1517.8400 720.0400 ;
        RECT 1516.2400 708.6800 1517.8400 709.1600 ;
        RECT 1516.2400 703.2400 1517.8400 703.7200 ;
        RECT 1516.2400 725.0000 1517.8400 725.4800 ;
        RECT 1572.7800 686.9200 1575.7800 687.4000 ;
        RECT 1572.7800 692.3600 1575.7800 692.8400 ;
        RECT 1561.2400 686.9200 1562.8400 687.4000 ;
        RECT 1561.2400 692.3600 1562.8400 692.8400 ;
        RECT 1572.7800 670.6000 1575.7800 671.0800 ;
        RECT 1572.7800 676.0400 1575.7800 676.5200 ;
        RECT 1572.7800 681.4800 1575.7800 681.9600 ;
        RECT 1561.2400 670.6000 1562.8400 671.0800 ;
        RECT 1561.2400 676.0400 1562.8400 676.5200 ;
        RECT 1561.2400 681.4800 1562.8400 681.9600 ;
        RECT 1572.7800 659.7200 1575.7800 660.2000 ;
        RECT 1572.7800 665.1600 1575.7800 665.6400 ;
        RECT 1561.2400 659.7200 1562.8400 660.2000 ;
        RECT 1561.2400 665.1600 1562.8400 665.6400 ;
        RECT 1572.7800 643.4000 1575.7800 643.8800 ;
        RECT 1572.7800 648.8400 1575.7800 649.3200 ;
        RECT 1572.7800 654.2800 1575.7800 654.7600 ;
        RECT 1561.2400 643.4000 1562.8400 643.8800 ;
        RECT 1561.2400 648.8400 1562.8400 649.3200 ;
        RECT 1561.2400 654.2800 1562.8400 654.7600 ;
        RECT 1516.2400 686.9200 1517.8400 687.4000 ;
        RECT 1516.2400 692.3600 1517.8400 692.8400 ;
        RECT 1516.2400 670.6000 1517.8400 671.0800 ;
        RECT 1516.2400 676.0400 1517.8400 676.5200 ;
        RECT 1516.2400 681.4800 1517.8400 681.9600 ;
        RECT 1516.2400 659.7200 1517.8400 660.2000 ;
        RECT 1516.2400 665.1600 1517.8400 665.6400 ;
        RECT 1516.2400 643.4000 1517.8400 643.8800 ;
        RECT 1516.2400 648.8400 1517.8400 649.3200 ;
        RECT 1516.2400 654.2800 1517.8400 654.7600 ;
        RECT 1572.7800 697.8000 1575.7800 698.2800 ;
        RECT 1516.2400 697.8000 1517.8400 698.2800 ;
        RECT 1561.2400 697.8000 1562.8400 698.2800 ;
        RECT 1471.2400 730.4400 1472.8400 730.9200 ;
        RECT 1471.2400 735.8800 1472.8400 736.3600 ;
        RECT 1471.2400 741.3200 1472.8400 741.8000 ;
        RECT 1426.2400 730.4400 1427.8400 730.9200 ;
        RECT 1426.2400 735.8800 1427.8400 736.3600 ;
        RECT 1426.2400 741.3200 1427.8400 741.8000 ;
        RECT 1471.2400 714.1200 1472.8400 714.6000 ;
        RECT 1471.2400 719.5600 1472.8400 720.0400 ;
        RECT 1471.2400 703.2400 1472.8400 703.7200 ;
        RECT 1471.2400 708.6800 1472.8400 709.1600 ;
        RECT 1426.2400 714.1200 1427.8400 714.6000 ;
        RECT 1426.2400 719.5600 1427.8400 720.0400 ;
        RECT 1426.2400 703.2400 1427.8400 703.7200 ;
        RECT 1426.2400 708.6800 1427.8400 709.1600 ;
        RECT 1426.2400 725.0000 1427.8400 725.4800 ;
        RECT 1471.2400 725.0000 1472.8400 725.4800 ;
        RECT 1376.6800 741.3200 1379.6800 741.8000 ;
        RECT 1376.6800 735.8800 1379.6800 736.3600 ;
        RECT 1376.6800 730.4400 1379.6800 730.9200 ;
        RECT 1376.6800 719.5600 1379.6800 720.0400 ;
        RECT 1376.6800 714.1200 1379.6800 714.6000 ;
        RECT 1376.6800 708.6800 1379.6800 709.1600 ;
        RECT 1376.6800 703.2400 1379.6800 703.7200 ;
        RECT 1376.6800 725.0000 1379.6800 725.4800 ;
        RECT 1471.2400 686.9200 1472.8400 687.4000 ;
        RECT 1471.2400 692.3600 1472.8400 692.8400 ;
        RECT 1471.2400 670.6000 1472.8400 671.0800 ;
        RECT 1471.2400 676.0400 1472.8400 676.5200 ;
        RECT 1471.2400 681.4800 1472.8400 681.9600 ;
        RECT 1426.2400 686.9200 1427.8400 687.4000 ;
        RECT 1426.2400 692.3600 1427.8400 692.8400 ;
        RECT 1426.2400 670.6000 1427.8400 671.0800 ;
        RECT 1426.2400 676.0400 1427.8400 676.5200 ;
        RECT 1426.2400 681.4800 1427.8400 681.9600 ;
        RECT 1471.2400 659.7200 1472.8400 660.2000 ;
        RECT 1471.2400 665.1600 1472.8400 665.6400 ;
        RECT 1471.2400 643.4000 1472.8400 643.8800 ;
        RECT 1471.2400 648.8400 1472.8400 649.3200 ;
        RECT 1471.2400 654.2800 1472.8400 654.7600 ;
        RECT 1426.2400 659.7200 1427.8400 660.2000 ;
        RECT 1426.2400 665.1600 1427.8400 665.6400 ;
        RECT 1426.2400 643.4000 1427.8400 643.8800 ;
        RECT 1426.2400 648.8400 1427.8400 649.3200 ;
        RECT 1426.2400 654.2800 1427.8400 654.7600 ;
        RECT 1376.6800 686.9200 1379.6800 687.4000 ;
        RECT 1376.6800 692.3600 1379.6800 692.8400 ;
        RECT 1376.6800 676.0400 1379.6800 676.5200 ;
        RECT 1376.6800 670.6000 1379.6800 671.0800 ;
        RECT 1376.6800 681.4800 1379.6800 681.9600 ;
        RECT 1376.6800 659.7200 1379.6800 660.2000 ;
        RECT 1376.6800 665.1600 1379.6800 665.6400 ;
        RECT 1376.6800 648.8400 1379.6800 649.3200 ;
        RECT 1376.6800 643.4000 1379.6800 643.8800 ;
        RECT 1376.6800 654.2800 1379.6800 654.7600 ;
        RECT 1376.6800 697.8000 1379.6800 698.2800 ;
        RECT 1426.2400 697.8000 1427.8400 698.2800 ;
        RECT 1471.2400 697.8000 1472.8400 698.2800 ;
        RECT 1572.7800 632.5200 1575.7800 633.0000 ;
        RECT 1572.7800 637.9600 1575.7800 638.4400 ;
        RECT 1561.2400 632.5200 1562.8400 633.0000 ;
        RECT 1561.2400 637.9600 1562.8400 638.4400 ;
        RECT 1572.7800 616.2000 1575.7800 616.6800 ;
        RECT 1572.7800 621.6400 1575.7800 622.1200 ;
        RECT 1572.7800 627.0800 1575.7800 627.5600 ;
        RECT 1561.2400 616.2000 1562.8400 616.6800 ;
        RECT 1561.2400 621.6400 1562.8400 622.1200 ;
        RECT 1561.2400 627.0800 1562.8400 627.5600 ;
        RECT 1572.7800 605.3200 1575.7800 605.8000 ;
        RECT 1572.7800 610.7600 1575.7800 611.2400 ;
        RECT 1561.2400 605.3200 1562.8400 605.8000 ;
        RECT 1561.2400 610.7600 1562.8400 611.2400 ;
        RECT 1572.7800 589.0000 1575.7800 589.4800 ;
        RECT 1572.7800 594.4400 1575.7800 594.9200 ;
        RECT 1572.7800 599.8800 1575.7800 600.3600 ;
        RECT 1561.2400 589.0000 1562.8400 589.4800 ;
        RECT 1561.2400 594.4400 1562.8400 594.9200 ;
        RECT 1561.2400 599.8800 1562.8400 600.3600 ;
        RECT 1516.2400 632.5200 1517.8400 633.0000 ;
        RECT 1516.2400 637.9600 1517.8400 638.4400 ;
        RECT 1516.2400 616.2000 1517.8400 616.6800 ;
        RECT 1516.2400 621.6400 1517.8400 622.1200 ;
        RECT 1516.2400 627.0800 1517.8400 627.5600 ;
        RECT 1516.2400 605.3200 1517.8400 605.8000 ;
        RECT 1516.2400 610.7600 1517.8400 611.2400 ;
        RECT 1516.2400 589.0000 1517.8400 589.4800 ;
        RECT 1516.2400 594.4400 1517.8400 594.9200 ;
        RECT 1516.2400 599.8800 1517.8400 600.3600 ;
        RECT 1572.7800 578.1200 1575.7800 578.6000 ;
        RECT 1572.7800 583.5600 1575.7800 584.0400 ;
        RECT 1561.2400 578.1200 1562.8400 578.6000 ;
        RECT 1561.2400 583.5600 1562.8400 584.0400 ;
        RECT 1572.7800 561.8000 1575.7800 562.2800 ;
        RECT 1572.7800 567.2400 1575.7800 567.7200 ;
        RECT 1572.7800 572.6800 1575.7800 573.1600 ;
        RECT 1561.2400 561.8000 1562.8400 562.2800 ;
        RECT 1561.2400 567.2400 1562.8400 567.7200 ;
        RECT 1561.2400 572.6800 1562.8400 573.1600 ;
        RECT 1572.7800 550.9200 1575.7800 551.4000 ;
        RECT 1572.7800 556.3600 1575.7800 556.8400 ;
        RECT 1561.2400 550.9200 1562.8400 551.4000 ;
        RECT 1561.2400 556.3600 1562.8400 556.8400 ;
        RECT 1572.7800 545.4800 1575.7800 545.9600 ;
        RECT 1561.2400 545.4800 1562.8400 545.9600 ;
        RECT 1516.2400 578.1200 1517.8400 578.6000 ;
        RECT 1516.2400 583.5600 1517.8400 584.0400 ;
        RECT 1516.2400 561.8000 1517.8400 562.2800 ;
        RECT 1516.2400 567.2400 1517.8400 567.7200 ;
        RECT 1516.2400 572.6800 1517.8400 573.1600 ;
        RECT 1516.2400 550.9200 1517.8400 551.4000 ;
        RECT 1516.2400 556.3600 1517.8400 556.8400 ;
        RECT 1516.2400 545.4800 1517.8400 545.9600 ;
        RECT 1471.2400 632.5200 1472.8400 633.0000 ;
        RECT 1471.2400 637.9600 1472.8400 638.4400 ;
        RECT 1471.2400 616.2000 1472.8400 616.6800 ;
        RECT 1471.2400 621.6400 1472.8400 622.1200 ;
        RECT 1471.2400 627.0800 1472.8400 627.5600 ;
        RECT 1426.2400 632.5200 1427.8400 633.0000 ;
        RECT 1426.2400 637.9600 1427.8400 638.4400 ;
        RECT 1426.2400 616.2000 1427.8400 616.6800 ;
        RECT 1426.2400 621.6400 1427.8400 622.1200 ;
        RECT 1426.2400 627.0800 1427.8400 627.5600 ;
        RECT 1471.2400 605.3200 1472.8400 605.8000 ;
        RECT 1471.2400 610.7600 1472.8400 611.2400 ;
        RECT 1471.2400 589.0000 1472.8400 589.4800 ;
        RECT 1471.2400 594.4400 1472.8400 594.9200 ;
        RECT 1471.2400 599.8800 1472.8400 600.3600 ;
        RECT 1426.2400 605.3200 1427.8400 605.8000 ;
        RECT 1426.2400 610.7600 1427.8400 611.2400 ;
        RECT 1426.2400 589.0000 1427.8400 589.4800 ;
        RECT 1426.2400 594.4400 1427.8400 594.9200 ;
        RECT 1426.2400 599.8800 1427.8400 600.3600 ;
        RECT 1376.6800 632.5200 1379.6800 633.0000 ;
        RECT 1376.6800 637.9600 1379.6800 638.4400 ;
        RECT 1376.6800 621.6400 1379.6800 622.1200 ;
        RECT 1376.6800 616.2000 1379.6800 616.6800 ;
        RECT 1376.6800 627.0800 1379.6800 627.5600 ;
        RECT 1376.6800 605.3200 1379.6800 605.8000 ;
        RECT 1376.6800 610.7600 1379.6800 611.2400 ;
        RECT 1376.6800 594.4400 1379.6800 594.9200 ;
        RECT 1376.6800 589.0000 1379.6800 589.4800 ;
        RECT 1376.6800 599.8800 1379.6800 600.3600 ;
        RECT 1471.2400 578.1200 1472.8400 578.6000 ;
        RECT 1471.2400 583.5600 1472.8400 584.0400 ;
        RECT 1471.2400 561.8000 1472.8400 562.2800 ;
        RECT 1471.2400 567.2400 1472.8400 567.7200 ;
        RECT 1471.2400 572.6800 1472.8400 573.1600 ;
        RECT 1426.2400 578.1200 1427.8400 578.6000 ;
        RECT 1426.2400 583.5600 1427.8400 584.0400 ;
        RECT 1426.2400 561.8000 1427.8400 562.2800 ;
        RECT 1426.2400 567.2400 1427.8400 567.7200 ;
        RECT 1426.2400 572.6800 1427.8400 573.1600 ;
        RECT 1471.2400 556.3600 1472.8400 556.8400 ;
        RECT 1471.2400 550.9200 1472.8400 551.4000 ;
        RECT 1471.2400 545.4800 1472.8400 545.9600 ;
        RECT 1426.2400 556.3600 1427.8400 556.8400 ;
        RECT 1426.2400 550.9200 1427.8400 551.4000 ;
        RECT 1426.2400 545.4800 1427.8400 545.9600 ;
        RECT 1376.6800 578.1200 1379.6800 578.6000 ;
        RECT 1376.6800 583.5600 1379.6800 584.0400 ;
        RECT 1376.6800 567.2400 1379.6800 567.7200 ;
        RECT 1376.6800 561.8000 1379.6800 562.2800 ;
        RECT 1376.6800 572.6800 1379.6800 573.1600 ;
        RECT 1376.6800 550.9200 1379.6800 551.4000 ;
        RECT 1376.6800 556.3600 1379.6800 556.8400 ;
        RECT 1376.6800 545.4800 1379.6800 545.9600 ;
        RECT 1376.6800 743.6700 1575.7800 746.6700 ;
        RECT 1376.6800 538.5700 1575.7800 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 308.9300 1562.8400 517.0300 ;
        RECT 1516.2400 308.9300 1517.8400 517.0300 ;
        RECT 1471.2400 308.9300 1472.8400 517.0300 ;
        RECT 1426.2400 308.9300 1427.8400 517.0300 ;
        RECT 1572.7800 308.9300 1575.7800 517.0300 ;
        RECT 1376.6800 308.9300 1379.6800 517.0300 ;
      LAYER met3 ;
        RECT 1572.7800 511.6800 1575.7800 512.1600 ;
        RECT 1561.2400 511.6800 1562.8400 512.1600 ;
        RECT 1572.7800 500.8000 1575.7800 501.2800 ;
        RECT 1572.7800 506.2400 1575.7800 506.7200 ;
        RECT 1561.2400 500.8000 1562.8400 501.2800 ;
        RECT 1561.2400 506.2400 1562.8400 506.7200 ;
        RECT 1572.7800 484.4800 1575.7800 484.9600 ;
        RECT 1572.7800 489.9200 1575.7800 490.4000 ;
        RECT 1561.2400 484.4800 1562.8400 484.9600 ;
        RECT 1561.2400 489.9200 1562.8400 490.4000 ;
        RECT 1572.7800 473.6000 1575.7800 474.0800 ;
        RECT 1572.7800 479.0400 1575.7800 479.5200 ;
        RECT 1561.2400 473.6000 1562.8400 474.0800 ;
        RECT 1561.2400 479.0400 1562.8400 479.5200 ;
        RECT 1572.7800 495.3600 1575.7800 495.8400 ;
        RECT 1561.2400 495.3600 1562.8400 495.8400 ;
        RECT 1516.2400 500.8000 1517.8400 501.2800 ;
        RECT 1516.2400 506.2400 1517.8400 506.7200 ;
        RECT 1516.2400 511.6800 1517.8400 512.1600 ;
        RECT 1516.2400 484.4800 1517.8400 484.9600 ;
        RECT 1516.2400 489.9200 1517.8400 490.4000 ;
        RECT 1516.2400 479.0400 1517.8400 479.5200 ;
        RECT 1516.2400 473.6000 1517.8400 474.0800 ;
        RECT 1516.2400 495.3600 1517.8400 495.8400 ;
        RECT 1572.7800 457.2800 1575.7800 457.7600 ;
        RECT 1572.7800 462.7200 1575.7800 463.2000 ;
        RECT 1561.2400 457.2800 1562.8400 457.7600 ;
        RECT 1561.2400 462.7200 1562.8400 463.2000 ;
        RECT 1572.7800 440.9600 1575.7800 441.4400 ;
        RECT 1572.7800 446.4000 1575.7800 446.8800 ;
        RECT 1572.7800 451.8400 1575.7800 452.3200 ;
        RECT 1561.2400 440.9600 1562.8400 441.4400 ;
        RECT 1561.2400 446.4000 1562.8400 446.8800 ;
        RECT 1561.2400 451.8400 1562.8400 452.3200 ;
        RECT 1572.7800 430.0800 1575.7800 430.5600 ;
        RECT 1572.7800 435.5200 1575.7800 436.0000 ;
        RECT 1561.2400 430.0800 1562.8400 430.5600 ;
        RECT 1561.2400 435.5200 1562.8400 436.0000 ;
        RECT 1572.7800 413.7600 1575.7800 414.2400 ;
        RECT 1572.7800 419.2000 1575.7800 419.6800 ;
        RECT 1572.7800 424.6400 1575.7800 425.1200 ;
        RECT 1561.2400 413.7600 1562.8400 414.2400 ;
        RECT 1561.2400 419.2000 1562.8400 419.6800 ;
        RECT 1561.2400 424.6400 1562.8400 425.1200 ;
        RECT 1516.2400 457.2800 1517.8400 457.7600 ;
        RECT 1516.2400 462.7200 1517.8400 463.2000 ;
        RECT 1516.2400 440.9600 1517.8400 441.4400 ;
        RECT 1516.2400 446.4000 1517.8400 446.8800 ;
        RECT 1516.2400 451.8400 1517.8400 452.3200 ;
        RECT 1516.2400 430.0800 1517.8400 430.5600 ;
        RECT 1516.2400 435.5200 1517.8400 436.0000 ;
        RECT 1516.2400 413.7600 1517.8400 414.2400 ;
        RECT 1516.2400 419.2000 1517.8400 419.6800 ;
        RECT 1516.2400 424.6400 1517.8400 425.1200 ;
        RECT 1572.7800 468.1600 1575.7800 468.6400 ;
        RECT 1516.2400 468.1600 1517.8400 468.6400 ;
        RECT 1561.2400 468.1600 1562.8400 468.6400 ;
        RECT 1471.2400 500.8000 1472.8400 501.2800 ;
        RECT 1471.2400 506.2400 1472.8400 506.7200 ;
        RECT 1471.2400 511.6800 1472.8400 512.1600 ;
        RECT 1426.2400 500.8000 1427.8400 501.2800 ;
        RECT 1426.2400 506.2400 1427.8400 506.7200 ;
        RECT 1426.2400 511.6800 1427.8400 512.1600 ;
        RECT 1471.2400 484.4800 1472.8400 484.9600 ;
        RECT 1471.2400 489.9200 1472.8400 490.4000 ;
        RECT 1471.2400 473.6000 1472.8400 474.0800 ;
        RECT 1471.2400 479.0400 1472.8400 479.5200 ;
        RECT 1426.2400 484.4800 1427.8400 484.9600 ;
        RECT 1426.2400 489.9200 1427.8400 490.4000 ;
        RECT 1426.2400 473.6000 1427.8400 474.0800 ;
        RECT 1426.2400 479.0400 1427.8400 479.5200 ;
        RECT 1426.2400 495.3600 1427.8400 495.8400 ;
        RECT 1471.2400 495.3600 1472.8400 495.8400 ;
        RECT 1376.6800 511.6800 1379.6800 512.1600 ;
        RECT 1376.6800 506.2400 1379.6800 506.7200 ;
        RECT 1376.6800 500.8000 1379.6800 501.2800 ;
        RECT 1376.6800 489.9200 1379.6800 490.4000 ;
        RECT 1376.6800 484.4800 1379.6800 484.9600 ;
        RECT 1376.6800 479.0400 1379.6800 479.5200 ;
        RECT 1376.6800 473.6000 1379.6800 474.0800 ;
        RECT 1376.6800 495.3600 1379.6800 495.8400 ;
        RECT 1471.2400 457.2800 1472.8400 457.7600 ;
        RECT 1471.2400 462.7200 1472.8400 463.2000 ;
        RECT 1471.2400 440.9600 1472.8400 441.4400 ;
        RECT 1471.2400 446.4000 1472.8400 446.8800 ;
        RECT 1471.2400 451.8400 1472.8400 452.3200 ;
        RECT 1426.2400 457.2800 1427.8400 457.7600 ;
        RECT 1426.2400 462.7200 1427.8400 463.2000 ;
        RECT 1426.2400 440.9600 1427.8400 441.4400 ;
        RECT 1426.2400 446.4000 1427.8400 446.8800 ;
        RECT 1426.2400 451.8400 1427.8400 452.3200 ;
        RECT 1471.2400 430.0800 1472.8400 430.5600 ;
        RECT 1471.2400 435.5200 1472.8400 436.0000 ;
        RECT 1471.2400 413.7600 1472.8400 414.2400 ;
        RECT 1471.2400 419.2000 1472.8400 419.6800 ;
        RECT 1471.2400 424.6400 1472.8400 425.1200 ;
        RECT 1426.2400 430.0800 1427.8400 430.5600 ;
        RECT 1426.2400 435.5200 1427.8400 436.0000 ;
        RECT 1426.2400 413.7600 1427.8400 414.2400 ;
        RECT 1426.2400 419.2000 1427.8400 419.6800 ;
        RECT 1426.2400 424.6400 1427.8400 425.1200 ;
        RECT 1376.6800 457.2800 1379.6800 457.7600 ;
        RECT 1376.6800 462.7200 1379.6800 463.2000 ;
        RECT 1376.6800 446.4000 1379.6800 446.8800 ;
        RECT 1376.6800 440.9600 1379.6800 441.4400 ;
        RECT 1376.6800 451.8400 1379.6800 452.3200 ;
        RECT 1376.6800 430.0800 1379.6800 430.5600 ;
        RECT 1376.6800 435.5200 1379.6800 436.0000 ;
        RECT 1376.6800 419.2000 1379.6800 419.6800 ;
        RECT 1376.6800 413.7600 1379.6800 414.2400 ;
        RECT 1376.6800 424.6400 1379.6800 425.1200 ;
        RECT 1376.6800 468.1600 1379.6800 468.6400 ;
        RECT 1426.2400 468.1600 1427.8400 468.6400 ;
        RECT 1471.2400 468.1600 1472.8400 468.6400 ;
        RECT 1572.7800 402.8800 1575.7800 403.3600 ;
        RECT 1572.7800 408.3200 1575.7800 408.8000 ;
        RECT 1561.2400 402.8800 1562.8400 403.3600 ;
        RECT 1561.2400 408.3200 1562.8400 408.8000 ;
        RECT 1572.7800 386.5600 1575.7800 387.0400 ;
        RECT 1572.7800 392.0000 1575.7800 392.4800 ;
        RECT 1572.7800 397.4400 1575.7800 397.9200 ;
        RECT 1561.2400 386.5600 1562.8400 387.0400 ;
        RECT 1561.2400 392.0000 1562.8400 392.4800 ;
        RECT 1561.2400 397.4400 1562.8400 397.9200 ;
        RECT 1572.7800 375.6800 1575.7800 376.1600 ;
        RECT 1572.7800 381.1200 1575.7800 381.6000 ;
        RECT 1561.2400 375.6800 1562.8400 376.1600 ;
        RECT 1561.2400 381.1200 1562.8400 381.6000 ;
        RECT 1572.7800 359.3600 1575.7800 359.8400 ;
        RECT 1572.7800 364.8000 1575.7800 365.2800 ;
        RECT 1572.7800 370.2400 1575.7800 370.7200 ;
        RECT 1561.2400 359.3600 1562.8400 359.8400 ;
        RECT 1561.2400 364.8000 1562.8400 365.2800 ;
        RECT 1561.2400 370.2400 1562.8400 370.7200 ;
        RECT 1516.2400 402.8800 1517.8400 403.3600 ;
        RECT 1516.2400 408.3200 1517.8400 408.8000 ;
        RECT 1516.2400 386.5600 1517.8400 387.0400 ;
        RECT 1516.2400 392.0000 1517.8400 392.4800 ;
        RECT 1516.2400 397.4400 1517.8400 397.9200 ;
        RECT 1516.2400 375.6800 1517.8400 376.1600 ;
        RECT 1516.2400 381.1200 1517.8400 381.6000 ;
        RECT 1516.2400 359.3600 1517.8400 359.8400 ;
        RECT 1516.2400 364.8000 1517.8400 365.2800 ;
        RECT 1516.2400 370.2400 1517.8400 370.7200 ;
        RECT 1572.7800 348.4800 1575.7800 348.9600 ;
        RECT 1572.7800 353.9200 1575.7800 354.4000 ;
        RECT 1561.2400 348.4800 1562.8400 348.9600 ;
        RECT 1561.2400 353.9200 1562.8400 354.4000 ;
        RECT 1572.7800 332.1600 1575.7800 332.6400 ;
        RECT 1572.7800 337.6000 1575.7800 338.0800 ;
        RECT 1572.7800 343.0400 1575.7800 343.5200 ;
        RECT 1561.2400 332.1600 1562.8400 332.6400 ;
        RECT 1561.2400 337.6000 1562.8400 338.0800 ;
        RECT 1561.2400 343.0400 1562.8400 343.5200 ;
        RECT 1572.7800 321.2800 1575.7800 321.7600 ;
        RECT 1572.7800 326.7200 1575.7800 327.2000 ;
        RECT 1561.2400 321.2800 1562.8400 321.7600 ;
        RECT 1561.2400 326.7200 1562.8400 327.2000 ;
        RECT 1572.7800 315.8400 1575.7800 316.3200 ;
        RECT 1561.2400 315.8400 1562.8400 316.3200 ;
        RECT 1516.2400 348.4800 1517.8400 348.9600 ;
        RECT 1516.2400 353.9200 1517.8400 354.4000 ;
        RECT 1516.2400 332.1600 1517.8400 332.6400 ;
        RECT 1516.2400 337.6000 1517.8400 338.0800 ;
        RECT 1516.2400 343.0400 1517.8400 343.5200 ;
        RECT 1516.2400 321.2800 1517.8400 321.7600 ;
        RECT 1516.2400 326.7200 1517.8400 327.2000 ;
        RECT 1516.2400 315.8400 1517.8400 316.3200 ;
        RECT 1471.2400 402.8800 1472.8400 403.3600 ;
        RECT 1471.2400 408.3200 1472.8400 408.8000 ;
        RECT 1471.2400 386.5600 1472.8400 387.0400 ;
        RECT 1471.2400 392.0000 1472.8400 392.4800 ;
        RECT 1471.2400 397.4400 1472.8400 397.9200 ;
        RECT 1426.2400 402.8800 1427.8400 403.3600 ;
        RECT 1426.2400 408.3200 1427.8400 408.8000 ;
        RECT 1426.2400 386.5600 1427.8400 387.0400 ;
        RECT 1426.2400 392.0000 1427.8400 392.4800 ;
        RECT 1426.2400 397.4400 1427.8400 397.9200 ;
        RECT 1471.2400 375.6800 1472.8400 376.1600 ;
        RECT 1471.2400 381.1200 1472.8400 381.6000 ;
        RECT 1471.2400 359.3600 1472.8400 359.8400 ;
        RECT 1471.2400 364.8000 1472.8400 365.2800 ;
        RECT 1471.2400 370.2400 1472.8400 370.7200 ;
        RECT 1426.2400 375.6800 1427.8400 376.1600 ;
        RECT 1426.2400 381.1200 1427.8400 381.6000 ;
        RECT 1426.2400 359.3600 1427.8400 359.8400 ;
        RECT 1426.2400 364.8000 1427.8400 365.2800 ;
        RECT 1426.2400 370.2400 1427.8400 370.7200 ;
        RECT 1376.6800 402.8800 1379.6800 403.3600 ;
        RECT 1376.6800 408.3200 1379.6800 408.8000 ;
        RECT 1376.6800 392.0000 1379.6800 392.4800 ;
        RECT 1376.6800 386.5600 1379.6800 387.0400 ;
        RECT 1376.6800 397.4400 1379.6800 397.9200 ;
        RECT 1376.6800 375.6800 1379.6800 376.1600 ;
        RECT 1376.6800 381.1200 1379.6800 381.6000 ;
        RECT 1376.6800 364.8000 1379.6800 365.2800 ;
        RECT 1376.6800 359.3600 1379.6800 359.8400 ;
        RECT 1376.6800 370.2400 1379.6800 370.7200 ;
        RECT 1471.2400 348.4800 1472.8400 348.9600 ;
        RECT 1471.2400 353.9200 1472.8400 354.4000 ;
        RECT 1471.2400 332.1600 1472.8400 332.6400 ;
        RECT 1471.2400 337.6000 1472.8400 338.0800 ;
        RECT 1471.2400 343.0400 1472.8400 343.5200 ;
        RECT 1426.2400 348.4800 1427.8400 348.9600 ;
        RECT 1426.2400 353.9200 1427.8400 354.4000 ;
        RECT 1426.2400 332.1600 1427.8400 332.6400 ;
        RECT 1426.2400 337.6000 1427.8400 338.0800 ;
        RECT 1426.2400 343.0400 1427.8400 343.5200 ;
        RECT 1471.2400 326.7200 1472.8400 327.2000 ;
        RECT 1471.2400 321.2800 1472.8400 321.7600 ;
        RECT 1471.2400 315.8400 1472.8400 316.3200 ;
        RECT 1426.2400 326.7200 1427.8400 327.2000 ;
        RECT 1426.2400 321.2800 1427.8400 321.7600 ;
        RECT 1426.2400 315.8400 1427.8400 316.3200 ;
        RECT 1376.6800 348.4800 1379.6800 348.9600 ;
        RECT 1376.6800 353.9200 1379.6800 354.4000 ;
        RECT 1376.6800 337.6000 1379.6800 338.0800 ;
        RECT 1376.6800 332.1600 1379.6800 332.6400 ;
        RECT 1376.6800 343.0400 1379.6800 343.5200 ;
        RECT 1376.6800 321.2800 1379.6800 321.7600 ;
        RECT 1376.6800 326.7200 1379.6800 327.2000 ;
        RECT 1376.6800 315.8400 1379.6800 316.3200 ;
        RECT 1376.6800 514.0300 1575.7800 517.0300 ;
        RECT 1376.6800 308.9300 1575.7800 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 79.2900 1562.8400 287.3900 ;
        RECT 1516.2400 79.2900 1517.8400 287.3900 ;
        RECT 1471.2400 79.2900 1472.8400 287.3900 ;
        RECT 1426.2400 79.2900 1427.8400 287.3900 ;
        RECT 1572.7800 79.2900 1575.7800 287.3900 ;
        RECT 1376.6800 79.2900 1379.6800 287.3900 ;
      LAYER met3 ;
        RECT 1572.7800 282.0400 1575.7800 282.5200 ;
        RECT 1561.2400 282.0400 1562.8400 282.5200 ;
        RECT 1572.7800 271.1600 1575.7800 271.6400 ;
        RECT 1572.7800 276.6000 1575.7800 277.0800 ;
        RECT 1561.2400 271.1600 1562.8400 271.6400 ;
        RECT 1561.2400 276.6000 1562.8400 277.0800 ;
        RECT 1572.7800 254.8400 1575.7800 255.3200 ;
        RECT 1572.7800 260.2800 1575.7800 260.7600 ;
        RECT 1561.2400 254.8400 1562.8400 255.3200 ;
        RECT 1561.2400 260.2800 1562.8400 260.7600 ;
        RECT 1572.7800 243.9600 1575.7800 244.4400 ;
        RECT 1572.7800 249.4000 1575.7800 249.8800 ;
        RECT 1561.2400 243.9600 1562.8400 244.4400 ;
        RECT 1561.2400 249.4000 1562.8400 249.8800 ;
        RECT 1572.7800 265.7200 1575.7800 266.2000 ;
        RECT 1561.2400 265.7200 1562.8400 266.2000 ;
        RECT 1516.2400 271.1600 1517.8400 271.6400 ;
        RECT 1516.2400 276.6000 1517.8400 277.0800 ;
        RECT 1516.2400 282.0400 1517.8400 282.5200 ;
        RECT 1516.2400 254.8400 1517.8400 255.3200 ;
        RECT 1516.2400 260.2800 1517.8400 260.7600 ;
        RECT 1516.2400 249.4000 1517.8400 249.8800 ;
        RECT 1516.2400 243.9600 1517.8400 244.4400 ;
        RECT 1516.2400 265.7200 1517.8400 266.2000 ;
        RECT 1572.7800 227.6400 1575.7800 228.1200 ;
        RECT 1572.7800 233.0800 1575.7800 233.5600 ;
        RECT 1561.2400 227.6400 1562.8400 228.1200 ;
        RECT 1561.2400 233.0800 1562.8400 233.5600 ;
        RECT 1572.7800 211.3200 1575.7800 211.8000 ;
        RECT 1572.7800 216.7600 1575.7800 217.2400 ;
        RECT 1572.7800 222.2000 1575.7800 222.6800 ;
        RECT 1561.2400 211.3200 1562.8400 211.8000 ;
        RECT 1561.2400 216.7600 1562.8400 217.2400 ;
        RECT 1561.2400 222.2000 1562.8400 222.6800 ;
        RECT 1572.7800 200.4400 1575.7800 200.9200 ;
        RECT 1572.7800 205.8800 1575.7800 206.3600 ;
        RECT 1561.2400 200.4400 1562.8400 200.9200 ;
        RECT 1561.2400 205.8800 1562.8400 206.3600 ;
        RECT 1572.7800 184.1200 1575.7800 184.6000 ;
        RECT 1572.7800 189.5600 1575.7800 190.0400 ;
        RECT 1572.7800 195.0000 1575.7800 195.4800 ;
        RECT 1561.2400 184.1200 1562.8400 184.6000 ;
        RECT 1561.2400 189.5600 1562.8400 190.0400 ;
        RECT 1561.2400 195.0000 1562.8400 195.4800 ;
        RECT 1516.2400 227.6400 1517.8400 228.1200 ;
        RECT 1516.2400 233.0800 1517.8400 233.5600 ;
        RECT 1516.2400 211.3200 1517.8400 211.8000 ;
        RECT 1516.2400 216.7600 1517.8400 217.2400 ;
        RECT 1516.2400 222.2000 1517.8400 222.6800 ;
        RECT 1516.2400 200.4400 1517.8400 200.9200 ;
        RECT 1516.2400 205.8800 1517.8400 206.3600 ;
        RECT 1516.2400 184.1200 1517.8400 184.6000 ;
        RECT 1516.2400 189.5600 1517.8400 190.0400 ;
        RECT 1516.2400 195.0000 1517.8400 195.4800 ;
        RECT 1572.7800 238.5200 1575.7800 239.0000 ;
        RECT 1516.2400 238.5200 1517.8400 239.0000 ;
        RECT 1561.2400 238.5200 1562.8400 239.0000 ;
        RECT 1471.2400 271.1600 1472.8400 271.6400 ;
        RECT 1471.2400 276.6000 1472.8400 277.0800 ;
        RECT 1471.2400 282.0400 1472.8400 282.5200 ;
        RECT 1426.2400 271.1600 1427.8400 271.6400 ;
        RECT 1426.2400 276.6000 1427.8400 277.0800 ;
        RECT 1426.2400 282.0400 1427.8400 282.5200 ;
        RECT 1471.2400 254.8400 1472.8400 255.3200 ;
        RECT 1471.2400 260.2800 1472.8400 260.7600 ;
        RECT 1471.2400 243.9600 1472.8400 244.4400 ;
        RECT 1471.2400 249.4000 1472.8400 249.8800 ;
        RECT 1426.2400 254.8400 1427.8400 255.3200 ;
        RECT 1426.2400 260.2800 1427.8400 260.7600 ;
        RECT 1426.2400 243.9600 1427.8400 244.4400 ;
        RECT 1426.2400 249.4000 1427.8400 249.8800 ;
        RECT 1426.2400 265.7200 1427.8400 266.2000 ;
        RECT 1471.2400 265.7200 1472.8400 266.2000 ;
        RECT 1376.6800 282.0400 1379.6800 282.5200 ;
        RECT 1376.6800 276.6000 1379.6800 277.0800 ;
        RECT 1376.6800 271.1600 1379.6800 271.6400 ;
        RECT 1376.6800 260.2800 1379.6800 260.7600 ;
        RECT 1376.6800 254.8400 1379.6800 255.3200 ;
        RECT 1376.6800 249.4000 1379.6800 249.8800 ;
        RECT 1376.6800 243.9600 1379.6800 244.4400 ;
        RECT 1376.6800 265.7200 1379.6800 266.2000 ;
        RECT 1471.2400 227.6400 1472.8400 228.1200 ;
        RECT 1471.2400 233.0800 1472.8400 233.5600 ;
        RECT 1471.2400 211.3200 1472.8400 211.8000 ;
        RECT 1471.2400 216.7600 1472.8400 217.2400 ;
        RECT 1471.2400 222.2000 1472.8400 222.6800 ;
        RECT 1426.2400 227.6400 1427.8400 228.1200 ;
        RECT 1426.2400 233.0800 1427.8400 233.5600 ;
        RECT 1426.2400 211.3200 1427.8400 211.8000 ;
        RECT 1426.2400 216.7600 1427.8400 217.2400 ;
        RECT 1426.2400 222.2000 1427.8400 222.6800 ;
        RECT 1471.2400 200.4400 1472.8400 200.9200 ;
        RECT 1471.2400 205.8800 1472.8400 206.3600 ;
        RECT 1471.2400 184.1200 1472.8400 184.6000 ;
        RECT 1471.2400 189.5600 1472.8400 190.0400 ;
        RECT 1471.2400 195.0000 1472.8400 195.4800 ;
        RECT 1426.2400 200.4400 1427.8400 200.9200 ;
        RECT 1426.2400 205.8800 1427.8400 206.3600 ;
        RECT 1426.2400 184.1200 1427.8400 184.6000 ;
        RECT 1426.2400 189.5600 1427.8400 190.0400 ;
        RECT 1426.2400 195.0000 1427.8400 195.4800 ;
        RECT 1376.6800 227.6400 1379.6800 228.1200 ;
        RECT 1376.6800 233.0800 1379.6800 233.5600 ;
        RECT 1376.6800 216.7600 1379.6800 217.2400 ;
        RECT 1376.6800 211.3200 1379.6800 211.8000 ;
        RECT 1376.6800 222.2000 1379.6800 222.6800 ;
        RECT 1376.6800 200.4400 1379.6800 200.9200 ;
        RECT 1376.6800 205.8800 1379.6800 206.3600 ;
        RECT 1376.6800 189.5600 1379.6800 190.0400 ;
        RECT 1376.6800 184.1200 1379.6800 184.6000 ;
        RECT 1376.6800 195.0000 1379.6800 195.4800 ;
        RECT 1376.6800 238.5200 1379.6800 239.0000 ;
        RECT 1426.2400 238.5200 1427.8400 239.0000 ;
        RECT 1471.2400 238.5200 1472.8400 239.0000 ;
        RECT 1572.7800 173.2400 1575.7800 173.7200 ;
        RECT 1572.7800 178.6800 1575.7800 179.1600 ;
        RECT 1561.2400 173.2400 1562.8400 173.7200 ;
        RECT 1561.2400 178.6800 1562.8400 179.1600 ;
        RECT 1572.7800 156.9200 1575.7800 157.4000 ;
        RECT 1572.7800 162.3600 1575.7800 162.8400 ;
        RECT 1572.7800 167.8000 1575.7800 168.2800 ;
        RECT 1561.2400 156.9200 1562.8400 157.4000 ;
        RECT 1561.2400 162.3600 1562.8400 162.8400 ;
        RECT 1561.2400 167.8000 1562.8400 168.2800 ;
        RECT 1572.7800 146.0400 1575.7800 146.5200 ;
        RECT 1572.7800 151.4800 1575.7800 151.9600 ;
        RECT 1561.2400 146.0400 1562.8400 146.5200 ;
        RECT 1561.2400 151.4800 1562.8400 151.9600 ;
        RECT 1572.7800 129.7200 1575.7800 130.2000 ;
        RECT 1572.7800 135.1600 1575.7800 135.6400 ;
        RECT 1572.7800 140.6000 1575.7800 141.0800 ;
        RECT 1561.2400 129.7200 1562.8400 130.2000 ;
        RECT 1561.2400 135.1600 1562.8400 135.6400 ;
        RECT 1561.2400 140.6000 1562.8400 141.0800 ;
        RECT 1516.2400 173.2400 1517.8400 173.7200 ;
        RECT 1516.2400 178.6800 1517.8400 179.1600 ;
        RECT 1516.2400 156.9200 1517.8400 157.4000 ;
        RECT 1516.2400 162.3600 1517.8400 162.8400 ;
        RECT 1516.2400 167.8000 1517.8400 168.2800 ;
        RECT 1516.2400 146.0400 1517.8400 146.5200 ;
        RECT 1516.2400 151.4800 1517.8400 151.9600 ;
        RECT 1516.2400 129.7200 1517.8400 130.2000 ;
        RECT 1516.2400 135.1600 1517.8400 135.6400 ;
        RECT 1516.2400 140.6000 1517.8400 141.0800 ;
        RECT 1572.7800 118.8400 1575.7800 119.3200 ;
        RECT 1572.7800 124.2800 1575.7800 124.7600 ;
        RECT 1561.2400 118.8400 1562.8400 119.3200 ;
        RECT 1561.2400 124.2800 1562.8400 124.7600 ;
        RECT 1572.7800 102.5200 1575.7800 103.0000 ;
        RECT 1572.7800 107.9600 1575.7800 108.4400 ;
        RECT 1572.7800 113.4000 1575.7800 113.8800 ;
        RECT 1561.2400 102.5200 1562.8400 103.0000 ;
        RECT 1561.2400 107.9600 1562.8400 108.4400 ;
        RECT 1561.2400 113.4000 1562.8400 113.8800 ;
        RECT 1572.7800 91.6400 1575.7800 92.1200 ;
        RECT 1572.7800 97.0800 1575.7800 97.5600 ;
        RECT 1561.2400 91.6400 1562.8400 92.1200 ;
        RECT 1561.2400 97.0800 1562.8400 97.5600 ;
        RECT 1572.7800 86.2000 1575.7800 86.6800 ;
        RECT 1561.2400 86.2000 1562.8400 86.6800 ;
        RECT 1516.2400 118.8400 1517.8400 119.3200 ;
        RECT 1516.2400 124.2800 1517.8400 124.7600 ;
        RECT 1516.2400 102.5200 1517.8400 103.0000 ;
        RECT 1516.2400 107.9600 1517.8400 108.4400 ;
        RECT 1516.2400 113.4000 1517.8400 113.8800 ;
        RECT 1516.2400 91.6400 1517.8400 92.1200 ;
        RECT 1516.2400 97.0800 1517.8400 97.5600 ;
        RECT 1516.2400 86.2000 1517.8400 86.6800 ;
        RECT 1471.2400 173.2400 1472.8400 173.7200 ;
        RECT 1471.2400 178.6800 1472.8400 179.1600 ;
        RECT 1471.2400 156.9200 1472.8400 157.4000 ;
        RECT 1471.2400 162.3600 1472.8400 162.8400 ;
        RECT 1471.2400 167.8000 1472.8400 168.2800 ;
        RECT 1426.2400 173.2400 1427.8400 173.7200 ;
        RECT 1426.2400 178.6800 1427.8400 179.1600 ;
        RECT 1426.2400 156.9200 1427.8400 157.4000 ;
        RECT 1426.2400 162.3600 1427.8400 162.8400 ;
        RECT 1426.2400 167.8000 1427.8400 168.2800 ;
        RECT 1471.2400 146.0400 1472.8400 146.5200 ;
        RECT 1471.2400 151.4800 1472.8400 151.9600 ;
        RECT 1471.2400 129.7200 1472.8400 130.2000 ;
        RECT 1471.2400 135.1600 1472.8400 135.6400 ;
        RECT 1471.2400 140.6000 1472.8400 141.0800 ;
        RECT 1426.2400 146.0400 1427.8400 146.5200 ;
        RECT 1426.2400 151.4800 1427.8400 151.9600 ;
        RECT 1426.2400 129.7200 1427.8400 130.2000 ;
        RECT 1426.2400 135.1600 1427.8400 135.6400 ;
        RECT 1426.2400 140.6000 1427.8400 141.0800 ;
        RECT 1376.6800 173.2400 1379.6800 173.7200 ;
        RECT 1376.6800 178.6800 1379.6800 179.1600 ;
        RECT 1376.6800 162.3600 1379.6800 162.8400 ;
        RECT 1376.6800 156.9200 1379.6800 157.4000 ;
        RECT 1376.6800 167.8000 1379.6800 168.2800 ;
        RECT 1376.6800 146.0400 1379.6800 146.5200 ;
        RECT 1376.6800 151.4800 1379.6800 151.9600 ;
        RECT 1376.6800 135.1600 1379.6800 135.6400 ;
        RECT 1376.6800 129.7200 1379.6800 130.2000 ;
        RECT 1376.6800 140.6000 1379.6800 141.0800 ;
        RECT 1471.2400 118.8400 1472.8400 119.3200 ;
        RECT 1471.2400 124.2800 1472.8400 124.7600 ;
        RECT 1471.2400 102.5200 1472.8400 103.0000 ;
        RECT 1471.2400 107.9600 1472.8400 108.4400 ;
        RECT 1471.2400 113.4000 1472.8400 113.8800 ;
        RECT 1426.2400 118.8400 1427.8400 119.3200 ;
        RECT 1426.2400 124.2800 1427.8400 124.7600 ;
        RECT 1426.2400 102.5200 1427.8400 103.0000 ;
        RECT 1426.2400 107.9600 1427.8400 108.4400 ;
        RECT 1426.2400 113.4000 1427.8400 113.8800 ;
        RECT 1471.2400 97.0800 1472.8400 97.5600 ;
        RECT 1471.2400 91.6400 1472.8400 92.1200 ;
        RECT 1471.2400 86.2000 1472.8400 86.6800 ;
        RECT 1426.2400 97.0800 1427.8400 97.5600 ;
        RECT 1426.2400 91.6400 1427.8400 92.1200 ;
        RECT 1426.2400 86.2000 1427.8400 86.6800 ;
        RECT 1376.6800 118.8400 1379.6800 119.3200 ;
        RECT 1376.6800 124.2800 1379.6800 124.7600 ;
        RECT 1376.6800 107.9600 1379.6800 108.4400 ;
        RECT 1376.6800 102.5200 1379.6800 103.0000 ;
        RECT 1376.6800 113.4000 1379.6800 113.8800 ;
        RECT 1376.6800 91.6400 1379.6800 92.1200 ;
        RECT 1376.6800 97.0800 1379.6800 97.5600 ;
        RECT 1376.6800 86.2000 1379.6800 86.6800 ;
        RECT 1376.6800 284.3900 1575.7800 287.3900 ;
        RECT 1376.6800 79.2900 1575.7800 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1376.6800 37.6700 1378.6800 58.6000 ;
        RECT 1573.7800 37.6700 1575.7800 58.6000 ;
      LAYER met3 ;
        RECT 1573.7800 54.1000 1575.7800 54.5800 ;
        RECT 1376.6800 54.1000 1378.6800 54.5800 ;
        RECT 1573.7800 43.2200 1575.7800 43.7000 ;
        RECT 1376.6800 43.2200 1378.6800 43.7000 ;
        RECT 1573.7800 48.6600 1575.7800 49.1400 ;
        RECT 1376.6800 48.6600 1378.6800 49.1400 ;
        RECT 1376.6800 56.6000 1575.7800 58.6000 ;
        RECT 1376.6800 37.6700 1575.7800 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 2605.3300 1562.8400 2813.4300 ;
        RECT 1516.2400 2605.3300 1517.8400 2813.4300 ;
        RECT 1471.2400 2605.3300 1472.8400 2813.4300 ;
        RECT 1426.2400 2605.3300 1427.8400 2813.4300 ;
        RECT 1572.7800 2605.3300 1575.7800 2813.4300 ;
        RECT 1376.6800 2605.3300 1379.6800 2813.4300 ;
      LAYER met3 ;
        RECT 1572.7800 2808.0800 1575.7800 2808.5600 ;
        RECT 1561.2400 2808.0800 1562.8400 2808.5600 ;
        RECT 1572.7800 2797.2000 1575.7800 2797.6800 ;
        RECT 1572.7800 2802.6400 1575.7800 2803.1200 ;
        RECT 1561.2400 2797.2000 1562.8400 2797.6800 ;
        RECT 1561.2400 2802.6400 1562.8400 2803.1200 ;
        RECT 1572.7800 2780.8800 1575.7800 2781.3600 ;
        RECT 1572.7800 2786.3200 1575.7800 2786.8000 ;
        RECT 1561.2400 2780.8800 1562.8400 2781.3600 ;
        RECT 1561.2400 2786.3200 1562.8400 2786.8000 ;
        RECT 1572.7800 2770.0000 1575.7800 2770.4800 ;
        RECT 1572.7800 2775.4400 1575.7800 2775.9200 ;
        RECT 1561.2400 2770.0000 1562.8400 2770.4800 ;
        RECT 1561.2400 2775.4400 1562.8400 2775.9200 ;
        RECT 1572.7800 2791.7600 1575.7800 2792.2400 ;
        RECT 1561.2400 2791.7600 1562.8400 2792.2400 ;
        RECT 1516.2400 2797.2000 1517.8400 2797.6800 ;
        RECT 1516.2400 2802.6400 1517.8400 2803.1200 ;
        RECT 1516.2400 2808.0800 1517.8400 2808.5600 ;
        RECT 1516.2400 2780.8800 1517.8400 2781.3600 ;
        RECT 1516.2400 2786.3200 1517.8400 2786.8000 ;
        RECT 1516.2400 2775.4400 1517.8400 2775.9200 ;
        RECT 1516.2400 2770.0000 1517.8400 2770.4800 ;
        RECT 1516.2400 2791.7600 1517.8400 2792.2400 ;
        RECT 1572.7800 2753.6800 1575.7800 2754.1600 ;
        RECT 1572.7800 2759.1200 1575.7800 2759.6000 ;
        RECT 1561.2400 2753.6800 1562.8400 2754.1600 ;
        RECT 1561.2400 2759.1200 1562.8400 2759.6000 ;
        RECT 1572.7800 2737.3600 1575.7800 2737.8400 ;
        RECT 1572.7800 2742.8000 1575.7800 2743.2800 ;
        RECT 1572.7800 2748.2400 1575.7800 2748.7200 ;
        RECT 1561.2400 2737.3600 1562.8400 2737.8400 ;
        RECT 1561.2400 2742.8000 1562.8400 2743.2800 ;
        RECT 1561.2400 2748.2400 1562.8400 2748.7200 ;
        RECT 1572.7800 2726.4800 1575.7800 2726.9600 ;
        RECT 1572.7800 2731.9200 1575.7800 2732.4000 ;
        RECT 1561.2400 2726.4800 1562.8400 2726.9600 ;
        RECT 1561.2400 2731.9200 1562.8400 2732.4000 ;
        RECT 1572.7800 2710.1600 1575.7800 2710.6400 ;
        RECT 1572.7800 2715.6000 1575.7800 2716.0800 ;
        RECT 1572.7800 2721.0400 1575.7800 2721.5200 ;
        RECT 1561.2400 2710.1600 1562.8400 2710.6400 ;
        RECT 1561.2400 2715.6000 1562.8400 2716.0800 ;
        RECT 1561.2400 2721.0400 1562.8400 2721.5200 ;
        RECT 1516.2400 2753.6800 1517.8400 2754.1600 ;
        RECT 1516.2400 2759.1200 1517.8400 2759.6000 ;
        RECT 1516.2400 2737.3600 1517.8400 2737.8400 ;
        RECT 1516.2400 2742.8000 1517.8400 2743.2800 ;
        RECT 1516.2400 2748.2400 1517.8400 2748.7200 ;
        RECT 1516.2400 2726.4800 1517.8400 2726.9600 ;
        RECT 1516.2400 2731.9200 1517.8400 2732.4000 ;
        RECT 1516.2400 2710.1600 1517.8400 2710.6400 ;
        RECT 1516.2400 2715.6000 1517.8400 2716.0800 ;
        RECT 1516.2400 2721.0400 1517.8400 2721.5200 ;
        RECT 1572.7800 2764.5600 1575.7800 2765.0400 ;
        RECT 1516.2400 2764.5600 1517.8400 2765.0400 ;
        RECT 1561.2400 2764.5600 1562.8400 2765.0400 ;
        RECT 1471.2400 2797.2000 1472.8400 2797.6800 ;
        RECT 1471.2400 2802.6400 1472.8400 2803.1200 ;
        RECT 1471.2400 2808.0800 1472.8400 2808.5600 ;
        RECT 1426.2400 2797.2000 1427.8400 2797.6800 ;
        RECT 1426.2400 2802.6400 1427.8400 2803.1200 ;
        RECT 1426.2400 2808.0800 1427.8400 2808.5600 ;
        RECT 1471.2400 2780.8800 1472.8400 2781.3600 ;
        RECT 1471.2400 2786.3200 1472.8400 2786.8000 ;
        RECT 1471.2400 2770.0000 1472.8400 2770.4800 ;
        RECT 1471.2400 2775.4400 1472.8400 2775.9200 ;
        RECT 1426.2400 2780.8800 1427.8400 2781.3600 ;
        RECT 1426.2400 2786.3200 1427.8400 2786.8000 ;
        RECT 1426.2400 2770.0000 1427.8400 2770.4800 ;
        RECT 1426.2400 2775.4400 1427.8400 2775.9200 ;
        RECT 1426.2400 2791.7600 1427.8400 2792.2400 ;
        RECT 1471.2400 2791.7600 1472.8400 2792.2400 ;
        RECT 1376.6800 2808.0800 1379.6800 2808.5600 ;
        RECT 1376.6800 2802.6400 1379.6800 2803.1200 ;
        RECT 1376.6800 2797.2000 1379.6800 2797.6800 ;
        RECT 1376.6800 2786.3200 1379.6800 2786.8000 ;
        RECT 1376.6800 2780.8800 1379.6800 2781.3600 ;
        RECT 1376.6800 2775.4400 1379.6800 2775.9200 ;
        RECT 1376.6800 2770.0000 1379.6800 2770.4800 ;
        RECT 1376.6800 2791.7600 1379.6800 2792.2400 ;
        RECT 1471.2400 2753.6800 1472.8400 2754.1600 ;
        RECT 1471.2400 2759.1200 1472.8400 2759.6000 ;
        RECT 1471.2400 2737.3600 1472.8400 2737.8400 ;
        RECT 1471.2400 2742.8000 1472.8400 2743.2800 ;
        RECT 1471.2400 2748.2400 1472.8400 2748.7200 ;
        RECT 1426.2400 2753.6800 1427.8400 2754.1600 ;
        RECT 1426.2400 2759.1200 1427.8400 2759.6000 ;
        RECT 1426.2400 2737.3600 1427.8400 2737.8400 ;
        RECT 1426.2400 2742.8000 1427.8400 2743.2800 ;
        RECT 1426.2400 2748.2400 1427.8400 2748.7200 ;
        RECT 1471.2400 2726.4800 1472.8400 2726.9600 ;
        RECT 1471.2400 2731.9200 1472.8400 2732.4000 ;
        RECT 1471.2400 2710.1600 1472.8400 2710.6400 ;
        RECT 1471.2400 2715.6000 1472.8400 2716.0800 ;
        RECT 1471.2400 2721.0400 1472.8400 2721.5200 ;
        RECT 1426.2400 2726.4800 1427.8400 2726.9600 ;
        RECT 1426.2400 2731.9200 1427.8400 2732.4000 ;
        RECT 1426.2400 2710.1600 1427.8400 2710.6400 ;
        RECT 1426.2400 2715.6000 1427.8400 2716.0800 ;
        RECT 1426.2400 2721.0400 1427.8400 2721.5200 ;
        RECT 1376.6800 2753.6800 1379.6800 2754.1600 ;
        RECT 1376.6800 2759.1200 1379.6800 2759.6000 ;
        RECT 1376.6800 2742.8000 1379.6800 2743.2800 ;
        RECT 1376.6800 2737.3600 1379.6800 2737.8400 ;
        RECT 1376.6800 2748.2400 1379.6800 2748.7200 ;
        RECT 1376.6800 2726.4800 1379.6800 2726.9600 ;
        RECT 1376.6800 2731.9200 1379.6800 2732.4000 ;
        RECT 1376.6800 2715.6000 1379.6800 2716.0800 ;
        RECT 1376.6800 2710.1600 1379.6800 2710.6400 ;
        RECT 1376.6800 2721.0400 1379.6800 2721.5200 ;
        RECT 1376.6800 2764.5600 1379.6800 2765.0400 ;
        RECT 1426.2400 2764.5600 1427.8400 2765.0400 ;
        RECT 1471.2400 2764.5600 1472.8400 2765.0400 ;
        RECT 1572.7800 2699.2800 1575.7800 2699.7600 ;
        RECT 1572.7800 2704.7200 1575.7800 2705.2000 ;
        RECT 1561.2400 2699.2800 1562.8400 2699.7600 ;
        RECT 1561.2400 2704.7200 1562.8400 2705.2000 ;
        RECT 1572.7800 2682.9600 1575.7800 2683.4400 ;
        RECT 1572.7800 2688.4000 1575.7800 2688.8800 ;
        RECT 1572.7800 2693.8400 1575.7800 2694.3200 ;
        RECT 1561.2400 2682.9600 1562.8400 2683.4400 ;
        RECT 1561.2400 2688.4000 1562.8400 2688.8800 ;
        RECT 1561.2400 2693.8400 1562.8400 2694.3200 ;
        RECT 1572.7800 2672.0800 1575.7800 2672.5600 ;
        RECT 1572.7800 2677.5200 1575.7800 2678.0000 ;
        RECT 1561.2400 2672.0800 1562.8400 2672.5600 ;
        RECT 1561.2400 2677.5200 1562.8400 2678.0000 ;
        RECT 1572.7800 2655.7600 1575.7800 2656.2400 ;
        RECT 1572.7800 2661.2000 1575.7800 2661.6800 ;
        RECT 1572.7800 2666.6400 1575.7800 2667.1200 ;
        RECT 1561.2400 2655.7600 1562.8400 2656.2400 ;
        RECT 1561.2400 2661.2000 1562.8400 2661.6800 ;
        RECT 1561.2400 2666.6400 1562.8400 2667.1200 ;
        RECT 1516.2400 2699.2800 1517.8400 2699.7600 ;
        RECT 1516.2400 2704.7200 1517.8400 2705.2000 ;
        RECT 1516.2400 2682.9600 1517.8400 2683.4400 ;
        RECT 1516.2400 2688.4000 1517.8400 2688.8800 ;
        RECT 1516.2400 2693.8400 1517.8400 2694.3200 ;
        RECT 1516.2400 2672.0800 1517.8400 2672.5600 ;
        RECT 1516.2400 2677.5200 1517.8400 2678.0000 ;
        RECT 1516.2400 2655.7600 1517.8400 2656.2400 ;
        RECT 1516.2400 2661.2000 1517.8400 2661.6800 ;
        RECT 1516.2400 2666.6400 1517.8400 2667.1200 ;
        RECT 1572.7800 2644.8800 1575.7800 2645.3600 ;
        RECT 1572.7800 2650.3200 1575.7800 2650.8000 ;
        RECT 1561.2400 2644.8800 1562.8400 2645.3600 ;
        RECT 1561.2400 2650.3200 1562.8400 2650.8000 ;
        RECT 1572.7800 2628.5600 1575.7800 2629.0400 ;
        RECT 1572.7800 2634.0000 1575.7800 2634.4800 ;
        RECT 1572.7800 2639.4400 1575.7800 2639.9200 ;
        RECT 1561.2400 2628.5600 1562.8400 2629.0400 ;
        RECT 1561.2400 2634.0000 1562.8400 2634.4800 ;
        RECT 1561.2400 2639.4400 1562.8400 2639.9200 ;
        RECT 1572.7800 2617.6800 1575.7800 2618.1600 ;
        RECT 1572.7800 2623.1200 1575.7800 2623.6000 ;
        RECT 1561.2400 2617.6800 1562.8400 2618.1600 ;
        RECT 1561.2400 2623.1200 1562.8400 2623.6000 ;
        RECT 1572.7800 2612.2400 1575.7800 2612.7200 ;
        RECT 1561.2400 2612.2400 1562.8400 2612.7200 ;
        RECT 1516.2400 2644.8800 1517.8400 2645.3600 ;
        RECT 1516.2400 2650.3200 1517.8400 2650.8000 ;
        RECT 1516.2400 2628.5600 1517.8400 2629.0400 ;
        RECT 1516.2400 2634.0000 1517.8400 2634.4800 ;
        RECT 1516.2400 2639.4400 1517.8400 2639.9200 ;
        RECT 1516.2400 2617.6800 1517.8400 2618.1600 ;
        RECT 1516.2400 2623.1200 1517.8400 2623.6000 ;
        RECT 1516.2400 2612.2400 1517.8400 2612.7200 ;
        RECT 1471.2400 2699.2800 1472.8400 2699.7600 ;
        RECT 1471.2400 2704.7200 1472.8400 2705.2000 ;
        RECT 1471.2400 2682.9600 1472.8400 2683.4400 ;
        RECT 1471.2400 2688.4000 1472.8400 2688.8800 ;
        RECT 1471.2400 2693.8400 1472.8400 2694.3200 ;
        RECT 1426.2400 2699.2800 1427.8400 2699.7600 ;
        RECT 1426.2400 2704.7200 1427.8400 2705.2000 ;
        RECT 1426.2400 2682.9600 1427.8400 2683.4400 ;
        RECT 1426.2400 2688.4000 1427.8400 2688.8800 ;
        RECT 1426.2400 2693.8400 1427.8400 2694.3200 ;
        RECT 1471.2400 2672.0800 1472.8400 2672.5600 ;
        RECT 1471.2400 2677.5200 1472.8400 2678.0000 ;
        RECT 1471.2400 2655.7600 1472.8400 2656.2400 ;
        RECT 1471.2400 2661.2000 1472.8400 2661.6800 ;
        RECT 1471.2400 2666.6400 1472.8400 2667.1200 ;
        RECT 1426.2400 2672.0800 1427.8400 2672.5600 ;
        RECT 1426.2400 2677.5200 1427.8400 2678.0000 ;
        RECT 1426.2400 2655.7600 1427.8400 2656.2400 ;
        RECT 1426.2400 2661.2000 1427.8400 2661.6800 ;
        RECT 1426.2400 2666.6400 1427.8400 2667.1200 ;
        RECT 1376.6800 2699.2800 1379.6800 2699.7600 ;
        RECT 1376.6800 2704.7200 1379.6800 2705.2000 ;
        RECT 1376.6800 2688.4000 1379.6800 2688.8800 ;
        RECT 1376.6800 2682.9600 1379.6800 2683.4400 ;
        RECT 1376.6800 2693.8400 1379.6800 2694.3200 ;
        RECT 1376.6800 2672.0800 1379.6800 2672.5600 ;
        RECT 1376.6800 2677.5200 1379.6800 2678.0000 ;
        RECT 1376.6800 2661.2000 1379.6800 2661.6800 ;
        RECT 1376.6800 2655.7600 1379.6800 2656.2400 ;
        RECT 1376.6800 2666.6400 1379.6800 2667.1200 ;
        RECT 1471.2400 2644.8800 1472.8400 2645.3600 ;
        RECT 1471.2400 2650.3200 1472.8400 2650.8000 ;
        RECT 1471.2400 2628.5600 1472.8400 2629.0400 ;
        RECT 1471.2400 2634.0000 1472.8400 2634.4800 ;
        RECT 1471.2400 2639.4400 1472.8400 2639.9200 ;
        RECT 1426.2400 2644.8800 1427.8400 2645.3600 ;
        RECT 1426.2400 2650.3200 1427.8400 2650.8000 ;
        RECT 1426.2400 2628.5600 1427.8400 2629.0400 ;
        RECT 1426.2400 2634.0000 1427.8400 2634.4800 ;
        RECT 1426.2400 2639.4400 1427.8400 2639.9200 ;
        RECT 1471.2400 2623.1200 1472.8400 2623.6000 ;
        RECT 1471.2400 2617.6800 1472.8400 2618.1600 ;
        RECT 1471.2400 2612.2400 1472.8400 2612.7200 ;
        RECT 1426.2400 2623.1200 1427.8400 2623.6000 ;
        RECT 1426.2400 2617.6800 1427.8400 2618.1600 ;
        RECT 1426.2400 2612.2400 1427.8400 2612.7200 ;
        RECT 1376.6800 2644.8800 1379.6800 2645.3600 ;
        RECT 1376.6800 2650.3200 1379.6800 2650.8000 ;
        RECT 1376.6800 2634.0000 1379.6800 2634.4800 ;
        RECT 1376.6800 2628.5600 1379.6800 2629.0400 ;
        RECT 1376.6800 2639.4400 1379.6800 2639.9200 ;
        RECT 1376.6800 2617.6800 1379.6800 2618.1600 ;
        RECT 1376.6800 2623.1200 1379.6800 2623.6000 ;
        RECT 1376.6800 2612.2400 1379.6800 2612.7200 ;
        RECT 1376.6800 2810.4300 1575.7800 2813.4300 ;
        RECT 1376.6800 2605.3300 1575.7800 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 2375.6900 1562.8400 2583.7900 ;
        RECT 1516.2400 2375.6900 1517.8400 2583.7900 ;
        RECT 1471.2400 2375.6900 1472.8400 2583.7900 ;
        RECT 1426.2400 2375.6900 1427.8400 2583.7900 ;
        RECT 1572.7800 2375.6900 1575.7800 2583.7900 ;
        RECT 1376.6800 2375.6900 1379.6800 2583.7900 ;
      LAYER met3 ;
        RECT 1572.7800 2578.4400 1575.7800 2578.9200 ;
        RECT 1561.2400 2578.4400 1562.8400 2578.9200 ;
        RECT 1572.7800 2567.5600 1575.7800 2568.0400 ;
        RECT 1572.7800 2573.0000 1575.7800 2573.4800 ;
        RECT 1561.2400 2567.5600 1562.8400 2568.0400 ;
        RECT 1561.2400 2573.0000 1562.8400 2573.4800 ;
        RECT 1572.7800 2551.2400 1575.7800 2551.7200 ;
        RECT 1572.7800 2556.6800 1575.7800 2557.1600 ;
        RECT 1561.2400 2551.2400 1562.8400 2551.7200 ;
        RECT 1561.2400 2556.6800 1562.8400 2557.1600 ;
        RECT 1572.7800 2540.3600 1575.7800 2540.8400 ;
        RECT 1572.7800 2545.8000 1575.7800 2546.2800 ;
        RECT 1561.2400 2540.3600 1562.8400 2540.8400 ;
        RECT 1561.2400 2545.8000 1562.8400 2546.2800 ;
        RECT 1572.7800 2562.1200 1575.7800 2562.6000 ;
        RECT 1561.2400 2562.1200 1562.8400 2562.6000 ;
        RECT 1516.2400 2567.5600 1517.8400 2568.0400 ;
        RECT 1516.2400 2573.0000 1517.8400 2573.4800 ;
        RECT 1516.2400 2578.4400 1517.8400 2578.9200 ;
        RECT 1516.2400 2551.2400 1517.8400 2551.7200 ;
        RECT 1516.2400 2556.6800 1517.8400 2557.1600 ;
        RECT 1516.2400 2545.8000 1517.8400 2546.2800 ;
        RECT 1516.2400 2540.3600 1517.8400 2540.8400 ;
        RECT 1516.2400 2562.1200 1517.8400 2562.6000 ;
        RECT 1572.7800 2524.0400 1575.7800 2524.5200 ;
        RECT 1572.7800 2529.4800 1575.7800 2529.9600 ;
        RECT 1561.2400 2524.0400 1562.8400 2524.5200 ;
        RECT 1561.2400 2529.4800 1562.8400 2529.9600 ;
        RECT 1572.7800 2507.7200 1575.7800 2508.2000 ;
        RECT 1572.7800 2513.1600 1575.7800 2513.6400 ;
        RECT 1572.7800 2518.6000 1575.7800 2519.0800 ;
        RECT 1561.2400 2507.7200 1562.8400 2508.2000 ;
        RECT 1561.2400 2513.1600 1562.8400 2513.6400 ;
        RECT 1561.2400 2518.6000 1562.8400 2519.0800 ;
        RECT 1572.7800 2496.8400 1575.7800 2497.3200 ;
        RECT 1572.7800 2502.2800 1575.7800 2502.7600 ;
        RECT 1561.2400 2496.8400 1562.8400 2497.3200 ;
        RECT 1561.2400 2502.2800 1562.8400 2502.7600 ;
        RECT 1572.7800 2480.5200 1575.7800 2481.0000 ;
        RECT 1572.7800 2485.9600 1575.7800 2486.4400 ;
        RECT 1572.7800 2491.4000 1575.7800 2491.8800 ;
        RECT 1561.2400 2480.5200 1562.8400 2481.0000 ;
        RECT 1561.2400 2485.9600 1562.8400 2486.4400 ;
        RECT 1561.2400 2491.4000 1562.8400 2491.8800 ;
        RECT 1516.2400 2524.0400 1517.8400 2524.5200 ;
        RECT 1516.2400 2529.4800 1517.8400 2529.9600 ;
        RECT 1516.2400 2507.7200 1517.8400 2508.2000 ;
        RECT 1516.2400 2513.1600 1517.8400 2513.6400 ;
        RECT 1516.2400 2518.6000 1517.8400 2519.0800 ;
        RECT 1516.2400 2496.8400 1517.8400 2497.3200 ;
        RECT 1516.2400 2502.2800 1517.8400 2502.7600 ;
        RECT 1516.2400 2480.5200 1517.8400 2481.0000 ;
        RECT 1516.2400 2485.9600 1517.8400 2486.4400 ;
        RECT 1516.2400 2491.4000 1517.8400 2491.8800 ;
        RECT 1572.7800 2534.9200 1575.7800 2535.4000 ;
        RECT 1516.2400 2534.9200 1517.8400 2535.4000 ;
        RECT 1561.2400 2534.9200 1562.8400 2535.4000 ;
        RECT 1471.2400 2567.5600 1472.8400 2568.0400 ;
        RECT 1471.2400 2573.0000 1472.8400 2573.4800 ;
        RECT 1471.2400 2578.4400 1472.8400 2578.9200 ;
        RECT 1426.2400 2567.5600 1427.8400 2568.0400 ;
        RECT 1426.2400 2573.0000 1427.8400 2573.4800 ;
        RECT 1426.2400 2578.4400 1427.8400 2578.9200 ;
        RECT 1471.2400 2551.2400 1472.8400 2551.7200 ;
        RECT 1471.2400 2556.6800 1472.8400 2557.1600 ;
        RECT 1471.2400 2540.3600 1472.8400 2540.8400 ;
        RECT 1471.2400 2545.8000 1472.8400 2546.2800 ;
        RECT 1426.2400 2551.2400 1427.8400 2551.7200 ;
        RECT 1426.2400 2556.6800 1427.8400 2557.1600 ;
        RECT 1426.2400 2540.3600 1427.8400 2540.8400 ;
        RECT 1426.2400 2545.8000 1427.8400 2546.2800 ;
        RECT 1426.2400 2562.1200 1427.8400 2562.6000 ;
        RECT 1471.2400 2562.1200 1472.8400 2562.6000 ;
        RECT 1376.6800 2578.4400 1379.6800 2578.9200 ;
        RECT 1376.6800 2573.0000 1379.6800 2573.4800 ;
        RECT 1376.6800 2567.5600 1379.6800 2568.0400 ;
        RECT 1376.6800 2556.6800 1379.6800 2557.1600 ;
        RECT 1376.6800 2551.2400 1379.6800 2551.7200 ;
        RECT 1376.6800 2545.8000 1379.6800 2546.2800 ;
        RECT 1376.6800 2540.3600 1379.6800 2540.8400 ;
        RECT 1376.6800 2562.1200 1379.6800 2562.6000 ;
        RECT 1471.2400 2524.0400 1472.8400 2524.5200 ;
        RECT 1471.2400 2529.4800 1472.8400 2529.9600 ;
        RECT 1471.2400 2507.7200 1472.8400 2508.2000 ;
        RECT 1471.2400 2513.1600 1472.8400 2513.6400 ;
        RECT 1471.2400 2518.6000 1472.8400 2519.0800 ;
        RECT 1426.2400 2524.0400 1427.8400 2524.5200 ;
        RECT 1426.2400 2529.4800 1427.8400 2529.9600 ;
        RECT 1426.2400 2507.7200 1427.8400 2508.2000 ;
        RECT 1426.2400 2513.1600 1427.8400 2513.6400 ;
        RECT 1426.2400 2518.6000 1427.8400 2519.0800 ;
        RECT 1471.2400 2496.8400 1472.8400 2497.3200 ;
        RECT 1471.2400 2502.2800 1472.8400 2502.7600 ;
        RECT 1471.2400 2480.5200 1472.8400 2481.0000 ;
        RECT 1471.2400 2485.9600 1472.8400 2486.4400 ;
        RECT 1471.2400 2491.4000 1472.8400 2491.8800 ;
        RECT 1426.2400 2496.8400 1427.8400 2497.3200 ;
        RECT 1426.2400 2502.2800 1427.8400 2502.7600 ;
        RECT 1426.2400 2480.5200 1427.8400 2481.0000 ;
        RECT 1426.2400 2485.9600 1427.8400 2486.4400 ;
        RECT 1426.2400 2491.4000 1427.8400 2491.8800 ;
        RECT 1376.6800 2524.0400 1379.6800 2524.5200 ;
        RECT 1376.6800 2529.4800 1379.6800 2529.9600 ;
        RECT 1376.6800 2513.1600 1379.6800 2513.6400 ;
        RECT 1376.6800 2507.7200 1379.6800 2508.2000 ;
        RECT 1376.6800 2518.6000 1379.6800 2519.0800 ;
        RECT 1376.6800 2496.8400 1379.6800 2497.3200 ;
        RECT 1376.6800 2502.2800 1379.6800 2502.7600 ;
        RECT 1376.6800 2485.9600 1379.6800 2486.4400 ;
        RECT 1376.6800 2480.5200 1379.6800 2481.0000 ;
        RECT 1376.6800 2491.4000 1379.6800 2491.8800 ;
        RECT 1376.6800 2534.9200 1379.6800 2535.4000 ;
        RECT 1426.2400 2534.9200 1427.8400 2535.4000 ;
        RECT 1471.2400 2534.9200 1472.8400 2535.4000 ;
        RECT 1572.7800 2469.6400 1575.7800 2470.1200 ;
        RECT 1572.7800 2475.0800 1575.7800 2475.5600 ;
        RECT 1561.2400 2469.6400 1562.8400 2470.1200 ;
        RECT 1561.2400 2475.0800 1562.8400 2475.5600 ;
        RECT 1572.7800 2453.3200 1575.7800 2453.8000 ;
        RECT 1572.7800 2458.7600 1575.7800 2459.2400 ;
        RECT 1572.7800 2464.2000 1575.7800 2464.6800 ;
        RECT 1561.2400 2453.3200 1562.8400 2453.8000 ;
        RECT 1561.2400 2458.7600 1562.8400 2459.2400 ;
        RECT 1561.2400 2464.2000 1562.8400 2464.6800 ;
        RECT 1572.7800 2442.4400 1575.7800 2442.9200 ;
        RECT 1572.7800 2447.8800 1575.7800 2448.3600 ;
        RECT 1561.2400 2442.4400 1562.8400 2442.9200 ;
        RECT 1561.2400 2447.8800 1562.8400 2448.3600 ;
        RECT 1572.7800 2426.1200 1575.7800 2426.6000 ;
        RECT 1572.7800 2431.5600 1575.7800 2432.0400 ;
        RECT 1572.7800 2437.0000 1575.7800 2437.4800 ;
        RECT 1561.2400 2426.1200 1562.8400 2426.6000 ;
        RECT 1561.2400 2431.5600 1562.8400 2432.0400 ;
        RECT 1561.2400 2437.0000 1562.8400 2437.4800 ;
        RECT 1516.2400 2469.6400 1517.8400 2470.1200 ;
        RECT 1516.2400 2475.0800 1517.8400 2475.5600 ;
        RECT 1516.2400 2453.3200 1517.8400 2453.8000 ;
        RECT 1516.2400 2458.7600 1517.8400 2459.2400 ;
        RECT 1516.2400 2464.2000 1517.8400 2464.6800 ;
        RECT 1516.2400 2442.4400 1517.8400 2442.9200 ;
        RECT 1516.2400 2447.8800 1517.8400 2448.3600 ;
        RECT 1516.2400 2426.1200 1517.8400 2426.6000 ;
        RECT 1516.2400 2431.5600 1517.8400 2432.0400 ;
        RECT 1516.2400 2437.0000 1517.8400 2437.4800 ;
        RECT 1572.7800 2415.2400 1575.7800 2415.7200 ;
        RECT 1572.7800 2420.6800 1575.7800 2421.1600 ;
        RECT 1561.2400 2415.2400 1562.8400 2415.7200 ;
        RECT 1561.2400 2420.6800 1562.8400 2421.1600 ;
        RECT 1572.7800 2398.9200 1575.7800 2399.4000 ;
        RECT 1572.7800 2404.3600 1575.7800 2404.8400 ;
        RECT 1572.7800 2409.8000 1575.7800 2410.2800 ;
        RECT 1561.2400 2398.9200 1562.8400 2399.4000 ;
        RECT 1561.2400 2404.3600 1562.8400 2404.8400 ;
        RECT 1561.2400 2409.8000 1562.8400 2410.2800 ;
        RECT 1572.7800 2388.0400 1575.7800 2388.5200 ;
        RECT 1572.7800 2393.4800 1575.7800 2393.9600 ;
        RECT 1561.2400 2388.0400 1562.8400 2388.5200 ;
        RECT 1561.2400 2393.4800 1562.8400 2393.9600 ;
        RECT 1572.7800 2382.6000 1575.7800 2383.0800 ;
        RECT 1561.2400 2382.6000 1562.8400 2383.0800 ;
        RECT 1516.2400 2415.2400 1517.8400 2415.7200 ;
        RECT 1516.2400 2420.6800 1517.8400 2421.1600 ;
        RECT 1516.2400 2398.9200 1517.8400 2399.4000 ;
        RECT 1516.2400 2404.3600 1517.8400 2404.8400 ;
        RECT 1516.2400 2409.8000 1517.8400 2410.2800 ;
        RECT 1516.2400 2388.0400 1517.8400 2388.5200 ;
        RECT 1516.2400 2393.4800 1517.8400 2393.9600 ;
        RECT 1516.2400 2382.6000 1517.8400 2383.0800 ;
        RECT 1471.2400 2469.6400 1472.8400 2470.1200 ;
        RECT 1471.2400 2475.0800 1472.8400 2475.5600 ;
        RECT 1471.2400 2453.3200 1472.8400 2453.8000 ;
        RECT 1471.2400 2458.7600 1472.8400 2459.2400 ;
        RECT 1471.2400 2464.2000 1472.8400 2464.6800 ;
        RECT 1426.2400 2469.6400 1427.8400 2470.1200 ;
        RECT 1426.2400 2475.0800 1427.8400 2475.5600 ;
        RECT 1426.2400 2453.3200 1427.8400 2453.8000 ;
        RECT 1426.2400 2458.7600 1427.8400 2459.2400 ;
        RECT 1426.2400 2464.2000 1427.8400 2464.6800 ;
        RECT 1471.2400 2442.4400 1472.8400 2442.9200 ;
        RECT 1471.2400 2447.8800 1472.8400 2448.3600 ;
        RECT 1471.2400 2426.1200 1472.8400 2426.6000 ;
        RECT 1471.2400 2431.5600 1472.8400 2432.0400 ;
        RECT 1471.2400 2437.0000 1472.8400 2437.4800 ;
        RECT 1426.2400 2442.4400 1427.8400 2442.9200 ;
        RECT 1426.2400 2447.8800 1427.8400 2448.3600 ;
        RECT 1426.2400 2426.1200 1427.8400 2426.6000 ;
        RECT 1426.2400 2431.5600 1427.8400 2432.0400 ;
        RECT 1426.2400 2437.0000 1427.8400 2437.4800 ;
        RECT 1376.6800 2469.6400 1379.6800 2470.1200 ;
        RECT 1376.6800 2475.0800 1379.6800 2475.5600 ;
        RECT 1376.6800 2458.7600 1379.6800 2459.2400 ;
        RECT 1376.6800 2453.3200 1379.6800 2453.8000 ;
        RECT 1376.6800 2464.2000 1379.6800 2464.6800 ;
        RECT 1376.6800 2442.4400 1379.6800 2442.9200 ;
        RECT 1376.6800 2447.8800 1379.6800 2448.3600 ;
        RECT 1376.6800 2431.5600 1379.6800 2432.0400 ;
        RECT 1376.6800 2426.1200 1379.6800 2426.6000 ;
        RECT 1376.6800 2437.0000 1379.6800 2437.4800 ;
        RECT 1471.2400 2415.2400 1472.8400 2415.7200 ;
        RECT 1471.2400 2420.6800 1472.8400 2421.1600 ;
        RECT 1471.2400 2398.9200 1472.8400 2399.4000 ;
        RECT 1471.2400 2404.3600 1472.8400 2404.8400 ;
        RECT 1471.2400 2409.8000 1472.8400 2410.2800 ;
        RECT 1426.2400 2415.2400 1427.8400 2415.7200 ;
        RECT 1426.2400 2420.6800 1427.8400 2421.1600 ;
        RECT 1426.2400 2398.9200 1427.8400 2399.4000 ;
        RECT 1426.2400 2404.3600 1427.8400 2404.8400 ;
        RECT 1426.2400 2409.8000 1427.8400 2410.2800 ;
        RECT 1471.2400 2393.4800 1472.8400 2393.9600 ;
        RECT 1471.2400 2388.0400 1472.8400 2388.5200 ;
        RECT 1471.2400 2382.6000 1472.8400 2383.0800 ;
        RECT 1426.2400 2393.4800 1427.8400 2393.9600 ;
        RECT 1426.2400 2388.0400 1427.8400 2388.5200 ;
        RECT 1426.2400 2382.6000 1427.8400 2383.0800 ;
        RECT 1376.6800 2415.2400 1379.6800 2415.7200 ;
        RECT 1376.6800 2420.6800 1379.6800 2421.1600 ;
        RECT 1376.6800 2404.3600 1379.6800 2404.8400 ;
        RECT 1376.6800 2398.9200 1379.6800 2399.4000 ;
        RECT 1376.6800 2409.8000 1379.6800 2410.2800 ;
        RECT 1376.6800 2388.0400 1379.6800 2388.5200 ;
        RECT 1376.6800 2393.4800 1379.6800 2393.9600 ;
        RECT 1376.6800 2382.6000 1379.6800 2383.0800 ;
        RECT 1376.6800 2580.7900 1575.7800 2583.7900 ;
        RECT 1376.6800 2375.6900 1575.7800 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 2146.0500 1562.8400 2354.1500 ;
        RECT 1516.2400 2146.0500 1517.8400 2354.1500 ;
        RECT 1471.2400 2146.0500 1472.8400 2354.1500 ;
        RECT 1426.2400 2146.0500 1427.8400 2354.1500 ;
        RECT 1572.7800 2146.0500 1575.7800 2354.1500 ;
        RECT 1376.6800 2146.0500 1379.6800 2354.1500 ;
      LAYER met3 ;
        RECT 1572.7800 2348.8000 1575.7800 2349.2800 ;
        RECT 1561.2400 2348.8000 1562.8400 2349.2800 ;
        RECT 1572.7800 2337.9200 1575.7800 2338.4000 ;
        RECT 1572.7800 2343.3600 1575.7800 2343.8400 ;
        RECT 1561.2400 2337.9200 1562.8400 2338.4000 ;
        RECT 1561.2400 2343.3600 1562.8400 2343.8400 ;
        RECT 1572.7800 2321.6000 1575.7800 2322.0800 ;
        RECT 1572.7800 2327.0400 1575.7800 2327.5200 ;
        RECT 1561.2400 2321.6000 1562.8400 2322.0800 ;
        RECT 1561.2400 2327.0400 1562.8400 2327.5200 ;
        RECT 1572.7800 2310.7200 1575.7800 2311.2000 ;
        RECT 1572.7800 2316.1600 1575.7800 2316.6400 ;
        RECT 1561.2400 2310.7200 1562.8400 2311.2000 ;
        RECT 1561.2400 2316.1600 1562.8400 2316.6400 ;
        RECT 1572.7800 2332.4800 1575.7800 2332.9600 ;
        RECT 1561.2400 2332.4800 1562.8400 2332.9600 ;
        RECT 1516.2400 2337.9200 1517.8400 2338.4000 ;
        RECT 1516.2400 2343.3600 1517.8400 2343.8400 ;
        RECT 1516.2400 2348.8000 1517.8400 2349.2800 ;
        RECT 1516.2400 2321.6000 1517.8400 2322.0800 ;
        RECT 1516.2400 2327.0400 1517.8400 2327.5200 ;
        RECT 1516.2400 2316.1600 1517.8400 2316.6400 ;
        RECT 1516.2400 2310.7200 1517.8400 2311.2000 ;
        RECT 1516.2400 2332.4800 1517.8400 2332.9600 ;
        RECT 1572.7800 2294.4000 1575.7800 2294.8800 ;
        RECT 1572.7800 2299.8400 1575.7800 2300.3200 ;
        RECT 1561.2400 2294.4000 1562.8400 2294.8800 ;
        RECT 1561.2400 2299.8400 1562.8400 2300.3200 ;
        RECT 1572.7800 2278.0800 1575.7800 2278.5600 ;
        RECT 1572.7800 2283.5200 1575.7800 2284.0000 ;
        RECT 1572.7800 2288.9600 1575.7800 2289.4400 ;
        RECT 1561.2400 2278.0800 1562.8400 2278.5600 ;
        RECT 1561.2400 2283.5200 1562.8400 2284.0000 ;
        RECT 1561.2400 2288.9600 1562.8400 2289.4400 ;
        RECT 1572.7800 2267.2000 1575.7800 2267.6800 ;
        RECT 1572.7800 2272.6400 1575.7800 2273.1200 ;
        RECT 1561.2400 2267.2000 1562.8400 2267.6800 ;
        RECT 1561.2400 2272.6400 1562.8400 2273.1200 ;
        RECT 1572.7800 2250.8800 1575.7800 2251.3600 ;
        RECT 1572.7800 2256.3200 1575.7800 2256.8000 ;
        RECT 1572.7800 2261.7600 1575.7800 2262.2400 ;
        RECT 1561.2400 2250.8800 1562.8400 2251.3600 ;
        RECT 1561.2400 2256.3200 1562.8400 2256.8000 ;
        RECT 1561.2400 2261.7600 1562.8400 2262.2400 ;
        RECT 1516.2400 2294.4000 1517.8400 2294.8800 ;
        RECT 1516.2400 2299.8400 1517.8400 2300.3200 ;
        RECT 1516.2400 2278.0800 1517.8400 2278.5600 ;
        RECT 1516.2400 2283.5200 1517.8400 2284.0000 ;
        RECT 1516.2400 2288.9600 1517.8400 2289.4400 ;
        RECT 1516.2400 2267.2000 1517.8400 2267.6800 ;
        RECT 1516.2400 2272.6400 1517.8400 2273.1200 ;
        RECT 1516.2400 2250.8800 1517.8400 2251.3600 ;
        RECT 1516.2400 2256.3200 1517.8400 2256.8000 ;
        RECT 1516.2400 2261.7600 1517.8400 2262.2400 ;
        RECT 1572.7800 2305.2800 1575.7800 2305.7600 ;
        RECT 1516.2400 2305.2800 1517.8400 2305.7600 ;
        RECT 1561.2400 2305.2800 1562.8400 2305.7600 ;
        RECT 1471.2400 2337.9200 1472.8400 2338.4000 ;
        RECT 1471.2400 2343.3600 1472.8400 2343.8400 ;
        RECT 1471.2400 2348.8000 1472.8400 2349.2800 ;
        RECT 1426.2400 2337.9200 1427.8400 2338.4000 ;
        RECT 1426.2400 2343.3600 1427.8400 2343.8400 ;
        RECT 1426.2400 2348.8000 1427.8400 2349.2800 ;
        RECT 1471.2400 2321.6000 1472.8400 2322.0800 ;
        RECT 1471.2400 2327.0400 1472.8400 2327.5200 ;
        RECT 1471.2400 2310.7200 1472.8400 2311.2000 ;
        RECT 1471.2400 2316.1600 1472.8400 2316.6400 ;
        RECT 1426.2400 2321.6000 1427.8400 2322.0800 ;
        RECT 1426.2400 2327.0400 1427.8400 2327.5200 ;
        RECT 1426.2400 2310.7200 1427.8400 2311.2000 ;
        RECT 1426.2400 2316.1600 1427.8400 2316.6400 ;
        RECT 1426.2400 2332.4800 1427.8400 2332.9600 ;
        RECT 1471.2400 2332.4800 1472.8400 2332.9600 ;
        RECT 1376.6800 2348.8000 1379.6800 2349.2800 ;
        RECT 1376.6800 2343.3600 1379.6800 2343.8400 ;
        RECT 1376.6800 2337.9200 1379.6800 2338.4000 ;
        RECT 1376.6800 2327.0400 1379.6800 2327.5200 ;
        RECT 1376.6800 2321.6000 1379.6800 2322.0800 ;
        RECT 1376.6800 2316.1600 1379.6800 2316.6400 ;
        RECT 1376.6800 2310.7200 1379.6800 2311.2000 ;
        RECT 1376.6800 2332.4800 1379.6800 2332.9600 ;
        RECT 1471.2400 2294.4000 1472.8400 2294.8800 ;
        RECT 1471.2400 2299.8400 1472.8400 2300.3200 ;
        RECT 1471.2400 2278.0800 1472.8400 2278.5600 ;
        RECT 1471.2400 2283.5200 1472.8400 2284.0000 ;
        RECT 1471.2400 2288.9600 1472.8400 2289.4400 ;
        RECT 1426.2400 2294.4000 1427.8400 2294.8800 ;
        RECT 1426.2400 2299.8400 1427.8400 2300.3200 ;
        RECT 1426.2400 2278.0800 1427.8400 2278.5600 ;
        RECT 1426.2400 2283.5200 1427.8400 2284.0000 ;
        RECT 1426.2400 2288.9600 1427.8400 2289.4400 ;
        RECT 1471.2400 2267.2000 1472.8400 2267.6800 ;
        RECT 1471.2400 2272.6400 1472.8400 2273.1200 ;
        RECT 1471.2400 2250.8800 1472.8400 2251.3600 ;
        RECT 1471.2400 2256.3200 1472.8400 2256.8000 ;
        RECT 1471.2400 2261.7600 1472.8400 2262.2400 ;
        RECT 1426.2400 2267.2000 1427.8400 2267.6800 ;
        RECT 1426.2400 2272.6400 1427.8400 2273.1200 ;
        RECT 1426.2400 2250.8800 1427.8400 2251.3600 ;
        RECT 1426.2400 2256.3200 1427.8400 2256.8000 ;
        RECT 1426.2400 2261.7600 1427.8400 2262.2400 ;
        RECT 1376.6800 2294.4000 1379.6800 2294.8800 ;
        RECT 1376.6800 2299.8400 1379.6800 2300.3200 ;
        RECT 1376.6800 2283.5200 1379.6800 2284.0000 ;
        RECT 1376.6800 2278.0800 1379.6800 2278.5600 ;
        RECT 1376.6800 2288.9600 1379.6800 2289.4400 ;
        RECT 1376.6800 2267.2000 1379.6800 2267.6800 ;
        RECT 1376.6800 2272.6400 1379.6800 2273.1200 ;
        RECT 1376.6800 2256.3200 1379.6800 2256.8000 ;
        RECT 1376.6800 2250.8800 1379.6800 2251.3600 ;
        RECT 1376.6800 2261.7600 1379.6800 2262.2400 ;
        RECT 1376.6800 2305.2800 1379.6800 2305.7600 ;
        RECT 1426.2400 2305.2800 1427.8400 2305.7600 ;
        RECT 1471.2400 2305.2800 1472.8400 2305.7600 ;
        RECT 1572.7800 2240.0000 1575.7800 2240.4800 ;
        RECT 1572.7800 2245.4400 1575.7800 2245.9200 ;
        RECT 1561.2400 2240.0000 1562.8400 2240.4800 ;
        RECT 1561.2400 2245.4400 1562.8400 2245.9200 ;
        RECT 1572.7800 2223.6800 1575.7800 2224.1600 ;
        RECT 1572.7800 2229.1200 1575.7800 2229.6000 ;
        RECT 1572.7800 2234.5600 1575.7800 2235.0400 ;
        RECT 1561.2400 2223.6800 1562.8400 2224.1600 ;
        RECT 1561.2400 2229.1200 1562.8400 2229.6000 ;
        RECT 1561.2400 2234.5600 1562.8400 2235.0400 ;
        RECT 1572.7800 2212.8000 1575.7800 2213.2800 ;
        RECT 1572.7800 2218.2400 1575.7800 2218.7200 ;
        RECT 1561.2400 2212.8000 1562.8400 2213.2800 ;
        RECT 1561.2400 2218.2400 1562.8400 2218.7200 ;
        RECT 1572.7800 2196.4800 1575.7800 2196.9600 ;
        RECT 1572.7800 2201.9200 1575.7800 2202.4000 ;
        RECT 1572.7800 2207.3600 1575.7800 2207.8400 ;
        RECT 1561.2400 2196.4800 1562.8400 2196.9600 ;
        RECT 1561.2400 2201.9200 1562.8400 2202.4000 ;
        RECT 1561.2400 2207.3600 1562.8400 2207.8400 ;
        RECT 1516.2400 2240.0000 1517.8400 2240.4800 ;
        RECT 1516.2400 2245.4400 1517.8400 2245.9200 ;
        RECT 1516.2400 2223.6800 1517.8400 2224.1600 ;
        RECT 1516.2400 2229.1200 1517.8400 2229.6000 ;
        RECT 1516.2400 2234.5600 1517.8400 2235.0400 ;
        RECT 1516.2400 2212.8000 1517.8400 2213.2800 ;
        RECT 1516.2400 2218.2400 1517.8400 2218.7200 ;
        RECT 1516.2400 2196.4800 1517.8400 2196.9600 ;
        RECT 1516.2400 2201.9200 1517.8400 2202.4000 ;
        RECT 1516.2400 2207.3600 1517.8400 2207.8400 ;
        RECT 1572.7800 2185.6000 1575.7800 2186.0800 ;
        RECT 1572.7800 2191.0400 1575.7800 2191.5200 ;
        RECT 1561.2400 2185.6000 1562.8400 2186.0800 ;
        RECT 1561.2400 2191.0400 1562.8400 2191.5200 ;
        RECT 1572.7800 2169.2800 1575.7800 2169.7600 ;
        RECT 1572.7800 2174.7200 1575.7800 2175.2000 ;
        RECT 1572.7800 2180.1600 1575.7800 2180.6400 ;
        RECT 1561.2400 2169.2800 1562.8400 2169.7600 ;
        RECT 1561.2400 2174.7200 1562.8400 2175.2000 ;
        RECT 1561.2400 2180.1600 1562.8400 2180.6400 ;
        RECT 1572.7800 2158.4000 1575.7800 2158.8800 ;
        RECT 1572.7800 2163.8400 1575.7800 2164.3200 ;
        RECT 1561.2400 2158.4000 1562.8400 2158.8800 ;
        RECT 1561.2400 2163.8400 1562.8400 2164.3200 ;
        RECT 1572.7800 2152.9600 1575.7800 2153.4400 ;
        RECT 1561.2400 2152.9600 1562.8400 2153.4400 ;
        RECT 1516.2400 2185.6000 1517.8400 2186.0800 ;
        RECT 1516.2400 2191.0400 1517.8400 2191.5200 ;
        RECT 1516.2400 2169.2800 1517.8400 2169.7600 ;
        RECT 1516.2400 2174.7200 1517.8400 2175.2000 ;
        RECT 1516.2400 2180.1600 1517.8400 2180.6400 ;
        RECT 1516.2400 2158.4000 1517.8400 2158.8800 ;
        RECT 1516.2400 2163.8400 1517.8400 2164.3200 ;
        RECT 1516.2400 2152.9600 1517.8400 2153.4400 ;
        RECT 1471.2400 2240.0000 1472.8400 2240.4800 ;
        RECT 1471.2400 2245.4400 1472.8400 2245.9200 ;
        RECT 1471.2400 2223.6800 1472.8400 2224.1600 ;
        RECT 1471.2400 2229.1200 1472.8400 2229.6000 ;
        RECT 1471.2400 2234.5600 1472.8400 2235.0400 ;
        RECT 1426.2400 2240.0000 1427.8400 2240.4800 ;
        RECT 1426.2400 2245.4400 1427.8400 2245.9200 ;
        RECT 1426.2400 2223.6800 1427.8400 2224.1600 ;
        RECT 1426.2400 2229.1200 1427.8400 2229.6000 ;
        RECT 1426.2400 2234.5600 1427.8400 2235.0400 ;
        RECT 1471.2400 2212.8000 1472.8400 2213.2800 ;
        RECT 1471.2400 2218.2400 1472.8400 2218.7200 ;
        RECT 1471.2400 2196.4800 1472.8400 2196.9600 ;
        RECT 1471.2400 2201.9200 1472.8400 2202.4000 ;
        RECT 1471.2400 2207.3600 1472.8400 2207.8400 ;
        RECT 1426.2400 2212.8000 1427.8400 2213.2800 ;
        RECT 1426.2400 2218.2400 1427.8400 2218.7200 ;
        RECT 1426.2400 2196.4800 1427.8400 2196.9600 ;
        RECT 1426.2400 2201.9200 1427.8400 2202.4000 ;
        RECT 1426.2400 2207.3600 1427.8400 2207.8400 ;
        RECT 1376.6800 2240.0000 1379.6800 2240.4800 ;
        RECT 1376.6800 2245.4400 1379.6800 2245.9200 ;
        RECT 1376.6800 2229.1200 1379.6800 2229.6000 ;
        RECT 1376.6800 2223.6800 1379.6800 2224.1600 ;
        RECT 1376.6800 2234.5600 1379.6800 2235.0400 ;
        RECT 1376.6800 2212.8000 1379.6800 2213.2800 ;
        RECT 1376.6800 2218.2400 1379.6800 2218.7200 ;
        RECT 1376.6800 2201.9200 1379.6800 2202.4000 ;
        RECT 1376.6800 2196.4800 1379.6800 2196.9600 ;
        RECT 1376.6800 2207.3600 1379.6800 2207.8400 ;
        RECT 1471.2400 2185.6000 1472.8400 2186.0800 ;
        RECT 1471.2400 2191.0400 1472.8400 2191.5200 ;
        RECT 1471.2400 2169.2800 1472.8400 2169.7600 ;
        RECT 1471.2400 2174.7200 1472.8400 2175.2000 ;
        RECT 1471.2400 2180.1600 1472.8400 2180.6400 ;
        RECT 1426.2400 2185.6000 1427.8400 2186.0800 ;
        RECT 1426.2400 2191.0400 1427.8400 2191.5200 ;
        RECT 1426.2400 2169.2800 1427.8400 2169.7600 ;
        RECT 1426.2400 2174.7200 1427.8400 2175.2000 ;
        RECT 1426.2400 2180.1600 1427.8400 2180.6400 ;
        RECT 1471.2400 2163.8400 1472.8400 2164.3200 ;
        RECT 1471.2400 2158.4000 1472.8400 2158.8800 ;
        RECT 1471.2400 2152.9600 1472.8400 2153.4400 ;
        RECT 1426.2400 2163.8400 1427.8400 2164.3200 ;
        RECT 1426.2400 2158.4000 1427.8400 2158.8800 ;
        RECT 1426.2400 2152.9600 1427.8400 2153.4400 ;
        RECT 1376.6800 2185.6000 1379.6800 2186.0800 ;
        RECT 1376.6800 2191.0400 1379.6800 2191.5200 ;
        RECT 1376.6800 2174.7200 1379.6800 2175.2000 ;
        RECT 1376.6800 2169.2800 1379.6800 2169.7600 ;
        RECT 1376.6800 2180.1600 1379.6800 2180.6400 ;
        RECT 1376.6800 2158.4000 1379.6800 2158.8800 ;
        RECT 1376.6800 2163.8400 1379.6800 2164.3200 ;
        RECT 1376.6800 2152.9600 1379.6800 2153.4400 ;
        RECT 1376.6800 2351.1500 1575.7800 2354.1500 ;
        RECT 1376.6800 2146.0500 1575.7800 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 1916.4100 1562.8400 2124.5100 ;
        RECT 1516.2400 1916.4100 1517.8400 2124.5100 ;
        RECT 1471.2400 1916.4100 1472.8400 2124.5100 ;
        RECT 1426.2400 1916.4100 1427.8400 2124.5100 ;
        RECT 1572.7800 1916.4100 1575.7800 2124.5100 ;
        RECT 1376.6800 1916.4100 1379.6800 2124.5100 ;
      LAYER met3 ;
        RECT 1572.7800 2119.1600 1575.7800 2119.6400 ;
        RECT 1561.2400 2119.1600 1562.8400 2119.6400 ;
        RECT 1572.7800 2108.2800 1575.7800 2108.7600 ;
        RECT 1572.7800 2113.7200 1575.7800 2114.2000 ;
        RECT 1561.2400 2108.2800 1562.8400 2108.7600 ;
        RECT 1561.2400 2113.7200 1562.8400 2114.2000 ;
        RECT 1572.7800 2091.9600 1575.7800 2092.4400 ;
        RECT 1572.7800 2097.4000 1575.7800 2097.8800 ;
        RECT 1561.2400 2091.9600 1562.8400 2092.4400 ;
        RECT 1561.2400 2097.4000 1562.8400 2097.8800 ;
        RECT 1572.7800 2081.0800 1575.7800 2081.5600 ;
        RECT 1572.7800 2086.5200 1575.7800 2087.0000 ;
        RECT 1561.2400 2081.0800 1562.8400 2081.5600 ;
        RECT 1561.2400 2086.5200 1562.8400 2087.0000 ;
        RECT 1572.7800 2102.8400 1575.7800 2103.3200 ;
        RECT 1561.2400 2102.8400 1562.8400 2103.3200 ;
        RECT 1516.2400 2108.2800 1517.8400 2108.7600 ;
        RECT 1516.2400 2113.7200 1517.8400 2114.2000 ;
        RECT 1516.2400 2119.1600 1517.8400 2119.6400 ;
        RECT 1516.2400 2091.9600 1517.8400 2092.4400 ;
        RECT 1516.2400 2097.4000 1517.8400 2097.8800 ;
        RECT 1516.2400 2086.5200 1517.8400 2087.0000 ;
        RECT 1516.2400 2081.0800 1517.8400 2081.5600 ;
        RECT 1516.2400 2102.8400 1517.8400 2103.3200 ;
        RECT 1572.7800 2064.7600 1575.7800 2065.2400 ;
        RECT 1572.7800 2070.2000 1575.7800 2070.6800 ;
        RECT 1561.2400 2064.7600 1562.8400 2065.2400 ;
        RECT 1561.2400 2070.2000 1562.8400 2070.6800 ;
        RECT 1572.7800 2048.4400 1575.7800 2048.9200 ;
        RECT 1572.7800 2053.8800 1575.7800 2054.3600 ;
        RECT 1572.7800 2059.3200 1575.7800 2059.8000 ;
        RECT 1561.2400 2048.4400 1562.8400 2048.9200 ;
        RECT 1561.2400 2053.8800 1562.8400 2054.3600 ;
        RECT 1561.2400 2059.3200 1562.8400 2059.8000 ;
        RECT 1572.7800 2037.5600 1575.7800 2038.0400 ;
        RECT 1572.7800 2043.0000 1575.7800 2043.4800 ;
        RECT 1561.2400 2037.5600 1562.8400 2038.0400 ;
        RECT 1561.2400 2043.0000 1562.8400 2043.4800 ;
        RECT 1572.7800 2021.2400 1575.7800 2021.7200 ;
        RECT 1572.7800 2026.6800 1575.7800 2027.1600 ;
        RECT 1572.7800 2032.1200 1575.7800 2032.6000 ;
        RECT 1561.2400 2021.2400 1562.8400 2021.7200 ;
        RECT 1561.2400 2026.6800 1562.8400 2027.1600 ;
        RECT 1561.2400 2032.1200 1562.8400 2032.6000 ;
        RECT 1516.2400 2064.7600 1517.8400 2065.2400 ;
        RECT 1516.2400 2070.2000 1517.8400 2070.6800 ;
        RECT 1516.2400 2048.4400 1517.8400 2048.9200 ;
        RECT 1516.2400 2053.8800 1517.8400 2054.3600 ;
        RECT 1516.2400 2059.3200 1517.8400 2059.8000 ;
        RECT 1516.2400 2037.5600 1517.8400 2038.0400 ;
        RECT 1516.2400 2043.0000 1517.8400 2043.4800 ;
        RECT 1516.2400 2021.2400 1517.8400 2021.7200 ;
        RECT 1516.2400 2026.6800 1517.8400 2027.1600 ;
        RECT 1516.2400 2032.1200 1517.8400 2032.6000 ;
        RECT 1572.7800 2075.6400 1575.7800 2076.1200 ;
        RECT 1516.2400 2075.6400 1517.8400 2076.1200 ;
        RECT 1561.2400 2075.6400 1562.8400 2076.1200 ;
        RECT 1471.2400 2108.2800 1472.8400 2108.7600 ;
        RECT 1471.2400 2113.7200 1472.8400 2114.2000 ;
        RECT 1471.2400 2119.1600 1472.8400 2119.6400 ;
        RECT 1426.2400 2108.2800 1427.8400 2108.7600 ;
        RECT 1426.2400 2113.7200 1427.8400 2114.2000 ;
        RECT 1426.2400 2119.1600 1427.8400 2119.6400 ;
        RECT 1471.2400 2091.9600 1472.8400 2092.4400 ;
        RECT 1471.2400 2097.4000 1472.8400 2097.8800 ;
        RECT 1471.2400 2081.0800 1472.8400 2081.5600 ;
        RECT 1471.2400 2086.5200 1472.8400 2087.0000 ;
        RECT 1426.2400 2091.9600 1427.8400 2092.4400 ;
        RECT 1426.2400 2097.4000 1427.8400 2097.8800 ;
        RECT 1426.2400 2081.0800 1427.8400 2081.5600 ;
        RECT 1426.2400 2086.5200 1427.8400 2087.0000 ;
        RECT 1426.2400 2102.8400 1427.8400 2103.3200 ;
        RECT 1471.2400 2102.8400 1472.8400 2103.3200 ;
        RECT 1376.6800 2119.1600 1379.6800 2119.6400 ;
        RECT 1376.6800 2113.7200 1379.6800 2114.2000 ;
        RECT 1376.6800 2108.2800 1379.6800 2108.7600 ;
        RECT 1376.6800 2097.4000 1379.6800 2097.8800 ;
        RECT 1376.6800 2091.9600 1379.6800 2092.4400 ;
        RECT 1376.6800 2086.5200 1379.6800 2087.0000 ;
        RECT 1376.6800 2081.0800 1379.6800 2081.5600 ;
        RECT 1376.6800 2102.8400 1379.6800 2103.3200 ;
        RECT 1471.2400 2064.7600 1472.8400 2065.2400 ;
        RECT 1471.2400 2070.2000 1472.8400 2070.6800 ;
        RECT 1471.2400 2048.4400 1472.8400 2048.9200 ;
        RECT 1471.2400 2053.8800 1472.8400 2054.3600 ;
        RECT 1471.2400 2059.3200 1472.8400 2059.8000 ;
        RECT 1426.2400 2064.7600 1427.8400 2065.2400 ;
        RECT 1426.2400 2070.2000 1427.8400 2070.6800 ;
        RECT 1426.2400 2048.4400 1427.8400 2048.9200 ;
        RECT 1426.2400 2053.8800 1427.8400 2054.3600 ;
        RECT 1426.2400 2059.3200 1427.8400 2059.8000 ;
        RECT 1471.2400 2037.5600 1472.8400 2038.0400 ;
        RECT 1471.2400 2043.0000 1472.8400 2043.4800 ;
        RECT 1471.2400 2021.2400 1472.8400 2021.7200 ;
        RECT 1471.2400 2026.6800 1472.8400 2027.1600 ;
        RECT 1471.2400 2032.1200 1472.8400 2032.6000 ;
        RECT 1426.2400 2037.5600 1427.8400 2038.0400 ;
        RECT 1426.2400 2043.0000 1427.8400 2043.4800 ;
        RECT 1426.2400 2021.2400 1427.8400 2021.7200 ;
        RECT 1426.2400 2026.6800 1427.8400 2027.1600 ;
        RECT 1426.2400 2032.1200 1427.8400 2032.6000 ;
        RECT 1376.6800 2064.7600 1379.6800 2065.2400 ;
        RECT 1376.6800 2070.2000 1379.6800 2070.6800 ;
        RECT 1376.6800 2053.8800 1379.6800 2054.3600 ;
        RECT 1376.6800 2048.4400 1379.6800 2048.9200 ;
        RECT 1376.6800 2059.3200 1379.6800 2059.8000 ;
        RECT 1376.6800 2037.5600 1379.6800 2038.0400 ;
        RECT 1376.6800 2043.0000 1379.6800 2043.4800 ;
        RECT 1376.6800 2026.6800 1379.6800 2027.1600 ;
        RECT 1376.6800 2021.2400 1379.6800 2021.7200 ;
        RECT 1376.6800 2032.1200 1379.6800 2032.6000 ;
        RECT 1376.6800 2075.6400 1379.6800 2076.1200 ;
        RECT 1426.2400 2075.6400 1427.8400 2076.1200 ;
        RECT 1471.2400 2075.6400 1472.8400 2076.1200 ;
        RECT 1572.7800 2010.3600 1575.7800 2010.8400 ;
        RECT 1572.7800 2015.8000 1575.7800 2016.2800 ;
        RECT 1561.2400 2010.3600 1562.8400 2010.8400 ;
        RECT 1561.2400 2015.8000 1562.8400 2016.2800 ;
        RECT 1572.7800 1994.0400 1575.7800 1994.5200 ;
        RECT 1572.7800 1999.4800 1575.7800 1999.9600 ;
        RECT 1572.7800 2004.9200 1575.7800 2005.4000 ;
        RECT 1561.2400 1994.0400 1562.8400 1994.5200 ;
        RECT 1561.2400 1999.4800 1562.8400 1999.9600 ;
        RECT 1561.2400 2004.9200 1562.8400 2005.4000 ;
        RECT 1572.7800 1983.1600 1575.7800 1983.6400 ;
        RECT 1572.7800 1988.6000 1575.7800 1989.0800 ;
        RECT 1561.2400 1983.1600 1562.8400 1983.6400 ;
        RECT 1561.2400 1988.6000 1562.8400 1989.0800 ;
        RECT 1572.7800 1966.8400 1575.7800 1967.3200 ;
        RECT 1572.7800 1972.2800 1575.7800 1972.7600 ;
        RECT 1572.7800 1977.7200 1575.7800 1978.2000 ;
        RECT 1561.2400 1966.8400 1562.8400 1967.3200 ;
        RECT 1561.2400 1972.2800 1562.8400 1972.7600 ;
        RECT 1561.2400 1977.7200 1562.8400 1978.2000 ;
        RECT 1516.2400 2010.3600 1517.8400 2010.8400 ;
        RECT 1516.2400 2015.8000 1517.8400 2016.2800 ;
        RECT 1516.2400 1994.0400 1517.8400 1994.5200 ;
        RECT 1516.2400 1999.4800 1517.8400 1999.9600 ;
        RECT 1516.2400 2004.9200 1517.8400 2005.4000 ;
        RECT 1516.2400 1983.1600 1517.8400 1983.6400 ;
        RECT 1516.2400 1988.6000 1517.8400 1989.0800 ;
        RECT 1516.2400 1966.8400 1517.8400 1967.3200 ;
        RECT 1516.2400 1972.2800 1517.8400 1972.7600 ;
        RECT 1516.2400 1977.7200 1517.8400 1978.2000 ;
        RECT 1572.7800 1955.9600 1575.7800 1956.4400 ;
        RECT 1572.7800 1961.4000 1575.7800 1961.8800 ;
        RECT 1561.2400 1955.9600 1562.8400 1956.4400 ;
        RECT 1561.2400 1961.4000 1562.8400 1961.8800 ;
        RECT 1572.7800 1939.6400 1575.7800 1940.1200 ;
        RECT 1572.7800 1945.0800 1575.7800 1945.5600 ;
        RECT 1572.7800 1950.5200 1575.7800 1951.0000 ;
        RECT 1561.2400 1939.6400 1562.8400 1940.1200 ;
        RECT 1561.2400 1945.0800 1562.8400 1945.5600 ;
        RECT 1561.2400 1950.5200 1562.8400 1951.0000 ;
        RECT 1572.7800 1928.7600 1575.7800 1929.2400 ;
        RECT 1572.7800 1934.2000 1575.7800 1934.6800 ;
        RECT 1561.2400 1928.7600 1562.8400 1929.2400 ;
        RECT 1561.2400 1934.2000 1562.8400 1934.6800 ;
        RECT 1572.7800 1923.3200 1575.7800 1923.8000 ;
        RECT 1561.2400 1923.3200 1562.8400 1923.8000 ;
        RECT 1516.2400 1955.9600 1517.8400 1956.4400 ;
        RECT 1516.2400 1961.4000 1517.8400 1961.8800 ;
        RECT 1516.2400 1939.6400 1517.8400 1940.1200 ;
        RECT 1516.2400 1945.0800 1517.8400 1945.5600 ;
        RECT 1516.2400 1950.5200 1517.8400 1951.0000 ;
        RECT 1516.2400 1928.7600 1517.8400 1929.2400 ;
        RECT 1516.2400 1934.2000 1517.8400 1934.6800 ;
        RECT 1516.2400 1923.3200 1517.8400 1923.8000 ;
        RECT 1471.2400 2010.3600 1472.8400 2010.8400 ;
        RECT 1471.2400 2015.8000 1472.8400 2016.2800 ;
        RECT 1471.2400 1994.0400 1472.8400 1994.5200 ;
        RECT 1471.2400 1999.4800 1472.8400 1999.9600 ;
        RECT 1471.2400 2004.9200 1472.8400 2005.4000 ;
        RECT 1426.2400 2010.3600 1427.8400 2010.8400 ;
        RECT 1426.2400 2015.8000 1427.8400 2016.2800 ;
        RECT 1426.2400 1994.0400 1427.8400 1994.5200 ;
        RECT 1426.2400 1999.4800 1427.8400 1999.9600 ;
        RECT 1426.2400 2004.9200 1427.8400 2005.4000 ;
        RECT 1471.2400 1983.1600 1472.8400 1983.6400 ;
        RECT 1471.2400 1988.6000 1472.8400 1989.0800 ;
        RECT 1471.2400 1966.8400 1472.8400 1967.3200 ;
        RECT 1471.2400 1972.2800 1472.8400 1972.7600 ;
        RECT 1471.2400 1977.7200 1472.8400 1978.2000 ;
        RECT 1426.2400 1983.1600 1427.8400 1983.6400 ;
        RECT 1426.2400 1988.6000 1427.8400 1989.0800 ;
        RECT 1426.2400 1966.8400 1427.8400 1967.3200 ;
        RECT 1426.2400 1972.2800 1427.8400 1972.7600 ;
        RECT 1426.2400 1977.7200 1427.8400 1978.2000 ;
        RECT 1376.6800 2010.3600 1379.6800 2010.8400 ;
        RECT 1376.6800 2015.8000 1379.6800 2016.2800 ;
        RECT 1376.6800 1999.4800 1379.6800 1999.9600 ;
        RECT 1376.6800 1994.0400 1379.6800 1994.5200 ;
        RECT 1376.6800 2004.9200 1379.6800 2005.4000 ;
        RECT 1376.6800 1983.1600 1379.6800 1983.6400 ;
        RECT 1376.6800 1988.6000 1379.6800 1989.0800 ;
        RECT 1376.6800 1972.2800 1379.6800 1972.7600 ;
        RECT 1376.6800 1966.8400 1379.6800 1967.3200 ;
        RECT 1376.6800 1977.7200 1379.6800 1978.2000 ;
        RECT 1471.2400 1955.9600 1472.8400 1956.4400 ;
        RECT 1471.2400 1961.4000 1472.8400 1961.8800 ;
        RECT 1471.2400 1939.6400 1472.8400 1940.1200 ;
        RECT 1471.2400 1945.0800 1472.8400 1945.5600 ;
        RECT 1471.2400 1950.5200 1472.8400 1951.0000 ;
        RECT 1426.2400 1955.9600 1427.8400 1956.4400 ;
        RECT 1426.2400 1961.4000 1427.8400 1961.8800 ;
        RECT 1426.2400 1939.6400 1427.8400 1940.1200 ;
        RECT 1426.2400 1945.0800 1427.8400 1945.5600 ;
        RECT 1426.2400 1950.5200 1427.8400 1951.0000 ;
        RECT 1471.2400 1934.2000 1472.8400 1934.6800 ;
        RECT 1471.2400 1928.7600 1472.8400 1929.2400 ;
        RECT 1471.2400 1923.3200 1472.8400 1923.8000 ;
        RECT 1426.2400 1934.2000 1427.8400 1934.6800 ;
        RECT 1426.2400 1928.7600 1427.8400 1929.2400 ;
        RECT 1426.2400 1923.3200 1427.8400 1923.8000 ;
        RECT 1376.6800 1955.9600 1379.6800 1956.4400 ;
        RECT 1376.6800 1961.4000 1379.6800 1961.8800 ;
        RECT 1376.6800 1945.0800 1379.6800 1945.5600 ;
        RECT 1376.6800 1939.6400 1379.6800 1940.1200 ;
        RECT 1376.6800 1950.5200 1379.6800 1951.0000 ;
        RECT 1376.6800 1928.7600 1379.6800 1929.2400 ;
        RECT 1376.6800 1934.2000 1379.6800 1934.6800 ;
        RECT 1376.6800 1923.3200 1379.6800 1923.8000 ;
        RECT 1376.6800 2121.5100 1575.7800 2124.5100 ;
        RECT 1376.6800 1916.4100 1575.7800 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 1686.7700 1562.8400 1894.8700 ;
        RECT 1516.2400 1686.7700 1517.8400 1894.8700 ;
        RECT 1471.2400 1686.7700 1472.8400 1894.8700 ;
        RECT 1426.2400 1686.7700 1427.8400 1894.8700 ;
        RECT 1572.7800 1686.7700 1575.7800 1894.8700 ;
        RECT 1376.6800 1686.7700 1379.6800 1894.8700 ;
      LAYER met3 ;
        RECT 1572.7800 1889.5200 1575.7800 1890.0000 ;
        RECT 1561.2400 1889.5200 1562.8400 1890.0000 ;
        RECT 1572.7800 1878.6400 1575.7800 1879.1200 ;
        RECT 1572.7800 1884.0800 1575.7800 1884.5600 ;
        RECT 1561.2400 1878.6400 1562.8400 1879.1200 ;
        RECT 1561.2400 1884.0800 1562.8400 1884.5600 ;
        RECT 1572.7800 1862.3200 1575.7800 1862.8000 ;
        RECT 1572.7800 1867.7600 1575.7800 1868.2400 ;
        RECT 1561.2400 1862.3200 1562.8400 1862.8000 ;
        RECT 1561.2400 1867.7600 1562.8400 1868.2400 ;
        RECT 1572.7800 1851.4400 1575.7800 1851.9200 ;
        RECT 1572.7800 1856.8800 1575.7800 1857.3600 ;
        RECT 1561.2400 1851.4400 1562.8400 1851.9200 ;
        RECT 1561.2400 1856.8800 1562.8400 1857.3600 ;
        RECT 1572.7800 1873.2000 1575.7800 1873.6800 ;
        RECT 1561.2400 1873.2000 1562.8400 1873.6800 ;
        RECT 1516.2400 1878.6400 1517.8400 1879.1200 ;
        RECT 1516.2400 1884.0800 1517.8400 1884.5600 ;
        RECT 1516.2400 1889.5200 1517.8400 1890.0000 ;
        RECT 1516.2400 1862.3200 1517.8400 1862.8000 ;
        RECT 1516.2400 1867.7600 1517.8400 1868.2400 ;
        RECT 1516.2400 1856.8800 1517.8400 1857.3600 ;
        RECT 1516.2400 1851.4400 1517.8400 1851.9200 ;
        RECT 1516.2400 1873.2000 1517.8400 1873.6800 ;
        RECT 1572.7800 1835.1200 1575.7800 1835.6000 ;
        RECT 1572.7800 1840.5600 1575.7800 1841.0400 ;
        RECT 1561.2400 1835.1200 1562.8400 1835.6000 ;
        RECT 1561.2400 1840.5600 1562.8400 1841.0400 ;
        RECT 1572.7800 1818.8000 1575.7800 1819.2800 ;
        RECT 1572.7800 1824.2400 1575.7800 1824.7200 ;
        RECT 1572.7800 1829.6800 1575.7800 1830.1600 ;
        RECT 1561.2400 1818.8000 1562.8400 1819.2800 ;
        RECT 1561.2400 1824.2400 1562.8400 1824.7200 ;
        RECT 1561.2400 1829.6800 1562.8400 1830.1600 ;
        RECT 1572.7800 1807.9200 1575.7800 1808.4000 ;
        RECT 1572.7800 1813.3600 1575.7800 1813.8400 ;
        RECT 1561.2400 1807.9200 1562.8400 1808.4000 ;
        RECT 1561.2400 1813.3600 1562.8400 1813.8400 ;
        RECT 1572.7800 1791.6000 1575.7800 1792.0800 ;
        RECT 1572.7800 1797.0400 1575.7800 1797.5200 ;
        RECT 1572.7800 1802.4800 1575.7800 1802.9600 ;
        RECT 1561.2400 1791.6000 1562.8400 1792.0800 ;
        RECT 1561.2400 1797.0400 1562.8400 1797.5200 ;
        RECT 1561.2400 1802.4800 1562.8400 1802.9600 ;
        RECT 1516.2400 1835.1200 1517.8400 1835.6000 ;
        RECT 1516.2400 1840.5600 1517.8400 1841.0400 ;
        RECT 1516.2400 1818.8000 1517.8400 1819.2800 ;
        RECT 1516.2400 1824.2400 1517.8400 1824.7200 ;
        RECT 1516.2400 1829.6800 1517.8400 1830.1600 ;
        RECT 1516.2400 1807.9200 1517.8400 1808.4000 ;
        RECT 1516.2400 1813.3600 1517.8400 1813.8400 ;
        RECT 1516.2400 1791.6000 1517.8400 1792.0800 ;
        RECT 1516.2400 1797.0400 1517.8400 1797.5200 ;
        RECT 1516.2400 1802.4800 1517.8400 1802.9600 ;
        RECT 1572.7800 1846.0000 1575.7800 1846.4800 ;
        RECT 1516.2400 1846.0000 1517.8400 1846.4800 ;
        RECT 1561.2400 1846.0000 1562.8400 1846.4800 ;
        RECT 1471.2400 1878.6400 1472.8400 1879.1200 ;
        RECT 1471.2400 1884.0800 1472.8400 1884.5600 ;
        RECT 1471.2400 1889.5200 1472.8400 1890.0000 ;
        RECT 1426.2400 1878.6400 1427.8400 1879.1200 ;
        RECT 1426.2400 1884.0800 1427.8400 1884.5600 ;
        RECT 1426.2400 1889.5200 1427.8400 1890.0000 ;
        RECT 1471.2400 1862.3200 1472.8400 1862.8000 ;
        RECT 1471.2400 1867.7600 1472.8400 1868.2400 ;
        RECT 1471.2400 1851.4400 1472.8400 1851.9200 ;
        RECT 1471.2400 1856.8800 1472.8400 1857.3600 ;
        RECT 1426.2400 1862.3200 1427.8400 1862.8000 ;
        RECT 1426.2400 1867.7600 1427.8400 1868.2400 ;
        RECT 1426.2400 1851.4400 1427.8400 1851.9200 ;
        RECT 1426.2400 1856.8800 1427.8400 1857.3600 ;
        RECT 1426.2400 1873.2000 1427.8400 1873.6800 ;
        RECT 1471.2400 1873.2000 1472.8400 1873.6800 ;
        RECT 1376.6800 1889.5200 1379.6800 1890.0000 ;
        RECT 1376.6800 1884.0800 1379.6800 1884.5600 ;
        RECT 1376.6800 1878.6400 1379.6800 1879.1200 ;
        RECT 1376.6800 1867.7600 1379.6800 1868.2400 ;
        RECT 1376.6800 1862.3200 1379.6800 1862.8000 ;
        RECT 1376.6800 1856.8800 1379.6800 1857.3600 ;
        RECT 1376.6800 1851.4400 1379.6800 1851.9200 ;
        RECT 1376.6800 1873.2000 1379.6800 1873.6800 ;
        RECT 1471.2400 1835.1200 1472.8400 1835.6000 ;
        RECT 1471.2400 1840.5600 1472.8400 1841.0400 ;
        RECT 1471.2400 1818.8000 1472.8400 1819.2800 ;
        RECT 1471.2400 1824.2400 1472.8400 1824.7200 ;
        RECT 1471.2400 1829.6800 1472.8400 1830.1600 ;
        RECT 1426.2400 1835.1200 1427.8400 1835.6000 ;
        RECT 1426.2400 1840.5600 1427.8400 1841.0400 ;
        RECT 1426.2400 1818.8000 1427.8400 1819.2800 ;
        RECT 1426.2400 1824.2400 1427.8400 1824.7200 ;
        RECT 1426.2400 1829.6800 1427.8400 1830.1600 ;
        RECT 1471.2400 1807.9200 1472.8400 1808.4000 ;
        RECT 1471.2400 1813.3600 1472.8400 1813.8400 ;
        RECT 1471.2400 1791.6000 1472.8400 1792.0800 ;
        RECT 1471.2400 1797.0400 1472.8400 1797.5200 ;
        RECT 1471.2400 1802.4800 1472.8400 1802.9600 ;
        RECT 1426.2400 1807.9200 1427.8400 1808.4000 ;
        RECT 1426.2400 1813.3600 1427.8400 1813.8400 ;
        RECT 1426.2400 1791.6000 1427.8400 1792.0800 ;
        RECT 1426.2400 1797.0400 1427.8400 1797.5200 ;
        RECT 1426.2400 1802.4800 1427.8400 1802.9600 ;
        RECT 1376.6800 1835.1200 1379.6800 1835.6000 ;
        RECT 1376.6800 1840.5600 1379.6800 1841.0400 ;
        RECT 1376.6800 1824.2400 1379.6800 1824.7200 ;
        RECT 1376.6800 1818.8000 1379.6800 1819.2800 ;
        RECT 1376.6800 1829.6800 1379.6800 1830.1600 ;
        RECT 1376.6800 1807.9200 1379.6800 1808.4000 ;
        RECT 1376.6800 1813.3600 1379.6800 1813.8400 ;
        RECT 1376.6800 1797.0400 1379.6800 1797.5200 ;
        RECT 1376.6800 1791.6000 1379.6800 1792.0800 ;
        RECT 1376.6800 1802.4800 1379.6800 1802.9600 ;
        RECT 1376.6800 1846.0000 1379.6800 1846.4800 ;
        RECT 1426.2400 1846.0000 1427.8400 1846.4800 ;
        RECT 1471.2400 1846.0000 1472.8400 1846.4800 ;
        RECT 1572.7800 1780.7200 1575.7800 1781.2000 ;
        RECT 1572.7800 1786.1600 1575.7800 1786.6400 ;
        RECT 1561.2400 1780.7200 1562.8400 1781.2000 ;
        RECT 1561.2400 1786.1600 1562.8400 1786.6400 ;
        RECT 1572.7800 1764.4000 1575.7800 1764.8800 ;
        RECT 1572.7800 1769.8400 1575.7800 1770.3200 ;
        RECT 1572.7800 1775.2800 1575.7800 1775.7600 ;
        RECT 1561.2400 1764.4000 1562.8400 1764.8800 ;
        RECT 1561.2400 1769.8400 1562.8400 1770.3200 ;
        RECT 1561.2400 1775.2800 1562.8400 1775.7600 ;
        RECT 1572.7800 1753.5200 1575.7800 1754.0000 ;
        RECT 1572.7800 1758.9600 1575.7800 1759.4400 ;
        RECT 1561.2400 1753.5200 1562.8400 1754.0000 ;
        RECT 1561.2400 1758.9600 1562.8400 1759.4400 ;
        RECT 1572.7800 1737.2000 1575.7800 1737.6800 ;
        RECT 1572.7800 1742.6400 1575.7800 1743.1200 ;
        RECT 1572.7800 1748.0800 1575.7800 1748.5600 ;
        RECT 1561.2400 1737.2000 1562.8400 1737.6800 ;
        RECT 1561.2400 1742.6400 1562.8400 1743.1200 ;
        RECT 1561.2400 1748.0800 1562.8400 1748.5600 ;
        RECT 1516.2400 1780.7200 1517.8400 1781.2000 ;
        RECT 1516.2400 1786.1600 1517.8400 1786.6400 ;
        RECT 1516.2400 1764.4000 1517.8400 1764.8800 ;
        RECT 1516.2400 1769.8400 1517.8400 1770.3200 ;
        RECT 1516.2400 1775.2800 1517.8400 1775.7600 ;
        RECT 1516.2400 1753.5200 1517.8400 1754.0000 ;
        RECT 1516.2400 1758.9600 1517.8400 1759.4400 ;
        RECT 1516.2400 1737.2000 1517.8400 1737.6800 ;
        RECT 1516.2400 1742.6400 1517.8400 1743.1200 ;
        RECT 1516.2400 1748.0800 1517.8400 1748.5600 ;
        RECT 1572.7800 1726.3200 1575.7800 1726.8000 ;
        RECT 1572.7800 1731.7600 1575.7800 1732.2400 ;
        RECT 1561.2400 1726.3200 1562.8400 1726.8000 ;
        RECT 1561.2400 1731.7600 1562.8400 1732.2400 ;
        RECT 1572.7800 1710.0000 1575.7800 1710.4800 ;
        RECT 1572.7800 1715.4400 1575.7800 1715.9200 ;
        RECT 1572.7800 1720.8800 1575.7800 1721.3600 ;
        RECT 1561.2400 1710.0000 1562.8400 1710.4800 ;
        RECT 1561.2400 1715.4400 1562.8400 1715.9200 ;
        RECT 1561.2400 1720.8800 1562.8400 1721.3600 ;
        RECT 1572.7800 1699.1200 1575.7800 1699.6000 ;
        RECT 1572.7800 1704.5600 1575.7800 1705.0400 ;
        RECT 1561.2400 1699.1200 1562.8400 1699.6000 ;
        RECT 1561.2400 1704.5600 1562.8400 1705.0400 ;
        RECT 1572.7800 1693.6800 1575.7800 1694.1600 ;
        RECT 1561.2400 1693.6800 1562.8400 1694.1600 ;
        RECT 1516.2400 1726.3200 1517.8400 1726.8000 ;
        RECT 1516.2400 1731.7600 1517.8400 1732.2400 ;
        RECT 1516.2400 1710.0000 1517.8400 1710.4800 ;
        RECT 1516.2400 1715.4400 1517.8400 1715.9200 ;
        RECT 1516.2400 1720.8800 1517.8400 1721.3600 ;
        RECT 1516.2400 1699.1200 1517.8400 1699.6000 ;
        RECT 1516.2400 1704.5600 1517.8400 1705.0400 ;
        RECT 1516.2400 1693.6800 1517.8400 1694.1600 ;
        RECT 1471.2400 1780.7200 1472.8400 1781.2000 ;
        RECT 1471.2400 1786.1600 1472.8400 1786.6400 ;
        RECT 1471.2400 1764.4000 1472.8400 1764.8800 ;
        RECT 1471.2400 1769.8400 1472.8400 1770.3200 ;
        RECT 1471.2400 1775.2800 1472.8400 1775.7600 ;
        RECT 1426.2400 1780.7200 1427.8400 1781.2000 ;
        RECT 1426.2400 1786.1600 1427.8400 1786.6400 ;
        RECT 1426.2400 1764.4000 1427.8400 1764.8800 ;
        RECT 1426.2400 1769.8400 1427.8400 1770.3200 ;
        RECT 1426.2400 1775.2800 1427.8400 1775.7600 ;
        RECT 1471.2400 1753.5200 1472.8400 1754.0000 ;
        RECT 1471.2400 1758.9600 1472.8400 1759.4400 ;
        RECT 1471.2400 1737.2000 1472.8400 1737.6800 ;
        RECT 1471.2400 1742.6400 1472.8400 1743.1200 ;
        RECT 1471.2400 1748.0800 1472.8400 1748.5600 ;
        RECT 1426.2400 1753.5200 1427.8400 1754.0000 ;
        RECT 1426.2400 1758.9600 1427.8400 1759.4400 ;
        RECT 1426.2400 1737.2000 1427.8400 1737.6800 ;
        RECT 1426.2400 1742.6400 1427.8400 1743.1200 ;
        RECT 1426.2400 1748.0800 1427.8400 1748.5600 ;
        RECT 1376.6800 1780.7200 1379.6800 1781.2000 ;
        RECT 1376.6800 1786.1600 1379.6800 1786.6400 ;
        RECT 1376.6800 1769.8400 1379.6800 1770.3200 ;
        RECT 1376.6800 1764.4000 1379.6800 1764.8800 ;
        RECT 1376.6800 1775.2800 1379.6800 1775.7600 ;
        RECT 1376.6800 1753.5200 1379.6800 1754.0000 ;
        RECT 1376.6800 1758.9600 1379.6800 1759.4400 ;
        RECT 1376.6800 1742.6400 1379.6800 1743.1200 ;
        RECT 1376.6800 1737.2000 1379.6800 1737.6800 ;
        RECT 1376.6800 1748.0800 1379.6800 1748.5600 ;
        RECT 1471.2400 1726.3200 1472.8400 1726.8000 ;
        RECT 1471.2400 1731.7600 1472.8400 1732.2400 ;
        RECT 1471.2400 1710.0000 1472.8400 1710.4800 ;
        RECT 1471.2400 1715.4400 1472.8400 1715.9200 ;
        RECT 1471.2400 1720.8800 1472.8400 1721.3600 ;
        RECT 1426.2400 1726.3200 1427.8400 1726.8000 ;
        RECT 1426.2400 1731.7600 1427.8400 1732.2400 ;
        RECT 1426.2400 1710.0000 1427.8400 1710.4800 ;
        RECT 1426.2400 1715.4400 1427.8400 1715.9200 ;
        RECT 1426.2400 1720.8800 1427.8400 1721.3600 ;
        RECT 1471.2400 1704.5600 1472.8400 1705.0400 ;
        RECT 1471.2400 1699.1200 1472.8400 1699.6000 ;
        RECT 1471.2400 1693.6800 1472.8400 1694.1600 ;
        RECT 1426.2400 1704.5600 1427.8400 1705.0400 ;
        RECT 1426.2400 1699.1200 1427.8400 1699.6000 ;
        RECT 1426.2400 1693.6800 1427.8400 1694.1600 ;
        RECT 1376.6800 1726.3200 1379.6800 1726.8000 ;
        RECT 1376.6800 1731.7600 1379.6800 1732.2400 ;
        RECT 1376.6800 1715.4400 1379.6800 1715.9200 ;
        RECT 1376.6800 1710.0000 1379.6800 1710.4800 ;
        RECT 1376.6800 1720.8800 1379.6800 1721.3600 ;
        RECT 1376.6800 1699.1200 1379.6800 1699.6000 ;
        RECT 1376.6800 1704.5600 1379.6800 1705.0400 ;
        RECT 1376.6800 1693.6800 1379.6800 1694.1600 ;
        RECT 1376.6800 1891.8700 1575.7800 1894.8700 ;
        RECT 1376.6800 1686.7700 1575.7800 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 1457.1300 1562.8400 1665.2300 ;
        RECT 1516.2400 1457.1300 1517.8400 1665.2300 ;
        RECT 1471.2400 1457.1300 1472.8400 1665.2300 ;
        RECT 1426.2400 1457.1300 1427.8400 1665.2300 ;
        RECT 1572.7800 1457.1300 1575.7800 1665.2300 ;
        RECT 1376.6800 1457.1300 1379.6800 1665.2300 ;
      LAYER met3 ;
        RECT 1572.7800 1659.8800 1575.7800 1660.3600 ;
        RECT 1561.2400 1659.8800 1562.8400 1660.3600 ;
        RECT 1572.7800 1649.0000 1575.7800 1649.4800 ;
        RECT 1572.7800 1654.4400 1575.7800 1654.9200 ;
        RECT 1561.2400 1649.0000 1562.8400 1649.4800 ;
        RECT 1561.2400 1654.4400 1562.8400 1654.9200 ;
        RECT 1572.7800 1632.6800 1575.7800 1633.1600 ;
        RECT 1572.7800 1638.1200 1575.7800 1638.6000 ;
        RECT 1561.2400 1632.6800 1562.8400 1633.1600 ;
        RECT 1561.2400 1638.1200 1562.8400 1638.6000 ;
        RECT 1572.7800 1621.8000 1575.7800 1622.2800 ;
        RECT 1572.7800 1627.2400 1575.7800 1627.7200 ;
        RECT 1561.2400 1621.8000 1562.8400 1622.2800 ;
        RECT 1561.2400 1627.2400 1562.8400 1627.7200 ;
        RECT 1572.7800 1643.5600 1575.7800 1644.0400 ;
        RECT 1561.2400 1643.5600 1562.8400 1644.0400 ;
        RECT 1516.2400 1649.0000 1517.8400 1649.4800 ;
        RECT 1516.2400 1654.4400 1517.8400 1654.9200 ;
        RECT 1516.2400 1659.8800 1517.8400 1660.3600 ;
        RECT 1516.2400 1632.6800 1517.8400 1633.1600 ;
        RECT 1516.2400 1638.1200 1517.8400 1638.6000 ;
        RECT 1516.2400 1627.2400 1517.8400 1627.7200 ;
        RECT 1516.2400 1621.8000 1517.8400 1622.2800 ;
        RECT 1516.2400 1643.5600 1517.8400 1644.0400 ;
        RECT 1572.7800 1605.4800 1575.7800 1605.9600 ;
        RECT 1572.7800 1610.9200 1575.7800 1611.4000 ;
        RECT 1561.2400 1605.4800 1562.8400 1605.9600 ;
        RECT 1561.2400 1610.9200 1562.8400 1611.4000 ;
        RECT 1572.7800 1589.1600 1575.7800 1589.6400 ;
        RECT 1572.7800 1594.6000 1575.7800 1595.0800 ;
        RECT 1572.7800 1600.0400 1575.7800 1600.5200 ;
        RECT 1561.2400 1589.1600 1562.8400 1589.6400 ;
        RECT 1561.2400 1594.6000 1562.8400 1595.0800 ;
        RECT 1561.2400 1600.0400 1562.8400 1600.5200 ;
        RECT 1572.7800 1578.2800 1575.7800 1578.7600 ;
        RECT 1572.7800 1583.7200 1575.7800 1584.2000 ;
        RECT 1561.2400 1578.2800 1562.8400 1578.7600 ;
        RECT 1561.2400 1583.7200 1562.8400 1584.2000 ;
        RECT 1572.7800 1561.9600 1575.7800 1562.4400 ;
        RECT 1572.7800 1567.4000 1575.7800 1567.8800 ;
        RECT 1572.7800 1572.8400 1575.7800 1573.3200 ;
        RECT 1561.2400 1561.9600 1562.8400 1562.4400 ;
        RECT 1561.2400 1567.4000 1562.8400 1567.8800 ;
        RECT 1561.2400 1572.8400 1562.8400 1573.3200 ;
        RECT 1516.2400 1605.4800 1517.8400 1605.9600 ;
        RECT 1516.2400 1610.9200 1517.8400 1611.4000 ;
        RECT 1516.2400 1589.1600 1517.8400 1589.6400 ;
        RECT 1516.2400 1594.6000 1517.8400 1595.0800 ;
        RECT 1516.2400 1600.0400 1517.8400 1600.5200 ;
        RECT 1516.2400 1578.2800 1517.8400 1578.7600 ;
        RECT 1516.2400 1583.7200 1517.8400 1584.2000 ;
        RECT 1516.2400 1561.9600 1517.8400 1562.4400 ;
        RECT 1516.2400 1567.4000 1517.8400 1567.8800 ;
        RECT 1516.2400 1572.8400 1517.8400 1573.3200 ;
        RECT 1572.7800 1616.3600 1575.7800 1616.8400 ;
        RECT 1516.2400 1616.3600 1517.8400 1616.8400 ;
        RECT 1561.2400 1616.3600 1562.8400 1616.8400 ;
        RECT 1471.2400 1649.0000 1472.8400 1649.4800 ;
        RECT 1471.2400 1654.4400 1472.8400 1654.9200 ;
        RECT 1471.2400 1659.8800 1472.8400 1660.3600 ;
        RECT 1426.2400 1649.0000 1427.8400 1649.4800 ;
        RECT 1426.2400 1654.4400 1427.8400 1654.9200 ;
        RECT 1426.2400 1659.8800 1427.8400 1660.3600 ;
        RECT 1471.2400 1632.6800 1472.8400 1633.1600 ;
        RECT 1471.2400 1638.1200 1472.8400 1638.6000 ;
        RECT 1471.2400 1621.8000 1472.8400 1622.2800 ;
        RECT 1471.2400 1627.2400 1472.8400 1627.7200 ;
        RECT 1426.2400 1632.6800 1427.8400 1633.1600 ;
        RECT 1426.2400 1638.1200 1427.8400 1638.6000 ;
        RECT 1426.2400 1621.8000 1427.8400 1622.2800 ;
        RECT 1426.2400 1627.2400 1427.8400 1627.7200 ;
        RECT 1426.2400 1643.5600 1427.8400 1644.0400 ;
        RECT 1471.2400 1643.5600 1472.8400 1644.0400 ;
        RECT 1376.6800 1659.8800 1379.6800 1660.3600 ;
        RECT 1376.6800 1654.4400 1379.6800 1654.9200 ;
        RECT 1376.6800 1649.0000 1379.6800 1649.4800 ;
        RECT 1376.6800 1638.1200 1379.6800 1638.6000 ;
        RECT 1376.6800 1632.6800 1379.6800 1633.1600 ;
        RECT 1376.6800 1627.2400 1379.6800 1627.7200 ;
        RECT 1376.6800 1621.8000 1379.6800 1622.2800 ;
        RECT 1376.6800 1643.5600 1379.6800 1644.0400 ;
        RECT 1471.2400 1605.4800 1472.8400 1605.9600 ;
        RECT 1471.2400 1610.9200 1472.8400 1611.4000 ;
        RECT 1471.2400 1589.1600 1472.8400 1589.6400 ;
        RECT 1471.2400 1594.6000 1472.8400 1595.0800 ;
        RECT 1471.2400 1600.0400 1472.8400 1600.5200 ;
        RECT 1426.2400 1605.4800 1427.8400 1605.9600 ;
        RECT 1426.2400 1610.9200 1427.8400 1611.4000 ;
        RECT 1426.2400 1589.1600 1427.8400 1589.6400 ;
        RECT 1426.2400 1594.6000 1427.8400 1595.0800 ;
        RECT 1426.2400 1600.0400 1427.8400 1600.5200 ;
        RECT 1471.2400 1578.2800 1472.8400 1578.7600 ;
        RECT 1471.2400 1583.7200 1472.8400 1584.2000 ;
        RECT 1471.2400 1561.9600 1472.8400 1562.4400 ;
        RECT 1471.2400 1567.4000 1472.8400 1567.8800 ;
        RECT 1471.2400 1572.8400 1472.8400 1573.3200 ;
        RECT 1426.2400 1578.2800 1427.8400 1578.7600 ;
        RECT 1426.2400 1583.7200 1427.8400 1584.2000 ;
        RECT 1426.2400 1561.9600 1427.8400 1562.4400 ;
        RECT 1426.2400 1567.4000 1427.8400 1567.8800 ;
        RECT 1426.2400 1572.8400 1427.8400 1573.3200 ;
        RECT 1376.6800 1605.4800 1379.6800 1605.9600 ;
        RECT 1376.6800 1610.9200 1379.6800 1611.4000 ;
        RECT 1376.6800 1594.6000 1379.6800 1595.0800 ;
        RECT 1376.6800 1589.1600 1379.6800 1589.6400 ;
        RECT 1376.6800 1600.0400 1379.6800 1600.5200 ;
        RECT 1376.6800 1578.2800 1379.6800 1578.7600 ;
        RECT 1376.6800 1583.7200 1379.6800 1584.2000 ;
        RECT 1376.6800 1567.4000 1379.6800 1567.8800 ;
        RECT 1376.6800 1561.9600 1379.6800 1562.4400 ;
        RECT 1376.6800 1572.8400 1379.6800 1573.3200 ;
        RECT 1376.6800 1616.3600 1379.6800 1616.8400 ;
        RECT 1426.2400 1616.3600 1427.8400 1616.8400 ;
        RECT 1471.2400 1616.3600 1472.8400 1616.8400 ;
        RECT 1572.7800 1551.0800 1575.7800 1551.5600 ;
        RECT 1572.7800 1556.5200 1575.7800 1557.0000 ;
        RECT 1561.2400 1551.0800 1562.8400 1551.5600 ;
        RECT 1561.2400 1556.5200 1562.8400 1557.0000 ;
        RECT 1572.7800 1534.7600 1575.7800 1535.2400 ;
        RECT 1572.7800 1540.2000 1575.7800 1540.6800 ;
        RECT 1572.7800 1545.6400 1575.7800 1546.1200 ;
        RECT 1561.2400 1534.7600 1562.8400 1535.2400 ;
        RECT 1561.2400 1540.2000 1562.8400 1540.6800 ;
        RECT 1561.2400 1545.6400 1562.8400 1546.1200 ;
        RECT 1572.7800 1523.8800 1575.7800 1524.3600 ;
        RECT 1572.7800 1529.3200 1575.7800 1529.8000 ;
        RECT 1561.2400 1523.8800 1562.8400 1524.3600 ;
        RECT 1561.2400 1529.3200 1562.8400 1529.8000 ;
        RECT 1572.7800 1507.5600 1575.7800 1508.0400 ;
        RECT 1572.7800 1513.0000 1575.7800 1513.4800 ;
        RECT 1572.7800 1518.4400 1575.7800 1518.9200 ;
        RECT 1561.2400 1507.5600 1562.8400 1508.0400 ;
        RECT 1561.2400 1513.0000 1562.8400 1513.4800 ;
        RECT 1561.2400 1518.4400 1562.8400 1518.9200 ;
        RECT 1516.2400 1551.0800 1517.8400 1551.5600 ;
        RECT 1516.2400 1556.5200 1517.8400 1557.0000 ;
        RECT 1516.2400 1534.7600 1517.8400 1535.2400 ;
        RECT 1516.2400 1540.2000 1517.8400 1540.6800 ;
        RECT 1516.2400 1545.6400 1517.8400 1546.1200 ;
        RECT 1516.2400 1523.8800 1517.8400 1524.3600 ;
        RECT 1516.2400 1529.3200 1517.8400 1529.8000 ;
        RECT 1516.2400 1507.5600 1517.8400 1508.0400 ;
        RECT 1516.2400 1513.0000 1517.8400 1513.4800 ;
        RECT 1516.2400 1518.4400 1517.8400 1518.9200 ;
        RECT 1572.7800 1496.6800 1575.7800 1497.1600 ;
        RECT 1572.7800 1502.1200 1575.7800 1502.6000 ;
        RECT 1561.2400 1496.6800 1562.8400 1497.1600 ;
        RECT 1561.2400 1502.1200 1562.8400 1502.6000 ;
        RECT 1572.7800 1480.3600 1575.7800 1480.8400 ;
        RECT 1572.7800 1485.8000 1575.7800 1486.2800 ;
        RECT 1572.7800 1491.2400 1575.7800 1491.7200 ;
        RECT 1561.2400 1480.3600 1562.8400 1480.8400 ;
        RECT 1561.2400 1485.8000 1562.8400 1486.2800 ;
        RECT 1561.2400 1491.2400 1562.8400 1491.7200 ;
        RECT 1572.7800 1469.4800 1575.7800 1469.9600 ;
        RECT 1572.7800 1474.9200 1575.7800 1475.4000 ;
        RECT 1561.2400 1469.4800 1562.8400 1469.9600 ;
        RECT 1561.2400 1474.9200 1562.8400 1475.4000 ;
        RECT 1572.7800 1464.0400 1575.7800 1464.5200 ;
        RECT 1561.2400 1464.0400 1562.8400 1464.5200 ;
        RECT 1516.2400 1496.6800 1517.8400 1497.1600 ;
        RECT 1516.2400 1502.1200 1517.8400 1502.6000 ;
        RECT 1516.2400 1480.3600 1517.8400 1480.8400 ;
        RECT 1516.2400 1485.8000 1517.8400 1486.2800 ;
        RECT 1516.2400 1491.2400 1517.8400 1491.7200 ;
        RECT 1516.2400 1469.4800 1517.8400 1469.9600 ;
        RECT 1516.2400 1474.9200 1517.8400 1475.4000 ;
        RECT 1516.2400 1464.0400 1517.8400 1464.5200 ;
        RECT 1471.2400 1551.0800 1472.8400 1551.5600 ;
        RECT 1471.2400 1556.5200 1472.8400 1557.0000 ;
        RECT 1471.2400 1534.7600 1472.8400 1535.2400 ;
        RECT 1471.2400 1540.2000 1472.8400 1540.6800 ;
        RECT 1471.2400 1545.6400 1472.8400 1546.1200 ;
        RECT 1426.2400 1551.0800 1427.8400 1551.5600 ;
        RECT 1426.2400 1556.5200 1427.8400 1557.0000 ;
        RECT 1426.2400 1534.7600 1427.8400 1535.2400 ;
        RECT 1426.2400 1540.2000 1427.8400 1540.6800 ;
        RECT 1426.2400 1545.6400 1427.8400 1546.1200 ;
        RECT 1471.2400 1523.8800 1472.8400 1524.3600 ;
        RECT 1471.2400 1529.3200 1472.8400 1529.8000 ;
        RECT 1471.2400 1507.5600 1472.8400 1508.0400 ;
        RECT 1471.2400 1513.0000 1472.8400 1513.4800 ;
        RECT 1471.2400 1518.4400 1472.8400 1518.9200 ;
        RECT 1426.2400 1523.8800 1427.8400 1524.3600 ;
        RECT 1426.2400 1529.3200 1427.8400 1529.8000 ;
        RECT 1426.2400 1507.5600 1427.8400 1508.0400 ;
        RECT 1426.2400 1513.0000 1427.8400 1513.4800 ;
        RECT 1426.2400 1518.4400 1427.8400 1518.9200 ;
        RECT 1376.6800 1551.0800 1379.6800 1551.5600 ;
        RECT 1376.6800 1556.5200 1379.6800 1557.0000 ;
        RECT 1376.6800 1540.2000 1379.6800 1540.6800 ;
        RECT 1376.6800 1534.7600 1379.6800 1535.2400 ;
        RECT 1376.6800 1545.6400 1379.6800 1546.1200 ;
        RECT 1376.6800 1523.8800 1379.6800 1524.3600 ;
        RECT 1376.6800 1529.3200 1379.6800 1529.8000 ;
        RECT 1376.6800 1513.0000 1379.6800 1513.4800 ;
        RECT 1376.6800 1507.5600 1379.6800 1508.0400 ;
        RECT 1376.6800 1518.4400 1379.6800 1518.9200 ;
        RECT 1471.2400 1496.6800 1472.8400 1497.1600 ;
        RECT 1471.2400 1502.1200 1472.8400 1502.6000 ;
        RECT 1471.2400 1480.3600 1472.8400 1480.8400 ;
        RECT 1471.2400 1485.8000 1472.8400 1486.2800 ;
        RECT 1471.2400 1491.2400 1472.8400 1491.7200 ;
        RECT 1426.2400 1496.6800 1427.8400 1497.1600 ;
        RECT 1426.2400 1502.1200 1427.8400 1502.6000 ;
        RECT 1426.2400 1480.3600 1427.8400 1480.8400 ;
        RECT 1426.2400 1485.8000 1427.8400 1486.2800 ;
        RECT 1426.2400 1491.2400 1427.8400 1491.7200 ;
        RECT 1471.2400 1474.9200 1472.8400 1475.4000 ;
        RECT 1471.2400 1469.4800 1472.8400 1469.9600 ;
        RECT 1471.2400 1464.0400 1472.8400 1464.5200 ;
        RECT 1426.2400 1474.9200 1427.8400 1475.4000 ;
        RECT 1426.2400 1469.4800 1427.8400 1469.9600 ;
        RECT 1426.2400 1464.0400 1427.8400 1464.5200 ;
        RECT 1376.6800 1496.6800 1379.6800 1497.1600 ;
        RECT 1376.6800 1502.1200 1379.6800 1502.6000 ;
        RECT 1376.6800 1485.8000 1379.6800 1486.2800 ;
        RECT 1376.6800 1480.3600 1379.6800 1480.8400 ;
        RECT 1376.6800 1491.2400 1379.6800 1491.7200 ;
        RECT 1376.6800 1469.4800 1379.6800 1469.9600 ;
        RECT 1376.6800 1474.9200 1379.6800 1475.4000 ;
        RECT 1376.6800 1464.0400 1379.6800 1464.5200 ;
        RECT 1376.6800 1662.2300 1575.7800 1665.2300 ;
        RECT 1376.6800 1457.1300 1575.7800 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 1227.4900 1562.8400 1435.5900 ;
        RECT 1516.2400 1227.4900 1517.8400 1435.5900 ;
        RECT 1471.2400 1227.4900 1472.8400 1435.5900 ;
        RECT 1426.2400 1227.4900 1427.8400 1435.5900 ;
        RECT 1572.7800 1227.4900 1575.7800 1435.5900 ;
        RECT 1376.6800 1227.4900 1379.6800 1435.5900 ;
      LAYER met3 ;
        RECT 1572.7800 1430.2400 1575.7800 1430.7200 ;
        RECT 1561.2400 1430.2400 1562.8400 1430.7200 ;
        RECT 1572.7800 1419.3600 1575.7800 1419.8400 ;
        RECT 1572.7800 1424.8000 1575.7800 1425.2800 ;
        RECT 1561.2400 1419.3600 1562.8400 1419.8400 ;
        RECT 1561.2400 1424.8000 1562.8400 1425.2800 ;
        RECT 1572.7800 1403.0400 1575.7800 1403.5200 ;
        RECT 1572.7800 1408.4800 1575.7800 1408.9600 ;
        RECT 1561.2400 1403.0400 1562.8400 1403.5200 ;
        RECT 1561.2400 1408.4800 1562.8400 1408.9600 ;
        RECT 1572.7800 1392.1600 1575.7800 1392.6400 ;
        RECT 1572.7800 1397.6000 1575.7800 1398.0800 ;
        RECT 1561.2400 1392.1600 1562.8400 1392.6400 ;
        RECT 1561.2400 1397.6000 1562.8400 1398.0800 ;
        RECT 1572.7800 1413.9200 1575.7800 1414.4000 ;
        RECT 1561.2400 1413.9200 1562.8400 1414.4000 ;
        RECT 1516.2400 1419.3600 1517.8400 1419.8400 ;
        RECT 1516.2400 1424.8000 1517.8400 1425.2800 ;
        RECT 1516.2400 1430.2400 1517.8400 1430.7200 ;
        RECT 1516.2400 1403.0400 1517.8400 1403.5200 ;
        RECT 1516.2400 1408.4800 1517.8400 1408.9600 ;
        RECT 1516.2400 1397.6000 1517.8400 1398.0800 ;
        RECT 1516.2400 1392.1600 1517.8400 1392.6400 ;
        RECT 1516.2400 1413.9200 1517.8400 1414.4000 ;
        RECT 1572.7800 1375.8400 1575.7800 1376.3200 ;
        RECT 1572.7800 1381.2800 1575.7800 1381.7600 ;
        RECT 1561.2400 1375.8400 1562.8400 1376.3200 ;
        RECT 1561.2400 1381.2800 1562.8400 1381.7600 ;
        RECT 1572.7800 1359.5200 1575.7800 1360.0000 ;
        RECT 1572.7800 1364.9600 1575.7800 1365.4400 ;
        RECT 1572.7800 1370.4000 1575.7800 1370.8800 ;
        RECT 1561.2400 1359.5200 1562.8400 1360.0000 ;
        RECT 1561.2400 1364.9600 1562.8400 1365.4400 ;
        RECT 1561.2400 1370.4000 1562.8400 1370.8800 ;
        RECT 1572.7800 1348.6400 1575.7800 1349.1200 ;
        RECT 1572.7800 1354.0800 1575.7800 1354.5600 ;
        RECT 1561.2400 1348.6400 1562.8400 1349.1200 ;
        RECT 1561.2400 1354.0800 1562.8400 1354.5600 ;
        RECT 1572.7800 1332.3200 1575.7800 1332.8000 ;
        RECT 1572.7800 1337.7600 1575.7800 1338.2400 ;
        RECT 1572.7800 1343.2000 1575.7800 1343.6800 ;
        RECT 1561.2400 1332.3200 1562.8400 1332.8000 ;
        RECT 1561.2400 1337.7600 1562.8400 1338.2400 ;
        RECT 1561.2400 1343.2000 1562.8400 1343.6800 ;
        RECT 1516.2400 1375.8400 1517.8400 1376.3200 ;
        RECT 1516.2400 1381.2800 1517.8400 1381.7600 ;
        RECT 1516.2400 1359.5200 1517.8400 1360.0000 ;
        RECT 1516.2400 1364.9600 1517.8400 1365.4400 ;
        RECT 1516.2400 1370.4000 1517.8400 1370.8800 ;
        RECT 1516.2400 1348.6400 1517.8400 1349.1200 ;
        RECT 1516.2400 1354.0800 1517.8400 1354.5600 ;
        RECT 1516.2400 1332.3200 1517.8400 1332.8000 ;
        RECT 1516.2400 1337.7600 1517.8400 1338.2400 ;
        RECT 1516.2400 1343.2000 1517.8400 1343.6800 ;
        RECT 1572.7800 1386.7200 1575.7800 1387.2000 ;
        RECT 1516.2400 1386.7200 1517.8400 1387.2000 ;
        RECT 1561.2400 1386.7200 1562.8400 1387.2000 ;
        RECT 1471.2400 1419.3600 1472.8400 1419.8400 ;
        RECT 1471.2400 1424.8000 1472.8400 1425.2800 ;
        RECT 1471.2400 1430.2400 1472.8400 1430.7200 ;
        RECT 1426.2400 1419.3600 1427.8400 1419.8400 ;
        RECT 1426.2400 1424.8000 1427.8400 1425.2800 ;
        RECT 1426.2400 1430.2400 1427.8400 1430.7200 ;
        RECT 1471.2400 1403.0400 1472.8400 1403.5200 ;
        RECT 1471.2400 1408.4800 1472.8400 1408.9600 ;
        RECT 1471.2400 1392.1600 1472.8400 1392.6400 ;
        RECT 1471.2400 1397.6000 1472.8400 1398.0800 ;
        RECT 1426.2400 1403.0400 1427.8400 1403.5200 ;
        RECT 1426.2400 1408.4800 1427.8400 1408.9600 ;
        RECT 1426.2400 1392.1600 1427.8400 1392.6400 ;
        RECT 1426.2400 1397.6000 1427.8400 1398.0800 ;
        RECT 1426.2400 1413.9200 1427.8400 1414.4000 ;
        RECT 1471.2400 1413.9200 1472.8400 1414.4000 ;
        RECT 1376.6800 1430.2400 1379.6800 1430.7200 ;
        RECT 1376.6800 1424.8000 1379.6800 1425.2800 ;
        RECT 1376.6800 1419.3600 1379.6800 1419.8400 ;
        RECT 1376.6800 1408.4800 1379.6800 1408.9600 ;
        RECT 1376.6800 1403.0400 1379.6800 1403.5200 ;
        RECT 1376.6800 1397.6000 1379.6800 1398.0800 ;
        RECT 1376.6800 1392.1600 1379.6800 1392.6400 ;
        RECT 1376.6800 1413.9200 1379.6800 1414.4000 ;
        RECT 1471.2400 1375.8400 1472.8400 1376.3200 ;
        RECT 1471.2400 1381.2800 1472.8400 1381.7600 ;
        RECT 1471.2400 1359.5200 1472.8400 1360.0000 ;
        RECT 1471.2400 1364.9600 1472.8400 1365.4400 ;
        RECT 1471.2400 1370.4000 1472.8400 1370.8800 ;
        RECT 1426.2400 1375.8400 1427.8400 1376.3200 ;
        RECT 1426.2400 1381.2800 1427.8400 1381.7600 ;
        RECT 1426.2400 1359.5200 1427.8400 1360.0000 ;
        RECT 1426.2400 1364.9600 1427.8400 1365.4400 ;
        RECT 1426.2400 1370.4000 1427.8400 1370.8800 ;
        RECT 1471.2400 1348.6400 1472.8400 1349.1200 ;
        RECT 1471.2400 1354.0800 1472.8400 1354.5600 ;
        RECT 1471.2400 1332.3200 1472.8400 1332.8000 ;
        RECT 1471.2400 1337.7600 1472.8400 1338.2400 ;
        RECT 1471.2400 1343.2000 1472.8400 1343.6800 ;
        RECT 1426.2400 1348.6400 1427.8400 1349.1200 ;
        RECT 1426.2400 1354.0800 1427.8400 1354.5600 ;
        RECT 1426.2400 1332.3200 1427.8400 1332.8000 ;
        RECT 1426.2400 1337.7600 1427.8400 1338.2400 ;
        RECT 1426.2400 1343.2000 1427.8400 1343.6800 ;
        RECT 1376.6800 1375.8400 1379.6800 1376.3200 ;
        RECT 1376.6800 1381.2800 1379.6800 1381.7600 ;
        RECT 1376.6800 1364.9600 1379.6800 1365.4400 ;
        RECT 1376.6800 1359.5200 1379.6800 1360.0000 ;
        RECT 1376.6800 1370.4000 1379.6800 1370.8800 ;
        RECT 1376.6800 1348.6400 1379.6800 1349.1200 ;
        RECT 1376.6800 1354.0800 1379.6800 1354.5600 ;
        RECT 1376.6800 1337.7600 1379.6800 1338.2400 ;
        RECT 1376.6800 1332.3200 1379.6800 1332.8000 ;
        RECT 1376.6800 1343.2000 1379.6800 1343.6800 ;
        RECT 1376.6800 1386.7200 1379.6800 1387.2000 ;
        RECT 1426.2400 1386.7200 1427.8400 1387.2000 ;
        RECT 1471.2400 1386.7200 1472.8400 1387.2000 ;
        RECT 1572.7800 1321.4400 1575.7800 1321.9200 ;
        RECT 1572.7800 1326.8800 1575.7800 1327.3600 ;
        RECT 1561.2400 1321.4400 1562.8400 1321.9200 ;
        RECT 1561.2400 1326.8800 1562.8400 1327.3600 ;
        RECT 1572.7800 1305.1200 1575.7800 1305.6000 ;
        RECT 1572.7800 1310.5600 1575.7800 1311.0400 ;
        RECT 1572.7800 1316.0000 1575.7800 1316.4800 ;
        RECT 1561.2400 1305.1200 1562.8400 1305.6000 ;
        RECT 1561.2400 1310.5600 1562.8400 1311.0400 ;
        RECT 1561.2400 1316.0000 1562.8400 1316.4800 ;
        RECT 1572.7800 1294.2400 1575.7800 1294.7200 ;
        RECT 1572.7800 1299.6800 1575.7800 1300.1600 ;
        RECT 1561.2400 1294.2400 1562.8400 1294.7200 ;
        RECT 1561.2400 1299.6800 1562.8400 1300.1600 ;
        RECT 1572.7800 1277.9200 1575.7800 1278.4000 ;
        RECT 1572.7800 1283.3600 1575.7800 1283.8400 ;
        RECT 1572.7800 1288.8000 1575.7800 1289.2800 ;
        RECT 1561.2400 1277.9200 1562.8400 1278.4000 ;
        RECT 1561.2400 1283.3600 1562.8400 1283.8400 ;
        RECT 1561.2400 1288.8000 1562.8400 1289.2800 ;
        RECT 1516.2400 1321.4400 1517.8400 1321.9200 ;
        RECT 1516.2400 1326.8800 1517.8400 1327.3600 ;
        RECT 1516.2400 1305.1200 1517.8400 1305.6000 ;
        RECT 1516.2400 1310.5600 1517.8400 1311.0400 ;
        RECT 1516.2400 1316.0000 1517.8400 1316.4800 ;
        RECT 1516.2400 1294.2400 1517.8400 1294.7200 ;
        RECT 1516.2400 1299.6800 1517.8400 1300.1600 ;
        RECT 1516.2400 1277.9200 1517.8400 1278.4000 ;
        RECT 1516.2400 1283.3600 1517.8400 1283.8400 ;
        RECT 1516.2400 1288.8000 1517.8400 1289.2800 ;
        RECT 1572.7800 1267.0400 1575.7800 1267.5200 ;
        RECT 1572.7800 1272.4800 1575.7800 1272.9600 ;
        RECT 1561.2400 1267.0400 1562.8400 1267.5200 ;
        RECT 1561.2400 1272.4800 1562.8400 1272.9600 ;
        RECT 1572.7800 1250.7200 1575.7800 1251.2000 ;
        RECT 1572.7800 1256.1600 1575.7800 1256.6400 ;
        RECT 1572.7800 1261.6000 1575.7800 1262.0800 ;
        RECT 1561.2400 1250.7200 1562.8400 1251.2000 ;
        RECT 1561.2400 1256.1600 1562.8400 1256.6400 ;
        RECT 1561.2400 1261.6000 1562.8400 1262.0800 ;
        RECT 1572.7800 1239.8400 1575.7800 1240.3200 ;
        RECT 1572.7800 1245.2800 1575.7800 1245.7600 ;
        RECT 1561.2400 1239.8400 1562.8400 1240.3200 ;
        RECT 1561.2400 1245.2800 1562.8400 1245.7600 ;
        RECT 1572.7800 1234.4000 1575.7800 1234.8800 ;
        RECT 1561.2400 1234.4000 1562.8400 1234.8800 ;
        RECT 1516.2400 1267.0400 1517.8400 1267.5200 ;
        RECT 1516.2400 1272.4800 1517.8400 1272.9600 ;
        RECT 1516.2400 1250.7200 1517.8400 1251.2000 ;
        RECT 1516.2400 1256.1600 1517.8400 1256.6400 ;
        RECT 1516.2400 1261.6000 1517.8400 1262.0800 ;
        RECT 1516.2400 1239.8400 1517.8400 1240.3200 ;
        RECT 1516.2400 1245.2800 1517.8400 1245.7600 ;
        RECT 1516.2400 1234.4000 1517.8400 1234.8800 ;
        RECT 1471.2400 1321.4400 1472.8400 1321.9200 ;
        RECT 1471.2400 1326.8800 1472.8400 1327.3600 ;
        RECT 1471.2400 1305.1200 1472.8400 1305.6000 ;
        RECT 1471.2400 1310.5600 1472.8400 1311.0400 ;
        RECT 1471.2400 1316.0000 1472.8400 1316.4800 ;
        RECT 1426.2400 1321.4400 1427.8400 1321.9200 ;
        RECT 1426.2400 1326.8800 1427.8400 1327.3600 ;
        RECT 1426.2400 1305.1200 1427.8400 1305.6000 ;
        RECT 1426.2400 1310.5600 1427.8400 1311.0400 ;
        RECT 1426.2400 1316.0000 1427.8400 1316.4800 ;
        RECT 1471.2400 1294.2400 1472.8400 1294.7200 ;
        RECT 1471.2400 1299.6800 1472.8400 1300.1600 ;
        RECT 1471.2400 1277.9200 1472.8400 1278.4000 ;
        RECT 1471.2400 1283.3600 1472.8400 1283.8400 ;
        RECT 1471.2400 1288.8000 1472.8400 1289.2800 ;
        RECT 1426.2400 1294.2400 1427.8400 1294.7200 ;
        RECT 1426.2400 1299.6800 1427.8400 1300.1600 ;
        RECT 1426.2400 1277.9200 1427.8400 1278.4000 ;
        RECT 1426.2400 1283.3600 1427.8400 1283.8400 ;
        RECT 1426.2400 1288.8000 1427.8400 1289.2800 ;
        RECT 1376.6800 1321.4400 1379.6800 1321.9200 ;
        RECT 1376.6800 1326.8800 1379.6800 1327.3600 ;
        RECT 1376.6800 1310.5600 1379.6800 1311.0400 ;
        RECT 1376.6800 1305.1200 1379.6800 1305.6000 ;
        RECT 1376.6800 1316.0000 1379.6800 1316.4800 ;
        RECT 1376.6800 1294.2400 1379.6800 1294.7200 ;
        RECT 1376.6800 1299.6800 1379.6800 1300.1600 ;
        RECT 1376.6800 1283.3600 1379.6800 1283.8400 ;
        RECT 1376.6800 1277.9200 1379.6800 1278.4000 ;
        RECT 1376.6800 1288.8000 1379.6800 1289.2800 ;
        RECT 1471.2400 1267.0400 1472.8400 1267.5200 ;
        RECT 1471.2400 1272.4800 1472.8400 1272.9600 ;
        RECT 1471.2400 1250.7200 1472.8400 1251.2000 ;
        RECT 1471.2400 1256.1600 1472.8400 1256.6400 ;
        RECT 1471.2400 1261.6000 1472.8400 1262.0800 ;
        RECT 1426.2400 1267.0400 1427.8400 1267.5200 ;
        RECT 1426.2400 1272.4800 1427.8400 1272.9600 ;
        RECT 1426.2400 1250.7200 1427.8400 1251.2000 ;
        RECT 1426.2400 1256.1600 1427.8400 1256.6400 ;
        RECT 1426.2400 1261.6000 1427.8400 1262.0800 ;
        RECT 1471.2400 1245.2800 1472.8400 1245.7600 ;
        RECT 1471.2400 1239.8400 1472.8400 1240.3200 ;
        RECT 1471.2400 1234.4000 1472.8400 1234.8800 ;
        RECT 1426.2400 1245.2800 1427.8400 1245.7600 ;
        RECT 1426.2400 1239.8400 1427.8400 1240.3200 ;
        RECT 1426.2400 1234.4000 1427.8400 1234.8800 ;
        RECT 1376.6800 1267.0400 1379.6800 1267.5200 ;
        RECT 1376.6800 1272.4800 1379.6800 1272.9600 ;
        RECT 1376.6800 1256.1600 1379.6800 1256.6400 ;
        RECT 1376.6800 1250.7200 1379.6800 1251.2000 ;
        RECT 1376.6800 1261.6000 1379.6800 1262.0800 ;
        RECT 1376.6800 1239.8400 1379.6800 1240.3200 ;
        RECT 1376.6800 1245.2800 1379.6800 1245.7600 ;
        RECT 1376.6800 1234.4000 1379.6800 1234.8800 ;
        RECT 1376.6800 1432.5900 1575.7800 1435.5900 ;
        RECT 1376.6800 1227.4900 1575.7800 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 997.8500 1562.8400 1205.9500 ;
        RECT 1516.2400 997.8500 1517.8400 1205.9500 ;
        RECT 1471.2400 997.8500 1472.8400 1205.9500 ;
        RECT 1426.2400 997.8500 1427.8400 1205.9500 ;
        RECT 1572.7800 997.8500 1575.7800 1205.9500 ;
        RECT 1376.6800 997.8500 1379.6800 1205.9500 ;
      LAYER met3 ;
        RECT 1572.7800 1200.6000 1575.7800 1201.0800 ;
        RECT 1561.2400 1200.6000 1562.8400 1201.0800 ;
        RECT 1572.7800 1189.7200 1575.7800 1190.2000 ;
        RECT 1572.7800 1195.1600 1575.7800 1195.6400 ;
        RECT 1561.2400 1189.7200 1562.8400 1190.2000 ;
        RECT 1561.2400 1195.1600 1562.8400 1195.6400 ;
        RECT 1572.7800 1173.4000 1575.7800 1173.8800 ;
        RECT 1572.7800 1178.8400 1575.7800 1179.3200 ;
        RECT 1561.2400 1173.4000 1562.8400 1173.8800 ;
        RECT 1561.2400 1178.8400 1562.8400 1179.3200 ;
        RECT 1572.7800 1162.5200 1575.7800 1163.0000 ;
        RECT 1572.7800 1167.9600 1575.7800 1168.4400 ;
        RECT 1561.2400 1162.5200 1562.8400 1163.0000 ;
        RECT 1561.2400 1167.9600 1562.8400 1168.4400 ;
        RECT 1572.7800 1184.2800 1575.7800 1184.7600 ;
        RECT 1561.2400 1184.2800 1562.8400 1184.7600 ;
        RECT 1516.2400 1189.7200 1517.8400 1190.2000 ;
        RECT 1516.2400 1195.1600 1517.8400 1195.6400 ;
        RECT 1516.2400 1200.6000 1517.8400 1201.0800 ;
        RECT 1516.2400 1173.4000 1517.8400 1173.8800 ;
        RECT 1516.2400 1178.8400 1517.8400 1179.3200 ;
        RECT 1516.2400 1167.9600 1517.8400 1168.4400 ;
        RECT 1516.2400 1162.5200 1517.8400 1163.0000 ;
        RECT 1516.2400 1184.2800 1517.8400 1184.7600 ;
        RECT 1572.7800 1146.2000 1575.7800 1146.6800 ;
        RECT 1572.7800 1151.6400 1575.7800 1152.1200 ;
        RECT 1561.2400 1146.2000 1562.8400 1146.6800 ;
        RECT 1561.2400 1151.6400 1562.8400 1152.1200 ;
        RECT 1572.7800 1129.8800 1575.7800 1130.3600 ;
        RECT 1572.7800 1135.3200 1575.7800 1135.8000 ;
        RECT 1572.7800 1140.7600 1575.7800 1141.2400 ;
        RECT 1561.2400 1129.8800 1562.8400 1130.3600 ;
        RECT 1561.2400 1135.3200 1562.8400 1135.8000 ;
        RECT 1561.2400 1140.7600 1562.8400 1141.2400 ;
        RECT 1572.7800 1119.0000 1575.7800 1119.4800 ;
        RECT 1572.7800 1124.4400 1575.7800 1124.9200 ;
        RECT 1561.2400 1119.0000 1562.8400 1119.4800 ;
        RECT 1561.2400 1124.4400 1562.8400 1124.9200 ;
        RECT 1572.7800 1102.6800 1575.7800 1103.1600 ;
        RECT 1572.7800 1108.1200 1575.7800 1108.6000 ;
        RECT 1572.7800 1113.5600 1575.7800 1114.0400 ;
        RECT 1561.2400 1102.6800 1562.8400 1103.1600 ;
        RECT 1561.2400 1108.1200 1562.8400 1108.6000 ;
        RECT 1561.2400 1113.5600 1562.8400 1114.0400 ;
        RECT 1516.2400 1146.2000 1517.8400 1146.6800 ;
        RECT 1516.2400 1151.6400 1517.8400 1152.1200 ;
        RECT 1516.2400 1129.8800 1517.8400 1130.3600 ;
        RECT 1516.2400 1135.3200 1517.8400 1135.8000 ;
        RECT 1516.2400 1140.7600 1517.8400 1141.2400 ;
        RECT 1516.2400 1119.0000 1517.8400 1119.4800 ;
        RECT 1516.2400 1124.4400 1517.8400 1124.9200 ;
        RECT 1516.2400 1102.6800 1517.8400 1103.1600 ;
        RECT 1516.2400 1108.1200 1517.8400 1108.6000 ;
        RECT 1516.2400 1113.5600 1517.8400 1114.0400 ;
        RECT 1572.7800 1157.0800 1575.7800 1157.5600 ;
        RECT 1516.2400 1157.0800 1517.8400 1157.5600 ;
        RECT 1561.2400 1157.0800 1562.8400 1157.5600 ;
        RECT 1471.2400 1189.7200 1472.8400 1190.2000 ;
        RECT 1471.2400 1195.1600 1472.8400 1195.6400 ;
        RECT 1471.2400 1200.6000 1472.8400 1201.0800 ;
        RECT 1426.2400 1189.7200 1427.8400 1190.2000 ;
        RECT 1426.2400 1195.1600 1427.8400 1195.6400 ;
        RECT 1426.2400 1200.6000 1427.8400 1201.0800 ;
        RECT 1471.2400 1173.4000 1472.8400 1173.8800 ;
        RECT 1471.2400 1178.8400 1472.8400 1179.3200 ;
        RECT 1471.2400 1162.5200 1472.8400 1163.0000 ;
        RECT 1471.2400 1167.9600 1472.8400 1168.4400 ;
        RECT 1426.2400 1173.4000 1427.8400 1173.8800 ;
        RECT 1426.2400 1178.8400 1427.8400 1179.3200 ;
        RECT 1426.2400 1162.5200 1427.8400 1163.0000 ;
        RECT 1426.2400 1167.9600 1427.8400 1168.4400 ;
        RECT 1426.2400 1184.2800 1427.8400 1184.7600 ;
        RECT 1471.2400 1184.2800 1472.8400 1184.7600 ;
        RECT 1376.6800 1200.6000 1379.6800 1201.0800 ;
        RECT 1376.6800 1195.1600 1379.6800 1195.6400 ;
        RECT 1376.6800 1189.7200 1379.6800 1190.2000 ;
        RECT 1376.6800 1178.8400 1379.6800 1179.3200 ;
        RECT 1376.6800 1173.4000 1379.6800 1173.8800 ;
        RECT 1376.6800 1167.9600 1379.6800 1168.4400 ;
        RECT 1376.6800 1162.5200 1379.6800 1163.0000 ;
        RECT 1376.6800 1184.2800 1379.6800 1184.7600 ;
        RECT 1471.2400 1146.2000 1472.8400 1146.6800 ;
        RECT 1471.2400 1151.6400 1472.8400 1152.1200 ;
        RECT 1471.2400 1129.8800 1472.8400 1130.3600 ;
        RECT 1471.2400 1135.3200 1472.8400 1135.8000 ;
        RECT 1471.2400 1140.7600 1472.8400 1141.2400 ;
        RECT 1426.2400 1146.2000 1427.8400 1146.6800 ;
        RECT 1426.2400 1151.6400 1427.8400 1152.1200 ;
        RECT 1426.2400 1129.8800 1427.8400 1130.3600 ;
        RECT 1426.2400 1135.3200 1427.8400 1135.8000 ;
        RECT 1426.2400 1140.7600 1427.8400 1141.2400 ;
        RECT 1471.2400 1119.0000 1472.8400 1119.4800 ;
        RECT 1471.2400 1124.4400 1472.8400 1124.9200 ;
        RECT 1471.2400 1102.6800 1472.8400 1103.1600 ;
        RECT 1471.2400 1108.1200 1472.8400 1108.6000 ;
        RECT 1471.2400 1113.5600 1472.8400 1114.0400 ;
        RECT 1426.2400 1119.0000 1427.8400 1119.4800 ;
        RECT 1426.2400 1124.4400 1427.8400 1124.9200 ;
        RECT 1426.2400 1102.6800 1427.8400 1103.1600 ;
        RECT 1426.2400 1108.1200 1427.8400 1108.6000 ;
        RECT 1426.2400 1113.5600 1427.8400 1114.0400 ;
        RECT 1376.6800 1146.2000 1379.6800 1146.6800 ;
        RECT 1376.6800 1151.6400 1379.6800 1152.1200 ;
        RECT 1376.6800 1135.3200 1379.6800 1135.8000 ;
        RECT 1376.6800 1129.8800 1379.6800 1130.3600 ;
        RECT 1376.6800 1140.7600 1379.6800 1141.2400 ;
        RECT 1376.6800 1119.0000 1379.6800 1119.4800 ;
        RECT 1376.6800 1124.4400 1379.6800 1124.9200 ;
        RECT 1376.6800 1108.1200 1379.6800 1108.6000 ;
        RECT 1376.6800 1102.6800 1379.6800 1103.1600 ;
        RECT 1376.6800 1113.5600 1379.6800 1114.0400 ;
        RECT 1376.6800 1157.0800 1379.6800 1157.5600 ;
        RECT 1426.2400 1157.0800 1427.8400 1157.5600 ;
        RECT 1471.2400 1157.0800 1472.8400 1157.5600 ;
        RECT 1572.7800 1091.8000 1575.7800 1092.2800 ;
        RECT 1572.7800 1097.2400 1575.7800 1097.7200 ;
        RECT 1561.2400 1091.8000 1562.8400 1092.2800 ;
        RECT 1561.2400 1097.2400 1562.8400 1097.7200 ;
        RECT 1572.7800 1075.4800 1575.7800 1075.9600 ;
        RECT 1572.7800 1080.9200 1575.7800 1081.4000 ;
        RECT 1572.7800 1086.3600 1575.7800 1086.8400 ;
        RECT 1561.2400 1075.4800 1562.8400 1075.9600 ;
        RECT 1561.2400 1080.9200 1562.8400 1081.4000 ;
        RECT 1561.2400 1086.3600 1562.8400 1086.8400 ;
        RECT 1572.7800 1064.6000 1575.7800 1065.0800 ;
        RECT 1572.7800 1070.0400 1575.7800 1070.5200 ;
        RECT 1561.2400 1064.6000 1562.8400 1065.0800 ;
        RECT 1561.2400 1070.0400 1562.8400 1070.5200 ;
        RECT 1572.7800 1048.2800 1575.7800 1048.7600 ;
        RECT 1572.7800 1053.7200 1575.7800 1054.2000 ;
        RECT 1572.7800 1059.1600 1575.7800 1059.6400 ;
        RECT 1561.2400 1048.2800 1562.8400 1048.7600 ;
        RECT 1561.2400 1053.7200 1562.8400 1054.2000 ;
        RECT 1561.2400 1059.1600 1562.8400 1059.6400 ;
        RECT 1516.2400 1091.8000 1517.8400 1092.2800 ;
        RECT 1516.2400 1097.2400 1517.8400 1097.7200 ;
        RECT 1516.2400 1075.4800 1517.8400 1075.9600 ;
        RECT 1516.2400 1080.9200 1517.8400 1081.4000 ;
        RECT 1516.2400 1086.3600 1517.8400 1086.8400 ;
        RECT 1516.2400 1064.6000 1517.8400 1065.0800 ;
        RECT 1516.2400 1070.0400 1517.8400 1070.5200 ;
        RECT 1516.2400 1048.2800 1517.8400 1048.7600 ;
        RECT 1516.2400 1053.7200 1517.8400 1054.2000 ;
        RECT 1516.2400 1059.1600 1517.8400 1059.6400 ;
        RECT 1572.7800 1037.4000 1575.7800 1037.8800 ;
        RECT 1572.7800 1042.8400 1575.7800 1043.3200 ;
        RECT 1561.2400 1037.4000 1562.8400 1037.8800 ;
        RECT 1561.2400 1042.8400 1562.8400 1043.3200 ;
        RECT 1572.7800 1021.0800 1575.7800 1021.5600 ;
        RECT 1572.7800 1026.5200 1575.7800 1027.0000 ;
        RECT 1572.7800 1031.9600 1575.7800 1032.4400 ;
        RECT 1561.2400 1021.0800 1562.8400 1021.5600 ;
        RECT 1561.2400 1026.5200 1562.8400 1027.0000 ;
        RECT 1561.2400 1031.9600 1562.8400 1032.4400 ;
        RECT 1572.7800 1010.2000 1575.7800 1010.6800 ;
        RECT 1572.7800 1015.6400 1575.7800 1016.1200 ;
        RECT 1561.2400 1010.2000 1562.8400 1010.6800 ;
        RECT 1561.2400 1015.6400 1562.8400 1016.1200 ;
        RECT 1572.7800 1004.7600 1575.7800 1005.2400 ;
        RECT 1561.2400 1004.7600 1562.8400 1005.2400 ;
        RECT 1516.2400 1037.4000 1517.8400 1037.8800 ;
        RECT 1516.2400 1042.8400 1517.8400 1043.3200 ;
        RECT 1516.2400 1021.0800 1517.8400 1021.5600 ;
        RECT 1516.2400 1026.5200 1517.8400 1027.0000 ;
        RECT 1516.2400 1031.9600 1517.8400 1032.4400 ;
        RECT 1516.2400 1010.2000 1517.8400 1010.6800 ;
        RECT 1516.2400 1015.6400 1517.8400 1016.1200 ;
        RECT 1516.2400 1004.7600 1517.8400 1005.2400 ;
        RECT 1471.2400 1091.8000 1472.8400 1092.2800 ;
        RECT 1471.2400 1097.2400 1472.8400 1097.7200 ;
        RECT 1471.2400 1075.4800 1472.8400 1075.9600 ;
        RECT 1471.2400 1080.9200 1472.8400 1081.4000 ;
        RECT 1471.2400 1086.3600 1472.8400 1086.8400 ;
        RECT 1426.2400 1091.8000 1427.8400 1092.2800 ;
        RECT 1426.2400 1097.2400 1427.8400 1097.7200 ;
        RECT 1426.2400 1075.4800 1427.8400 1075.9600 ;
        RECT 1426.2400 1080.9200 1427.8400 1081.4000 ;
        RECT 1426.2400 1086.3600 1427.8400 1086.8400 ;
        RECT 1471.2400 1064.6000 1472.8400 1065.0800 ;
        RECT 1471.2400 1070.0400 1472.8400 1070.5200 ;
        RECT 1471.2400 1048.2800 1472.8400 1048.7600 ;
        RECT 1471.2400 1053.7200 1472.8400 1054.2000 ;
        RECT 1471.2400 1059.1600 1472.8400 1059.6400 ;
        RECT 1426.2400 1064.6000 1427.8400 1065.0800 ;
        RECT 1426.2400 1070.0400 1427.8400 1070.5200 ;
        RECT 1426.2400 1048.2800 1427.8400 1048.7600 ;
        RECT 1426.2400 1053.7200 1427.8400 1054.2000 ;
        RECT 1426.2400 1059.1600 1427.8400 1059.6400 ;
        RECT 1376.6800 1091.8000 1379.6800 1092.2800 ;
        RECT 1376.6800 1097.2400 1379.6800 1097.7200 ;
        RECT 1376.6800 1080.9200 1379.6800 1081.4000 ;
        RECT 1376.6800 1075.4800 1379.6800 1075.9600 ;
        RECT 1376.6800 1086.3600 1379.6800 1086.8400 ;
        RECT 1376.6800 1064.6000 1379.6800 1065.0800 ;
        RECT 1376.6800 1070.0400 1379.6800 1070.5200 ;
        RECT 1376.6800 1053.7200 1379.6800 1054.2000 ;
        RECT 1376.6800 1048.2800 1379.6800 1048.7600 ;
        RECT 1376.6800 1059.1600 1379.6800 1059.6400 ;
        RECT 1471.2400 1037.4000 1472.8400 1037.8800 ;
        RECT 1471.2400 1042.8400 1472.8400 1043.3200 ;
        RECT 1471.2400 1021.0800 1472.8400 1021.5600 ;
        RECT 1471.2400 1026.5200 1472.8400 1027.0000 ;
        RECT 1471.2400 1031.9600 1472.8400 1032.4400 ;
        RECT 1426.2400 1037.4000 1427.8400 1037.8800 ;
        RECT 1426.2400 1042.8400 1427.8400 1043.3200 ;
        RECT 1426.2400 1021.0800 1427.8400 1021.5600 ;
        RECT 1426.2400 1026.5200 1427.8400 1027.0000 ;
        RECT 1426.2400 1031.9600 1427.8400 1032.4400 ;
        RECT 1471.2400 1015.6400 1472.8400 1016.1200 ;
        RECT 1471.2400 1010.2000 1472.8400 1010.6800 ;
        RECT 1471.2400 1004.7600 1472.8400 1005.2400 ;
        RECT 1426.2400 1015.6400 1427.8400 1016.1200 ;
        RECT 1426.2400 1010.2000 1427.8400 1010.6800 ;
        RECT 1426.2400 1004.7600 1427.8400 1005.2400 ;
        RECT 1376.6800 1037.4000 1379.6800 1037.8800 ;
        RECT 1376.6800 1042.8400 1379.6800 1043.3200 ;
        RECT 1376.6800 1026.5200 1379.6800 1027.0000 ;
        RECT 1376.6800 1021.0800 1379.6800 1021.5600 ;
        RECT 1376.6800 1031.9600 1379.6800 1032.4400 ;
        RECT 1376.6800 1010.2000 1379.6800 1010.6800 ;
        RECT 1376.6800 1015.6400 1379.6800 1016.1200 ;
        RECT 1376.6800 1004.7600 1379.6800 1005.2400 ;
        RECT 1376.6800 1202.9500 1575.7800 1205.9500 ;
        RECT 1376.6800 997.8500 1575.7800 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1561.2400 768.2100 1562.8400 976.3100 ;
        RECT 1516.2400 768.2100 1517.8400 976.3100 ;
        RECT 1471.2400 768.2100 1472.8400 976.3100 ;
        RECT 1426.2400 768.2100 1427.8400 976.3100 ;
        RECT 1572.7800 768.2100 1575.7800 976.3100 ;
        RECT 1376.6800 768.2100 1379.6800 976.3100 ;
      LAYER met3 ;
        RECT 1572.7800 970.9600 1575.7800 971.4400 ;
        RECT 1561.2400 970.9600 1562.8400 971.4400 ;
        RECT 1572.7800 960.0800 1575.7800 960.5600 ;
        RECT 1572.7800 965.5200 1575.7800 966.0000 ;
        RECT 1561.2400 960.0800 1562.8400 960.5600 ;
        RECT 1561.2400 965.5200 1562.8400 966.0000 ;
        RECT 1572.7800 943.7600 1575.7800 944.2400 ;
        RECT 1572.7800 949.2000 1575.7800 949.6800 ;
        RECT 1561.2400 943.7600 1562.8400 944.2400 ;
        RECT 1561.2400 949.2000 1562.8400 949.6800 ;
        RECT 1572.7800 932.8800 1575.7800 933.3600 ;
        RECT 1572.7800 938.3200 1575.7800 938.8000 ;
        RECT 1561.2400 932.8800 1562.8400 933.3600 ;
        RECT 1561.2400 938.3200 1562.8400 938.8000 ;
        RECT 1572.7800 954.6400 1575.7800 955.1200 ;
        RECT 1561.2400 954.6400 1562.8400 955.1200 ;
        RECT 1516.2400 960.0800 1517.8400 960.5600 ;
        RECT 1516.2400 965.5200 1517.8400 966.0000 ;
        RECT 1516.2400 970.9600 1517.8400 971.4400 ;
        RECT 1516.2400 943.7600 1517.8400 944.2400 ;
        RECT 1516.2400 949.2000 1517.8400 949.6800 ;
        RECT 1516.2400 938.3200 1517.8400 938.8000 ;
        RECT 1516.2400 932.8800 1517.8400 933.3600 ;
        RECT 1516.2400 954.6400 1517.8400 955.1200 ;
        RECT 1572.7800 916.5600 1575.7800 917.0400 ;
        RECT 1572.7800 922.0000 1575.7800 922.4800 ;
        RECT 1561.2400 916.5600 1562.8400 917.0400 ;
        RECT 1561.2400 922.0000 1562.8400 922.4800 ;
        RECT 1572.7800 900.2400 1575.7800 900.7200 ;
        RECT 1572.7800 905.6800 1575.7800 906.1600 ;
        RECT 1572.7800 911.1200 1575.7800 911.6000 ;
        RECT 1561.2400 900.2400 1562.8400 900.7200 ;
        RECT 1561.2400 905.6800 1562.8400 906.1600 ;
        RECT 1561.2400 911.1200 1562.8400 911.6000 ;
        RECT 1572.7800 889.3600 1575.7800 889.8400 ;
        RECT 1572.7800 894.8000 1575.7800 895.2800 ;
        RECT 1561.2400 889.3600 1562.8400 889.8400 ;
        RECT 1561.2400 894.8000 1562.8400 895.2800 ;
        RECT 1572.7800 873.0400 1575.7800 873.5200 ;
        RECT 1572.7800 878.4800 1575.7800 878.9600 ;
        RECT 1572.7800 883.9200 1575.7800 884.4000 ;
        RECT 1561.2400 873.0400 1562.8400 873.5200 ;
        RECT 1561.2400 878.4800 1562.8400 878.9600 ;
        RECT 1561.2400 883.9200 1562.8400 884.4000 ;
        RECT 1516.2400 916.5600 1517.8400 917.0400 ;
        RECT 1516.2400 922.0000 1517.8400 922.4800 ;
        RECT 1516.2400 900.2400 1517.8400 900.7200 ;
        RECT 1516.2400 905.6800 1517.8400 906.1600 ;
        RECT 1516.2400 911.1200 1517.8400 911.6000 ;
        RECT 1516.2400 889.3600 1517.8400 889.8400 ;
        RECT 1516.2400 894.8000 1517.8400 895.2800 ;
        RECT 1516.2400 873.0400 1517.8400 873.5200 ;
        RECT 1516.2400 878.4800 1517.8400 878.9600 ;
        RECT 1516.2400 883.9200 1517.8400 884.4000 ;
        RECT 1572.7800 927.4400 1575.7800 927.9200 ;
        RECT 1516.2400 927.4400 1517.8400 927.9200 ;
        RECT 1561.2400 927.4400 1562.8400 927.9200 ;
        RECT 1471.2400 960.0800 1472.8400 960.5600 ;
        RECT 1471.2400 965.5200 1472.8400 966.0000 ;
        RECT 1471.2400 970.9600 1472.8400 971.4400 ;
        RECT 1426.2400 960.0800 1427.8400 960.5600 ;
        RECT 1426.2400 965.5200 1427.8400 966.0000 ;
        RECT 1426.2400 970.9600 1427.8400 971.4400 ;
        RECT 1471.2400 943.7600 1472.8400 944.2400 ;
        RECT 1471.2400 949.2000 1472.8400 949.6800 ;
        RECT 1471.2400 932.8800 1472.8400 933.3600 ;
        RECT 1471.2400 938.3200 1472.8400 938.8000 ;
        RECT 1426.2400 943.7600 1427.8400 944.2400 ;
        RECT 1426.2400 949.2000 1427.8400 949.6800 ;
        RECT 1426.2400 932.8800 1427.8400 933.3600 ;
        RECT 1426.2400 938.3200 1427.8400 938.8000 ;
        RECT 1426.2400 954.6400 1427.8400 955.1200 ;
        RECT 1471.2400 954.6400 1472.8400 955.1200 ;
        RECT 1376.6800 970.9600 1379.6800 971.4400 ;
        RECT 1376.6800 965.5200 1379.6800 966.0000 ;
        RECT 1376.6800 960.0800 1379.6800 960.5600 ;
        RECT 1376.6800 949.2000 1379.6800 949.6800 ;
        RECT 1376.6800 943.7600 1379.6800 944.2400 ;
        RECT 1376.6800 938.3200 1379.6800 938.8000 ;
        RECT 1376.6800 932.8800 1379.6800 933.3600 ;
        RECT 1376.6800 954.6400 1379.6800 955.1200 ;
        RECT 1471.2400 916.5600 1472.8400 917.0400 ;
        RECT 1471.2400 922.0000 1472.8400 922.4800 ;
        RECT 1471.2400 900.2400 1472.8400 900.7200 ;
        RECT 1471.2400 905.6800 1472.8400 906.1600 ;
        RECT 1471.2400 911.1200 1472.8400 911.6000 ;
        RECT 1426.2400 916.5600 1427.8400 917.0400 ;
        RECT 1426.2400 922.0000 1427.8400 922.4800 ;
        RECT 1426.2400 900.2400 1427.8400 900.7200 ;
        RECT 1426.2400 905.6800 1427.8400 906.1600 ;
        RECT 1426.2400 911.1200 1427.8400 911.6000 ;
        RECT 1471.2400 889.3600 1472.8400 889.8400 ;
        RECT 1471.2400 894.8000 1472.8400 895.2800 ;
        RECT 1471.2400 873.0400 1472.8400 873.5200 ;
        RECT 1471.2400 878.4800 1472.8400 878.9600 ;
        RECT 1471.2400 883.9200 1472.8400 884.4000 ;
        RECT 1426.2400 889.3600 1427.8400 889.8400 ;
        RECT 1426.2400 894.8000 1427.8400 895.2800 ;
        RECT 1426.2400 873.0400 1427.8400 873.5200 ;
        RECT 1426.2400 878.4800 1427.8400 878.9600 ;
        RECT 1426.2400 883.9200 1427.8400 884.4000 ;
        RECT 1376.6800 916.5600 1379.6800 917.0400 ;
        RECT 1376.6800 922.0000 1379.6800 922.4800 ;
        RECT 1376.6800 905.6800 1379.6800 906.1600 ;
        RECT 1376.6800 900.2400 1379.6800 900.7200 ;
        RECT 1376.6800 911.1200 1379.6800 911.6000 ;
        RECT 1376.6800 889.3600 1379.6800 889.8400 ;
        RECT 1376.6800 894.8000 1379.6800 895.2800 ;
        RECT 1376.6800 878.4800 1379.6800 878.9600 ;
        RECT 1376.6800 873.0400 1379.6800 873.5200 ;
        RECT 1376.6800 883.9200 1379.6800 884.4000 ;
        RECT 1376.6800 927.4400 1379.6800 927.9200 ;
        RECT 1426.2400 927.4400 1427.8400 927.9200 ;
        RECT 1471.2400 927.4400 1472.8400 927.9200 ;
        RECT 1572.7800 862.1600 1575.7800 862.6400 ;
        RECT 1572.7800 867.6000 1575.7800 868.0800 ;
        RECT 1561.2400 862.1600 1562.8400 862.6400 ;
        RECT 1561.2400 867.6000 1562.8400 868.0800 ;
        RECT 1572.7800 845.8400 1575.7800 846.3200 ;
        RECT 1572.7800 851.2800 1575.7800 851.7600 ;
        RECT 1572.7800 856.7200 1575.7800 857.2000 ;
        RECT 1561.2400 845.8400 1562.8400 846.3200 ;
        RECT 1561.2400 851.2800 1562.8400 851.7600 ;
        RECT 1561.2400 856.7200 1562.8400 857.2000 ;
        RECT 1572.7800 834.9600 1575.7800 835.4400 ;
        RECT 1572.7800 840.4000 1575.7800 840.8800 ;
        RECT 1561.2400 834.9600 1562.8400 835.4400 ;
        RECT 1561.2400 840.4000 1562.8400 840.8800 ;
        RECT 1572.7800 818.6400 1575.7800 819.1200 ;
        RECT 1572.7800 824.0800 1575.7800 824.5600 ;
        RECT 1572.7800 829.5200 1575.7800 830.0000 ;
        RECT 1561.2400 818.6400 1562.8400 819.1200 ;
        RECT 1561.2400 824.0800 1562.8400 824.5600 ;
        RECT 1561.2400 829.5200 1562.8400 830.0000 ;
        RECT 1516.2400 862.1600 1517.8400 862.6400 ;
        RECT 1516.2400 867.6000 1517.8400 868.0800 ;
        RECT 1516.2400 845.8400 1517.8400 846.3200 ;
        RECT 1516.2400 851.2800 1517.8400 851.7600 ;
        RECT 1516.2400 856.7200 1517.8400 857.2000 ;
        RECT 1516.2400 834.9600 1517.8400 835.4400 ;
        RECT 1516.2400 840.4000 1517.8400 840.8800 ;
        RECT 1516.2400 818.6400 1517.8400 819.1200 ;
        RECT 1516.2400 824.0800 1517.8400 824.5600 ;
        RECT 1516.2400 829.5200 1517.8400 830.0000 ;
        RECT 1572.7800 807.7600 1575.7800 808.2400 ;
        RECT 1572.7800 813.2000 1575.7800 813.6800 ;
        RECT 1561.2400 807.7600 1562.8400 808.2400 ;
        RECT 1561.2400 813.2000 1562.8400 813.6800 ;
        RECT 1572.7800 791.4400 1575.7800 791.9200 ;
        RECT 1572.7800 796.8800 1575.7800 797.3600 ;
        RECT 1572.7800 802.3200 1575.7800 802.8000 ;
        RECT 1561.2400 791.4400 1562.8400 791.9200 ;
        RECT 1561.2400 796.8800 1562.8400 797.3600 ;
        RECT 1561.2400 802.3200 1562.8400 802.8000 ;
        RECT 1572.7800 780.5600 1575.7800 781.0400 ;
        RECT 1572.7800 786.0000 1575.7800 786.4800 ;
        RECT 1561.2400 780.5600 1562.8400 781.0400 ;
        RECT 1561.2400 786.0000 1562.8400 786.4800 ;
        RECT 1572.7800 775.1200 1575.7800 775.6000 ;
        RECT 1561.2400 775.1200 1562.8400 775.6000 ;
        RECT 1516.2400 807.7600 1517.8400 808.2400 ;
        RECT 1516.2400 813.2000 1517.8400 813.6800 ;
        RECT 1516.2400 791.4400 1517.8400 791.9200 ;
        RECT 1516.2400 796.8800 1517.8400 797.3600 ;
        RECT 1516.2400 802.3200 1517.8400 802.8000 ;
        RECT 1516.2400 780.5600 1517.8400 781.0400 ;
        RECT 1516.2400 786.0000 1517.8400 786.4800 ;
        RECT 1516.2400 775.1200 1517.8400 775.6000 ;
        RECT 1471.2400 862.1600 1472.8400 862.6400 ;
        RECT 1471.2400 867.6000 1472.8400 868.0800 ;
        RECT 1471.2400 845.8400 1472.8400 846.3200 ;
        RECT 1471.2400 851.2800 1472.8400 851.7600 ;
        RECT 1471.2400 856.7200 1472.8400 857.2000 ;
        RECT 1426.2400 862.1600 1427.8400 862.6400 ;
        RECT 1426.2400 867.6000 1427.8400 868.0800 ;
        RECT 1426.2400 845.8400 1427.8400 846.3200 ;
        RECT 1426.2400 851.2800 1427.8400 851.7600 ;
        RECT 1426.2400 856.7200 1427.8400 857.2000 ;
        RECT 1471.2400 834.9600 1472.8400 835.4400 ;
        RECT 1471.2400 840.4000 1472.8400 840.8800 ;
        RECT 1471.2400 818.6400 1472.8400 819.1200 ;
        RECT 1471.2400 824.0800 1472.8400 824.5600 ;
        RECT 1471.2400 829.5200 1472.8400 830.0000 ;
        RECT 1426.2400 834.9600 1427.8400 835.4400 ;
        RECT 1426.2400 840.4000 1427.8400 840.8800 ;
        RECT 1426.2400 818.6400 1427.8400 819.1200 ;
        RECT 1426.2400 824.0800 1427.8400 824.5600 ;
        RECT 1426.2400 829.5200 1427.8400 830.0000 ;
        RECT 1376.6800 862.1600 1379.6800 862.6400 ;
        RECT 1376.6800 867.6000 1379.6800 868.0800 ;
        RECT 1376.6800 851.2800 1379.6800 851.7600 ;
        RECT 1376.6800 845.8400 1379.6800 846.3200 ;
        RECT 1376.6800 856.7200 1379.6800 857.2000 ;
        RECT 1376.6800 834.9600 1379.6800 835.4400 ;
        RECT 1376.6800 840.4000 1379.6800 840.8800 ;
        RECT 1376.6800 824.0800 1379.6800 824.5600 ;
        RECT 1376.6800 818.6400 1379.6800 819.1200 ;
        RECT 1376.6800 829.5200 1379.6800 830.0000 ;
        RECT 1471.2400 807.7600 1472.8400 808.2400 ;
        RECT 1471.2400 813.2000 1472.8400 813.6800 ;
        RECT 1471.2400 791.4400 1472.8400 791.9200 ;
        RECT 1471.2400 796.8800 1472.8400 797.3600 ;
        RECT 1471.2400 802.3200 1472.8400 802.8000 ;
        RECT 1426.2400 807.7600 1427.8400 808.2400 ;
        RECT 1426.2400 813.2000 1427.8400 813.6800 ;
        RECT 1426.2400 791.4400 1427.8400 791.9200 ;
        RECT 1426.2400 796.8800 1427.8400 797.3600 ;
        RECT 1426.2400 802.3200 1427.8400 802.8000 ;
        RECT 1471.2400 786.0000 1472.8400 786.4800 ;
        RECT 1471.2400 780.5600 1472.8400 781.0400 ;
        RECT 1471.2400 775.1200 1472.8400 775.6000 ;
        RECT 1426.2400 786.0000 1427.8400 786.4800 ;
        RECT 1426.2400 780.5600 1427.8400 781.0400 ;
        RECT 1426.2400 775.1200 1427.8400 775.6000 ;
        RECT 1376.6800 807.7600 1379.6800 808.2400 ;
        RECT 1376.6800 813.2000 1379.6800 813.6800 ;
        RECT 1376.6800 796.8800 1379.6800 797.3600 ;
        RECT 1376.6800 791.4400 1379.6800 791.9200 ;
        RECT 1376.6800 802.3200 1379.6800 802.8000 ;
        RECT 1376.6800 780.5600 1379.6800 781.0400 ;
        RECT 1376.6800 786.0000 1379.6800 786.4800 ;
        RECT 1376.6800 775.1200 1379.6800 775.6000 ;
        RECT 1376.6800 973.3100 1575.7800 976.3100 ;
        RECT 1376.6800 768.2100 1575.7800 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1596.9000 2833.6100 1598.9000 2854.5400 ;
        RECT 1794.0000 2833.6100 1796.0000 2854.5400 ;
      LAYER met3 ;
        RECT 1794.0000 2850.0400 1796.0000 2850.5200 ;
        RECT 1596.9000 2850.0400 1598.9000 2850.5200 ;
        RECT 1794.0000 2839.1600 1796.0000 2839.6400 ;
        RECT 1596.9000 2839.1600 1598.9000 2839.6400 ;
        RECT 1794.0000 2844.6000 1796.0000 2845.0800 ;
        RECT 1596.9000 2844.6000 1598.9000 2845.0800 ;
        RECT 1596.9000 2852.5400 1796.0000 2854.5400 ;
        RECT 1596.9000 2833.6100 1796.0000 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 538.5700 1783.0600 746.6700 ;
        RECT 1736.4600 538.5700 1738.0600 746.6700 ;
        RECT 1691.4600 538.5700 1693.0600 746.6700 ;
        RECT 1646.4600 538.5700 1648.0600 746.6700 ;
        RECT 1793.0000 538.5700 1796.0000 746.6700 ;
        RECT 1596.9000 538.5700 1599.9000 746.6700 ;
      LAYER met3 ;
        RECT 1793.0000 741.3200 1796.0000 741.8000 ;
        RECT 1781.4600 741.3200 1783.0600 741.8000 ;
        RECT 1793.0000 730.4400 1796.0000 730.9200 ;
        RECT 1793.0000 735.8800 1796.0000 736.3600 ;
        RECT 1781.4600 730.4400 1783.0600 730.9200 ;
        RECT 1781.4600 735.8800 1783.0600 736.3600 ;
        RECT 1793.0000 714.1200 1796.0000 714.6000 ;
        RECT 1793.0000 719.5600 1796.0000 720.0400 ;
        RECT 1781.4600 714.1200 1783.0600 714.6000 ;
        RECT 1781.4600 719.5600 1783.0600 720.0400 ;
        RECT 1793.0000 703.2400 1796.0000 703.7200 ;
        RECT 1793.0000 708.6800 1796.0000 709.1600 ;
        RECT 1781.4600 703.2400 1783.0600 703.7200 ;
        RECT 1781.4600 708.6800 1783.0600 709.1600 ;
        RECT 1793.0000 725.0000 1796.0000 725.4800 ;
        RECT 1781.4600 725.0000 1783.0600 725.4800 ;
        RECT 1736.4600 730.4400 1738.0600 730.9200 ;
        RECT 1736.4600 735.8800 1738.0600 736.3600 ;
        RECT 1736.4600 741.3200 1738.0600 741.8000 ;
        RECT 1736.4600 714.1200 1738.0600 714.6000 ;
        RECT 1736.4600 719.5600 1738.0600 720.0400 ;
        RECT 1736.4600 708.6800 1738.0600 709.1600 ;
        RECT 1736.4600 703.2400 1738.0600 703.7200 ;
        RECT 1736.4600 725.0000 1738.0600 725.4800 ;
        RECT 1793.0000 686.9200 1796.0000 687.4000 ;
        RECT 1793.0000 692.3600 1796.0000 692.8400 ;
        RECT 1781.4600 686.9200 1783.0600 687.4000 ;
        RECT 1781.4600 692.3600 1783.0600 692.8400 ;
        RECT 1793.0000 670.6000 1796.0000 671.0800 ;
        RECT 1793.0000 676.0400 1796.0000 676.5200 ;
        RECT 1793.0000 681.4800 1796.0000 681.9600 ;
        RECT 1781.4600 670.6000 1783.0600 671.0800 ;
        RECT 1781.4600 676.0400 1783.0600 676.5200 ;
        RECT 1781.4600 681.4800 1783.0600 681.9600 ;
        RECT 1793.0000 659.7200 1796.0000 660.2000 ;
        RECT 1793.0000 665.1600 1796.0000 665.6400 ;
        RECT 1781.4600 659.7200 1783.0600 660.2000 ;
        RECT 1781.4600 665.1600 1783.0600 665.6400 ;
        RECT 1793.0000 643.4000 1796.0000 643.8800 ;
        RECT 1793.0000 648.8400 1796.0000 649.3200 ;
        RECT 1793.0000 654.2800 1796.0000 654.7600 ;
        RECT 1781.4600 643.4000 1783.0600 643.8800 ;
        RECT 1781.4600 648.8400 1783.0600 649.3200 ;
        RECT 1781.4600 654.2800 1783.0600 654.7600 ;
        RECT 1736.4600 686.9200 1738.0600 687.4000 ;
        RECT 1736.4600 692.3600 1738.0600 692.8400 ;
        RECT 1736.4600 670.6000 1738.0600 671.0800 ;
        RECT 1736.4600 676.0400 1738.0600 676.5200 ;
        RECT 1736.4600 681.4800 1738.0600 681.9600 ;
        RECT 1736.4600 659.7200 1738.0600 660.2000 ;
        RECT 1736.4600 665.1600 1738.0600 665.6400 ;
        RECT 1736.4600 643.4000 1738.0600 643.8800 ;
        RECT 1736.4600 648.8400 1738.0600 649.3200 ;
        RECT 1736.4600 654.2800 1738.0600 654.7600 ;
        RECT 1793.0000 697.8000 1796.0000 698.2800 ;
        RECT 1736.4600 697.8000 1738.0600 698.2800 ;
        RECT 1781.4600 697.8000 1783.0600 698.2800 ;
        RECT 1691.4600 730.4400 1693.0600 730.9200 ;
        RECT 1691.4600 735.8800 1693.0600 736.3600 ;
        RECT 1691.4600 741.3200 1693.0600 741.8000 ;
        RECT 1646.4600 730.4400 1648.0600 730.9200 ;
        RECT 1646.4600 735.8800 1648.0600 736.3600 ;
        RECT 1646.4600 741.3200 1648.0600 741.8000 ;
        RECT 1691.4600 714.1200 1693.0600 714.6000 ;
        RECT 1691.4600 719.5600 1693.0600 720.0400 ;
        RECT 1691.4600 703.2400 1693.0600 703.7200 ;
        RECT 1691.4600 708.6800 1693.0600 709.1600 ;
        RECT 1646.4600 714.1200 1648.0600 714.6000 ;
        RECT 1646.4600 719.5600 1648.0600 720.0400 ;
        RECT 1646.4600 703.2400 1648.0600 703.7200 ;
        RECT 1646.4600 708.6800 1648.0600 709.1600 ;
        RECT 1646.4600 725.0000 1648.0600 725.4800 ;
        RECT 1691.4600 725.0000 1693.0600 725.4800 ;
        RECT 1596.9000 741.3200 1599.9000 741.8000 ;
        RECT 1596.9000 735.8800 1599.9000 736.3600 ;
        RECT 1596.9000 730.4400 1599.9000 730.9200 ;
        RECT 1596.9000 719.5600 1599.9000 720.0400 ;
        RECT 1596.9000 714.1200 1599.9000 714.6000 ;
        RECT 1596.9000 708.6800 1599.9000 709.1600 ;
        RECT 1596.9000 703.2400 1599.9000 703.7200 ;
        RECT 1596.9000 725.0000 1599.9000 725.4800 ;
        RECT 1691.4600 686.9200 1693.0600 687.4000 ;
        RECT 1691.4600 692.3600 1693.0600 692.8400 ;
        RECT 1691.4600 670.6000 1693.0600 671.0800 ;
        RECT 1691.4600 676.0400 1693.0600 676.5200 ;
        RECT 1691.4600 681.4800 1693.0600 681.9600 ;
        RECT 1646.4600 686.9200 1648.0600 687.4000 ;
        RECT 1646.4600 692.3600 1648.0600 692.8400 ;
        RECT 1646.4600 670.6000 1648.0600 671.0800 ;
        RECT 1646.4600 676.0400 1648.0600 676.5200 ;
        RECT 1646.4600 681.4800 1648.0600 681.9600 ;
        RECT 1691.4600 659.7200 1693.0600 660.2000 ;
        RECT 1691.4600 665.1600 1693.0600 665.6400 ;
        RECT 1691.4600 643.4000 1693.0600 643.8800 ;
        RECT 1691.4600 648.8400 1693.0600 649.3200 ;
        RECT 1691.4600 654.2800 1693.0600 654.7600 ;
        RECT 1646.4600 659.7200 1648.0600 660.2000 ;
        RECT 1646.4600 665.1600 1648.0600 665.6400 ;
        RECT 1646.4600 643.4000 1648.0600 643.8800 ;
        RECT 1646.4600 648.8400 1648.0600 649.3200 ;
        RECT 1646.4600 654.2800 1648.0600 654.7600 ;
        RECT 1596.9000 686.9200 1599.9000 687.4000 ;
        RECT 1596.9000 692.3600 1599.9000 692.8400 ;
        RECT 1596.9000 676.0400 1599.9000 676.5200 ;
        RECT 1596.9000 670.6000 1599.9000 671.0800 ;
        RECT 1596.9000 681.4800 1599.9000 681.9600 ;
        RECT 1596.9000 659.7200 1599.9000 660.2000 ;
        RECT 1596.9000 665.1600 1599.9000 665.6400 ;
        RECT 1596.9000 648.8400 1599.9000 649.3200 ;
        RECT 1596.9000 643.4000 1599.9000 643.8800 ;
        RECT 1596.9000 654.2800 1599.9000 654.7600 ;
        RECT 1596.9000 697.8000 1599.9000 698.2800 ;
        RECT 1646.4600 697.8000 1648.0600 698.2800 ;
        RECT 1691.4600 697.8000 1693.0600 698.2800 ;
        RECT 1793.0000 632.5200 1796.0000 633.0000 ;
        RECT 1793.0000 637.9600 1796.0000 638.4400 ;
        RECT 1781.4600 632.5200 1783.0600 633.0000 ;
        RECT 1781.4600 637.9600 1783.0600 638.4400 ;
        RECT 1793.0000 616.2000 1796.0000 616.6800 ;
        RECT 1793.0000 621.6400 1796.0000 622.1200 ;
        RECT 1793.0000 627.0800 1796.0000 627.5600 ;
        RECT 1781.4600 616.2000 1783.0600 616.6800 ;
        RECT 1781.4600 621.6400 1783.0600 622.1200 ;
        RECT 1781.4600 627.0800 1783.0600 627.5600 ;
        RECT 1793.0000 605.3200 1796.0000 605.8000 ;
        RECT 1793.0000 610.7600 1796.0000 611.2400 ;
        RECT 1781.4600 605.3200 1783.0600 605.8000 ;
        RECT 1781.4600 610.7600 1783.0600 611.2400 ;
        RECT 1793.0000 589.0000 1796.0000 589.4800 ;
        RECT 1793.0000 594.4400 1796.0000 594.9200 ;
        RECT 1793.0000 599.8800 1796.0000 600.3600 ;
        RECT 1781.4600 589.0000 1783.0600 589.4800 ;
        RECT 1781.4600 594.4400 1783.0600 594.9200 ;
        RECT 1781.4600 599.8800 1783.0600 600.3600 ;
        RECT 1736.4600 632.5200 1738.0600 633.0000 ;
        RECT 1736.4600 637.9600 1738.0600 638.4400 ;
        RECT 1736.4600 616.2000 1738.0600 616.6800 ;
        RECT 1736.4600 621.6400 1738.0600 622.1200 ;
        RECT 1736.4600 627.0800 1738.0600 627.5600 ;
        RECT 1736.4600 605.3200 1738.0600 605.8000 ;
        RECT 1736.4600 610.7600 1738.0600 611.2400 ;
        RECT 1736.4600 589.0000 1738.0600 589.4800 ;
        RECT 1736.4600 594.4400 1738.0600 594.9200 ;
        RECT 1736.4600 599.8800 1738.0600 600.3600 ;
        RECT 1793.0000 578.1200 1796.0000 578.6000 ;
        RECT 1793.0000 583.5600 1796.0000 584.0400 ;
        RECT 1781.4600 578.1200 1783.0600 578.6000 ;
        RECT 1781.4600 583.5600 1783.0600 584.0400 ;
        RECT 1793.0000 561.8000 1796.0000 562.2800 ;
        RECT 1793.0000 567.2400 1796.0000 567.7200 ;
        RECT 1793.0000 572.6800 1796.0000 573.1600 ;
        RECT 1781.4600 561.8000 1783.0600 562.2800 ;
        RECT 1781.4600 567.2400 1783.0600 567.7200 ;
        RECT 1781.4600 572.6800 1783.0600 573.1600 ;
        RECT 1793.0000 550.9200 1796.0000 551.4000 ;
        RECT 1793.0000 556.3600 1796.0000 556.8400 ;
        RECT 1781.4600 550.9200 1783.0600 551.4000 ;
        RECT 1781.4600 556.3600 1783.0600 556.8400 ;
        RECT 1793.0000 545.4800 1796.0000 545.9600 ;
        RECT 1781.4600 545.4800 1783.0600 545.9600 ;
        RECT 1736.4600 578.1200 1738.0600 578.6000 ;
        RECT 1736.4600 583.5600 1738.0600 584.0400 ;
        RECT 1736.4600 561.8000 1738.0600 562.2800 ;
        RECT 1736.4600 567.2400 1738.0600 567.7200 ;
        RECT 1736.4600 572.6800 1738.0600 573.1600 ;
        RECT 1736.4600 550.9200 1738.0600 551.4000 ;
        RECT 1736.4600 556.3600 1738.0600 556.8400 ;
        RECT 1736.4600 545.4800 1738.0600 545.9600 ;
        RECT 1691.4600 632.5200 1693.0600 633.0000 ;
        RECT 1691.4600 637.9600 1693.0600 638.4400 ;
        RECT 1691.4600 616.2000 1693.0600 616.6800 ;
        RECT 1691.4600 621.6400 1693.0600 622.1200 ;
        RECT 1691.4600 627.0800 1693.0600 627.5600 ;
        RECT 1646.4600 632.5200 1648.0600 633.0000 ;
        RECT 1646.4600 637.9600 1648.0600 638.4400 ;
        RECT 1646.4600 616.2000 1648.0600 616.6800 ;
        RECT 1646.4600 621.6400 1648.0600 622.1200 ;
        RECT 1646.4600 627.0800 1648.0600 627.5600 ;
        RECT 1691.4600 605.3200 1693.0600 605.8000 ;
        RECT 1691.4600 610.7600 1693.0600 611.2400 ;
        RECT 1691.4600 589.0000 1693.0600 589.4800 ;
        RECT 1691.4600 594.4400 1693.0600 594.9200 ;
        RECT 1691.4600 599.8800 1693.0600 600.3600 ;
        RECT 1646.4600 605.3200 1648.0600 605.8000 ;
        RECT 1646.4600 610.7600 1648.0600 611.2400 ;
        RECT 1646.4600 589.0000 1648.0600 589.4800 ;
        RECT 1646.4600 594.4400 1648.0600 594.9200 ;
        RECT 1646.4600 599.8800 1648.0600 600.3600 ;
        RECT 1596.9000 632.5200 1599.9000 633.0000 ;
        RECT 1596.9000 637.9600 1599.9000 638.4400 ;
        RECT 1596.9000 621.6400 1599.9000 622.1200 ;
        RECT 1596.9000 616.2000 1599.9000 616.6800 ;
        RECT 1596.9000 627.0800 1599.9000 627.5600 ;
        RECT 1596.9000 605.3200 1599.9000 605.8000 ;
        RECT 1596.9000 610.7600 1599.9000 611.2400 ;
        RECT 1596.9000 594.4400 1599.9000 594.9200 ;
        RECT 1596.9000 589.0000 1599.9000 589.4800 ;
        RECT 1596.9000 599.8800 1599.9000 600.3600 ;
        RECT 1691.4600 578.1200 1693.0600 578.6000 ;
        RECT 1691.4600 583.5600 1693.0600 584.0400 ;
        RECT 1691.4600 561.8000 1693.0600 562.2800 ;
        RECT 1691.4600 567.2400 1693.0600 567.7200 ;
        RECT 1691.4600 572.6800 1693.0600 573.1600 ;
        RECT 1646.4600 578.1200 1648.0600 578.6000 ;
        RECT 1646.4600 583.5600 1648.0600 584.0400 ;
        RECT 1646.4600 561.8000 1648.0600 562.2800 ;
        RECT 1646.4600 567.2400 1648.0600 567.7200 ;
        RECT 1646.4600 572.6800 1648.0600 573.1600 ;
        RECT 1691.4600 556.3600 1693.0600 556.8400 ;
        RECT 1691.4600 550.9200 1693.0600 551.4000 ;
        RECT 1691.4600 545.4800 1693.0600 545.9600 ;
        RECT 1646.4600 556.3600 1648.0600 556.8400 ;
        RECT 1646.4600 550.9200 1648.0600 551.4000 ;
        RECT 1646.4600 545.4800 1648.0600 545.9600 ;
        RECT 1596.9000 578.1200 1599.9000 578.6000 ;
        RECT 1596.9000 583.5600 1599.9000 584.0400 ;
        RECT 1596.9000 567.2400 1599.9000 567.7200 ;
        RECT 1596.9000 561.8000 1599.9000 562.2800 ;
        RECT 1596.9000 572.6800 1599.9000 573.1600 ;
        RECT 1596.9000 550.9200 1599.9000 551.4000 ;
        RECT 1596.9000 556.3600 1599.9000 556.8400 ;
        RECT 1596.9000 545.4800 1599.9000 545.9600 ;
        RECT 1596.9000 743.6700 1796.0000 746.6700 ;
        RECT 1596.9000 538.5700 1796.0000 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 308.9300 1783.0600 517.0300 ;
        RECT 1736.4600 308.9300 1738.0600 517.0300 ;
        RECT 1691.4600 308.9300 1693.0600 517.0300 ;
        RECT 1646.4600 308.9300 1648.0600 517.0300 ;
        RECT 1793.0000 308.9300 1796.0000 517.0300 ;
        RECT 1596.9000 308.9300 1599.9000 517.0300 ;
      LAYER met3 ;
        RECT 1793.0000 511.6800 1796.0000 512.1600 ;
        RECT 1781.4600 511.6800 1783.0600 512.1600 ;
        RECT 1793.0000 500.8000 1796.0000 501.2800 ;
        RECT 1793.0000 506.2400 1796.0000 506.7200 ;
        RECT 1781.4600 500.8000 1783.0600 501.2800 ;
        RECT 1781.4600 506.2400 1783.0600 506.7200 ;
        RECT 1793.0000 484.4800 1796.0000 484.9600 ;
        RECT 1793.0000 489.9200 1796.0000 490.4000 ;
        RECT 1781.4600 484.4800 1783.0600 484.9600 ;
        RECT 1781.4600 489.9200 1783.0600 490.4000 ;
        RECT 1793.0000 473.6000 1796.0000 474.0800 ;
        RECT 1793.0000 479.0400 1796.0000 479.5200 ;
        RECT 1781.4600 473.6000 1783.0600 474.0800 ;
        RECT 1781.4600 479.0400 1783.0600 479.5200 ;
        RECT 1793.0000 495.3600 1796.0000 495.8400 ;
        RECT 1781.4600 495.3600 1783.0600 495.8400 ;
        RECT 1736.4600 500.8000 1738.0600 501.2800 ;
        RECT 1736.4600 506.2400 1738.0600 506.7200 ;
        RECT 1736.4600 511.6800 1738.0600 512.1600 ;
        RECT 1736.4600 484.4800 1738.0600 484.9600 ;
        RECT 1736.4600 489.9200 1738.0600 490.4000 ;
        RECT 1736.4600 479.0400 1738.0600 479.5200 ;
        RECT 1736.4600 473.6000 1738.0600 474.0800 ;
        RECT 1736.4600 495.3600 1738.0600 495.8400 ;
        RECT 1793.0000 457.2800 1796.0000 457.7600 ;
        RECT 1793.0000 462.7200 1796.0000 463.2000 ;
        RECT 1781.4600 457.2800 1783.0600 457.7600 ;
        RECT 1781.4600 462.7200 1783.0600 463.2000 ;
        RECT 1793.0000 440.9600 1796.0000 441.4400 ;
        RECT 1793.0000 446.4000 1796.0000 446.8800 ;
        RECT 1793.0000 451.8400 1796.0000 452.3200 ;
        RECT 1781.4600 440.9600 1783.0600 441.4400 ;
        RECT 1781.4600 446.4000 1783.0600 446.8800 ;
        RECT 1781.4600 451.8400 1783.0600 452.3200 ;
        RECT 1793.0000 430.0800 1796.0000 430.5600 ;
        RECT 1793.0000 435.5200 1796.0000 436.0000 ;
        RECT 1781.4600 430.0800 1783.0600 430.5600 ;
        RECT 1781.4600 435.5200 1783.0600 436.0000 ;
        RECT 1793.0000 413.7600 1796.0000 414.2400 ;
        RECT 1793.0000 419.2000 1796.0000 419.6800 ;
        RECT 1793.0000 424.6400 1796.0000 425.1200 ;
        RECT 1781.4600 413.7600 1783.0600 414.2400 ;
        RECT 1781.4600 419.2000 1783.0600 419.6800 ;
        RECT 1781.4600 424.6400 1783.0600 425.1200 ;
        RECT 1736.4600 457.2800 1738.0600 457.7600 ;
        RECT 1736.4600 462.7200 1738.0600 463.2000 ;
        RECT 1736.4600 440.9600 1738.0600 441.4400 ;
        RECT 1736.4600 446.4000 1738.0600 446.8800 ;
        RECT 1736.4600 451.8400 1738.0600 452.3200 ;
        RECT 1736.4600 430.0800 1738.0600 430.5600 ;
        RECT 1736.4600 435.5200 1738.0600 436.0000 ;
        RECT 1736.4600 413.7600 1738.0600 414.2400 ;
        RECT 1736.4600 419.2000 1738.0600 419.6800 ;
        RECT 1736.4600 424.6400 1738.0600 425.1200 ;
        RECT 1793.0000 468.1600 1796.0000 468.6400 ;
        RECT 1736.4600 468.1600 1738.0600 468.6400 ;
        RECT 1781.4600 468.1600 1783.0600 468.6400 ;
        RECT 1691.4600 500.8000 1693.0600 501.2800 ;
        RECT 1691.4600 506.2400 1693.0600 506.7200 ;
        RECT 1691.4600 511.6800 1693.0600 512.1600 ;
        RECT 1646.4600 500.8000 1648.0600 501.2800 ;
        RECT 1646.4600 506.2400 1648.0600 506.7200 ;
        RECT 1646.4600 511.6800 1648.0600 512.1600 ;
        RECT 1691.4600 484.4800 1693.0600 484.9600 ;
        RECT 1691.4600 489.9200 1693.0600 490.4000 ;
        RECT 1691.4600 473.6000 1693.0600 474.0800 ;
        RECT 1691.4600 479.0400 1693.0600 479.5200 ;
        RECT 1646.4600 484.4800 1648.0600 484.9600 ;
        RECT 1646.4600 489.9200 1648.0600 490.4000 ;
        RECT 1646.4600 473.6000 1648.0600 474.0800 ;
        RECT 1646.4600 479.0400 1648.0600 479.5200 ;
        RECT 1646.4600 495.3600 1648.0600 495.8400 ;
        RECT 1691.4600 495.3600 1693.0600 495.8400 ;
        RECT 1596.9000 511.6800 1599.9000 512.1600 ;
        RECT 1596.9000 506.2400 1599.9000 506.7200 ;
        RECT 1596.9000 500.8000 1599.9000 501.2800 ;
        RECT 1596.9000 489.9200 1599.9000 490.4000 ;
        RECT 1596.9000 484.4800 1599.9000 484.9600 ;
        RECT 1596.9000 479.0400 1599.9000 479.5200 ;
        RECT 1596.9000 473.6000 1599.9000 474.0800 ;
        RECT 1596.9000 495.3600 1599.9000 495.8400 ;
        RECT 1691.4600 457.2800 1693.0600 457.7600 ;
        RECT 1691.4600 462.7200 1693.0600 463.2000 ;
        RECT 1691.4600 440.9600 1693.0600 441.4400 ;
        RECT 1691.4600 446.4000 1693.0600 446.8800 ;
        RECT 1691.4600 451.8400 1693.0600 452.3200 ;
        RECT 1646.4600 457.2800 1648.0600 457.7600 ;
        RECT 1646.4600 462.7200 1648.0600 463.2000 ;
        RECT 1646.4600 440.9600 1648.0600 441.4400 ;
        RECT 1646.4600 446.4000 1648.0600 446.8800 ;
        RECT 1646.4600 451.8400 1648.0600 452.3200 ;
        RECT 1691.4600 430.0800 1693.0600 430.5600 ;
        RECT 1691.4600 435.5200 1693.0600 436.0000 ;
        RECT 1691.4600 413.7600 1693.0600 414.2400 ;
        RECT 1691.4600 419.2000 1693.0600 419.6800 ;
        RECT 1691.4600 424.6400 1693.0600 425.1200 ;
        RECT 1646.4600 430.0800 1648.0600 430.5600 ;
        RECT 1646.4600 435.5200 1648.0600 436.0000 ;
        RECT 1646.4600 413.7600 1648.0600 414.2400 ;
        RECT 1646.4600 419.2000 1648.0600 419.6800 ;
        RECT 1646.4600 424.6400 1648.0600 425.1200 ;
        RECT 1596.9000 457.2800 1599.9000 457.7600 ;
        RECT 1596.9000 462.7200 1599.9000 463.2000 ;
        RECT 1596.9000 446.4000 1599.9000 446.8800 ;
        RECT 1596.9000 440.9600 1599.9000 441.4400 ;
        RECT 1596.9000 451.8400 1599.9000 452.3200 ;
        RECT 1596.9000 430.0800 1599.9000 430.5600 ;
        RECT 1596.9000 435.5200 1599.9000 436.0000 ;
        RECT 1596.9000 419.2000 1599.9000 419.6800 ;
        RECT 1596.9000 413.7600 1599.9000 414.2400 ;
        RECT 1596.9000 424.6400 1599.9000 425.1200 ;
        RECT 1596.9000 468.1600 1599.9000 468.6400 ;
        RECT 1646.4600 468.1600 1648.0600 468.6400 ;
        RECT 1691.4600 468.1600 1693.0600 468.6400 ;
        RECT 1793.0000 402.8800 1796.0000 403.3600 ;
        RECT 1793.0000 408.3200 1796.0000 408.8000 ;
        RECT 1781.4600 402.8800 1783.0600 403.3600 ;
        RECT 1781.4600 408.3200 1783.0600 408.8000 ;
        RECT 1793.0000 386.5600 1796.0000 387.0400 ;
        RECT 1793.0000 392.0000 1796.0000 392.4800 ;
        RECT 1793.0000 397.4400 1796.0000 397.9200 ;
        RECT 1781.4600 386.5600 1783.0600 387.0400 ;
        RECT 1781.4600 392.0000 1783.0600 392.4800 ;
        RECT 1781.4600 397.4400 1783.0600 397.9200 ;
        RECT 1793.0000 375.6800 1796.0000 376.1600 ;
        RECT 1793.0000 381.1200 1796.0000 381.6000 ;
        RECT 1781.4600 375.6800 1783.0600 376.1600 ;
        RECT 1781.4600 381.1200 1783.0600 381.6000 ;
        RECT 1793.0000 359.3600 1796.0000 359.8400 ;
        RECT 1793.0000 364.8000 1796.0000 365.2800 ;
        RECT 1793.0000 370.2400 1796.0000 370.7200 ;
        RECT 1781.4600 359.3600 1783.0600 359.8400 ;
        RECT 1781.4600 364.8000 1783.0600 365.2800 ;
        RECT 1781.4600 370.2400 1783.0600 370.7200 ;
        RECT 1736.4600 402.8800 1738.0600 403.3600 ;
        RECT 1736.4600 408.3200 1738.0600 408.8000 ;
        RECT 1736.4600 386.5600 1738.0600 387.0400 ;
        RECT 1736.4600 392.0000 1738.0600 392.4800 ;
        RECT 1736.4600 397.4400 1738.0600 397.9200 ;
        RECT 1736.4600 375.6800 1738.0600 376.1600 ;
        RECT 1736.4600 381.1200 1738.0600 381.6000 ;
        RECT 1736.4600 359.3600 1738.0600 359.8400 ;
        RECT 1736.4600 364.8000 1738.0600 365.2800 ;
        RECT 1736.4600 370.2400 1738.0600 370.7200 ;
        RECT 1793.0000 348.4800 1796.0000 348.9600 ;
        RECT 1793.0000 353.9200 1796.0000 354.4000 ;
        RECT 1781.4600 348.4800 1783.0600 348.9600 ;
        RECT 1781.4600 353.9200 1783.0600 354.4000 ;
        RECT 1793.0000 332.1600 1796.0000 332.6400 ;
        RECT 1793.0000 337.6000 1796.0000 338.0800 ;
        RECT 1793.0000 343.0400 1796.0000 343.5200 ;
        RECT 1781.4600 332.1600 1783.0600 332.6400 ;
        RECT 1781.4600 337.6000 1783.0600 338.0800 ;
        RECT 1781.4600 343.0400 1783.0600 343.5200 ;
        RECT 1793.0000 321.2800 1796.0000 321.7600 ;
        RECT 1793.0000 326.7200 1796.0000 327.2000 ;
        RECT 1781.4600 321.2800 1783.0600 321.7600 ;
        RECT 1781.4600 326.7200 1783.0600 327.2000 ;
        RECT 1793.0000 315.8400 1796.0000 316.3200 ;
        RECT 1781.4600 315.8400 1783.0600 316.3200 ;
        RECT 1736.4600 348.4800 1738.0600 348.9600 ;
        RECT 1736.4600 353.9200 1738.0600 354.4000 ;
        RECT 1736.4600 332.1600 1738.0600 332.6400 ;
        RECT 1736.4600 337.6000 1738.0600 338.0800 ;
        RECT 1736.4600 343.0400 1738.0600 343.5200 ;
        RECT 1736.4600 321.2800 1738.0600 321.7600 ;
        RECT 1736.4600 326.7200 1738.0600 327.2000 ;
        RECT 1736.4600 315.8400 1738.0600 316.3200 ;
        RECT 1691.4600 402.8800 1693.0600 403.3600 ;
        RECT 1691.4600 408.3200 1693.0600 408.8000 ;
        RECT 1691.4600 386.5600 1693.0600 387.0400 ;
        RECT 1691.4600 392.0000 1693.0600 392.4800 ;
        RECT 1691.4600 397.4400 1693.0600 397.9200 ;
        RECT 1646.4600 402.8800 1648.0600 403.3600 ;
        RECT 1646.4600 408.3200 1648.0600 408.8000 ;
        RECT 1646.4600 386.5600 1648.0600 387.0400 ;
        RECT 1646.4600 392.0000 1648.0600 392.4800 ;
        RECT 1646.4600 397.4400 1648.0600 397.9200 ;
        RECT 1691.4600 375.6800 1693.0600 376.1600 ;
        RECT 1691.4600 381.1200 1693.0600 381.6000 ;
        RECT 1691.4600 359.3600 1693.0600 359.8400 ;
        RECT 1691.4600 364.8000 1693.0600 365.2800 ;
        RECT 1691.4600 370.2400 1693.0600 370.7200 ;
        RECT 1646.4600 375.6800 1648.0600 376.1600 ;
        RECT 1646.4600 381.1200 1648.0600 381.6000 ;
        RECT 1646.4600 359.3600 1648.0600 359.8400 ;
        RECT 1646.4600 364.8000 1648.0600 365.2800 ;
        RECT 1646.4600 370.2400 1648.0600 370.7200 ;
        RECT 1596.9000 402.8800 1599.9000 403.3600 ;
        RECT 1596.9000 408.3200 1599.9000 408.8000 ;
        RECT 1596.9000 392.0000 1599.9000 392.4800 ;
        RECT 1596.9000 386.5600 1599.9000 387.0400 ;
        RECT 1596.9000 397.4400 1599.9000 397.9200 ;
        RECT 1596.9000 375.6800 1599.9000 376.1600 ;
        RECT 1596.9000 381.1200 1599.9000 381.6000 ;
        RECT 1596.9000 364.8000 1599.9000 365.2800 ;
        RECT 1596.9000 359.3600 1599.9000 359.8400 ;
        RECT 1596.9000 370.2400 1599.9000 370.7200 ;
        RECT 1691.4600 348.4800 1693.0600 348.9600 ;
        RECT 1691.4600 353.9200 1693.0600 354.4000 ;
        RECT 1691.4600 332.1600 1693.0600 332.6400 ;
        RECT 1691.4600 337.6000 1693.0600 338.0800 ;
        RECT 1691.4600 343.0400 1693.0600 343.5200 ;
        RECT 1646.4600 348.4800 1648.0600 348.9600 ;
        RECT 1646.4600 353.9200 1648.0600 354.4000 ;
        RECT 1646.4600 332.1600 1648.0600 332.6400 ;
        RECT 1646.4600 337.6000 1648.0600 338.0800 ;
        RECT 1646.4600 343.0400 1648.0600 343.5200 ;
        RECT 1691.4600 326.7200 1693.0600 327.2000 ;
        RECT 1691.4600 321.2800 1693.0600 321.7600 ;
        RECT 1691.4600 315.8400 1693.0600 316.3200 ;
        RECT 1646.4600 326.7200 1648.0600 327.2000 ;
        RECT 1646.4600 321.2800 1648.0600 321.7600 ;
        RECT 1646.4600 315.8400 1648.0600 316.3200 ;
        RECT 1596.9000 348.4800 1599.9000 348.9600 ;
        RECT 1596.9000 353.9200 1599.9000 354.4000 ;
        RECT 1596.9000 337.6000 1599.9000 338.0800 ;
        RECT 1596.9000 332.1600 1599.9000 332.6400 ;
        RECT 1596.9000 343.0400 1599.9000 343.5200 ;
        RECT 1596.9000 321.2800 1599.9000 321.7600 ;
        RECT 1596.9000 326.7200 1599.9000 327.2000 ;
        RECT 1596.9000 315.8400 1599.9000 316.3200 ;
        RECT 1596.9000 514.0300 1796.0000 517.0300 ;
        RECT 1596.9000 308.9300 1796.0000 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 79.2900 1783.0600 287.3900 ;
        RECT 1736.4600 79.2900 1738.0600 287.3900 ;
        RECT 1691.4600 79.2900 1693.0600 287.3900 ;
        RECT 1646.4600 79.2900 1648.0600 287.3900 ;
        RECT 1793.0000 79.2900 1796.0000 287.3900 ;
        RECT 1596.9000 79.2900 1599.9000 287.3900 ;
      LAYER met3 ;
        RECT 1793.0000 282.0400 1796.0000 282.5200 ;
        RECT 1781.4600 282.0400 1783.0600 282.5200 ;
        RECT 1793.0000 271.1600 1796.0000 271.6400 ;
        RECT 1793.0000 276.6000 1796.0000 277.0800 ;
        RECT 1781.4600 271.1600 1783.0600 271.6400 ;
        RECT 1781.4600 276.6000 1783.0600 277.0800 ;
        RECT 1793.0000 254.8400 1796.0000 255.3200 ;
        RECT 1793.0000 260.2800 1796.0000 260.7600 ;
        RECT 1781.4600 254.8400 1783.0600 255.3200 ;
        RECT 1781.4600 260.2800 1783.0600 260.7600 ;
        RECT 1793.0000 243.9600 1796.0000 244.4400 ;
        RECT 1793.0000 249.4000 1796.0000 249.8800 ;
        RECT 1781.4600 243.9600 1783.0600 244.4400 ;
        RECT 1781.4600 249.4000 1783.0600 249.8800 ;
        RECT 1793.0000 265.7200 1796.0000 266.2000 ;
        RECT 1781.4600 265.7200 1783.0600 266.2000 ;
        RECT 1736.4600 271.1600 1738.0600 271.6400 ;
        RECT 1736.4600 276.6000 1738.0600 277.0800 ;
        RECT 1736.4600 282.0400 1738.0600 282.5200 ;
        RECT 1736.4600 254.8400 1738.0600 255.3200 ;
        RECT 1736.4600 260.2800 1738.0600 260.7600 ;
        RECT 1736.4600 249.4000 1738.0600 249.8800 ;
        RECT 1736.4600 243.9600 1738.0600 244.4400 ;
        RECT 1736.4600 265.7200 1738.0600 266.2000 ;
        RECT 1793.0000 227.6400 1796.0000 228.1200 ;
        RECT 1793.0000 233.0800 1796.0000 233.5600 ;
        RECT 1781.4600 227.6400 1783.0600 228.1200 ;
        RECT 1781.4600 233.0800 1783.0600 233.5600 ;
        RECT 1793.0000 211.3200 1796.0000 211.8000 ;
        RECT 1793.0000 216.7600 1796.0000 217.2400 ;
        RECT 1793.0000 222.2000 1796.0000 222.6800 ;
        RECT 1781.4600 211.3200 1783.0600 211.8000 ;
        RECT 1781.4600 216.7600 1783.0600 217.2400 ;
        RECT 1781.4600 222.2000 1783.0600 222.6800 ;
        RECT 1793.0000 200.4400 1796.0000 200.9200 ;
        RECT 1793.0000 205.8800 1796.0000 206.3600 ;
        RECT 1781.4600 200.4400 1783.0600 200.9200 ;
        RECT 1781.4600 205.8800 1783.0600 206.3600 ;
        RECT 1793.0000 184.1200 1796.0000 184.6000 ;
        RECT 1793.0000 189.5600 1796.0000 190.0400 ;
        RECT 1793.0000 195.0000 1796.0000 195.4800 ;
        RECT 1781.4600 184.1200 1783.0600 184.6000 ;
        RECT 1781.4600 189.5600 1783.0600 190.0400 ;
        RECT 1781.4600 195.0000 1783.0600 195.4800 ;
        RECT 1736.4600 227.6400 1738.0600 228.1200 ;
        RECT 1736.4600 233.0800 1738.0600 233.5600 ;
        RECT 1736.4600 211.3200 1738.0600 211.8000 ;
        RECT 1736.4600 216.7600 1738.0600 217.2400 ;
        RECT 1736.4600 222.2000 1738.0600 222.6800 ;
        RECT 1736.4600 200.4400 1738.0600 200.9200 ;
        RECT 1736.4600 205.8800 1738.0600 206.3600 ;
        RECT 1736.4600 184.1200 1738.0600 184.6000 ;
        RECT 1736.4600 189.5600 1738.0600 190.0400 ;
        RECT 1736.4600 195.0000 1738.0600 195.4800 ;
        RECT 1793.0000 238.5200 1796.0000 239.0000 ;
        RECT 1736.4600 238.5200 1738.0600 239.0000 ;
        RECT 1781.4600 238.5200 1783.0600 239.0000 ;
        RECT 1691.4600 271.1600 1693.0600 271.6400 ;
        RECT 1691.4600 276.6000 1693.0600 277.0800 ;
        RECT 1691.4600 282.0400 1693.0600 282.5200 ;
        RECT 1646.4600 271.1600 1648.0600 271.6400 ;
        RECT 1646.4600 276.6000 1648.0600 277.0800 ;
        RECT 1646.4600 282.0400 1648.0600 282.5200 ;
        RECT 1691.4600 254.8400 1693.0600 255.3200 ;
        RECT 1691.4600 260.2800 1693.0600 260.7600 ;
        RECT 1691.4600 243.9600 1693.0600 244.4400 ;
        RECT 1691.4600 249.4000 1693.0600 249.8800 ;
        RECT 1646.4600 254.8400 1648.0600 255.3200 ;
        RECT 1646.4600 260.2800 1648.0600 260.7600 ;
        RECT 1646.4600 243.9600 1648.0600 244.4400 ;
        RECT 1646.4600 249.4000 1648.0600 249.8800 ;
        RECT 1646.4600 265.7200 1648.0600 266.2000 ;
        RECT 1691.4600 265.7200 1693.0600 266.2000 ;
        RECT 1596.9000 282.0400 1599.9000 282.5200 ;
        RECT 1596.9000 276.6000 1599.9000 277.0800 ;
        RECT 1596.9000 271.1600 1599.9000 271.6400 ;
        RECT 1596.9000 260.2800 1599.9000 260.7600 ;
        RECT 1596.9000 254.8400 1599.9000 255.3200 ;
        RECT 1596.9000 249.4000 1599.9000 249.8800 ;
        RECT 1596.9000 243.9600 1599.9000 244.4400 ;
        RECT 1596.9000 265.7200 1599.9000 266.2000 ;
        RECT 1691.4600 227.6400 1693.0600 228.1200 ;
        RECT 1691.4600 233.0800 1693.0600 233.5600 ;
        RECT 1691.4600 211.3200 1693.0600 211.8000 ;
        RECT 1691.4600 216.7600 1693.0600 217.2400 ;
        RECT 1691.4600 222.2000 1693.0600 222.6800 ;
        RECT 1646.4600 227.6400 1648.0600 228.1200 ;
        RECT 1646.4600 233.0800 1648.0600 233.5600 ;
        RECT 1646.4600 211.3200 1648.0600 211.8000 ;
        RECT 1646.4600 216.7600 1648.0600 217.2400 ;
        RECT 1646.4600 222.2000 1648.0600 222.6800 ;
        RECT 1691.4600 200.4400 1693.0600 200.9200 ;
        RECT 1691.4600 205.8800 1693.0600 206.3600 ;
        RECT 1691.4600 184.1200 1693.0600 184.6000 ;
        RECT 1691.4600 189.5600 1693.0600 190.0400 ;
        RECT 1691.4600 195.0000 1693.0600 195.4800 ;
        RECT 1646.4600 200.4400 1648.0600 200.9200 ;
        RECT 1646.4600 205.8800 1648.0600 206.3600 ;
        RECT 1646.4600 184.1200 1648.0600 184.6000 ;
        RECT 1646.4600 189.5600 1648.0600 190.0400 ;
        RECT 1646.4600 195.0000 1648.0600 195.4800 ;
        RECT 1596.9000 227.6400 1599.9000 228.1200 ;
        RECT 1596.9000 233.0800 1599.9000 233.5600 ;
        RECT 1596.9000 216.7600 1599.9000 217.2400 ;
        RECT 1596.9000 211.3200 1599.9000 211.8000 ;
        RECT 1596.9000 222.2000 1599.9000 222.6800 ;
        RECT 1596.9000 200.4400 1599.9000 200.9200 ;
        RECT 1596.9000 205.8800 1599.9000 206.3600 ;
        RECT 1596.9000 189.5600 1599.9000 190.0400 ;
        RECT 1596.9000 184.1200 1599.9000 184.6000 ;
        RECT 1596.9000 195.0000 1599.9000 195.4800 ;
        RECT 1596.9000 238.5200 1599.9000 239.0000 ;
        RECT 1646.4600 238.5200 1648.0600 239.0000 ;
        RECT 1691.4600 238.5200 1693.0600 239.0000 ;
        RECT 1793.0000 173.2400 1796.0000 173.7200 ;
        RECT 1793.0000 178.6800 1796.0000 179.1600 ;
        RECT 1781.4600 173.2400 1783.0600 173.7200 ;
        RECT 1781.4600 178.6800 1783.0600 179.1600 ;
        RECT 1793.0000 156.9200 1796.0000 157.4000 ;
        RECT 1793.0000 162.3600 1796.0000 162.8400 ;
        RECT 1793.0000 167.8000 1796.0000 168.2800 ;
        RECT 1781.4600 156.9200 1783.0600 157.4000 ;
        RECT 1781.4600 162.3600 1783.0600 162.8400 ;
        RECT 1781.4600 167.8000 1783.0600 168.2800 ;
        RECT 1793.0000 146.0400 1796.0000 146.5200 ;
        RECT 1793.0000 151.4800 1796.0000 151.9600 ;
        RECT 1781.4600 146.0400 1783.0600 146.5200 ;
        RECT 1781.4600 151.4800 1783.0600 151.9600 ;
        RECT 1793.0000 129.7200 1796.0000 130.2000 ;
        RECT 1793.0000 135.1600 1796.0000 135.6400 ;
        RECT 1793.0000 140.6000 1796.0000 141.0800 ;
        RECT 1781.4600 129.7200 1783.0600 130.2000 ;
        RECT 1781.4600 135.1600 1783.0600 135.6400 ;
        RECT 1781.4600 140.6000 1783.0600 141.0800 ;
        RECT 1736.4600 173.2400 1738.0600 173.7200 ;
        RECT 1736.4600 178.6800 1738.0600 179.1600 ;
        RECT 1736.4600 156.9200 1738.0600 157.4000 ;
        RECT 1736.4600 162.3600 1738.0600 162.8400 ;
        RECT 1736.4600 167.8000 1738.0600 168.2800 ;
        RECT 1736.4600 146.0400 1738.0600 146.5200 ;
        RECT 1736.4600 151.4800 1738.0600 151.9600 ;
        RECT 1736.4600 129.7200 1738.0600 130.2000 ;
        RECT 1736.4600 135.1600 1738.0600 135.6400 ;
        RECT 1736.4600 140.6000 1738.0600 141.0800 ;
        RECT 1793.0000 118.8400 1796.0000 119.3200 ;
        RECT 1793.0000 124.2800 1796.0000 124.7600 ;
        RECT 1781.4600 118.8400 1783.0600 119.3200 ;
        RECT 1781.4600 124.2800 1783.0600 124.7600 ;
        RECT 1793.0000 102.5200 1796.0000 103.0000 ;
        RECT 1793.0000 107.9600 1796.0000 108.4400 ;
        RECT 1793.0000 113.4000 1796.0000 113.8800 ;
        RECT 1781.4600 102.5200 1783.0600 103.0000 ;
        RECT 1781.4600 107.9600 1783.0600 108.4400 ;
        RECT 1781.4600 113.4000 1783.0600 113.8800 ;
        RECT 1793.0000 91.6400 1796.0000 92.1200 ;
        RECT 1793.0000 97.0800 1796.0000 97.5600 ;
        RECT 1781.4600 91.6400 1783.0600 92.1200 ;
        RECT 1781.4600 97.0800 1783.0600 97.5600 ;
        RECT 1793.0000 86.2000 1796.0000 86.6800 ;
        RECT 1781.4600 86.2000 1783.0600 86.6800 ;
        RECT 1736.4600 118.8400 1738.0600 119.3200 ;
        RECT 1736.4600 124.2800 1738.0600 124.7600 ;
        RECT 1736.4600 102.5200 1738.0600 103.0000 ;
        RECT 1736.4600 107.9600 1738.0600 108.4400 ;
        RECT 1736.4600 113.4000 1738.0600 113.8800 ;
        RECT 1736.4600 91.6400 1738.0600 92.1200 ;
        RECT 1736.4600 97.0800 1738.0600 97.5600 ;
        RECT 1736.4600 86.2000 1738.0600 86.6800 ;
        RECT 1691.4600 173.2400 1693.0600 173.7200 ;
        RECT 1691.4600 178.6800 1693.0600 179.1600 ;
        RECT 1691.4600 156.9200 1693.0600 157.4000 ;
        RECT 1691.4600 162.3600 1693.0600 162.8400 ;
        RECT 1691.4600 167.8000 1693.0600 168.2800 ;
        RECT 1646.4600 173.2400 1648.0600 173.7200 ;
        RECT 1646.4600 178.6800 1648.0600 179.1600 ;
        RECT 1646.4600 156.9200 1648.0600 157.4000 ;
        RECT 1646.4600 162.3600 1648.0600 162.8400 ;
        RECT 1646.4600 167.8000 1648.0600 168.2800 ;
        RECT 1691.4600 146.0400 1693.0600 146.5200 ;
        RECT 1691.4600 151.4800 1693.0600 151.9600 ;
        RECT 1691.4600 129.7200 1693.0600 130.2000 ;
        RECT 1691.4600 135.1600 1693.0600 135.6400 ;
        RECT 1691.4600 140.6000 1693.0600 141.0800 ;
        RECT 1646.4600 146.0400 1648.0600 146.5200 ;
        RECT 1646.4600 151.4800 1648.0600 151.9600 ;
        RECT 1646.4600 129.7200 1648.0600 130.2000 ;
        RECT 1646.4600 135.1600 1648.0600 135.6400 ;
        RECT 1646.4600 140.6000 1648.0600 141.0800 ;
        RECT 1596.9000 173.2400 1599.9000 173.7200 ;
        RECT 1596.9000 178.6800 1599.9000 179.1600 ;
        RECT 1596.9000 162.3600 1599.9000 162.8400 ;
        RECT 1596.9000 156.9200 1599.9000 157.4000 ;
        RECT 1596.9000 167.8000 1599.9000 168.2800 ;
        RECT 1596.9000 146.0400 1599.9000 146.5200 ;
        RECT 1596.9000 151.4800 1599.9000 151.9600 ;
        RECT 1596.9000 135.1600 1599.9000 135.6400 ;
        RECT 1596.9000 129.7200 1599.9000 130.2000 ;
        RECT 1596.9000 140.6000 1599.9000 141.0800 ;
        RECT 1691.4600 118.8400 1693.0600 119.3200 ;
        RECT 1691.4600 124.2800 1693.0600 124.7600 ;
        RECT 1691.4600 102.5200 1693.0600 103.0000 ;
        RECT 1691.4600 107.9600 1693.0600 108.4400 ;
        RECT 1691.4600 113.4000 1693.0600 113.8800 ;
        RECT 1646.4600 118.8400 1648.0600 119.3200 ;
        RECT 1646.4600 124.2800 1648.0600 124.7600 ;
        RECT 1646.4600 102.5200 1648.0600 103.0000 ;
        RECT 1646.4600 107.9600 1648.0600 108.4400 ;
        RECT 1646.4600 113.4000 1648.0600 113.8800 ;
        RECT 1691.4600 97.0800 1693.0600 97.5600 ;
        RECT 1691.4600 91.6400 1693.0600 92.1200 ;
        RECT 1691.4600 86.2000 1693.0600 86.6800 ;
        RECT 1646.4600 97.0800 1648.0600 97.5600 ;
        RECT 1646.4600 91.6400 1648.0600 92.1200 ;
        RECT 1646.4600 86.2000 1648.0600 86.6800 ;
        RECT 1596.9000 118.8400 1599.9000 119.3200 ;
        RECT 1596.9000 124.2800 1599.9000 124.7600 ;
        RECT 1596.9000 107.9600 1599.9000 108.4400 ;
        RECT 1596.9000 102.5200 1599.9000 103.0000 ;
        RECT 1596.9000 113.4000 1599.9000 113.8800 ;
        RECT 1596.9000 91.6400 1599.9000 92.1200 ;
        RECT 1596.9000 97.0800 1599.9000 97.5600 ;
        RECT 1596.9000 86.2000 1599.9000 86.6800 ;
        RECT 1596.9000 284.3900 1796.0000 287.3900 ;
        RECT 1596.9000 79.2900 1796.0000 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1596.9000 37.6700 1598.9000 58.6000 ;
        RECT 1794.0000 37.6700 1796.0000 58.6000 ;
      LAYER met3 ;
        RECT 1794.0000 54.1000 1796.0000 54.5800 ;
        RECT 1596.9000 54.1000 1598.9000 54.5800 ;
        RECT 1794.0000 43.2200 1796.0000 43.7000 ;
        RECT 1596.9000 43.2200 1598.9000 43.7000 ;
        RECT 1794.0000 48.6600 1796.0000 49.1400 ;
        RECT 1596.9000 48.6600 1598.9000 49.1400 ;
        RECT 1596.9000 56.6000 1796.0000 58.6000 ;
        RECT 1596.9000 37.6700 1796.0000 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 2605.3300 1783.0600 2813.4300 ;
        RECT 1736.4600 2605.3300 1738.0600 2813.4300 ;
        RECT 1691.4600 2605.3300 1693.0600 2813.4300 ;
        RECT 1646.4600 2605.3300 1648.0600 2813.4300 ;
        RECT 1793.0000 2605.3300 1796.0000 2813.4300 ;
        RECT 1596.9000 2605.3300 1599.9000 2813.4300 ;
      LAYER met3 ;
        RECT 1793.0000 2808.0800 1796.0000 2808.5600 ;
        RECT 1781.4600 2808.0800 1783.0600 2808.5600 ;
        RECT 1793.0000 2797.2000 1796.0000 2797.6800 ;
        RECT 1793.0000 2802.6400 1796.0000 2803.1200 ;
        RECT 1781.4600 2797.2000 1783.0600 2797.6800 ;
        RECT 1781.4600 2802.6400 1783.0600 2803.1200 ;
        RECT 1793.0000 2780.8800 1796.0000 2781.3600 ;
        RECT 1793.0000 2786.3200 1796.0000 2786.8000 ;
        RECT 1781.4600 2780.8800 1783.0600 2781.3600 ;
        RECT 1781.4600 2786.3200 1783.0600 2786.8000 ;
        RECT 1793.0000 2770.0000 1796.0000 2770.4800 ;
        RECT 1793.0000 2775.4400 1796.0000 2775.9200 ;
        RECT 1781.4600 2770.0000 1783.0600 2770.4800 ;
        RECT 1781.4600 2775.4400 1783.0600 2775.9200 ;
        RECT 1793.0000 2791.7600 1796.0000 2792.2400 ;
        RECT 1781.4600 2791.7600 1783.0600 2792.2400 ;
        RECT 1736.4600 2797.2000 1738.0600 2797.6800 ;
        RECT 1736.4600 2802.6400 1738.0600 2803.1200 ;
        RECT 1736.4600 2808.0800 1738.0600 2808.5600 ;
        RECT 1736.4600 2780.8800 1738.0600 2781.3600 ;
        RECT 1736.4600 2786.3200 1738.0600 2786.8000 ;
        RECT 1736.4600 2775.4400 1738.0600 2775.9200 ;
        RECT 1736.4600 2770.0000 1738.0600 2770.4800 ;
        RECT 1736.4600 2791.7600 1738.0600 2792.2400 ;
        RECT 1793.0000 2753.6800 1796.0000 2754.1600 ;
        RECT 1793.0000 2759.1200 1796.0000 2759.6000 ;
        RECT 1781.4600 2753.6800 1783.0600 2754.1600 ;
        RECT 1781.4600 2759.1200 1783.0600 2759.6000 ;
        RECT 1793.0000 2737.3600 1796.0000 2737.8400 ;
        RECT 1793.0000 2742.8000 1796.0000 2743.2800 ;
        RECT 1793.0000 2748.2400 1796.0000 2748.7200 ;
        RECT 1781.4600 2737.3600 1783.0600 2737.8400 ;
        RECT 1781.4600 2742.8000 1783.0600 2743.2800 ;
        RECT 1781.4600 2748.2400 1783.0600 2748.7200 ;
        RECT 1793.0000 2726.4800 1796.0000 2726.9600 ;
        RECT 1793.0000 2731.9200 1796.0000 2732.4000 ;
        RECT 1781.4600 2726.4800 1783.0600 2726.9600 ;
        RECT 1781.4600 2731.9200 1783.0600 2732.4000 ;
        RECT 1793.0000 2710.1600 1796.0000 2710.6400 ;
        RECT 1793.0000 2715.6000 1796.0000 2716.0800 ;
        RECT 1793.0000 2721.0400 1796.0000 2721.5200 ;
        RECT 1781.4600 2710.1600 1783.0600 2710.6400 ;
        RECT 1781.4600 2715.6000 1783.0600 2716.0800 ;
        RECT 1781.4600 2721.0400 1783.0600 2721.5200 ;
        RECT 1736.4600 2753.6800 1738.0600 2754.1600 ;
        RECT 1736.4600 2759.1200 1738.0600 2759.6000 ;
        RECT 1736.4600 2737.3600 1738.0600 2737.8400 ;
        RECT 1736.4600 2742.8000 1738.0600 2743.2800 ;
        RECT 1736.4600 2748.2400 1738.0600 2748.7200 ;
        RECT 1736.4600 2726.4800 1738.0600 2726.9600 ;
        RECT 1736.4600 2731.9200 1738.0600 2732.4000 ;
        RECT 1736.4600 2710.1600 1738.0600 2710.6400 ;
        RECT 1736.4600 2715.6000 1738.0600 2716.0800 ;
        RECT 1736.4600 2721.0400 1738.0600 2721.5200 ;
        RECT 1793.0000 2764.5600 1796.0000 2765.0400 ;
        RECT 1736.4600 2764.5600 1738.0600 2765.0400 ;
        RECT 1781.4600 2764.5600 1783.0600 2765.0400 ;
        RECT 1691.4600 2797.2000 1693.0600 2797.6800 ;
        RECT 1691.4600 2802.6400 1693.0600 2803.1200 ;
        RECT 1691.4600 2808.0800 1693.0600 2808.5600 ;
        RECT 1646.4600 2797.2000 1648.0600 2797.6800 ;
        RECT 1646.4600 2802.6400 1648.0600 2803.1200 ;
        RECT 1646.4600 2808.0800 1648.0600 2808.5600 ;
        RECT 1691.4600 2780.8800 1693.0600 2781.3600 ;
        RECT 1691.4600 2786.3200 1693.0600 2786.8000 ;
        RECT 1691.4600 2770.0000 1693.0600 2770.4800 ;
        RECT 1691.4600 2775.4400 1693.0600 2775.9200 ;
        RECT 1646.4600 2780.8800 1648.0600 2781.3600 ;
        RECT 1646.4600 2786.3200 1648.0600 2786.8000 ;
        RECT 1646.4600 2770.0000 1648.0600 2770.4800 ;
        RECT 1646.4600 2775.4400 1648.0600 2775.9200 ;
        RECT 1646.4600 2791.7600 1648.0600 2792.2400 ;
        RECT 1691.4600 2791.7600 1693.0600 2792.2400 ;
        RECT 1596.9000 2808.0800 1599.9000 2808.5600 ;
        RECT 1596.9000 2802.6400 1599.9000 2803.1200 ;
        RECT 1596.9000 2797.2000 1599.9000 2797.6800 ;
        RECT 1596.9000 2786.3200 1599.9000 2786.8000 ;
        RECT 1596.9000 2780.8800 1599.9000 2781.3600 ;
        RECT 1596.9000 2775.4400 1599.9000 2775.9200 ;
        RECT 1596.9000 2770.0000 1599.9000 2770.4800 ;
        RECT 1596.9000 2791.7600 1599.9000 2792.2400 ;
        RECT 1691.4600 2753.6800 1693.0600 2754.1600 ;
        RECT 1691.4600 2759.1200 1693.0600 2759.6000 ;
        RECT 1691.4600 2737.3600 1693.0600 2737.8400 ;
        RECT 1691.4600 2742.8000 1693.0600 2743.2800 ;
        RECT 1691.4600 2748.2400 1693.0600 2748.7200 ;
        RECT 1646.4600 2753.6800 1648.0600 2754.1600 ;
        RECT 1646.4600 2759.1200 1648.0600 2759.6000 ;
        RECT 1646.4600 2737.3600 1648.0600 2737.8400 ;
        RECT 1646.4600 2742.8000 1648.0600 2743.2800 ;
        RECT 1646.4600 2748.2400 1648.0600 2748.7200 ;
        RECT 1691.4600 2726.4800 1693.0600 2726.9600 ;
        RECT 1691.4600 2731.9200 1693.0600 2732.4000 ;
        RECT 1691.4600 2710.1600 1693.0600 2710.6400 ;
        RECT 1691.4600 2715.6000 1693.0600 2716.0800 ;
        RECT 1691.4600 2721.0400 1693.0600 2721.5200 ;
        RECT 1646.4600 2726.4800 1648.0600 2726.9600 ;
        RECT 1646.4600 2731.9200 1648.0600 2732.4000 ;
        RECT 1646.4600 2710.1600 1648.0600 2710.6400 ;
        RECT 1646.4600 2715.6000 1648.0600 2716.0800 ;
        RECT 1646.4600 2721.0400 1648.0600 2721.5200 ;
        RECT 1596.9000 2753.6800 1599.9000 2754.1600 ;
        RECT 1596.9000 2759.1200 1599.9000 2759.6000 ;
        RECT 1596.9000 2742.8000 1599.9000 2743.2800 ;
        RECT 1596.9000 2737.3600 1599.9000 2737.8400 ;
        RECT 1596.9000 2748.2400 1599.9000 2748.7200 ;
        RECT 1596.9000 2726.4800 1599.9000 2726.9600 ;
        RECT 1596.9000 2731.9200 1599.9000 2732.4000 ;
        RECT 1596.9000 2715.6000 1599.9000 2716.0800 ;
        RECT 1596.9000 2710.1600 1599.9000 2710.6400 ;
        RECT 1596.9000 2721.0400 1599.9000 2721.5200 ;
        RECT 1596.9000 2764.5600 1599.9000 2765.0400 ;
        RECT 1646.4600 2764.5600 1648.0600 2765.0400 ;
        RECT 1691.4600 2764.5600 1693.0600 2765.0400 ;
        RECT 1793.0000 2699.2800 1796.0000 2699.7600 ;
        RECT 1793.0000 2704.7200 1796.0000 2705.2000 ;
        RECT 1781.4600 2699.2800 1783.0600 2699.7600 ;
        RECT 1781.4600 2704.7200 1783.0600 2705.2000 ;
        RECT 1793.0000 2682.9600 1796.0000 2683.4400 ;
        RECT 1793.0000 2688.4000 1796.0000 2688.8800 ;
        RECT 1793.0000 2693.8400 1796.0000 2694.3200 ;
        RECT 1781.4600 2682.9600 1783.0600 2683.4400 ;
        RECT 1781.4600 2688.4000 1783.0600 2688.8800 ;
        RECT 1781.4600 2693.8400 1783.0600 2694.3200 ;
        RECT 1793.0000 2672.0800 1796.0000 2672.5600 ;
        RECT 1793.0000 2677.5200 1796.0000 2678.0000 ;
        RECT 1781.4600 2672.0800 1783.0600 2672.5600 ;
        RECT 1781.4600 2677.5200 1783.0600 2678.0000 ;
        RECT 1793.0000 2655.7600 1796.0000 2656.2400 ;
        RECT 1793.0000 2661.2000 1796.0000 2661.6800 ;
        RECT 1793.0000 2666.6400 1796.0000 2667.1200 ;
        RECT 1781.4600 2655.7600 1783.0600 2656.2400 ;
        RECT 1781.4600 2661.2000 1783.0600 2661.6800 ;
        RECT 1781.4600 2666.6400 1783.0600 2667.1200 ;
        RECT 1736.4600 2699.2800 1738.0600 2699.7600 ;
        RECT 1736.4600 2704.7200 1738.0600 2705.2000 ;
        RECT 1736.4600 2682.9600 1738.0600 2683.4400 ;
        RECT 1736.4600 2688.4000 1738.0600 2688.8800 ;
        RECT 1736.4600 2693.8400 1738.0600 2694.3200 ;
        RECT 1736.4600 2672.0800 1738.0600 2672.5600 ;
        RECT 1736.4600 2677.5200 1738.0600 2678.0000 ;
        RECT 1736.4600 2655.7600 1738.0600 2656.2400 ;
        RECT 1736.4600 2661.2000 1738.0600 2661.6800 ;
        RECT 1736.4600 2666.6400 1738.0600 2667.1200 ;
        RECT 1793.0000 2644.8800 1796.0000 2645.3600 ;
        RECT 1793.0000 2650.3200 1796.0000 2650.8000 ;
        RECT 1781.4600 2644.8800 1783.0600 2645.3600 ;
        RECT 1781.4600 2650.3200 1783.0600 2650.8000 ;
        RECT 1793.0000 2628.5600 1796.0000 2629.0400 ;
        RECT 1793.0000 2634.0000 1796.0000 2634.4800 ;
        RECT 1793.0000 2639.4400 1796.0000 2639.9200 ;
        RECT 1781.4600 2628.5600 1783.0600 2629.0400 ;
        RECT 1781.4600 2634.0000 1783.0600 2634.4800 ;
        RECT 1781.4600 2639.4400 1783.0600 2639.9200 ;
        RECT 1793.0000 2617.6800 1796.0000 2618.1600 ;
        RECT 1793.0000 2623.1200 1796.0000 2623.6000 ;
        RECT 1781.4600 2617.6800 1783.0600 2618.1600 ;
        RECT 1781.4600 2623.1200 1783.0600 2623.6000 ;
        RECT 1793.0000 2612.2400 1796.0000 2612.7200 ;
        RECT 1781.4600 2612.2400 1783.0600 2612.7200 ;
        RECT 1736.4600 2644.8800 1738.0600 2645.3600 ;
        RECT 1736.4600 2650.3200 1738.0600 2650.8000 ;
        RECT 1736.4600 2628.5600 1738.0600 2629.0400 ;
        RECT 1736.4600 2634.0000 1738.0600 2634.4800 ;
        RECT 1736.4600 2639.4400 1738.0600 2639.9200 ;
        RECT 1736.4600 2617.6800 1738.0600 2618.1600 ;
        RECT 1736.4600 2623.1200 1738.0600 2623.6000 ;
        RECT 1736.4600 2612.2400 1738.0600 2612.7200 ;
        RECT 1691.4600 2699.2800 1693.0600 2699.7600 ;
        RECT 1691.4600 2704.7200 1693.0600 2705.2000 ;
        RECT 1691.4600 2682.9600 1693.0600 2683.4400 ;
        RECT 1691.4600 2688.4000 1693.0600 2688.8800 ;
        RECT 1691.4600 2693.8400 1693.0600 2694.3200 ;
        RECT 1646.4600 2699.2800 1648.0600 2699.7600 ;
        RECT 1646.4600 2704.7200 1648.0600 2705.2000 ;
        RECT 1646.4600 2682.9600 1648.0600 2683.4400 ;
        RECT 1646.4600 2688.4000 1648.0600 2688.8800 ;
        RECT 1646.4600 2693.8400 1648.0600 2694.3200 ;
        RECT 1691.4600 2672.0800 1693.0600 2672.5600 ;
        RECT 1691.4600 2677.5200 1693.0600 2678.0000 ;
        RECT 1691.4600 2655.7600 1693.0600 2656.2400 ;
        RECT 1691.4600 2661.2000 1693.0600 2661.6800 ;
        RECT 1691.4600 2666.6400 1693.0600 2667.1200 ;
        RECT 1646.4600 2672.0800 1648.0600 2672.5600 ;
        RECT 1646.4600 2677.5200 1648.0600 2678.0000 ;
        RECT 1646.4600 2655.7600 1648.0600 2656.2400 ;
        RECT 1646.4600 2661.2000 1648.0600 2661.6800 ;
        RECT 1646.4600 2666.6400 1648.0600 2667.1200 ;
        RECT 1596.9000 2699.2800 1599.9000 2699.7600 ;
        RECT 1596.9000 2704.7200 1599.9000 2705.2000 ;
        RECT 1596.9000 2688.4000 1599.9000 2688.8800 ;
        RECT 1596.9000 2682.9600 1599.9000 2683.4400 ;
        RECT 1596.9000 2693.8400 1599.9000 2694.3200 ;
        RECT 1596.9000 2672.0800 1599.9000 2672.5600 ;
        RECT 1596.9000 2677.5200 1599.9000 2678.0000 ;
        RECT 1596.9000 2661.2000 1599.9000 2661.6800 ;
        RECT 1596.9000 2655.7600 1599.9000 2656.2400 ;
        RECT 1596.9000 2666.6400 1599.9000 2667.1200 ;
        RECT 1691.4600 2644.8800 1693.0600 2645.3600 ;
        RECT 1691.4600 2650.3200 1693.0600 2650.8000 ;
        RECT 1691.4600 2628.5600 1693.0600 2629.0400 ;
        RECT 1691.4600 2634.0000 1693.0600 2634.4800 ;
        RECT 1691.4600 2639.4400 1693.0600 2639.9200 ;
        RECT 1646.4600 2644.8800 1648.0600 2645.3600 ;
        RECT 1646.4600 2650.3200 1648.0600 2650.8000 ;
        RECT 1646.4600 2628.5600 1648.0600 2629.0400 ;
        RECT 1646.4600 2634.0000 1648.0600 2634.4800 ;
        RECT 1646.4600 2639.4400 1648.0600 2639.9200 ;
        RECT 1691.4600 2623.1200 1693.0600 2623.6000 ;
        RECT 1691.4600 2617.6800 1693.0600 2618.1600 ;
        RECT 1691.4600 2612.2400 1693.0600 2612.7200 ;
        RECT 1646.4600 2623.1200 1648.0600 2623.6000 ;
        RECT 1646.4600 2617.6800 1648.0600 2618.1600 ;
        RECT 1646.4600 2612.2400 1648.0600 2612.7200 ;
        RECT 1596.9000 2644.8800 1599.9000 2645.3600 ;
        RECT 1596.9000 2650.3200 1599.9000 2650.8000 ;
        RECT 1596.9000 2634.0000 1599.9000 2634.4800 ;
        RECT 1596.9000 2628.5600 1599.9000 2629.0400 ;
        RECT 1596.9000 2639.4400 1599.9000 2639.9200 ;
        RECT 1596.9000 2617.6800 1599.9000 2618.1600 ;
        RECT 1596.9000 2623.1200 1599.9000 2623.6000 ;
        RECT 1596.9000 2612.2400 1599.9000 2612.7200 ;
        RECT 1596.9000 2810.4300 1796.0000 2813.4300 ;
        RECT 1596.9000 2605.3300 1796.0000 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 2375.6900 1783.0600 2583.7900 ;
        RECT 1736.4600 2375.6900 1738.0600 2583.7900 ;
        RECT 1691.4600 2375.6900 1693.0600 2583.7900 ;
        RECT 1646.4600 2375.6900 1648.0600 2583.7900 ;
        RECT 1793.0000 2375.6900 1796.0000 2583.7900 ;
        RECT 1596.9000 2375.6900 1599.9000 2583.7900 ;
      LAYER met3 ;
        RECT 1793.0000 2578.4400 1796.0000 2578.9200 ;
        RECT 1781.4600 2578.4400 1783.0600 2578.9200 ;
        RECT 1793.0000 2567.5600 1796.0000 2568.0400 ;
        RECT 1793.0000 2573.0000 1796.0000 2573.4800 ;
        RECT 1781.4600 2567.5600 1783.0600 2568.0400 ;
        RECT 1781.4600 2573.0000 1783.0600 2573.4800 ;
        RECT 1793.0000 2551.2400 1796.0000 2551.7200 ;
        RECT 1793.0000 2556.6800 1796.0000 2557.1600 ;
        RECT 1781.4600 2551.2400 1783.0600 2551.7200 ;
        RECT 1781.4600 2556.6800 1783.0600 2557.1600 ;
        RECT 1793.0000 2540.3600 1796.0000 2540.8400 ;
        RECT 1793.0000 2545.8000 1796.0000 2546.2800 ;
        RECT 1781.4600 2540.3600 1783.0600 2540.8400 ;
        RECT 1781.4600 2545.8000 1783.0600 2546.2800 ;
        RECT 1793.0000 2562.1200 1796.0000 2562.6000 ;
        RECT 1781.4600 2562.1200 1783.0600 2562.6000 ;
        RECT 1736.4600 2567.5600 1738.0600 2568.0400 ;
        RECT 1736.4600 2573.0000 1738.0600 2573.4800 ;
        RECT 1736.4600 2578.4400 1738.0600 2578.9200 ;
        RECT 1736.4600 2551.2400 1738.0600 2551.7200 ;
        RECT 1736.4600 2556.6800 1738.0600 2557.1600 ;
        RECT 1736.4600 2545.8000 1738.0600 2546.2800 ;
        RECT 1736.4600 2540.3600 1738.0600 2540.8400 ;
        RECT 1736.4600 2562.1200 1738.0600 2562.6000 ;
        RECT 1793.0000 2524.0400 1796.0000 2524.5200 ;
        RECT 1793.0000 2529.4800 1796.0000 2529.9600 ;
        RECT 1781.4600 2524.0400 1783.0600 2524.5200 ;
        RECT 1781.4600 2529.4800 1783.0600 2529.9600 ;
        RECT 1793.0000 2507.7200 1796.0000 2508.2000 ;
        RECT 1793.0000 2513.1600 1796.0000 2513.6400 ;
        RECT 1793.0000 2518.6000 1796.0000 2519.0800 ;
        RECT 1781.4600 2507.7200 1783.0600 2508.2000 ;
        RECT 1781.4600 2513.1600 1783.0600 2513.6400 ;
        RECT 1781.4600 2518.6000 1783.0600 2519.0800 ;
        RECT 1793.0000 2496.8400 1796.0000 2497.3200 ;
        RECT 1793.0000 2502.2800 1796.0000 2502.7600 ;
        RECT 1781.4600 2496.8400 1783.0600 2497.3200 ;
        RECT 1781.4600 2502.2800 1783.0600 2502.7600 ;
        RECT 1793.0000 2480.5200 1796.0000 2481.0000 ;
        RECT 1793.0000 2485.9600 1796.0000 2486.4400 ;
        RECT 1793.0000 2491.4000 1796.0000 2491.8800 ;
        RECT 1781.4600 2480.5200 1783.0600 2481.0000 ;
        RECT 1781.4600 2485.9600 1783.0600 2486.4400 ;
        RECT 1781.4600 2491.4000 1783.0600 2491.8800 ;
        RECT 1736.4600 2524.0400 1738.0600 2524.5200 ;
        RECT 1736.4600 2529.4800 1738.0600 2529.9600 ;
        RECT 1736.4600 2507.7200 1738.0600 2508.2000 ;
        RECT 1736.4600 2513.1600 1738.0600 2513.6400 ;
        RECT 1736.4600 2518.6000 1738.0600 2519.0800 ;
        RECT 1736.4600 2496.8400 1738.0600 2497.3200 ;
        RECT 1736.4600 2502.2800 1738.0600 2502.7600 ;
        RECT 1736.4600 2480.5200 1738.0600 2481.0000 ;
        RECT 1736.4600 2485.9600 1738.0600 2486.4400 ;
        RECT 1736.4600 2491.4000 1738.0600 2491.8800 ;
        RECT 1793.0000 2534.9200 1796.0000 2535.4000 ;
        RECT 1736.4600 2534.9200 1738.0600 2535.4000 ;
        RECT 1781.4600 2534.9200 1783.0600 2535.4000 ;
        RECT 1691.4600 2567.5600 1693.0600 2568.0400 ;
        RECT 1691.4600 2573.0000 1693.0600 2573.4800 ;
        RECT 1691.4600 2578.4400 1693.0600 2578.9200 ;
        RECT 1646.4600 2567.5600 1648.0600 2568.0400 ;
        RECT 1646.4600 2573.0000 1648.0600 2573.4800 ;
        RECT 1646.4600 2578.4400 1648.0600 2578.9200 ;
        RECT 1691.4600 2551.2400 1693.0600 2551.7200 ;
        RECT 1691.4600 2556.6800 1693.0600 2557.1600 ;
        RECT 1691.4600 2540.3600 1693.0600 2540.8400 ;
        RECT 1691.4600 2545.8000 1693.0600 2546.2800 ;
        RECT 1646.4600 2551.2400 1648.0600 2551.7200 ;
        RECT 1646.4600 2556.6800 1648.0600 2557.1600 ;
        RECT 1646.4600 2540.3600 1648.0600 2540.8400 ;
        RECT 1646.4600 2545.8000 1648.0600 2546.2800 ;
        RECT 1646.4600 2562.1200 1648.0600 2562.6000 ;
        RECT 1691.4600 2562.1200 1693.0600 2562.6000 ;
        RECT 1596.9000 2578.4400 1599.9000 2578.9200 ;
        RECT 1596.9000 2573.0000 1599.9000 2573.4800 ;
        RECT 1596.9000 2567.5600 1599.9000 2568.0400 ;
        RECT 1596.9000 2556.6800 1599.9000 2557.1600 ;
        RECT 1596.9000 2551.2400 1599.9000 2551.7200 ;
        RECT 1596.9000 2545.8000 1599.9000 2546.2800 ;
        RECT 1596.9000 2540.3600 1599.9000 2540.8400 ;
        RECT 1596.9000 2562.1200 1599.9000 2562.6000 ;
        RECT 1691.4600 2524.0400 1693.0600 2524.5200 ;
        RECT 1691.4600 2529.4800 1693.0600 2529.9600 ;
        RECT 1691.4600 2507.7200 1693.0600 2508.2000 ;
        RECT 1691.4600 2513.1600 1693.0600 2513.6400 ;
        RECT 1691.4600 2518.6000 1693.0600 2519.0800 ;
        RECT 1646.4600 2524.0400 1648.0600 2524.5200 ;
        RECT 1646.4600 2529.4800 1648.0600 2529.9600 ;
        RECT 1646.4600 2507.7200 1648.0600 2508.2000 ;
        RECT 1646.4600 2513.1600 1648.0600 2513.6400 ;
        RECT 1646.4600 2518.6000 1648.0600 2519.0800 ;
        RECT 1691.4600 2496.8400 1693.0600 2497.3200 ;
        RECT 1691.4600 2502.2800 1693.0600 2502.7600 ;
        RECT 1691.4600 2480.5200 1693.0600 2481.0000 ;
        RECT 1691.4600 2485.9600 1693.0600 2486.4400 ;
        RECT 1691.4600 2491.4000 1693.0600 2491.8800 ;
        RECT 1646.4600 2496.8400 1648.0600 2497.3200 ;
        RECT 1646.4600 2502.2800 1648.0600 2502.7600 ;
        RECT 1646.4600 2480.5200 1648.0600 2481.0000 ;
        RECT 1646.4600 2485.9600 1648.0600 2486.4400 ;
        RECT 1646.4600 2491.4000 1648.0600 2491.8800 ;
        RECT 1596.9000 2524.0400 1599.9000 2524.5200 ;
        RECT 1596.9000 2529.4800 1599.9000 2529.9600 ;
        RECT 1596.9000 2513.1600 1599.9000 2513.6400 ;
        RECT 1596.9000 2507.7200 1599.9000 2508.2000 ;
        RECT 1596.9000 2518.6000 1599.9000 2519.0800 ;
        RECT 1596.9000 2496.8400 1599.9000 2497.3200 ;
        RECT 1596.9000 2502.2800 1599.9000 2502.7600 ;
        RECT 1596.9000 2485.9600 1599.9000 2486.4400 ;
        RECT 1596.9000 2480.5200 1599.9000 2481.0000 ;
        RECT 1596.9000 2491.4000 1599.9000 2491.8800 ;
        RECT 1596.9000 2534.9200 1599.9000 2535.4000 ;
        RECT 1646.4600 2534.9200 1648.0600 2535.4000 ;
        RECT 1691.4600 2534.9200 1693.0600 2535.4000 ;
        RECT 1793.0000 2469.6400 1796.0000 2470.1200 ;
        RECT 1793.0000 2475.0800 1796.0000 2475.5600 ;
        RECT 1781.4600 2469.6400 1783.0600 2470.1200 ;
        RECT 1781.4600 2475.0800 1783.0600 2475.5600 ;
        RECT 1793.0000 2453.3200 1796.0000 2453.8000 ;
        RECT 1793.0000 2458.7600 1796.0000 2459.2400 ;
        RECT 1793.0000 2464.2000 1796.0000 2464.6800 ;
        RECT 1781.4600 2453.3200 1783.0600 2453.8000 ;
        RECT 1781.4600 2458.7600 1783.0600 2459.2400 ;
        RECT 1781.4600 2464.2000 1783.0600 2464.6800 ;
        RECT 1793.0000 2442.4400 1796.0000 2442.9200 ;
        RECT 1793.0000 2447.8800 1796.0000 2448.3600 ;
        RECT 1781.4600 2442.4400 1783.0600 2442.9200 ;
        RECT 1781.4600 2447.8800 1783.0600 2448.3600 ;
        RECT 1793.0000 2426.1200 1796.0000 2426.6000 ;
        RECT 1793.0000 2431.5600 1796.0000 2432.0400 ;
        RECT 1793.0000 2437.0000 1796.0000 2437.4800 ;
        RECT 1781.4600 2426.1200 1783.0600 2426.6000 ;
        RECT 1781.4600 2431.5600 1783.0600 2432.0400 ;
        RECT 1781.4600 2437.0000 1783.0600 2437.4800 ;
        RECT 1736.4600 2469.6400 1738.0600 2470.1200 ;
        RECT 1736.4600 2475.0800 1738.0600 2475.5600 ;
        RECT 1736.4600 2453.3200 1738.0600 2453.8000 ;
        RECT 1736.4600 2458.7600 1738.0600 2459.2400 ;
        RECT 1736.4600 2464.2000 1738.0600 2464.6800 ;
        RECT 1736.4600 2442.4400 1738.0600 2442.9200 ;
        RECT 1736.4600 2447.8800 1738.0600 2448.3600 ;
        RECT 1736.4600 2426.1200 1738.0600 2426.6000 ;
        RECT 1736.4600 2431.5600 1738.0600 2432.0400 ;
        RECT 1736.4600 2437.0000 1738.0600 2437.4800 ;
        RECT 1793.0000 2415.2400 1796.0000 2415.7200 ;
        RECT 1793.0000 2420.6800 1796.0000 2421.1600 ;
        RECT 1781.4600 2415.2400 1783.0600 2415.7200 ;
        RECT 1781.4600 2420.6800 1783.0600 2421.1600 ;
        RECT 1793.0000 2398.9200 1796.0000 2399.4000 ;
        RECT 1793.0000 2404.3600 1796.0000 2404.8400 ;
        RECT 1793.0000 2409.8000 1796.0000 2410.2800 ;
        RECT 1781.4600 2398.9200 1783.0600 2399.4000 ;
        RECT 1781.4600 2404.3600 1783.0600 2404.8400 ;
        RECT 1781.4600 2409.8000 1783.0600 2410.2800 ;
        RECT 1793.0000 2388.0400 1796.0000 2388.5200 ;
        RECT 1793.0000 2393.4800 1796.0000 2393.9600 ;
        RECT 1781.4600 2388.0400 1783.0600 2388.5200 ;
        RECT 1781.4600 2393.4800 1783.0600 2393.9600 ;
        RECT 1793.0000 2382.6000 1796.0000 2383.0800 ;
        RECT 1781.4600 2382.6000 1783.0600 2383.0800 ;
        RECT 1736.4600 2415.2400 1738.0600 2415.7200 ;
        RECT 1736.4600 2420.6800 1738.0600 2421.1600 ;
        RECT 1736.4600 2398.9200 1738.0600 2399.4000 ;
        RECT 1736.4600 2404.3600 1738.0600 2404.8400 ;
        RECT 1736.4600 2409.8000 1738.0600 2410.2800 ;
        RECT 1736.4600 2388.0400 1738.0600 2388.5200 ;
        RECT 1736.4600 2393.4800 1738.0600 2393.9600 ;
        RECT 1736.4600 2382.6000 1738.0600 2383.0800 ;
        RECT 1691.4600 2469.6400 1693.0600 2470.1200 ;
        RECT 1691.4600 2475.0800 1693.0600 2475.5600 ;
        RECT 1691.4600 2453.3200 1693.0600 2453.8000 ;
        RECT 1691.4600 2458.7600 1693.0600 2459.2400 ;
        RECT 1691.4600 2464.2000 1693.0600 2464.6800 ;
        RECT 1646.4600 2469.6400 1648.0600 2470.1200 ;
        RECT 1646.4600 2475.0800 1648.0600 2475.5600 ;
        RECT 1646.4600 2453.3200 1648.0600 2453.8000 ;
        RECT 1646.4600 2458.7600 1648.0600 2459.2400 ;
        RECT 1646.4600 2464.2000 1648.0600 2464.6800 ;
        RECT 1691.4600 2442.4400 1693.0600 2442.9200 ;
        RECT 1691.4600 2447.8800 1693.0600 2448.3600 ;
        RECT 1691.4600 2426.1200 1693.0600 2426.6000 ;
        RECT 1691.4600 2431.5600 1693.0600 2432.0400 ;
        RECT 1691.4600 2437.0000 1693.0600 2437.4800 ;
        RECT 1646.4600 2442.4400 1648.0600 2442.9200 ;
        RECT 1646.4600 2447.8800 1648.0600 2448.3600 ;
        RECT 1646.4600 2426.1200 1648.0600 2426.6000 ;
        RECT 1646.4600 2431.5600 1648.0600 2432.0400 ;
        RECT 1646.4600 2437.0000 1648.0600 2437.4800 ;
        RECT 1596.9000 2469.6400 1599.9000 2470.1200 ;
        RECT 1596.9000 2475.0800 1599.9000 2475.5600 ;
        RECT 1596.9000 2458.7600 1599.9000 2459.2400 ;
        RECT 1596.9000 2453.3200 1599.9000 2453.8000 ;
        RECT 1596.9000 2464.2000 1599.9000 2464.6800 ;
        RECT 1596.9000 2442.4400 1599.9000 2442.9200 ;
        RECT 1596.9000 2447.8800 1599.9000 2448.3600 ;
        RECT 1596.9000 2431.5600 1599.9000 2432.0400 ;
        RECT 1596.9000 2426.1200 1599.9000 2426.6000 ;
        RECT 1596.9000 2437.0000 1599.9000 2437.4800 ;
        RECT 1691.4600 2415.2400 1693.0600 2415.7200 ;
        RECT 1691.4600 2420.6800 1693.0600 2421.1600 ;
        RECT 1691.4600 2398.9200 1693.0600 2399.4000 ;
        RECT 1691.4600 2404.3600 1693.0600 2404.8400 ;
        RECT 1691.4600 2409.8000 1693.0600 2410.2800 ;
        RECT 1646.4600 2415.2400 1648.0600 2415.7200 ;
        RECT 1646.4600 2420.6800 1648.0600 2421.1600 ;
        RECT 1646.4600 2398.9200 1648.0600 2399.4000 ;
        RECT 1646.4600 2404.3600 1648.0600 2404.8400 ;
        RECT 1646.4600 2409.8000 1648.0600 2410.2800 ;
        RECT 1691.4600 2393.4800 1693.0600 2393.9600 ;
        RECT 1691.4600 2388.0400 1693.0600 2388.5200 ;
        RECT 1691.4600 2382.6000 1693.0600 2383.0800 ;
        RECT 1646.4600 2393.4800 1648.0600 2393.9600 ;
        RECT 1646.4600 2388.0400 1648.0600 2388.5200 ;
        RECT 1646.4600 2382.6000 1648.0600 2383.0800 ;
        RECT 1596.9000 2415.2400 1599.9000 2415.7200 ;
        RECT 1596.9000 2420.6800 1599.9000 2421.1600 ;
        RECT 1596.9000 2404.3600 1599.9000 2404.8400 ;
        RECT 1596.9000 2398.9200 1599.9000 2399.4000 ;
        RECT 1596.9000 2409.8000 1599.9000 2410.2800 ;
        RECT 1596.9000 2388.0400 1599.9000 2388.5200 ;
        RECT 1596.9000 2393.4800 1599.9000 2393.9600 ;
        RECT 1596.9000 2382.6000 1599.9000 2383.0800 ;
        RECT 1596.9000 2580.7900 1796.0000 2583.7900 ;
        RECT 1596.9000 2375.6900 1796.0000 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 2146.0500 1783.0600 2354.1500 ;
        RECT 1736.4600 2146.0500 1738.0600 2354.1500 ;
        RECT 1691.4600 2146.0500 1693.0600 2354.1500 ;
        RECT 1646.4600 2146.0500 1648.0600 2354.1500 ;
        RECT 1793.0000 2146.0500 1796.0000 2354.1500 ;
        RECT 1596.9000 2146.0500 1599.9000 2354.1500 ;
      LAYER met3 ;
        RECT 1793.0000 2348.8000 1796.0000 2349.2800 ;
        RECT 1781.4600 2348.8000 1783.0600 2349.2800 ;
        RECT 1793.0000 2337.9200 1796.0000 2338.4000 ;
        RECT 1793.0000 2343.3600 1796.0000 2343.8400 ;
        RECT 1781.4600 2337.9200 1783.0600 2338.4000 ;
        RECT 1781.4600 2343.3600 1783.0600 2343.8400 ;
        RECT 1793.0000 2321.6000 1796.0000 2322.0800 ;
        RECT 1793.0000 2327.0400 1796.0000 2327.5200 ;
        RECT 1781.4600 2321.6000 1783.0600 2322.0800 ;
        RECT 1781.4600 2327.0400 1783.0600 2327.5200 ;
        RECT 1793.0000 2310.7200 1796.0000 2311.2000 ;
        RECT 1793.0000 2316.1600 1796.0000 2316.6400 ;
        RECT 1781.4600 2310.7200 1783.0600 2311.2000 ;
        RECT 1781.4600 2316.1600 1783.0600 2316.6400 ;
        RECT 1793.0000 2332.4800 1796.0000 2332.9600 ;
        RECT 1781.4600 2332.4800 1783.0600 2332.9600 ;
        RECT 1736.4600 2337.9200 1738.0600 2338.4000 ;
        RECT 1736.4600 2343.3600 1738.0600 2343.8400 ;
        RECT 1736.4600 2348.8000 1738.0600 2349.2800 ;
        RECT 1736.4600 2321.6000 1738.0600 2322.0800 ;
        RECT 1736.4600 2327.0400 1738.0600 2327.5200 ;
        RECT 1736.4600 2316.1600 1738.0600 2316.6400 ;
        RECT 1736.4600 2310.7200 1738.0600 2311.2000 ;
        RECT 1736.4600 2332.4800 1738.0600 2332.9600 ;
        RECT 1793.0000 2294.4000 1796.0000 2294.8800 ;
        RECT 1793.0000 2299.8400 1796.0000 2300.3200 ;
        RECT 1781.4600 2294.4000 1783.0600 2294.8800 ;
        RECT 1781.4600 2299.8400 1783.0600 2300.3200 ;
        RECT 1793.0000 2278.0800 1796.0000 2278.5600 ;
        RECT 1793.0000 2283.5200 1796.0000 2284.0000 ;
        RECT 1793.0000 2288.9600 1796.0000 2289.4400 ;
        RECT 1781.4600 2278.0800 1783.0600 2278.5600 ;
        RECT 1781.4600 2283.5200 1783.0600 2284.0000 ;
        RECT 1781.4600 2288.9600 1783.0600 2289.4400 ;
        RECT 1793.0000 2267.2000 1796.0000 2267.6800 ;
        RECT 1793.0000 2272.6400 1796.0000 2273.1200 ;
        RECT 1781.4600 2267.2000 1783.0600 2267.6800 ;
        RECT 1781.4600 2272.6400 1783.0600 2273.1200 ;
        RECT 1793.0000 2250.8800 1796.0000 2251.3600 ;
        RECT 1793.0000 2256.3200 1796.0000 2256.8000 ;
        RECT 1793.0000 2261.7600 1796.0000 2262.2400 ;
        RECT 1781.4600 2250.8800 1783.0600 2251.3600 ;
        RECT 1781.4600 2256.3200 1783.0600 2256.8000 ;
        RECT 1781.4600 2261.7600 1783.0600 2262.2400 ;
        RECT 1736.4600 2294.4000 1738.0600 2294.8800 ;
        RECT 1736.4600 2299.8400 1738.0600 2300.3200 ;
        RECT 1736.4600 2278.0800 1738.0600 2278.5600 ;
        RECT 1736.4600 2283.5200 1738.0600 2284.0000 ;
        RECT 1736.4600 2288.9600 1738.0600 2289.4400 ;
        RECT 1736.4600 2267.2000 1738.0600 2267.6800 ;
        RECT 1736.4600 2272.6400 1738.0600 2273.1200 ;
        RECT 1736.4600 2250.8800 1738.0600 2251.3600 ;
        RECT 1736.4600 2256.3200 1738.0600 2256.8000 ;
        RECT 1736.4600 2261.7600 1738.0600 2262.2400 ;
        RECT 1793.0000 2305.2800 1796.0000 2305.7600 ;
        RECT 1736.4600 2305.2800 1738.0600 2305.7600 ;
        RECT 1781.4600 2305.2800 1783.0600 2305.7600 ;
        RECT 1691.4600 2337.9200 1693.0600 2338.4000 ;
        RECT 1691.4600 2343.3600 1693.0600 2343.8400 ;
        RECT 1691.4600 2348.8000 1693.0600 2349.2800 ;
        RECT 1646.4600 2337.9200 1648.0600 2338.4000 ;
        RECT 1646.4600 2343.3600 1648.0600 2343.8400 ;
        RECT 1646.4600 2348.8000 1648.0600 2349.2800 ;
        RECT 1691.4600 2321.6000 1693.0600 2322.0800 ;
        RECT 1691.4600 2327.0400 1693.0600 2327.5200 ;
        RECT 1691.4600 2310.7200 1693.0600 2311.2000 ;
        RECT 1691.4600 2316.1600 1693.0600 2316.6400 ;
        RECT 1646.4600 2321.6000 1648.0600 2322.0800 ;
        RECT 1646.4600 2327.0400 1648.0600 2327.5200 ;
        RECT 1646.4600 2310.7200 1648.0600 2311.2000 ;
        RECT 1646.4600 2316.1600 1648.0600 2316.6400 ;
        RECT 1646.4600 2332.4800 1648.0600 2332.9600 ;
        RECT 1691.4600 2332.4800 1693.0600 2332.9600 ;
        RECT 1596.9000 2348.8000 1599.9000 2349.2800 ;
        RECT 1596.9000 2343.3600 1599.9000 2343.8400 ;
        RECT 1596.9000 2337.9200 1599.9000 2338.4000 ;
        RECT 1596.9000 2327.0400 1599.9000 2327.5200 ;
        RECT 1596.9000 2321.6000 1599.9000 2322.0800 ;
        RECT 1596.9000 2316.1600 1599.9000 2316.6400 ;
        RECT 1596.9000 2310.7200 1599.9000 2311.2000 ;
        RECT 1596.9000 2332.4800 1599.9000 2332.9600 ;
        RECT 1691.4600 2294.4000 1693.0600 2294.8800 ;
        RECT 1691.4600 2299.8400 1693.0600 2300.3200 ;
        RECT 1691.4600 2278.0800 1693.0600 2278.5600 ;
        RECT 1691.4600 2283.5200 1693.0600 2284.0000 ;
        RECT 1691.4600 2288.9600 1693.0600 2289.4400 ;
        RECT 1646.4600 2294.4000 1648.0600 2294.8800 ;
        RECT 1646.4600 2299.8400 1648.0600 2300.3200 ;
        RECT 1646.4600 2278.0800 1648.0600 2278.5600 ;
        RECT 1646.4600 2283.5200 1648.0600 2284.0000 ;
        RECT 1646.4600 2288.9600 1648.0600 2289.4400 ;
        RECT 1691.4600 2267.2000 1693.0600 2267.6800 ;
        RECT 1691.4600 2272.6400 1693.0600 2273.1200 ;
        RECT 1691.4600 2250.8800 1693.0600 2251.3600 ;
        RECT 1691.4600 2256.3200 1693.0600 2256.8000 ;
        RECT 1691.4600 2261.7600 1693.0600 2262.2400 ;
        RECT 1646.4600 2267.2000 1648.0600 2267.6800 ;
        RECT 1646.4600 2272.6400 1648.0600 2273.1200 ;
        RECT 1646.4600 2250.8800 1648.0600 2251.3600 ;
        RECT 1646.4600 2256.3200 1648.0600 2256.8000 ;
        RECT 1646.4600 2261.7600 1648.0600 2262.2400 ;
        RECT 1596.9000 2294.4000 1599.9000 2294.8800 ;
        RECT 1596.9000 2299.8400 1599.9000 2300.3200 ;
        RECT 1596.9000 2283.5200 1599.9000 2284.0000 ;
        RECT 1596.9000 2278.0800 1599.9000 2278.5600 ;
        RECT 1596.9000 2288.9600 1599.9000 2289.4400 ;
        RECT 1596.9000 2267.2000 1599.9000 2267.6800 ;
        RECT 1596.9000 2272.6400 1599.9000 2273.1200 ;
        RECT 1596.9000 2256.3200 1599.9000 2256.8000 ;
        RECT 1596.9000 2250.8800 1599.9000 2251.3600 ;
        RECT 1596.9000 2261.7600 1599.9000 2262.2400 ;
        RECT 1596.9000 2305.2800 1599.9000 2305.7600 ;
        RECT 1646.4600 2305.2800 1648.0600 2305.7600 ;
        RECT 1691.4600 2305.2800 1693.0600 2305.7600 ;
        RECT 1793.0000 2240.0000 1796.0000 2240.4800 ;
        RECT 1793.0000 2245.4400 1796.0000 2245.9200 ;
        RECT 1781.4600 2240.0000 1783.0600 2240.4800 ;
        RECT 1781.4600 2245.4400 1783.0600 2245.9200 ;
        RECT 1793.0000 2223.6800 1796.0000 2224.1600 ;
        RECT 1793.0000 2229.1200 1796.0000 2229.6000 ;
        RECT 1793.0000 2234.5600 1796.0000 2235.0400 ;
        RECT 1781.4600 2223.6800 1783.0600 2224.1600 ;
        RECT 1781.4600 2229.1200 1783.0600 2229.6000 ;
        RECT 1781.4600 2234.5600 1783.0600 2235.0400 ;
        RECT 1793.0000 2212.8000 1796.0000 2213.2800 ;
        RECT 1793.0000 2218.2400 1796.0000 2218.7200 ;
        RECT 1781.4600 2212.8000 1783.0600 2213.2800 ;
        RECT 1781.4600 2218.2400 1783.0600 2218.7200 ;
        RECT 1793.0000 2196.4800 1796.0000 2196.9600 ;
        RECT 1793.0000 2201.9200 1796.0000 2202.4000 ;
        RECT 1793.0000 2207.3600 1796.0000 2207.8400 ;
        RECT 1781.4600 2196.4800 1783.0600 2196.9600 ;
        RECT 1781.4600 2201.9200 1783.0600 2202.4000 ;
        RECT 1781.4600 2207.3600 1783.0600 2207.8400 ;
        RECT 1736.4600 2240.0000 1738.0600 2240.4800 ;
        RECT 1736.4600 2245.4400 1738.0600 2245.9200 ;
        RECT 1736.4600 2223.6800 1738.0600 2224.1600 ;
        RECT 1736.4600 2229.1200 1738.0600 2229.6000 ;
        RECT 1736.4600 2234.5600 1738.0600 2235.0400 ;
        RECT 1736.4600 2212.8000 1738.0600 2213.2800 ;
        RECT 1736.4600 2218.2400 1738.0600 2218.7200 ;
        RECT 1736.4600 2196.4800 1738.0600 2196.9600 ;
        RECT 1736.4600 2201.9200 1738.0600 2202.4000 ;
        RECT 1736.4600 2207.3600 1738.0600 2207.8400 ;
        RECT 1793.0000 2185.6000 1796.0000 2186.0800 ;
        RECT 1793.0000 2191.0400 1796.0000 2191.5200 ;
        RECT 1781.4600 2185.6000 1783.0600 2186.0800 ;
        RECT 1781.4600 2191.0400 1783.0600 2191.5200 ;
        RECT 1793.0000 2169.2800 1796.0000 2169.7600 ;
        RECT 1793.0000 2174.7200 1796.0000 2175.2000 ;
        RECT 1793.0000 2180.1600 1796.0000 2180.6400 ;
        RECT 1781.4600 2169.2800 1783.0600 2169.7600 ;
        RECT 1781.4600 2174.7200 1783.0600 2175.2000 ;
        RECT 1781.4600 2180.1600 1783.0600 2180.6400 ;
        RECT 1793.0000 2158.4000 1796.0000 2158.8800 ;
        RECT 1793.0000 2163.8400 1796.0000 2164.3200 ;
        RECT 1781.4600 2158.4000 1783.0600 2158.8800 ;
        RECT 1781.4600 2163.8400 1783.0600 2164.3200 ;
        RECT 1793.0000 2152.9600 1796.0000 2153.4400 ;
        RECT 1781.4600 2152.9600 1783.0600 2153.4400 ;
        RECT 1736.4600 2185.6000 1738.0600 2186.0800 ;
        RECT 1736.4600 2191.0400 1738.0600 2191.5200 ;
        RECT 1736.4600 2169.2800 1738.0600 2169.7600 ;
        RECT 1736.4600 2174.7200 1738.0600 2175.2000 ;
        RECT 1736.4600 2180.1600 1738.0600 2180.6400 ;
        RECT 1736.4600 2158.4000 1738.0600 2158.8800 ;
        RECT 1736.4600 2163.8400 1738.0600 2164.3200 ;
        RECT 1736.4600 2152.9600 1738.0600 2153.4400 ;
        RECT 1691.4600 2240.0000 1693.0600 2240.4800 ;
        RECT 1691.4600 2245.4400 1693.0600 2245.9200 ;
        RECT 1691.4600 2223.6800 1693.0600 2224.1600 ;
        RECT 1691.4600 2229.1200 1693.0600 2229.6000 ;
        RECT 1691.4600 2234.5600 1693.0600 2235.0400 ;
        RECT 1646.4600 2240.0000 1648.0600 2240.4800 ;
        RECT 1646.4600 2245.4400 1648.0600 2245.9200 ;
        RECT 1646.4600 2223.6800 1648.0600 2224.1600 ;
        RECT 1646.4600 2229.1200 1648.0600 2229.6000 ;
        RECT 1646.4600 2234.5600 1648.0600 2235.0400 ;
        RECT 1691.4600 2212.8000 1693.0600 2213.2800 ;
        RECT 1691.4600 2218.2400 1693.0600 2218.7200 ;
        RECT 1691.4600 2196.4800 1693.0600 2196.9600 ;
        RECT 1691.4600 2201.9200 1693.0600 2202.4000 ;
        RECT 1691.4600 2207.3600 1693.0600 2207.8400 ;
        RECT 1646.4600 2212.8000 1648.0600 2213.2800 ;
        RECT 1646.4600 2218.2400 1648.0600 2218.7200 ;
        RECT 1646.4600 2196.4800 1648.0600 2196.9600 ;
        RECT 1646.4600 2201.9200 1648.0600 2202.4000 ;
        RECT 1646.4600 2207.3600 1648.0600 2207.8400 ;
        RECT 1596.9000 2240.0000 1599.9000 2240.4800 ;
        RECT 1596.9000 2245.4400 1599.9000 2245.9200 ;
        RECT 1596.9000 2229.1200 1599.9000 2229.6000 ;
        RECT 1596.9000 2223.6800 1599.9000 2224.1600 ;
        RECT 1596.9000 2234.5600 1599.9000 2235.0400 ;
        RECT 1596.9000 2212.8000 1599.9000 2213.2800 ;
        RECT 1596.9000 2218.2400 1599.9000 2218.7200 ;
        RECT 1596.9000 2201.9200 1599.9000 2202.4000 ;
        RECT 1596.9000 2196.4800 1599.9000 2196.9600 ;
        RECT 1596.9000 2207.3600 1599.9000 2207.8400 ;
        RECT 1691.4600 2185.6000 1693.0600 2186.0800 ;
        RECT 1691.4600 2191.0400 1693.0600 2191.5200 ;
        RECT 1691.4600 2169.2800 1693.0600 2169.7600 ;
        RECT 1691.4600 2174.7200 1693.0600 2175.2000 ;
        RECT 1691.4600 2180.1600 1693.0600 2180.6400 ;
        RECT 1646.4600 2185.6000 1648.0600 2186.0800 ;
        RECT 1646.4600 2191.0400 1648.0600 2191.5200 ;
        RECT 1646.4600 2169.2800 1648.0600 2169.7600 ;
        RECT 1646.4600 2174.7200 1648.0600 2175.2000 ;
        RECT 1646.4600 2180.1600 1648.0600 2180.6400 ;
        RECT 1691.4600 2163.8400 1693.0600 2164.3200 ;
        RECT 1691.4600 2158.4000 1693.0600 2158.8800 ;
        RECT 1691.4600 2152.9600 1693.0600 2153.4400 ;
        RECT 1646.4600 2163.8400 1648.0600 2164.3200 ;
        RECT 1646.4600 2158.4000 1648.0600 2158.8800 ;
        RECT 1646.4600 2152.9600 1648.0600 2153.4400 ;
        RECT 1596.9000 2185.6000 1599.9000 2186.0800 ;
        RECT 1596.9000 2191.0400 1599.9000 2191.5200 ;
        RECT 1596.9000 2174.7200 1599.9000 2175.2000 ;
        RECT 1596.9000 2169.2800 1599.9000 2169.7600 ;
        RECT 1596.9000 2180.1600 1599.9000 2180.6400 ;
        RECT 1596.9000 2158.4000 1599.9000 2158.8800 ;
        RECT 1596.9000 2163.8400 1599.9000 2164.3200 ;
        RECT 1596.9000 2152.9600 1599.9000 2153.4400 ;
        RECT 1596.9000 2351.1500 1796.0000 2354.1500 ;
        RECT 1596.9000 2146.0500 1796.0000 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 1916.4100 1783.0600 2124.5100 ;
        RECT 1736.4600 1916.4100 1738.0600 2124.5100 ;
        RECT 1691.4600 1916.4100 1693.0600 2124.5100 ;
        RECT 1646.4600 1916.4100 1648.0600 2124.5100 ;
        RECT 1793.0000 1916.4100 1796.0000 2124.5100 ;
        RECT 1596.9000 1916.4100 1599.9000 2124.5100 ;
      LAYER met3 ;
        RECT 1793.0000 2119.1600 1796.0000 2119.6400 ;
        RECT 1781.4600 2119.1600 1783.0600 2119.6400 ;
        RECT 1793.0000 2108.2800 1796.0000 2108.7600 ;
        RECT 1793.0000 2113.7200 1796.0000 2114.2000 ;
        RECT 1781.4600 2108.2800 1783.0600 2108.7600 ;
        RECT 1781.4600 2113.7200 1783.0600 2114.2000 ;
        RECT 1793.0000 2091.9600 1796.0000 2092.4400 ;
        RECT 1793.0000 2097.4000 1796.0000 2097.8800 ;
        RECT 1781.4600 2091.9600 1783.0600 2092.4400 ;
        RECT 1781.4600 2097.4000 1783.0600 2097.8800 ;
        RECT 1793.0000 2081.0800 1796.0000 2081.5600 ;
        RECT 1793.0000 2086.5200 1796.0000 2087.0000 ;
        RECT 1781.4600 2081.0800 1783.0600 2081.5600 ;
        RECT 1781.4600 2086.5200 1783.0600 2087.0000 ;
        RECT 1793.0000 2102.8400 1796.0000 2103.3200 ;
        RECT 1781.4600 2102.8400 1783.0600 2103.3200 ;
        RECT 1736.4600 2108.2800 1738.0600 2108.7600 ;
        RECT 1736.4600 2113.7200 1738.0600 2114.2000 ;
        RECT 1736.4600 2119.1600 1738.0600 2119.6400 ;
        RECT 1736.4600 2091.9600 1738.0600 2092.4400 ;
        RECT 1736.4600 2097.4000 1738.0600 2097.8800 ;
        RECT 1736.4600 2086.5200 1738.0600 2087.0000 ;
        RECT 1736.4600 2081.0800 1738.0600 2081.5600 ;
        RECT 1736.4600 2102.8400 1738.0600 2103.3200 ;
        RECT 1793.0000 2064.7600 1796.0000 2065.2400 ;
        RECT 1793.0000 2070.2000 1796.0000 2070.6800 ;
        RECT 1781.4600 2064.7600 1783.0600 2065.2400 ;
        RECT 1781.4600 2070.2000 1783.0600 2070.6800 ;
        RECT 1793.0000 2048.4400 1796.0000 2048.9200 ;
        RECT 1793.0000 2053.8800 1796.0000 2054.3600 ;
        RECT 1793.0000 2059.3200 1796.0000 2059.8000 ;
        RECT 1781.4600 2048.4400 1783.0600 2048.9200 ;
        RECT 1781.4600 2053.8800 1783.0600 2054.3600 ;
        RECT 1781.4600 2059.3200 1783.0600 2059.8000 ;
        RECT 1793.0000 2037.5600 1796.0000 2038.0400 ;
        RECT 1793.0000 2043.0000 1796.0000 2043.4800 ;
        RECT 1781.4600 2037.5600 1783.0600 2038.0400 ;
        RECT 1781.4600 2043.0000 1783.0600 2043.4800 ;
        RECT 1793.0000 2021.2400 1796.0000 2021.7200 ;
        RECT 1793.0000 2026.6800 1796.0000 2027.1600 ;
        RECT 1793.0000 2032.1200 1796.0000 2032.6000 ;
        RECT 1781.4600 2021.2400 1783.0600 2021.7200 ;
        RECT 1781.4600 2026.6800 1783.0600 2027.1600 ;
        RECT 1781.4600 2032.1200 1783.0600 2032.6000 ;
        RECT 1736.4600 2064.7600 1738.0600 2065.2400 ;
        RECT 1736.4600 2070.2000 1738.0600 2070.6800 ;
        RECT 1736.4600 2048.4400 1738.0600 2048.9200 ;
        RECT 1736.4600 2053.8800 1738.0600 2054.3600 ;
        RECT 1736.4600 2059.3200 1738.0600 2059.8000 ;
        RECT 1736.4600 2037.5600 1738.0600 2038.0400 ;
        RECT 1736.4600 2043.0000 1738.0600 2043.4800 ;
        RECT 1736.4600 2021.2400 1738.0600 2021.7200 ;
        RECT 1736.4600 2026.6800 1738.0600 2027.1600 ;
        RECT 1736.4600 2032.1200 1738.0600 2032.6000 ;
        RECT 1793.0000 2075.6400 1796.0000 2076.1200 ;
        RECT 1736.4600 2075.6400 1738.0600 2076.1200 ;
        RECT 1781.4600 2075.6400 1783.0600 2076.1200 ;
        RECT 1691.4600 2108.2800 1693.0600 2108.7600 ;
        RECT 1691.4600 2113.7200 1693.0600 2114.2000 ;
        RECT 1691.4600 2119.1600 1693.0600 2119.6400 ;
        RECT 1646.4600 2108.2800 1648.0600 2108.7600 ;
        RECT 1646.4600 2113.7200 1648.0600 2114.2000 ;
        RECT 1646.4600 2119.1600 1648.0600 2119.6400 ;
        RECT 1691.4600 2091.9600 1693.0600 2092.4400 ;
        RECT 1691.4600 2097.4000 1693.0600 2097.8800 ;
        RECT 1691.4600 2081.0800 1693.0600 2081.5600 ;
        RECT 1691.4600 2086.5200 1693.0600 2087.0000 ;
        RECT 1646.4600 2091.9600 1648.0600 2092.4400 ;
        RECT 1646.4600 2097.4000 1648.0600 2097.8800 ;
        RECT 1646.4600 2081.0800 1648.0600 2081.5600 ;
        RECT 1646.4600 2086.5200 1648.0600 2087.0000 ;
        RECT 1646.4600 2102.8400 1648.0600 2103.3200 ;
        RECT 1691.4600 2102.8400 1693.0600 2103.3200 ;
        RECT 1596.9000 2119.1600 1599.9000 2119.6400 ;
        RECT 1596.9000 2113.7200 1599.9000 2114.2000 ;
        RECT 1596.9000 2108.2800 1599.9000 2108.7600 ;
        RECT 1596.9000 2097.4000 1599.9000 2097.8800 ;
        RECT 1596.9000 2091.9600 1599.9000 2092.4400 ;
        RECT 1596.9000 2086.5200 1599.9000 2087.0000 ;
        RECT 1596.9000 2081.0800 1599.9000 2081.5600 ;
        RECT 1596.9000 2102.8400 1599.9000 2103.3200 ;
        RECT 1691.4600 2064.7600 1693.0600 2065.2400 ;
        RECT 1691.4600 2070.2000 1693.0600 2070.6800 ;
        RECT 1691.4600 2048.4400 1693.0600 2048.9200 ;
        RECT 1691.4600 2053.8800 1693.0600 2054.3600 ;
        RECT 1691.4600 2059.3200 1693.0600 2059.8000 ;
        RECT 1646.4600 2064.7600 1648.0600 2065.2400 ;
        RECT 1646.4600 2070.2000 1648.0600 2070.6800 ;
        RECT 1646.4600 2048.4400 1648.0600 2048.9200 ;
        RECT 1646.4600 2053.8800 1648.0600 2054.3600 ;
        RECT 1646.4600 2059.3200 1648.0600 2059.8000 ;
        RECT 1691.4600 2037.5600 1693.0600 2038.0400 ;
        RECT 1691.4600 2043.0000 1693.0600 2043.4800 ;
        RECT 1691.4600 2021.2400 1693.0600 2021.7200 ;
        RECT 1691.4600 2026.6800 1693.0600 2027.1600 ;
        RECT 1691.4600 2032.1200 1693.0600 2032.6000 ;
        RECT 1646.4600 2037.5600 1648.0600 2038.0400 ;
        RECT 1646.4600 2043.0000 1648.0600 2043.4800 ;
        RECT 1646.4600 2021.2400 1648.0600 2021.7200 ;
        RECT 1646.4600 2026.6800 1648.0600 2027.1600 ;
        RECT 1646.4600 2032.1200 1648.0600 2032.6000 ;
        RECT 1596.9000 2064.7600 1599.9000 2065.2400 ;
        RECT 1596.9000 2070.2000 1599.9000 2070.6800 ;
        RECT 1596.9000 2053.8800 1599.9000 2054.3600 ;
        RECT 1596.9000 2048.4400 1599.9000 2048.9200 ;
        RECT 1596.9000 2059.3200 1599.9000 2059.8000 ;
        RECT 1596.9000 2037.5600 1599.9000 2038.0400 ;
        RECT 1596.9000 2043.0000 1599.9000 2043.4800 ;
        RECT 1596.9000 2026.6800 1599.9000 2027.1600 ;
        RECT 1596.9000 2021.2400 1599.9000 2021.7200 ;
        RECT 1596.9000 2032.1200 1599.9000 2032.6000 ;
        RECT 1596.9000 2075.6400 1599.9000 2076.1200 ;
        RECT 1646.4600 2075.6400 1648.0600 2076.1200 ;
        RECT 1691.4600 2075.6400 1693.0600 2076.1200 ;
        RECT 1793.0000 2010.3600 1796.0000 2010.8400 ;
        RECT 1793.0000 2015.8000 1796.0000 2016.2800 ;
        RECT 1781.4600 2010.3600 1783.0600 2010.8400 ;
        RECT 1781.4600 2015.8000 1783.0600 2016.2800 ;
        RECT 1793.0000 1994.0400 1796.0000 1994.5200 ;
        RECT 1793.0000 1999.4800 1796.0000 1999.9600 ;
        RECT 1793.0000 2004.9200 1796.0000 2005.4000 ;
        RECT 1781.4600 1994.0400 1783.0600 1994.5200 ;
        RECT 1781.4600 1999.4800 1783.0600 1999.9600 ;
        RECT 1781.4600 2004.9200 1783.0600 2005.4000 ;
        RECT 1793.0000 1983.1600 1796.0000 1983.6400 ;
        RECT 1793.0000 1988.6000 1796.0000 1989.0800 ;
        RECT 1781.4600 1983.1600 1783.0600 1983.6400 ;
        RECT 1781.4600 1988.6000 1783.0600 1989.0800 ;
        RECT 1793.0000 1966.8400 1796.0000 1967.3200 ;
        RECT 1793.0000 1972.2800 1796.0000 1972.7600 ;
        RECT 1793.0000 1977.7200 1796.0000 1978.2000 ;
        RECT 1781.4600 1966.8400 1783.0600 1967.3200 ;
        RECT 1781.4600 1972.2800 1783.0600 1972.7600 ;
        RECT 1781.4600 1977.7200 1783.0600 1978.2000 ;
        RECT 1736.4600 2010.3600 1738.0600 2010.8400 ;
        RECT 1736.4600 2015.8000 1738.0600 2016.2800 ;
        RECT 1736.4600 1994.0400 1738.0600 1994.5200 ;
        RECT 1736.4600 1999.4800 1738.0600 1999.9600 ;
        RECT 1736.4600 2004.9200 1738.0600 2005.4000 ;
        RECT 1736.4600 1983.1600 1738.0600 1983.6400 ;
        RECT 1736.4600 1988.6000 1738.0600 1989.0800 ;
        RECT 1736.4600 1966.8400 1738.0600 1967.3200 ;
        RECT 1736.4600 1972.2800 1738.0600 1972.7600 ;
        RECT 1736.4600 1977.7200 1738.0600 1978.2000 ;
        RECT 1793.0000 1955.9600 1796.0000 1956.4400 ;
        RECT 1793.0000 1961.4000 1796.0000 1961.8800 ;
        RECT 1781.4600 1955.9600 1783.0600 1956.4400 ;
        RECT 1781.4600 1961.4000 1783.0600 1961.8800 ;
        RECT 1793.0000 1939.6400 1796.0000 1940.1200 ;
        RECT 1793.0000 1945.0800 1796.0000 1945.5600 ;
        RECT 1793.0000 1950.5200 1796.0000 1951.0000 ;
        RECT 1781.4600 1939.6400 1783.0600 1940.1200 ;
        RECT 1781.4600 1945.0800 1783.0600 1945.5600 ;
        RECT 1781.4600 1950.5200 1783.0600 1951.0000 ;
        RECT 1793.0000 1928.7600 1796.0000 1929.2400 ;
        RECT 1793.0000 1934.2000 1796.0000 1934.6800 ;
        RECT 1781.4600 1928.7600 1783.0600 1929.2400 ;
        RECT 1781.4600 1934.2000 1783.0600 1934.6800 ;
        RECT 1793.0000 1923.3200 1796.0000 1923.8000 ;
        RECT 1781.4600 1923.3200 1783.0600 1923.8000 ;
        RECT 1736.4600 1955.9600 1738.0600 1956.4400 ;
        RECT 1736.4600 1961.4000 1738.0600 1961.8800 ;
        RECT 1736.4600 1939.6400 1738.0600 1940.1200 ;
        RECT 1736.4600 1945.0800 1738.0600 1945.5600 ;
        RECT 1736.4600 1950.5200 1738.0600 1951.0000 ;
        RECT 1736.4600 1928.7600 1738.0600 1929.2400 ;
        RECT 1736.4600 1934.2000 1738.0600 1934.6800 ;
        RECT 1736.4600 1923.3200 1738.0600 1923.8000 ;
        RECT 1691.4600 2010.3600 1693.0600 2010.8400 ;
        RECT 1691.4600 2015.8000 1693.0600 2016.2800 ;
        RECT 1691.4600 1994.0400 1693.0600 1994.5200 ;
        RECT 1691.4600 1999.4800 1693.0600 1999.9600 ;
        RECT 1691.4600 2004.9200 1693.0600 2005.4000 ;
        RECT 1646.4600 2010.3600 1648.0600 2010.8400 ;
        RECT 1646.4600 2015.8000 1648.0600 2016.2800 ;
        RECT 1646.4600 1994.0400 1648.0600 1994.5200 ;
        RECT 1646.4600 1999.4800 1648.0600 1999.9600 ;
        RECT 1646.4600 2004.9200 1648.0600 2005.4000 ;
        RECT 1691.4600 1983.1600 1693.0600 1983.6400 ;
        RECT 1691.4600 1988.6000 1693.0600 1989.0800 ;
        RECT 1691.4600 1966.8400 1693.0600 1967.3200 ;
        RECT 1691.4600 1972.2800 1693.0600 1972.7600 ;
        RECT 1691.4600 1977.7200 1693.0600 1978.2000 ;
        RECT 1646.4600 1983.1600 1648.0600 1983.6400 ;
        RECT 1646.4600 1988.6000 1648.0600 1989.0800 ;
        RECT 1646.4600 1966.8400 1648.0600 1967.3200 ;
        RECT 1646.4600 1972.2800 1648.0600 1972.7600 ;
        RECT 1646.4600 1977.7200 1648.0600 1978.2000 ;
        RECT 1596.9000 2010.3600 1599.9000 2010.8400 ;
        RECT 1596.9000 2015.8000 1599.9000 2016.2800 ;
        RECT 1596.9000 1999.4800 1599.9000 1999.9600 ;
        RECT 1596.9000 1994.0400 1599.9000 1994.5200 ;
        RECT 1596.9000 2004.9200 1599.9000 2005.4000 ;
        RECT 1596.9000 1983.1600 1599.9000 1983.6400 ;
        RECT 1596.9000 1988.6000 1599.9000 1989.0800 ;
        RECT 1596.9000 1972.2800 1599.9000 1972.7600 ;
        RECT 1596.9000 1966.8400 1599.9000 1967.3200 ;
        RECT 1596.9000 1977.7200 1599.9000 1978.2000 ;
        RECT 1691.4600 1955.9600 1693.0600 1956.4400 ;
        RECT 1691.4600 1961.4000 1693.0600 1961.8800 ;
        RECT 1691.4600 1939.6400 1693.0600 1940.1200 ;
        RECT 1691.4600 1945.0800 1693.0600 1945.5600 ;
        RECT 1691.4600 1950.5200 1693.0600 1951.0000 ;
        RECT 1646.4600 1955.9600 1648.0600 1956.4400 ;
        RECT 1646.4600 1961.4000 1648.0600 1961.8800 ;
        RECT 1646.4600 1939.6400 1648.0600 1940.1200 ;
        RECT 1646.4600 1945.0800 1648.0600 1945.5600 ;
        RECT 1646.4600 1950.5200 1648.0600 1951.0000 ;
        RECT 1691.4600 1934.2000 1693.0600 1934.6800 ;
        RECT 1691.4600 1928.7600 1693.0600 1929.2400 ;
        RECT 1691.4600 1923.3200 1693.0600 1923.8000 ;
        RECT 1646.4600 1934.2000 1648.0600 1934.6800 ;
        RECT 1646.4600 1928.7600 1648.0600 1929.2400 ;
        RECT 1646.4600 1923.3200 1648.0600 1923.8000 ;
        RECT 1596.9000 1955.9600 1599.9000 1956.4400 ;
        RECT 1596.9000 1961.4000 1599.9000 1961.8800 ;
        RECT 1596.9000 1945.0800 1599.9000 1945.5600 ;
        RECT 1596.9000 1939.6400 1599.9000 1940.1200 ;
        RECT 1596.9000 1950.5200 1599.9000 1951.0000 ;
        RECT 1596.9000 1928.7600 1599.9000 1929.2400 ;
        RECT 1596.9000 1934.2000 1599.9000 1934.6800 ;
        RECT 1596.9000 1923.3200 1599.9000 1923.8000 ;
        RECT 1596.9000 2121.5100 1796.0000 2124.5100 ;
        RECT 1596.9000 1916.4100 1796.0000 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 1686.7700 1783.0600 1894.8700 ;
        RECT 1736.4600 1686.7700 1738.0600 1894.8700 ;
        RECT 1691.4600 1686.7700 1693.0600 1894.8700 ;
        RECT 1646.4600 1686.7700 1648.0600 1894.8700 ;
        RECT 1793.0000 1686.7700 1796.0000 1894.8700 ;
        RECT 1596.9000 1686.7700 1599.9000 1894.8700 ;
      LAYER met3 ;
        RECT 1793.0000 1889.5200 1796.0000 1890.0000 ;
        RECT 1781.4600 1889.5200 1783.0600 1890.0000 ;
        RECT 1793.0000 1878.6400 1796.0000 1879.1200 ;
        RECT 1793.0000 1884.0800 1796.0000 1884.5600 ;
        RECT 1781.4600 1878.6400 1783.0600 1879.1200 ;
        RECT 1781.4600 1884.0800 1783.0600 1884.5600 ;
        RECT 1793.0000 1862.3200 1796.0000 1862.8000 ;
        RECT 1793.0000 1867.7600 1796.0000 1868.2400 ;
        RECT 1781.4600 1862.3200 1783.0600 1862.8000 ;
        RECT 1781.4600 1867.7600 1783.0600 1868.2400 ;
        RECT 1793.0000 1851.4400 1796.0000 1851.9200 ;
        RECT 1793.0000 1856.8800 1796.0000 1857.3600 ;
        RECT 1781.4600 1851.4400 1783.0600 1851.9200 ;
        RECT 1781.4600 1856.8800 1783.0600 1857.3600 ;
        RECT 1793.0000 1873.2000 1796.0000 1873.6800 ;
        RECT 1781.4600 1873.2000 1783.0600 1873.6800 ;
        RECT 1736.4600 1878.6400 1738.0600 1879.1200 ;
        RECT 1736.4600 1884.0800 1738.0600 1884.5600 ;
        RECT 1736.4600 1889.5200 1738.0600 1890.0000 ;
        RECT 1736.4600 1862.3200 1738.0600 1862.8000 ;
        RECT 1736.4600 1867.7600 1738.0600 1868.2400 ;
        RECT 1736.4600 1856.8800 1738.0600 1857.3600 ;
        RECT 1736.4600 1851.4400 1738.0600 1851.9200 ;
        RECT 1736.4600 1873.2000 1738.0600 1873.6800 ;
        RECT 1793.0000 1835.1200 1796.0000 1835.6000 ;
        RECT 1793.0000 1840.5600 1796.0000 1841.0400 ;
        RECT 1781.4600 1835.1200 1783.0600 1835.6000 ;
        RECT 1781.4600 1840.5600 1783.0600 1841.0400 ;
        RECT 1793.0000 1818.8000 1796.0000 1819.2800 ;
        RECT 1793.0000 1824.2400 1796.0000 1824.7200 ;
        RECT 1793.0000 1829.6800 1796.0000 1830.1600 ;
        RECT 1781.4600 1818.8000 1783.0600 1819.2800 ;
        RECT 1781.4600 1824.2400 1783.0600 1824.7200 ;
        RECT 1781.4600 1829.6800 1783.0600 1830.1600 ;
        RECT 1793.0000 1807.9200 1796.0000 1808.4000 ;
        RECT 1793.0000 1813.3600 1796.0000 1813.8400 ;
        RECT 1781.4600 1807.9200 1783.0600 1808.4000 ;
        RECT 1781.4600 1813.3600 1783.0600 1813.8400 ;
        RECT 1793.0000 1791.6000 1796.0000 1792.0800 ;
        RECT 1793.0000 1797.0400 1796.0000 1797.5200 ;
        RECT 1793.0000 1802.4800 1796.0000 1802.9600 ;
        RECT 1781.4600 1791.6000 1783.0600 1792.0800 ;
        RECT 1781.4600 1797.0400 1783.0600 1797.5200 ;
        RECT 1781.4600 1802.4800 1783.0600 1802.9600 ;
        RECT 1736.4600 1835.1200 1738.0600 1835.6000 ;
        RECT 1736.4600 1840.5600 1738.0600 1841.0400 ;
        RECT 1736.4600 1818.8000 1738.0600 1819.2800 ;
        RECT 1736.4600 1824.2400 1738.0600 1824.7200 ;
        RECT 1736.4600 1829.6800 1738.0600 1830.1600 ;
        RECT 1736.4600 1807.9200 1738.0600 1808.4000 ;
        RECT 1736.4600 1813.3600 1738.0600 1813.8400 ;
        RECT 1736.4600 1791.6000 1738.0600 1792.0800 ;
        RECT 1736.4600 1797.0400 1738.0600 1797.5200 ;
        RECT 1736.4600 1802.4800 1738.0600 1802.9600 ;
        RECT 1793.0000 1846.0000 1796.0000 1846.4800 ;
        RECT 1736.4600 1846.0000 1738.0600 1846.4800 ;
        RECT 1781.4600 1846.0000 1783.0600 1846.4800 ;
        RECT 1691.4600 1878.6400 1693.0600 1879.1200 ;
        RECT 1691.4600 1884.0800 1693.0600 1884.5600 ;
        RECT 1691.4600 1889.5200 1693.0600 1890.0000 ;
        RECT 1646.4600 1878.6400 1648.0600 1879.1200 ;
        RECT 1646.4600 1884.0800 1648.0600 1884.5600 ;
        RECT 1646.4600 1889.5200 1648.0600 1890.0000 ;
        RECT 1691.4600 1862.3200 1693.0600 1862.8000 ;
        RECT 1691.4600 1867.7600 1693.0600 1868.2400 ;
        RECT 1691.4600 1851.4400 1693.0600 1851.9200 ;
        RECT 1691.4600 1856.8800 1693.0600 1857.3600 ;
        RECT 1646.4600 1862.3200 1648.0600 1862.8000 ;
        RECT 1646.4600 1867.7600 1648.0600 1868.2400 ;
        RECT 1646.4600 1851.4400 1648.0600 1851.9200 ;
        RECT 1646.4600 1856.8800 1648.0600 1857.3600 ;
        RECT 1646.4600 1873.2000 1648.0600 1873.6800 ;
        RECT 1691.4600 1873.2000 1693.0600 1873.6800 ;
        RECT 1596.9000 1889.5200 1599.9000 1890.0000 ;
        RECT 1596.9000 1884.0800 1599.9000 1884.5600 ;
        RECT 1596.9000 1878.6400 1599.9000 1879.1200 ;
        RECT 1596.9000 1867.7600 1599.9000 1868.2400 ;
        RECT 1596.9000 1862.3200 1599.9000 1862.8000 ;
        RECT 1596.9000 1856.8800 1599.9000 1857.3600 ;
        RECT 1596.9000 1851.4400 1599.9000 1851.9200 ;
        RECT 1596.9000 1873.2000 1599.9000 1873.6800 ;
        RECT 1691.4600 1835.1200 1693.0600 1835.6000 ;
        RECT 1691.4600 1840.5600 1693.0600 1841.0400 ;
        RECT 1691.4600 1818.8000 1693.0600 1819.2800 ;
        RECT 1691.4600 1824.2400 1693.0600 1824.7200 ;
        RECT 1691.4600 1829.6800 1693.0600 1830.1600 ;
        RECT 1646.4600 1835.1200 1648.0600 1835.6000 ;
        RECT 1646.4600 1840.5600 1648.0600 1841.0400 ;
        RECT 1646.4600 1818.8000 1648.0600 1819.2800 ;
        RECT 1646.4600 1824.2400 1648.0600 1824.7200 ;
        RECT 1646.4600 1829.6800 1648.0600 1830.1600 ;
        RECT 1691.4600 1807.9200 1693.0600 1808.4000 ;
        RECT 1691.4600 1813.3600 1693.0600 1813.8400 ;
        RECT 1691.4600 1791.6000 1693.0600 1792.0800 ;
        RECT 1691.4600 1797.0400 1693.0600 1797.5200 ;
        RECT 1691.4600 1802.4800 1693.0600 1802.9600 ;
        RECT 1646.4600 1807.9200 1648.0600 1808.4000 ;
        RECT 1646.4600 1813.3600 1648.0600 1813.8400 ;
        RECT 1646.4600 1791.6000 1648.0600 1792.0800 ;
        RECT 1646.4600 1797.0400 1648.0600 1797.5200 ;
        RECT 1646.4600 1802.4800 1648.0600 1802.9600 ;
        RECT 1596.9000 1835.1200 1599.9000 1835.6000 ;
        RECT 1596.9000 1840.5600 1599.9000 1841.0400 ;
        RECT 1596.9000 1824.2400 1599.9000 1824.7200 ;
        RECT 1596.9000 1818.8000 1599.9000 1819.2800 ;
        RECT 1596.9000 1829.6800 1599.9000 1830.1600 ;
        RECT 1596.9000 1807.9200 1599.9000 1808.4000 ;
        RECT 1596.9000 1813.3600 1599.9000 1813.8400 ;
        RECT 1596.9000 1797.0400 1599.9000 1797.5200 ;
        RECT 1596.9000 1791.6000 1599.9000 1792.0800 ;
        RECT 1596.9000 1802.4800 1599.9000 1802.9600 ;
        RECT 1596.9000 1846.0000 1599.9000 1846.4800 ;
        RECT 1646.4600 1846.0000 1648.0600 1846.4800 ;
        RECT 1691.4600 1846.0000 1693.0600 1846.4800 ;
        RECT 1793.0000 1780.7200 1796.0000 1781.2000 ;
        RECT 1793.0000 1786.1600 1796.0000 1786.6400 ;
        RECT 1781.4600 1780.7200 1783.0600 1781.2000 ;
        RECT 1781.4600 1786.1600 1783.0600 1786.6400 ;
        RECT 1793.0000 1764.4000 1796.0000 1764.8800 ;
        RECT 1793.0000 1769.8400 1796.0000 1770.3200 ;
        RECT 1793.0000 1775.2800 1796.0000 1775.7600 ;
        RECT 1781.4600 1764.4000 1783.0600 1764.8800 ;
        RECT 1781.4600 1769.8400 1783.0600 1770.3200 ;
        RECT 1781.4600 1775.2800 1783.0600 1775.7600 ;
        RECT 1793.0000 1753.5200 1796.0000 1754.0000 ;
        RECT 1793.0000 1758.9600 1796.0000 1759.4400 ;
        RECT 1781.4600 1753.5200 1783.0600 1754.0000 ;
        RECT 1781.4600 1758.9600 1783.0600 1759.4400 ;
        RECT 1793.0000 1737.2000 1796.0000 1737.6800 ;
        RECT 1793.0000 1742.6400 1796.0000 1743.1200 ;
        RECT 1793.0000 1748.0800 1796.0000 1748.5600 ;
        RECT 1781.4600 1737.2000 1783.0600 1737.6800 ;
        RECT 1781.4600 1742.6400 1783.0600 1743.1200 ;
        RECT 1781.4600 1748.0800 1783.0600 1748.5600 ;
        RECT 1736.4600 1780.7200 1738.0600 1781.2000 ;
        RECT 1736.4600 1786.1600 1738.0600 1786.6400 ;
        RECT 1736.4600 1764.4000 1738.0600 1764.8800 ;
        RECT 1736.4600 1769.8400 1738.0600 1770.3200 ;
        RECT 1736.4600 1775.2800 1738.0600 1775.7600 ;
        RECT 1736.4600 1753.5200 1738.0600 1754.0000 ;
        RECT 1736.4600 1758.9600 1738.0600 1759.4400 ;
        RECT 1736.4600 1737.2000 1738.0600 1737.6800 ;
        RECT 1736.4600 1742.6400 1738.0600 1743.1200 ;
        RECT 1736.4600 1748.0800 1738.0600 1748.5600 ;
        RECT 1793.0000 1726.3200 1796.0000 1726.8000 ;
        RECT 1793.0000 1731.7600 1796.0000 1732.2400 ;
        RECT 1781.4600 1726.3200 1783.0600 1726.8000 ;
        RECT 1781.4600 1731.7600 1783.0600 1732.2400 ;
        RECT 1793.0000 1710.0000 1796.0000 1710.4800 ;
        RECT 1793.0000 1715.4400 1796.0000 1715.9200 ;
        RECT 1793.0000 1720.8800 1796.0000 1721.3600 ;
        RECT 1781.4600 1710.0000 1783.0600 1710.4800 ;
        RECT 1781.4600 1715.4400 1783.0600 1715.9200 ;
        RECT 1781.4600 1720.8800 1783.0600 1721.3600 ;
        RECT 1793.0000 1699.1200 1796.0000 1699.6000 ;
        RECT 1793.0000 1704.5600 1796.0000 1705.0400 ;
        RECT 1781.4600 1699.1200 1783.0600 1699.6000 ;
        RECT 1781.4600 1704.5600 1783.0600 1705.0400 ;
        RECT 1793.0000 1693.6800 1796.0000 1694.1600 ;
        RECT 1781.4600 1693.6800 1783.0600 1694.1600 ;
        RECT 1736.4600 1726.3200 1738.0600 1726.8000 ;
        RECT 1736.4600 1731.7600 1738.0600 1732.2400 ;
        RECT 1736.4600 1710.0000 1738.0600 1710.4800 ;
        RECT 1736.4600 1715.4400 1738.0600 1715.9200 ;
        RECT 1736.4600 1720.8800 1738.0600 1721.3600 ;
        RECT 1736.4600 1699.1200 1738.0600 1699.6000 ;
        RECT 1736.4600 1704.5600 1738.0600 1705.0400 ;
        RECT 1736.4600 1693.6800 1738.0600 1694.1600 ;
        RECT 1691.4600 1780.7200 1693.0600 1781.2000 ;
        RECT 1691.4600 1786.1600 1693.0600 1786.6400 ;
        RECT 1691.4600 1764.4000 1693.0600 1764.8800 ;
        RECT 1691.4600 1769.8400 1693.0600 1770.3200 ;
        RECT 1691.4600 1775.2800 1693.0600 1775.7600 ;
        RECT 1646.4600 1780.7200 1648.0600 1781.2000 ;
        RECT 1646.4600 1786.1600 1648.0600 1786.6400 ;
        RECT 1646.4600 1764.4000 1648.0600 1764.8800 ;
        RECT 1646.4600 1769.8400 1648.0600 1770.3200 ;
        RECT 1646.4600 1775.2800 1648.0600 1775.7600 ;
        RECT 1691.4600 1753.5200 1693.0600 1754.0000 ;
        RECT 1691.4600 1758.9600 1693.0600 1759.4400 ;
        RECT 1691.4600 1737.2000 1693.0600 1737.6800 ;
        RECT 1691.4600 1742.6400 1693.0600 1743.1200 ;
        RECT 1691.4600 1748.0800 1693.0600 1748.5600 ;
        RECT 1646.4600 1753.5200 1648.0600 1754.0000 ;
        RECT 1646.4600 1758.9600 1648.0600 1759.4400 ;
        RECT 1646.4600 1737.2000 1648.0600 1737.6800 ;
        RECT 1646.4600 1742.6400 1648.0600 1743.1200 ;
        RECT 1646.4600 1748.0800 1648.0600 1748.5600 ;
        RECT 1596.9000 1780.7200 1599.9000 1781.2000 ;
        RECT 1596.9000 1786.1600 1599.9000 1786.6400 ;
        RECT 1596.9000 1769.8400 1599.9000 1770.3200 ;
        RECT 1596.9000 1764.4000 1599.9000 1764.8800 ;
        RECT 1596.9000 1775.2800 1599.9000 1775.7600 ;
        RECT 1596.9000 1753.5200 1599.9000 1754.0000 ;
        RECT 1596.9000 1758.9600 1599.9000 1759.4400 ;
        RECT 1596.9000 1742.6400 1599.9000 1743.1200 ;
        RECT 1596.9000 1737.2000 1599.9000 1737.6800 ;
        RECT 1596.9000 1748.0800 1599.9000 1748.5600 ;
        RECT 1691.4600 1726.3200 1693.0600 1726.8000 ;
        RECT 1691.4600 1731.7600 1693.0600 1732.2400 ;
        RECT 1691.4600 1710.0000 1693.0600 1710.4800 ;
        RECT 1691.4600 1715.4400 1693.0600 1715.9200 ;
        RECT 1691.4600 1720.8800 1693.0600 1721.3600 ;
        RECT 1646.4600 1726.3200 1648.0600 1726.8000 ;
        RECT 1646.4600 1731.7600 1648.0600 1732.2400 ;
        RECT 1646.4600 1710.0000 1648.0600 1710.4800 ;
        RECT 1646.4600 1715.4400 1648.0600 1715.9200 ;
        RECT 1646.4600 1720.8800 1648.0600 1721.3600 ;
        RECT 1691.4600 1704.5600 1693.0600 1705.0400 ;
        RECT 1691.4600 1699.1200 1693.0600 1699.6000 ;
        RECT 1691.4600 1693.6800 1693.0600 1694.1600 ;
        RECT 1646.4600 1704.5600 1648.0600 1705.0400 ;
        RECT 1646.4600 1699.1200 1648.0600 1699.6000 ;
        RECT 1646.4600 1693.6800 1648.0600 1694.1600 ;
        RECT 1596.9000 1726.3200 1599.9000 1726.8000 ;
        RECT 1596.9000 1731.7600 1599.9000 1732.2400 ;
        RECT 1596.9000 1715.4400 1599.9000 1715.9200 ;
        RECT 1596.9000 1710.0000 1599.9000 1710.4800 ;
        RECT 1596.9000 1720.8800 1599.9000 1721.3600 ;
        RECT 1596.9000 1699.1200 1599.9000 1699.6000 ;
        RECT 1596.9000 1704.5600 1599.9000 1705.0400 ;
        RECT 1596.9000 1693.6800 1599.9000 1694.1600 ;
        RECT 1596.9000 1891.8700 1796.0000 1894.8700 ;
        RECT 1596.9000 1686.7700 1796.0000 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 1457.1300 1783.0600 1665.2300 ;
        RECT 1736.4600 1457.1300 1738.0600 1665.2300 ;
        RECT 1691.4600 1457.1300 1693.0600 1665.2300 ;
        RECT 1646.4600 1457.1300 1648.0600 1665.2300 ;
        RECT 1793.0000 1457.1300 1796.0000 1665.2300 ;
        RECT 1596.9000 1457.1300 1599.9000 1665.2300 ;
      LAYER met3 ;
        RECT 1793.0000 1659.8800 1796.0000 1660.3600 ;
        RECT 1781.4600 1659.8800 1783.0600 1660.3600 ;
        RECT 1793.0000 1649.0000 1796.0000 1649.4800 ;
        RECT 1793.0000 1654.4400 1796.0000 1654.9200 ;
        RECT 1781.4600 1649.0000 1783.0600 1649.4800 ;
        RECT 1781.4600 1654.4400 1783.0600 1654.9200 ;
        RECT 1793.0000 1632.6800 1796.0000 1633.1600 ;
        RECT 1793.0000 1638.1200 1796.0000 1638.6000 ;
        RECT 1781.4600 1632.6800 1783.0600 1633.1600 ;
        RECT 1781.4600 1638.1200 1783.0600 1638.6000 ;
        RECT 1793.0000 1621.8000 1796.0000 1622.2800 ;
        RECT 1793.0000 1627.2400 1796.0000 1627.7200 ;
        RECT 1781.4600 1621.8000 1783.0600 1622.2800 ;
        RECT 1781.4600 1627.2400 1783.0600 1627.7200 ;
        RECT 1793.0000 1643.5600 1796.0000 1644.0400 ;
        RECT 1781.4600 1643.5600 1783.0600 1644.0400 ;
        RECT 1736.4600 1649.0000 1738.0600 1649.4800 ;
        RECT 1736.4600 1654.4400 1738.0600 1654.9200 ;
        RECT 1736.4600 1659.8800 1738.0600 1660.3600 ;
        RECT 1736.4600 1632.6800 1738.0600 1633.1600 ;
        RECT 1736.4600 1638.1200 1738.0600 1638.6000 ;
        RECT 1736.4600 1627.2400 1738.0600 1627.7200 ;
        RECT 1736.4600 1621.8000 1738.0600 1622.2800 ;
        RECT 1736.4600 1643.5600 1738.0600 1644.0400 ;
        RECT 1793.0000 1605.4800 1796.0000 1605.9600 ;
        RECT 1793.0000 1610.9200 1796.0000 1611.4000 ;
        RECT 1781.4600 1605.4800 1783.0600 1605.9600 ;
        RECT 1781.4600 1610.9200 1783.0600 1611.4000 ;
        RECT 1793.0000 1589.1600 1796.0000 1589.6400 ;
        RECT 1793.0000 1594.6000 1796.0000 1595.0800 ;
        RECT 1793.0000 1600.0400 1796.0000 1600.5200 ;
        RECT 1781.4600 1589.1600 1783.0600 1589.6400 ;
        RECT 1781.4600 1594.6000 1783.0600 1595.0800 ;
        RECT 1781.4600 1600.0400 1783.0600 1600.5200 ;
        RECT 1793.0000 1578.2800 1796.0000 1578.7600 ;
        RECT 1793.0000 1583.7200 1796.0000 1584.2000 ;
        RECT 1781.4600 1578.2800 1783.0600 1578.7600 ;
        RECT 1781.4600 1583.7200 1783.0600 1584.2000 ;
        RECT 1793.0000 1561.9600 1796.0000 1562.4400 ;
        RECT 1793.0000 1567.4000 1796.0000 1567.8800 ;
        RECT 1793.0000 1572.8400 1796.0000 1573.3200 ;
        RECT 1781.4600 1561.9600 1783.0600 1562.4400 ;
        RECT 1781.4600 1567.4000 1783.0600 1567.8800 ;
        RECT 1781.4600 1572.8400 1783.0600 1573.3200 ;
        RECT 1736.4600 1605.4800 1738.0600 1605.9600 ;
        RECT 1736.4600 1610.9200 1738.0600 1611.4000 ;
        RECT 1736.4600 1589.1600 1738.0600 1589.6400 ;
        RECT 1736.4600 1594.6000 1738.0600 1595.0800 ;
        RECT 1736.4600 1600.0400 1738.0600 1600.5200 ;
        RECT 1736.4600 1578.2800 1738.0600 1578.7600 ;
        RECT 1736.4600 1583.7200 1738.0600 1584.2000 ;
        RECT 1736.4600 1561.9600 1738.0600 1562.4400 ;
        RECT 1736.4600 1567.4000 1738.0600 1567.8800 ;
        RECT 1736.4600 1572.8400 1738.0600 1573.3200 ;
        RECT 1793.0000 1616.3600 1796.0000 1616.8400 ;
        RECT 1736.4600 1616.3600 1738.0600 1616.8400 ;
        RECT 1781.4600 1616.3600 1783.0600 1616.8400 ;
        RECT 1691.4600 1649.0000 1693.0600 1649.4800 ;
        RECT 1691.4600 1654.4400 1693.0600 1654.9200 ;
        RECT 1691.4600 1659.8800 1693.0600 1660.3600 ;
        RECT 1646.4600 1649.0000 1648.0600 1649.4800 ;
        RECT 1646.4600 1654.4400 1648.0600 1654.9200 ;
        RECT 1646.4600 1659.8800 1648.0600 1660.3600 ;
        RECT 1691.4600 1632.6800 1693.0600 1633.1600 ;
        RECT 1691.4600 1638.1200 1693.0600 1638.6000 ;
        RECT 1691.4600 1621.8000 1693.0600 1622.2800 ;
        RECT 1691.4600 1627.2400 1693.0600 1627.7200 ;
        RECT 1646.4600 1632.6800 1648.0600 1633.1600 ;
        RECT 1646.4600 1638.1200 1648.0600 1638.6000 ;
        RECT 1646.4600 1621.8000 1648.0600 1622.2800 ;
        RECT 1646.4600 1627.2400 1648.0600 1627.7200 ;
        RECT 1646.4600 1643.5600 1648.0600 1644.0400 ;
        RECT 1691.4600 1643.5600 1693.0600 1644.0400 ;
        RECT 1596.9000 1659.8800 1599.9000 1660.3600 ;
        RECT 1596.9000 1654.4400 1599.9000 1654.9200 ;
        RECT 1596.9000 1649.0000 1599.9000 1649.4800 ;
        RECT 1596.9000 1638.1200 1599.9000 1638.6000 ;
        RECT 1596.9000 1632.6800 1599.9000 1633.1600 ;
        RECT 1596.9000 1627.2400 1599.9000 1627.7200 ;
        RECT 1596.9000 1621.8000 1599.9000 1622.2800 ;
        RECT 1596.9000 1643.5600 1599.9000 1644.0400 ;
        RECT 1691.4600 1605.4800 1693.0600 1605.9600 ;
        RECT 1691.4600 1610.9200 1693.0600 1611.4000 ;
        RECT 1691.4600 1589.1600 1693.0600 1589.6400 ;
        RECT 1691.4600 1594.6000 1693.0600 1595.0800 ;
        RECT 1691.4600 1600.0400 1693.0600 1600.5200 ;
        RECT 1646.4600 1605.4800 1648.0600 1605.9600 ;
        RECT 1646.4600 1610.9200 1648.0600 1611.4000 ;
        RECT 1646.4600 1589.1600 1648.0600 1589.6400 ;
        RECT 1646.4600 1594.6000 1648.0600 1595.0800 ;
        RECT 1646.4600 1600.0400 1648.0600 1600.5200 ;
        RECT 1691.4600 1578.2800 1693.0600 1578.7600 ;
        RECT 1691.4600 1583.7200 1693.0600 1584.2000 ;
        RECT 1691.4600 1561.9600 1693.0600 1562.4400 ;
        RECT 1691.4600 1567.4000 1693.0600 1567.8800 ;
        RECT 1691.4600 1572.8400 1693.0600 1573.3200 ;
        RECT 1646.4600 1578.2800 1648.0600 1578.7600 ;
        RECT 1646.4600 1583.7200 1648.0600 1584.2000 ;
        RECT 1646.4600 1561.9600 1648.0600 1562.4400 ;
        RECT 1646.4600 1567.4000 1648.0600 1567.8800 ;
        RECT 1646.4600 1572.8400 1648.0600 1573.3200 ;
        RECT 1596.9000 1605.4800 1599.9000 1605.9600 ;
        RECT 1596.9000 1610.9200 1599.9000 1611.4000 ;
        RECT 1596.9000 1594.6000 1599.9000 1595.0800 ;
        RECT 1596.9000 1589.1600 1599.9000 1589.6400 ;
        RECT 1596.9000 1600.0400 1599.9000 1600.5200 ;
        RECT 1596.9000 1578.2800 1599.9000 1578.7600 ;
        RECT 1596.9000 1583.7200 1599.9000 1584.2000 ;
        RECT 1596.9000 1567.4000 1599.9000 1567.8800 ;
        RECT 1596.9000 1561.9600 1599.9000 1562.4400 ;
        RECT 1596.9000 1572.8400 1599.9000 1573.3200 ;
        RECT 1596.9000 1616.3600 1599.9000 1616.8400 ;
        RECT 1646.4600 1616.3600 1648.0600 1616.8400 ;
        RECT 1691.4600 1616.3600 1693.0600 1616.8400 ;
        RECT 1793.0000 1551.0800 1796.0000 1551.5600 ;
        RECT 1793.0000 1556.5200 1796.0000 1557.0000 ;
        RECT 1781.4600 1551.0800 1783.0600 1551.5600 ;
        RECT 1781.4600 1556.5200 1783.0600 1557.0000 ;
        RECT 1793.0000 1534.7600 1796.0000 1535.2400 ;
        RECT 1793.0000 1540.2000 1796.0000 1540.6800 ;
        RECT 1793.0000 1545.6400 1796.0000 1546.1200 ;
        RECT 1781.4600 1534.7600 1783.0600 1535.2400 ;
        RECT 1781.4600 1540.2000 1783.0600 1540.6800 ;
        RECT 1781.4600 1545.6400 1783.0600 1546.1200 ;
        RECT 1793.0000 1523.8800 1796.0000 1524.3600 ;
        RECT 1793.0000 1529.3200 1796.0000 1529.8000 ;
        RECT 1781.4600 1523.8800 1783.0600 1524.3600 ;
        RECT 1781.4600 1529.3200 1783.0600 1529.8000 ;
        RECT 1793.0000 1507.5600 1796.0000 1508.0400 ;
        RECT 1793.0000 1513.0000 1796.0000 1513.4800 ;
        RECT 1793.0000 1518.4400 1796.0000 1518.9200 ;
        RECT 1781.4600 1507.5600 1783.0600 1508.0400 ;
        RECT 1781.4600 1513.0000 1783.0600 1513.4800 ;
        RECT 1781.4600 1518.4400 1783.0600 1518.9200 ;
        RECT 1736.4600 1551.0800 1738.0600 1551.5600 ;
        RECT 1736.4600 1556.5200 1738.0600 1557.0000 ;
        RECT 1736.4600 1534.7600 1738.0600 1535.2400 ;
        RECT 1736.4600 1540.2000 1738.0600 1540.6800 ;
        RECT 1736.4600 1545.6400 1738.0600 1546.1200 ;
        RECT 1736.4600 1523.8800 1738.0600 1524.3600 ;
        RECT 1736.4600 1529.3200 1738.0600 1529.8000 ;
        RECT 1736.4600 1507.5600 1738.0600 1508.0400 ;
        RECT 1736.4600 1513.0000 1738.0600 1513.4800 ;
        RECT 1736.4600 1518.4400 1738.0600 1518.9200 ;
        RECT 1793.0000 1496.6800 1796.0000 1497.1600 ;
        RECT 1793.0000 1502.1200 1796.0000 1502.6000 ;
        RECT 1781.4600 1496.6800 1783.0600 1497.1600 ;
        RECT 1781.4600 1502.1200 1783.0600 1502.6000 ;
        RECT 1793.0000 1480.3600 1796.0000 1480.8400 ;
        RECT 1793.0000 1485.8000 1796.0000 1486.2800 ;
        RECT 1793.0000 1491.2400 1796.0000 1491.7200 ;
        RECT 1781.4600 1480.3600 1783.0600 1480.8400 ;
        RECT 1781.4600 1485.8000 1783.0600 1486.2800 ;
        RECT 1781.4600 1491.2400 1783.0600 1491.7200 ;
        RECT 1793.0000 1469.4800 1796.0000 1469.9600 ;
        RECT 1793.0000 1474.9200 1796.0000 1475.4000 ;
        RECT 1781.4600 1469.4800 1783.0600 1469.9600 ;
        RECT 1781.4600 1474.9200 1783.0600 1475.4000 ;
        RECT 1793.0000 1464.0400 1796.0000 1464.5200 ;
        RECT 1781.4600 1464.0400 1783.0600 1464.5200 ;
        RECT 1736.4600 1496.6800 1738.0600 1497.1600 ;
        RECT 1736.4600 1502.1200 1738.0600 1502.6000 ;
        RECT 1736.4600 1480.3600 1738.0600 1480.8400 ;
        RECT 1736.4600 1485.8000 1738.0600 1486.2800 ;
        RECT 1736.4600 1491.2400 1738.0600 1491.7200 ;
        RECT 1736.4600 1469.4800 1738.0600 1469.9600 ;
        RECT 1736.4600 1474.9200 1738.0600 1475.4000 ;
        RECT 1736.4600 1464.0400 1738.0600 1464.5200 ;
        RECT 1691.4600 1551.0800 1693.0600 1551.5600 ;
        RECT 1691.4600 1556.5200 1693.0600 1557.0000 ;
        RECT 1691.4600 1534.7600 1693.0600 1535.2400 ;
        RECT 1691.4600 1540.2000 1693.0600 1540.6800 ;
        RECT 1691.4600 1545.6400 1693.0600 1546.1200 ;
        RECT 1646.4600 1551.0800 1648.0600 1551.5600 ;
        RECT 1646.4600 1556.5200 1648.0600 1557.0000 ;
        RECT 1646.4600 1534.7600 1648.0600 1535.2400 ;
        RECT 1646.4600 1540.2000 1648.0600 1540.6800 ;
        RECT 1646.4600 1545.6400 1648.0600 1546.1200 ;
        RECT 1691.4600 1523.8800 1693.0600 1524.3600 ;
        RECT 1691.4600 1529.3200 1693.0600 1529.8000 ;
        RECT 1691.4600 1507.5600 1693.0600 1508.0400 ;
        RECT 1691.4600 1513.0000 1693.0600 1513.4800 ;
        RECT 1691.4600 1518.4400 1693.0600 1518.9200 ;
        RECT 1646.4600 1523.8800 1648.0600 1524.3600 ;
        RECT 1646.4600 1529.3200 1648.0600 1529.8000 ;
        RECT 1646.4600 1507.5600 1648.0600 1508.0400 ;
        RECT 1646.4600 1513.0000 1648.0600 1513.4800 ;
        RECT 1646.4600 1518.4400 1648.0600 1518.9200 ;
        RECT 1596.9000 1551.0800 1599.9000 1551.5600 ;
        RECT 1596.9000 1556.5200 1599.9000 1557.0000 ;
        RECT 1596.9000 1540.2000 1599.9000 1540.6800 ;
        RECT 1596.9000 1534.7600 1599.9000 1535.2400 ;
        RECT 1596.9000 1545.6400 1599.9000 1546.1200 ;
        RECT 1596.9000 1523.8800 1599.9000 1524.3600 ;
        RECT 1596.9000 1529.3200 1599.9000 1529.8000 ;
        RECT 1596.9000 1513.0000 1599.9000 1513.4800 ;
        RECT 1596.9000 1507.5600 1599.9000 1508.0400 ;
        RECT 1596.9000 1518.4400 1599.9000 1518.9200 ;
        RECT 1691.4600 1496.6800 1693.0600 1497.1600 ;
        RECT 1691.4600 1502.1200 1693.0600 1502.6000 ;
        RECT 1691.4600 1480.3600 1693.0600 1480.8400 ;
        RECT 1691.4600 1485.8000 1693.0600 1486.2800 ;
        RECT 1691.4600 1491.2400 1693.0600 1491.7200 ;
        RECT 1646.4600 1496.6800 1648.0600 1497.1600 ;
        RECT 1646.4600 1502.1200 1648.0600 1502.6000 ;
        RECT 1646.4600 1480.3600 1648.0600 1480.8400 ;
        RECT 1646.4600 1485.8000 1648.0600 1486.2800 ;
        RECT 1646.4600 1491.2400 1648.0600 1491.7200 ;
        RECT 1691.4600 1474.9200 1693.0600 1475.4000 ;
        RECT 1691.4600 1469.4800 1693.0600 1469.9600 ;
        RECT 1691.4600 1464.0400 1693.0600 1464.5200 ;
        RECT 1646.4600 1474.9200 1648.0600 1475.4000 ;
        RECT 1646.4600 1469.4800 1648.0600 1469.9600 ;
        RECT 1646.4600 1464.0400 1648.0600 1464.5200 ;
        RECT 1596.9000 1496.6800 1599.9000 1497.1600 ;
        RECT 1596.9000 1502.1200 1599.9000 1502.6000 ;
        RECT 1596.9000 1485.8000 1599.9000 1486.2800 ;
        RECT 1596.9000 1480.3600 1599.9000 1480.8400 ;
        RECT 1596.9000 1491.2400 1599.9000 1491.7200 ;
        RECT 1596.9000 1469.4800 1599.9000 1469.9600 ;
        RECT 1596.9000 1474.9200 1599.9000 1475.4000 ;
        RECT 1596.9000 1464.0400 1599.9000 1464.5200 ;
        RECT 1596.9000 1662.2300 1796.0000 1665.2300 ;
        RECT 1596.9000 1457.1300 1796.0000 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 1227.4900 1783.0600 1435.5900 ;
        RECT 1736.4600 1227.4900 1738.0600 1435.5900 ;
        RECT 1691.4600 1227.4900 1693.0600 1435.5900 ;
        RECT 1646.4600 1227.4900 1648.0600 1435.5900 ;
        RECT 1793.0000 1227.4900 1796.0000 1435.5900 ;
        RECT 1596.9000 1227.4900 1599.9000 1435.5900 ;
      LAYER met3 ;
        RECT 1793.0000 1430.2400 1796.0000 1430.7200 ;
        RECT 1781.4600 1430.2400 1783.0600 1430.7200 ;
        RECT 1793.0000 1419.3600 1796.0000 1419.8400 ;
        RECT 1793.0000 1424.8000 1796.0000 1425.2800 ;
        RECT 1781.4600 1419.3600 1783.0600 1419.8400 ;
        RECT 1781.4600 1424.8000 1783.0600 1425.2800 ;
        RECT 1793.0000 1403.0400 1796.0000 1403.5200 ;
        RECT 1793.0000 1408.4800 1796.0000 1408.9600 ;
        RECT 1781.4600 1403.0400 1783.0600 1403.5200 ;
        RECT 1781.4600 1408.4800 1783.0600 1408.9600 ;
        RECT 1793.0000 1392.1600 1796.0000 1392.6400 ;
        RECT 1793.0000 1397.6000 1796.0000 1398.0800 ;
        RECT 1781.4600 1392.1600 1783.0600 1392.6400 ;
        RECT 1781.4600 1397.6000 1783.0600 1398.0800 ;
        RECT 1793.0000 1413.9200 1796.0000 1414.4000 ;
        RECT 1781.4600 1413.9200 1783.0600 1414.4000 ;
        RECT 1736.4600 1419.3600 1738.0600 1419.8400 ;
        RECT 1736.4600 1424.8000 1738.0600 1425.2800 ;
        RECT 1736.4600 1430.2400 1738.0600 1430.7200 ;
        RECT 1736.4600 1403.0400 1738.0600 1403.5200 ;
        RECT 1736.4600 1408.4800 1738.0600 1408.9600 ;
        RECT 1736.4600 1397.6000 1738.0600 1398.0800 ;
        RECT 1736.4600 1392.1600 1738.0600 1392.6400 ;
        RECT 1736.4600 1413.9200 1738.0600 1414.4000 ;
        RECT 1793.0000 1375.8400 1796.0000 1376.3200 ;
        RECT 1793.0000 1381.2800 1796.0000 1381.7600 ;
        RECT 1781.4600 1375.8400 1783.0600 1376.3200 ;
        RECT 1781.4600 1381.2800 1783.0600 1381.7600 ;
        RECT 1793.0000 1359.5200 1796.0000 1360.0000 ;
        RECT 1793.0000 1364.9600 1796.0000 1365.4400 ;
        RECT 1793.0000 1370.4000 1796.0000 1370.8800 ;
        RECT 1781.4600 1359.5200 1783.0600 1360.0000 ;
        RECT 1781.4600 1364.9600 1783.0600 1365.4400 ;
        RECT 1781.4600 1370.4000 1783.0600 1370.8800 ;
        RECT 1793.0000 1348.6400 1796.0000 1349.1200 ;
        RECT 1793.0000 1354.0800 1796.0000 1354.5600 ;
        RECT 1781.4600 1348.6400 1783.0600 1349.1200 ;
        RECT 1781.4600 1354.0800 1783.0600 1354.5600 ;
        RECT 1793.0000 1332.3200 1796.0000 1332.8000 ;
        RECT 1793.0000 1337.7600 1796.0000 1338.2400 ;
        RECT 1793.0000 1343.2000 1796.0000 1343.6800 ;
        RECT 1781.4600 1332.3200 1783.0600 1332.8000 ;
        RECT 1781.4600 1337.7600 1783.0600 1338.2400 ;
        RECT 1781.4600 1343.2000 1783.0600 1343.6800 ;
        RECT 1736.4600 1375.8400 1738.0600 1376.3200 ;
        RECT 1736.4600 1381.2800 1738.0600 1381.7600 ;
        RECT 1736.4600 1359.5200 1738.0600 1360.0000 ;
        RECT 1736.4600 1364.9600 1738.0600 1365.4400 ;
        RECT 1736.4600 1370.4000 1738.0600 1370.8800 ;
        RECT 1736.4600 1348.6400 1738.0600 1349.1200 ;
        RECT 1736.4600 1354.0800 1738.0600 1354.5600 ;
        RECT 1736.4600 1332.3200 1738.0600 1332.8000 ;
        RECT 1736.4600 1337.7600 1738.0600 1338.2400 ;
        RECT 1736.4600 1343.2000 1738.0600 1343.6800 ;
        RECT 1793.0000 1386.7200 1796.0000 1387.2000 ;
        RECT 1736.4600 1386.7200 1738.0600 1387.2000 ;
        RECT 1781.4600 1386.7200 1783.0600 1387.2000 ;
        RECT 1691.4600 1419.3600 1693.0600 1419.8400 ;
        RECT 1691.4600 1424.8000 1693.0600 1425.2800 ;
        RECT 1691.4600 1430.2400 1693.0600 1430.7200 ;
        RECT 1646.4600 1419.3600 1648.0600 1419.8400 ;
        RECT 1646.4600 1424.8000 1648.0600 1425.2800 ;
        RECT 1646.4600 1430.2400 1648.0600 1430.7200 ;
        RECT 1691.4600 1403.0400 1693.0600 1403.5200 ;
        RECT 1691.4600 1408.4800 1693.0600 1408.9600 ;
        RECT 1691.4600 1392.1600 1693.0600 1392.6400 ;
        RECT 1691.4600 1397.6000 1693.0600 1398.0800 ;
        RECT 1646.4600 1403.0400 1648.0600 1403.5200 ;
        RECT 1646.4600 1408.4800 1648.0600 1408.9600 ;
        RECT 1646.4600 1392.1600 1648.0600 1392.6400 ;
        RECT 1646.4600 1397.6000 1648.0600 1398.0800 ;
        RECT 1646.4600 1413.9200 1648.0600 1414.4000 ;
        RECT 1691.4600 1413.9200 1693.0600 1414.4000 ;
        RECT 1596.9000 1430.2400 1599.9000 1430.7200 ;
        RECT 1596.9000 1424.8000 1599.9000 1425.2800 ;
        RECT 1596.9000 1419.3600 1599.9000 1419.8400 ;
        RECT 1596.9000 1408.4800 1599.9000 1408.9600 ;
        RECT 1596.9000 1403.0400 1599.9000 1403.5200 ;
        RECT 1596.9000 1397.6000 1599.9000 1398.0800 ;
        RECT 1596.9000 1392.1600 1599.9000 1392.6400 ;
        RECT 1596.9000 1413.9200 1599.9000 1414.4000 ;
        RECT 1691.4600 1375.8400 1693.0600 1376.3200 ;
        RECT 1691.4600 1381.2800 1693.0600 1381.7600 ;
        RECT 1691.4600 1359.5200 1693.0600 1360.0000 ;
        RECT 1691.4600 1364.9600 1693.0600 1365.4400 ;
        RECT 1691.4600 1370.4000 1693.0600 1370.8800 ;
        RECT 1646.4600 1375.8400 1648.0600 1376.3200 ;
        RECT 1646.4600 1381.2800 1648.0600 1381.7600 ;
        RECT 1646.4600 1359.5200 1648.0600 1360.0000 ;
        RECT 1646.4600 1364.9600 1648.0600 1365.4400 ;
        RECT 1646.4600 1370.4000 1648.0600 1370.8800 ;
        RECT 1691.4600 1348.6400 1693.0600 1349.1200 ;
        RECT 1691.4600 1354.0800 1693.0600 1354.5600 ;
        RECT 1691.4600 1332.3200 1693.0600 1332.8000 ;
        RECT 1691.4600 1337.7600 1693.0600 1338.2400 ;
        RECT 1691.4600 1343.2000 1693.0600 1343.6800 ;
        RECT 1646.4600 1348.6400 1648.0600 1349.1200 ;
        RECT 1646.4600 1354.0800 1648.0600 1354.5600 ;
        RECT 1646.4600 1332.3200 1648.0600 1332.8000 ;
        RECT 1646.4600 1337.7600 1648.0600 1338.2400 ;
        RECT 1646.4600 1343.2000 1648.0600 1343.6800 ;
        RECT 1596.9000 1375.8400 1599.9000 1376.3200 ;
        RECT 1596.9000 1381.2800 1599.9000 1381.7600 ;
        RECT 1596.9000 1364.9600 1599.9000 1365.4400 ;
        RECT 1596.9000 1359.5200 1599.9000 1360.0000 ;
        RECT 1596.9000 1370.4000 1599.9000 1370.8800 ;
        RECT 1596.9000 1348.6400 1599.9000 1349.1200 ;
        RECT 1596.9000 1354.0800 1599.9000 1354.5600 ;
        RECT 1596.9000 1337.7600 1599.9000 1338.2400 ;
        RECT 1596.9000 1332.3200 1599.9000 1332.8000 ;
        RECT 1596.9000 1343.2000 1599.9000 1343.6800 ;
        RECT 1596.9000 1386.7200 1599.9000 1387.2000 ;
        RECT 1646.4600 1386.7200 1648.0600 1387.2000 ;
        RECT 1691.4600 1386.7200 1693.0600 1387.2000 ;
        RECT 1793.0000 1321.4400 1796.0000 1321.9200 ;
        RECT 1793.0000 1326.8800 1796.0000 1327.3600 ;
        RECT 1781.4600 1321.4400 1783.0600 1321.9200 ;
        RECT 1781.4600 1326.8800 1783.0600 1327.3600 ;
        RECT 1793.0000 1305.1200 1796.0000 1305.6000 ;
        RECT 1793.0000 1310.5600 1796.0000 1311.0400 ;
        RECT 1793.0000 1316.0000 1796.0000 1316.4800 ;
        RECT 1781.4600 1305.1200 1783.0600 1305.6000 ;
        RECT 1781.4600 1310.5600 1783.0600 1311.0400 ;
        RECT 1781.4600 1316.0000 1783.0600 1316.4800 ;
        RECT 1793.0000 1294.2400 1796.0000 1294.7200 ;
        RECT 1793.0000 1299.6800 1796.0000 1300.1600 ;
        RECT 1781.4600 1294.2400 1783.0600 1294.7200 ;
        RECT 1781.4600 1299.6800 1783.0600 1300.1600 ;
        RECT 1793.0000 1277.9200 1796.0000 1278.4000 ;
        RECT 1793.0000 1283.3600 1796.0000 1283.8400 ;
        RECT 1793.0000 1288.8000 1796.0000 1289.2800 ;
        RECT 1781.4600 1277.9200 1783.0600 1278.4000 ;
        RECT 1781.4600 1283.3600 1783.0600 1283.8400 ;
        RECT 1781.4600 1288.8000 1783.0600 1289.2800 ;
        RECT 1736.4600 1321.4400 1738.0600 1321.9200 ;
        RECT 1736.4600 1326.8800 1738.0600 1327.3600 ;
        RECT 1736.4600 1305.1200 1738.0600 1305.6000 ;
        RECT 1736.4600 1310.5600 1738.0600 1311.0400 ;
        RECT 1736.4600 1316.0000 1738.0600 1316.4800 ;
        RECT 1736.4600 1294.2400 1738.0600 1294.7200 ;
        RECT 1736.4600 1299.6800 1738.0600 1300.1600 ;
        RECT 1736.4600 1277.9200 1738.0600 1278.4000 ;
        RECT 1736.4600 1283.3600 1738.0600 1283.8400 ;
        RECT 1736.4600 1288.8000 1738.0600 1289.2800 ;
        RECT 1793.0000 1267.0400 1796.0000 1267.5200 ;
        RECT 1793.0000 1272.4800 1796.0000 1272.9600 ;
        RECT 1781.4600 1267.0400 1783.0600 1267.5200 ;
        RECT 1781.4600 1272.4800 1783.0600 1272.9600 ;
        RECT 1793.0000 1250.7200 1796.0000 1251.2000 ;
        RECT 1793.0000 1256.1600 1796.0000 1256.6400 ;
        RECT 1793.0000 1261.6000 1796.0000 1262.0800 ;
        RECT 1781.4600 1250.7200 1783.0600 1251.2000 ;
        RECT 1781.4600 1256.1600 1783.0600 1256.6400 ;
        RECT 1781.4600 1261.6000 1783.0600 1262.0800 ;
        RECT 1793.0000 1239.8400 1796.0000 1240.3200 ;
        RECT 1793.0000 1245.2800 1796.0000 1245.7600 ;
        RECT 1781.4600 1239.8400 1783.0600 1240.3200 ;
        RECT 1781.4600 1245.2800 1783.0600 1245.7600 ;
        RECT 1793.0000 1234.4000 1796.0000 1234.8800 ;
        RECT 1781.4600 1234.4000 1783.0600 1234.8800 ;
        RECT 1736.4600 1267.0400 1738.0600 1267.5200 ;
        RECT 1736.4600 1272.4800 1738.0600 1272.9600 ;
        RECT 1736.4600 1250.7200 1738.0600 1251.2000 ;
        RECT 1736.4600 1256.1600 1738.0600 1256.6400 ;
        RECT 1736.4600 1261.6000 1738.0600 1262.0800 ;
        RECT 1736.4600 1239.8400 1738.0600 1240.3200 ;
        RECT 1736.4600 1245.2800 1738.0600 1245.7600 ;
        RECT 1736.4600 1234.4000 1738.0600 1234.8800 ;
        RECT 1691.4600 1321.4400 1693.0600 1321.9200 ;
        RECT 1691.4600 1326.8800 1693.0600 1327.3600 ;
        RECT 1691.4600 1305.1200 1693.0600 1305.6000 ;
        RECT 1691.4600 1310.5600 1693.0600 1311.0400 ;
        RECT 1691.4600 1316.0000 1693.0600 1316.4800 ;
        RECT 1646.4600 1321.4400 1648.0600 1321.9200 ;
        RECT 1646.4600 1326.8800 1648.0600 1327.3600 ;
        RECT 1646.4600 1305.1200 1648.0600 1305.6000 ;
        RECT 1646.4600 1310.5600 1648.0600 1311.0400 ;
        RECT 1646.4600 1316.0000 1648.0600 1316.4800 ;
        RECT 1691.4600 1294.2400 1693.0600 1294.7200 ;
        RECT 1691.4600 1299.6800 1693.0600 1300.1600 ;
        RECT 1691.4600 1277.9200 1693.0600 1278.4000 ;
        RECT 1691.4600 1283.3600 1693.0600 1283.8400 ;
        RECT 1691.4600 1288.8000 1693.0600 1289.2800 ;
        RECT 1646.4600 1294.2400 1648.0600 1294.7200 ;
        RECT 1646.4600 1299.6800 1648.0600 1300.1600 ;
        RECT 1646.4600 1277.9200 1648.0600 1278.4000 ;
        RECT 1646.4600 1283.3600 1648.0600 1283.8400 ;
        RECT 1646.4600 1288.8000 1648.0600 1289.2800 ;
        RECT 1596.9000 1321.4400 1599.9000 1321.9200 ;
        RECT 1596.9000 1326.8800 1599.9000 1327.3600 ;
        RECT 1596.9000 1310.5600 1599.9000 1311.0400 ;
        RECT 1596.9000 1305.1200 1599.9000 1305.6000 ;
        RECT 1596.9000 1316.0000 1599.9000 1316.4800 ;
        RECT 1596.9000 1294.2400 1599.9000 1294.7200 ;
        RECT 1596.9000 1299.6800 1599.9000 1300.1600 ;
        RECT 1596.9000 1283.3600 1599.9000 1283.8400 ;
        RECT 1596.9000 1277.9200 1599.9000 1278.4000 ;
        RECT 1596.9000 1288.8000 1599.9000 1289.2800 ;
        RECT 1691.4600 1267.0400 1693.0600 1267.5200 ;
        RECT 1691.4600 1272.4800 1693.0600 1272.9600 ;
        RECT 1691.4600 1250.7200 1693.0600 1251.2000 ;
        RECT 1691.4600 1256.1600 1693.0600 1256.6400 ;
        RECT 1691.4600 1261.6000 1693.0600 1262.0800 ;
        RECT 1646.4600 1267.0400 1648.0600 1267.5200 ;
        RECT 1646.4600 1272.4800 1648.0600 1272.9600 ;
        RECT 1646.4600 1250.7200 1648.0600 1251.2000 ;
        RECT 1646.4600 1256.1600 1648.0600 1256.6400 ;
        RECT 1646.4600 1261.6000 1648.0600 1262.0800 ;
        RECT 1691.4600 1245.2800 1693.0600 1245.7600 ;
        RECT 1691.4600 1239.8400 1693.0600 1240.3200 ;
        RECT 1691.4600 1234.4000 1693.0600 1234.8800 ;
        RECT 1646.4600 1245.2800 1648.0600 1245.7600 ;
        RECT 1646.4600 1239.8400 1648.0600 1240.3200 ;
        RECT 1646.4600 1234.4000 1648.0600 1234.8800 ;
        RECT 1596.9000 1267.0400 1599.9000 1267.5200 ;
        RECT 1596.9000 1272.4800 1599.9000 1272.9600 ;
        RECT 1596.9000 1256.1600 1599.9000 1256.6400 ;
        RECT 1596.9000 1250.7200 1599.9000 1251.2000 ;
        RECT 1596.9000 1261.6000 1599.9000 1262.0800 ;
        RECT 1596.9000 1239.8400 1599.9000 1240.3200 ;
        RECT 1596.9000 1245.2800 1599.9000 1245.7600 ;
        RECT 1596.9000 1234.4000 1599.9000 1234.8800 ;
        RECT 1596.9000 1432.5900 1796.0000 1435.5900 ;
        RECT 1596.9000 1227.4900 1796.0000 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 997.8500 1783.0600 1205.9500 ;
        RECT 1736.4600 997.8500 1738.0600 1205.9500 ;
        RECT 1691.4600 997.8500 1693.0600 1205.9500 ;
        RECT 1646.4600 997.8500 1648.0600 1205.9500 ;
        RECT 1793.0000 997.8500 1796.0000 1205.9500 ;
        RECT 1596.9000 997.8500 1599.9000 1205.9500 ;
      LAYER met3 ;
        RECT 1793.0000 1200.6000 1796.0000 1201.0800 ;
        RECT 1781.4600 1200.6000 1783.0600 1201.0800 ;
        RECT 1793.0000 1189.7200 1796.0000 1190.2000 ;
        RECT 1793.0000 1195.1600 1796.0000 1195.6400 ;
        RECT 1781.4600 1189.7200 1783.0600 1190.2000 ;
        RECT 1781.4600 1195.1600 1783.0600 1195.6400 ;
        RECT 1793.0000 1173.4000 1796.0000 1173.8800 ;
        RECT 1793.0000 1178.8400 1796.0000 1179.3200 ;
        RECT 1781.4600 1173.4000 1783.0600 1173.8800 ;
        RECT 1781.4600 1178.8400 1783.0600 1179.3200 ;
        RECT 1793.0000 1162.5200 1796.0000 1163.0000 ;
        RECT 1793.0000 1167.9600 1796.0000 1168.4400 ;
        RECT 1781.4600 1162.5200 1783.0600 1163.0000 ;
        RECT 1781.4600 1167.9600 1783.0600 1168.4400 ;
        RECT 1793.0000 1184.2800 1796.0000 1184.7600 ;
        RECT 1781.4600 1184.2800 1783.0600 1184.7600 ;
        RECT 1736.4600 1189.7200 1738.0600 1190.2000 ;
        RECT 1736.4600 1195.1600 1738.0600 1195.6400 ;
        RECT 1736.4600 1200.6000 1738.0600 1201.0800 ;
        RECT 1736.4600 1173.4000 1738.0600 1173.8800 ;
        RECT 1736.4600 1178.8400 1738.0600 1179.3200 ;
        RECT 1736.4600 1167.9600 1738.0600 1168.4400 ;
        RECT 1736.4600 1162.5200 1738.0600 1163.0000 ;
        RECT 1736.4600 1184.2800 1738.0600 1184.7600 ;
        RECT 1793.0000 1146.2000 1796.0000 1146.6800 ;
        RECT 1793.0000 1151.6400 1796.0000 1152.1200 ;
        RECT 1781.4600 1146.2000 1783.0600 1146.6800 ;
        RECT 1781.4600 1151.6400 1783.0600 1152.1200 ;
        RECT 1793.0000 1129.8800 1796.0000 1130.3600 ;
        RECT 1793.0000 1135.3200 1796.0000 1135.8000 ;
        RECT 1793.0000 1140.7600 1796.0000 1141.2400 ;
        RECT 1781.4600 1129.8800 1783.0600 1130.3600 ;
        RECT 1781.4600 1135.3200 1783.0600 1135.8000 ;
        RECT 1781.4600 1140.7600 1783.0600 1141.2400 ;
        RECT 1793.0000 1119.0000 1796.0000 1119.4800 ;
        RECT 1793.0000 1124.4400 1796.0000 1124.9200 ;
        RECT 1781.4600 1119.0000 1783.0600 1119.4800 ;
        RECT 1781.4600 1124.4400 1783.0600 1124.9200 ;
        RECT 1793.0000 1102.6800 1796.0000 1103.1600 ;
        RECT 1793.0000 1108.1200 1796.0000 1108.6000 ;
        RECT 1793.0000 1113.5600 1796.0000 1114.0400 ;
        RECT 1781.4600 1102.6800 1783.0600 1103.1600 ;
        RECT 1781.4600 1108.1200 1783.0600 1108.6000 ;
        RECT 1781.4600 1113.5600 1783.0600 1114.0400 ;
        RECT 1736.4600 1146.2000 1738.0600 1146.6800 ;
        RECT 1736.4600 1151.6400 1738.0600 1152.1200 ;
        RECT 1736.4600 1129.8800 1738.0600 1130.3600 ;
        RECT 1736.4600 1135.3200 1738.0600 1135.8000 ;
        RECT 1736.4600 1140.7600 1738.0600 1141.2400 ;
        RECT 1736.4600 1119.0000 1738.0600 1119.4800 ;
        RECT 1736.4600 1124.4400 1738.0600 1124.9200 ;
        RECT 1736.4600 1102.6800 1738.0600 1103.1600 ;
        RECT 1736.4600 1108.1200 1738.0600 1108.6000 ;
        RECT 1736.4600 1113.5600 1738.0600 1114.0400 ;
        RECT 1793.0000 1157.0800 1796.0000 1157.5600 ;
        RECT 1736.4600 1157.0800 1738.0600 1157.5600 ;
        RECT 1781.4600 1157.0800 1783.0600 1157.5600 ;
        RECT 1691.4600 1189.7200 1693.0600 1190.2000 ;
        RECT 1691.4600 1195.1600 1693.0600 1195.6400 ;
        RECT 1691.4600 1200.6000 1693.0600 1201.0800 ;
        RECT 1646.4600 1189.7200 1648.0600 1190.2000 ;
        RECT 1646.4600 1195.1600 1648.0600 1195.6400 ;
        RECT 1646.4600 1200.6000 1648.0600 1201.0800 ;
        RECT 1691.4600 1173.4000 1693.0600 1173.8800 ;
        RECT 1691.4600 1178.8400 1693.0600 1179.3200 ;
        RECT 1691.4600 1162.5200 1693.0600 1163.0000 ;
        RECT 1691.4600 1167.9600 1693.0600 1168.4400 ;
        RECT 1646.4600 1173.4000 1648.0600 1173.8800 ;
        RECT 1646.4600 1178.8400 1648.0600 1179.3200 ;
        RECT 1646.4600 1162.5200 1648.0600 1163.0000 ;
        RECT 1646.4600 1167.9600 1648.0600 1168.4400 ;
        RECT 1646.4600 1184.2800 1648.0600 1184.7600 ;
        RECT 1691.4600 1184.2800 1693.0600 1184.7600 ;
        RECT 1596.9000 1200.6000 1599.9000 1201.0800 ;
        RECT 1596.9000 1195.1600 1599.9000 1195.6400 ;
        RECT 1596.9000 1189.7200 1599.9000 1190.2000 ;
        RECT 1596.9000 1178.8400 1599.9000 1179.3200 ;
        RECT 1596.9000 1173.4000 1599.9000 1173.8800 ;
        RECT 1596.9000 1167.9600 1599.9000 1168.4400 ;
        RECT 1596.9000 1162.5200 1599.9000 1163.0000 ;
        RECT 1596.9000 1184.2800 1599.9000 1184.7600 ;
        RECT 1691.4600 1146.2000 1693.0600 1146.6800 ;
        RECT 1691.4600 1151.6400 1693.0600 1152.1200 ;
        RECT 1691.4600 1129.8800 1693.0600 1130.3600 ;
        RECT 1691.4600 1135.3200 1693.0600 1135.8000 ;
        RECT 1691.4600 1140.7600 1693.0600 1141.2400 ;
        RECT 1646.4600 1146.2000 1648.0600 1146.6800 ;
        RECT 1646.4600 1151.6400 1648.0600 1152.1200 ;
        RECT 1646.4600 1129.8800 1648.0600 1130.3600 ;
        RECT 1646.4600 1135.3200 1648.0600 1135.8000 ;
        RECT 1646.4600 1140.7600 1648.0600 1141.2400 ;
        RECT 1691.4600 1119.0000 1693.0600 1119.4800 ;
        RECT 1691.4600 1124.4400 1693.0600 1124.9200 ;
        RECT 1691.4600 1102.6800 1693.0600 1103.1600 ;
        RECT 1691.4600 1108.1200 1693.0600 1108.6000 ;
        RECT 1691.4600 1113.5600 1693.0600 1114.0400 ;
        RECT 1646.4600 1119.0000 1648.0600 1119.4800 ;
        RECT 1646.4600 1124.4400 1648.0600 1124.9200 ;
        RECT 1646.4600 1102.6800 1648.0600 1103.1600 ;
        RECT 1646.4600 1108.1200 1648.0600 1108.6000 ;
        RECT 1646.4600 1113.5600 1648.0600 1114.0400 ;
        RECT 1596.9000 1146.2000 1599.9000 1146.6800 ;
        RECT 1596.9000 1151.6400 1599.9000 1152.1200 ;
        RECT 1596.9000 1135.3200 1599.9000 1135.8000 ;
        RECT 1596.9000 1129.8800 1599.9000 1130.3600 ;
        RECT 1596.9000 1140.7600 1599.9000 1141.2400 ;
        RECT 1596.9000 1119.0000 1599.9000 1119.4800 ;
        RECT 1596.9000 1124.4400 1599.9000 1124.9200 ;
        RECT 1596.9000 1108.1200 1599.9000 1108.6000 ;
        RECT 1596.9000 1102.6800 1599.9000 1103.1600 ;
        RECT 1596.9000 1113.5600 1599.9000 1114.0400 ;
        RECT 1596.9000 1157.0800 1599.9000 1157.5600 ;
        RECT 1646.4600 1157.0800 1648.0600 1157.5600 ;
        RECT 1691.4600 1157.0800 1693.0600 1157.5600 ;
        RECT 1793.0000 1091.8000 1796.0000 1092.2800 ;
        RECT 1793.0000 1097.2400 1796.0000 1097.7200 ;
        RECT 1781.4600 1091.8000 1783.0600 1092.2800 ;
        RECT 1781.4600 1097.2400 1783.0600 1097.7200 ;
        RECT 1793.0000 1075.4800 1796.0000 1075.9600 ;
        RECT 1793.0000 1080.9200 1796.0000 1081.4000 ;
        RECT 1793.0000 1086.3600 1796.0000 1086.8400 ;
        RECT 1781.4600 1075.4800 1783.0600 1075.9600 ;
        RECT 1781.4600 1080.9200 1783.0600 1081.4000 ;
        RECT 1781.4600 1086.3600 1783.0600 1086.8400 ;
        RECT 1793.0000 1064.6000 1796.0000 1065.0800 ;
        RECT 1793.0000 1070.0400 1796.0000 1070.5200 ;
        RECT 1781.4600 1064.6000 1783.0600 1065.0800 ;
        RECT 1781.4600 1070.0400 1783.0600 1070.5200 ;
        RECT 1793.0000 1048.2800 1796.0000 1048.7600 ;
        RECT 1793.0000 1053.7200 1796.0000 1054.2000 ;
        RECT 1793.0000 1059.1600 1796.0000 1059.6400 ;
        RECT 1781.4600 1048.2800 1783.0600 1048.7600 ;
        RECT 1781.4600 1053.7200 1783.0600 1054.2000 ;
        RECT 1781.4600 1059.1600 1783.0600 1059.6400 ;
        RECT 1736.4600 1091.8000 1738.0600 1092.2800 ;
        RECT 1736.4600 1097.2400 1738.0600 1097.7200 ;
        RECT 1736.4600 1075.4800 1738.0600 1075.9600 ;
        RECT 1736.4600 1080.9200 1738.0600 1081.4000 ;
        RECT 1736.4600 1086.3600 1738.0600 1086.8400 ;
        RECT 1736.4600 1064.6000 1738.0600 1065.0800 ;
        RECT 1736.4600 1070.0400 1738.0600 1070.5200 ;
        RECT 1736.4600 1048.2800 1738.0600 1048.7600 ;
        RECT 1736.4600 1053.7200 1738.0600 1054.2000 ;
        RECT 1736.4600 1059.1600 1738.0600 1059.6400 ;
        RECT 1793.0000 1037.4000 1796.0000 1037.8800 ;
        RECT 1793.0000 1042.8400 1796.0000 1043.3200 ;
        RECT 1781.4600 1037.4000 1783.0600 1037.8800 ;
        RECT 1781.4600 1042.8400 1783.0600 1043.3200 ;
        RECT 1793.0000 1021.0800 1796.0000 1021.5600 ;
        RECT 1793.0000 1026.5200 1796.0000 1027.0000 ;
        RECT 1793.0000 1031.9600 1796.0000 1032.4400 ;
        RECT 1781.4600 1021.0800 1783.0600 1021.5600 ;
        RECT 1781.4600 1026.5200 1783.0600 1027.0000 ;
        RECT 1781.4600 1031.9600 1783.0600 1032.4400 ;
        RECT 1793.0000 1010.2000 1796.0000 1010.6800 ;
        RECT 1793.0000 1015.6400 1796.0000 1016.1200 ;
        RECT 1781.4600 1010.2000 1783.0600 1010.6800 ;
        RECT 1781.4600 1015.6400 1783.0600 1016.1200 ;
        RECT 1793.0000 1004.7600 1796.0000 1005.2400 ;
        RECT 1781.4600 1004.7600 1783.0600 1005.2400 ;
        RECT 1736.4600 1037.4000 1738.0600 1037.8800 ;
        RECT 1736.4600 1042.8400 1738.0600 1043.3200 ;
        RECT 1736.4600 1021.0800 1738.0600 1021.5600 ;
        RECT 1736.4600 1026.5200 1738.0600 1027.0000 ;
        RECT 1736.4600 1031.9600 1738.0600 1032.4400 ;
        RECT 1736.4600 1010.2000 1738.0600 1010.6800 ;
        RECT 1736.4600 1015.6400 1738.0600 1016.1200 ;
        RECT 1736.4600 1004.7600 1738.0600 1005.2400 ;
        RECT 1691.4600 1091.8000 1693.0600 1092.2800 ;
        RECT 1691.4600 1097.2400 1693.0600 1097.7200 ;
        RECT 1691.4600 1075.4800 1693.0600 1075.9600 ;
        RECT 1691.4600 1080.9200 1693.0600 1081.4000 ;
        RECT 1691.4600 1086.3600 1693.0600 1086.8400 ;
        RECT 1646.4600 1091.8000 1648.0600 1092.2800 ;
        RECT 1646.4600 1097.2400 1648.0600 1097.7200 ;
        RECT 1646.4600 1075.4800 1648.0600 1075.9600 ;
        RECT 1646.4600 1080.9200 1648.0600 1081.4000 ;
        RECT 1646.4600 1086.3600 1648.0600 1086.8400 ;
        RECT 1691.4600 1064.6000 1693.0600 1065.0800 ;
        RECT 1691.4600 1070.0400 1693.0600 1070.5200 ;
        RECT 1691.4600 1048.2800 1693.0600 1048.7600 ;
        RECT 1691.4600 1053.7200 1693.0600 1054.2000 ;
        RECT 1691.4600 1059.1600 1693.0600 1059.6400 ;
        RECT 1646.4600 1064.6000 1648.0600 1065.0800 ;
        RECT 1646.4600 1070.0400 1648.0600 1070.5200 ;
        RECT 1646.4600 1048.2800 1648.0600 1048.7600 ;
        RECT 1646.4600 1053.7200 1648.0600 1054.2000 ;
        RECT 1646.4600 1059.1600 1648.0600 1059.6400 ;
        RECT 1596.9000 1091.8000 1599.9000 1092.2800 ;
        RECT 1596.9000 1097.2400 1599.9000 1097.7200 ;
        RECT 1596.9000 1080.9200 1599.9000 1081.4000 ;
        RECT 1596.9000 1075.4800 1599.9000 1075.9600 ;
        RECT 1596.9000 1086.3600 1599.9000 1086.8400 ;
        RECT 1596.9000 1064.6000 1599.9000 1065.0800 ;
        RECT 1596.9000 1070.0400 1599.9000 1070.5200 ;
        RECT 1596.9000 1053.7200 1599.9000 1054.2000 ;
        RECT 1596.9000 1048.2800 1599.9000 1048.7600 ;
        RECT 1596.9000 1059.1600 1599.9000 1059.6400 ;
        RECT 1691.4600 1037.4000 1693.0600 1037.8800 ;
        RECT 1691.4600 1042.8400 1693.0600 1043.3200 ;
        RECT 1691.4600 1021.0800 1693.0600 1021.5600 ;
        RECT 1691.4600 1026.5200 1693.0600 1027.0000 ;
        RECT 1691.4600 1031.9600 1693.0600 1032.4400 ;
        RECT 1646.4600 1037.4000 1648.0600 1037.8800 ;
        RECT 1646.4600 1042.8400 1648.0600 1043.3200 ;
        RECT 1646.4600 1021.0800 1648.0600 1021.5600 ;
        RECT 1646.4600 1026.5200 1648.0600 1027.0000 ;
        RECT 1646.4600 1031.9600 1648.0600 1032.4400 ;
        RECT 1691.4600 1015.6400 1693.0600 1016.1200 ;
        RECT 1691.4600 1010.2000 1693.0600 1010.6800 ;
        RECT 1691.4600 1004.7600 1693.0600 1005.2400 ;
        RECT 1646.4600 1015.6400 1648.0600 1016.1200 ;
        RECT 1646.4600 1010.2000 1648.0600 1010.6800 ;
        RECT 1646.4600 1004.7600 1648.0600 1005.2400 ;
        RECT 1596.9000 1037.4000 1599.9000 1037.8800 ;
        RECT 1596.9000 1042.8400 1599.9000 1043.3200 ;
        RECT 1596.9000 1026.5200 1599.9000 1027.0000 ;
        RECT 1596.9000 1021.0800 1599.9000 1021.5600 ;
        RECT 1596.9000 1031.9600 1599.9000 1032.4400 ;
        RECT 1596.9000 1010.2000 1599.9000 1010.6800 ;
        RECT 1596.9000 1015.6400 1599.9000 1016.1200 ;
        RECT 1596.9000 1004.7600 1599.9000 1005.2400 ;
        RECT 1596.9000 1202.9500 1796.0000 1205.9500 ;
        RECT 1596.9000 997.8500 1796.0000 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1781.4600 768.2100 1783.0600 976.3100 ;
        RECT 1736.4600 768.2100 1738.0600 976.3100 ;
        RECT 1691.4600 768.2100 1693.0600 976.3100 ;
        RECT 1646.4600 768.2100 1648.0600 976.3100 ;
        RECT 1793.0000 768.2100 1796.0000 976.3100 ;
        RECT 1596.9000 768.2100 1599.9000 976.3100 ;
      LAYER met3 ;
        RECT 1793.0000 970.9600 1796.0000 971.4400 ;
        RECT 1781.4600 970.9600 1783.0600 971.4400 ;
        RECT 1793.0000 960.0800 1796.0000 960.5600 ;
        RECT 1793.0000 965.5200 1796.0000 966.0000 ;
        RECT 1781.4600 960.0800 1783.0600 960.5600 ;
        RECT 1781.4600 965.5200 1783.0600 966.0000 ;
        RECT 1793.0000 943.7600 1796.0000 944.2400 ;
        RECT 1793.0000 949.2000 1796.0000 949.6800 ;
        RECT 1781.4600 943.7600 1783.0600 944.2400 ;
        RECT 1781.4600 949.2000 1783.0600 949.6800 ;
        RECT 1793.0000 932.8800 1796.0000 933.3600 ;
        RECT 1793.0000 938.3200 1796.0000 938.8000 ;
        RECT 1781.4600 932.8800 1783.0600 933.3600 ;
        RECT 1781.4600 938.3200 1783.0600 938.8000 ;
        RECT 1793.0000 954.6400 1796.0000 955.1200 ;
        RECT 1781.4600 954.6400 1783.0600 955.1200 ;
        RECT 1736.4600 960.0800 1738.0600 960.5600 ;
        RECT 1736.4600 965.5200 1738.0600 966.0000 ;
        RECT 1736.4600 970.9600 1738.0600 971.4400 ;
        RECT 1736.4600 943.7600 1738.0600 944.2400 ;
        RECT 1736.4600 949.2000 1738.0600 949.6800 ;
        RECT 1736.4600 938.3200 1738.0600 938.8000 ;
        RECT 1736.4600 932.8800 1738.0600 933.3600 ;
        RECT 1736.4600 954.6400 1738.0600 955.1200 ;
        RECT 1793.0000 916.5600 1796.0000 917.0400 ;
        RECT 1793.0000 922.0000 1796.0000 922.4800 ;
        RECT 1781.4600 916.5600 1783.0600 917.0400 ;
        RECT 1781.4600 922.0000 1783.0600 922.4800 ;
        RECT 1793.0000 900.2400 1796.0000 900.7200 ;
        RECT 1793.0000 905.6800 1796.0000 906.1600 ;
        RECT 1793.0000 911.1200 1796.0000 911.6000 ;
        RECT 1781.4600 900.2400 1783.0600 900.7200 ;
        RECT 1781.4600 905.6800 1783.0600 906.1600 ;
        RECT 1781.4600 911.1200 1783.0600 911.6000 ;
        RECT 1793.0000 889.3600 1796.0000 889.8400 ;
        RECT 1793.0000 894.8000 1796.0000 895.2800 ;
        RECT 1781.4600 889.3600 1783.0600 889.8400 ;
        RECT 1781.4600 894.8000 1783.0600 895.2800 ;
        RECT 1793.0000 873.0400 1796.0000 873.5200 ;
        RECT 1793.0000 878.4800 1796.0000 878.9600 ;
        RECT 1793.0000 883.9200 1796.0000 884.4000 ;
        RECT 1781.4600 873.0400 1783.0600 873.5200 ;
        RECT 1781.4600 878.4800 1783.0600 878.9600 ;
        RECT 1781.4600 883.9200 1783.0600 884.4000 ;
        RECT 1736.4600 916.5600 1738.0600 917.0400 ;
        RECT 1736.4600 922.0000 1738.0600 922.4800 ;
        RECT 1736.4600 900.2400 1738.0600 900.7200 ;
        RECT 1736.4600 905.6800 1738.0600 906.1600 ;
        RECT 1736.4600 911.1200 1738.0600 911.6000 ;
        RECT 1736.4600 889.3600 1738.0600 889.8400 ;
        RECT 1736.4600 894.8000 1738.0600 895.2800 ;
        RECT 1736.4600 873.0400 1738.0600 873.5200 ;
        RECT 1736.4600 878.4800 1738.0600 878.9600 ;
        RECT 1736.4600 883.9200 1738.0600 884.4000 ;
        RECT 1793.0000 927.4400 1796.0000 927.9200 ;
        RECT 1736.4600 927.4400 1738.0600 927.9200 ;
        RECT 1781.4600 927.4400 1783.0600 927.9200 ;
        RECT 1691.4600 960.0800 1693.0600 960.5600 ;
        RECT 1691.4600 965.5200 1693.0600 966.0000 ;
        RECT 1691.4600 970.9600 1693.0600 971.4400 ;
        RECT 1646.4600 960.0800 1648.0600 960.5600 ;
        RECT 1646.4600 965.5200 1648.0600 966.0000 ;
        RECT 1646.4600 970.9600 1648.0600 971.4400 ;
        RECT 1691.4600 943.7600 1693.0600 944.2400 ;
        RECT 1691.4600 949.2000 1693.0600 949.6800 ;
        RECT 1691.4600 932.8800 1693.0600 933.3600 ;
        RECT 1691.4600 938.3200 1693.0600 938.8000 ;
        RECT 1646.4600 943.7600 1648.0600 944.2400 ;
        RECT 1646.4600 949.2000 1648.0600 949.6800 ;
        RECT 1646.4600 932.8800 1648.0600 933.3600 ;
        RECT 1646.4600 938.3200 1648.0600 938.8000 ;
        RECT 1646.4600 954.6400 1648.0600 955.1200 ;
        RECT 1691.4600 954.6400 1693.0600 955.1200 ;
        RECT 1596.9000 970.9600 1599.9000 971.4400 ;
        RECT 1596.9000 965.5200 1599.9000 966.0000 ;
        RECT 1596.9000 960.0800 1599.9000 960.5600 ;
        RECT 1596.9000 949.2000 1599.9000 949.6800 ;
        RECT 1596.9000 943.7600 1599.9000 944.2400 ;
        RECT 1596.9000 938.3200 1599.9000 938.8000 ;
        RECT 1596.9000 932.8800 1599.9000 933.3600 ;
        RECT 1596.9000 954.6400 1599.9000 955.1200 ;
        RECT 1691.4600 916.5600 1693.0600 917.0400 ;
        RECT 1691.4600 922.0000 1693.0600 922.4800 ;
        RECT 1691.4600 900.2400 1693.0600 900.7200 ;
        RECT 1691.4600 905.6800 1693.0600 906.1600 ;
        RECT 1691.4600 911.1200 1693.0600 911.6000 ;
        RECT 1646.4600 916.5600 1648.0600 917.0400 ;
        RECT 1646.4600 922.0000 1648.0600 922.4800 ;
        RECT 1646.4600 900.2400 1648.0600 900.7200 ;
        RECT 1646.4600 905.6800 1648.0600 906.1600 ;
        RECT 1646.4600 911.1200 1648.0600 911.6000 ;
        RECT 1691.4600 889.3600 1693.0600 889.8400 ;
        RECT 1691.4600 894.8000 1693.0600 895.2800 ;
        RECT 1691.4600 873.0400 1693.0600 873.5200 ;
        RECT 1691.4600 878.4800 1693.0600 878.9600 ;
        RECT 1691.4600 883.9200 1693.0600 884.4000 ;
        RECT 1646.4600 889.3600 1648.0600 889.8400 ;
        RECT 1646.4600 894.8000 1648.0600 895.2800 ;
        RECT 1646.4600 873.0400 1648.0600 873.5200 ;
        RECT 1646.4600 878.4800 1648.0600 878.9600 ;
        RECT 1646.4600 883.9200 1648.0600 884.4000 ;
        RECT 1596.9000 916.5600 1599.9000 917.0400 ;
        RECT 1596.9000 922.0000 1599.9000 922.4800 ;
        RECT 1596.9000 905.6800 1599.9000 906.1600 ;
        RECT 1596.9000 900.2400 1599.9000 900.7200 ;
        RECT 1596.9000 911.1200 1599.9000 911.6000 ;
        RECT 1596.9000 889.3600 1599.9000 889.8400 ;
        RECT 1596.9000 894.8000 1599.9000 895.2800 ;
        RECT 1596.9000 878.4800 1599.9000 878.9600 ;
        RECT 1596.9000 873.0400 1599.9000 873.5200 ;
        RECT 1596.9000 883.9200 1599.9000 884.4000 ;
        RECT 1596.9000 927.4400 1599.9000 927.9200 ;
        RECT 1646.4600 927.4400 1648.0600 927.9200 ;
        RECT 1691.4600 927.4400 1693.0600 927.9200 ;
        RECT 1793.0000 862.1600 1796.0000 862.6400 ;
        RECT 1793.0000 867.6000 1796.0000 868.0800 ;
        RECT 1781.4600 862.1600 1783.0600 862.6400 ;
        RECT 1781.4600 867.6000 1783.0600 868.0800 ;
        RECT 1793.0000 845.8400 1796.0000 846.3200 ;
        RECT 1793.0000 851.2800 1796.0000 851.7600 ;
        RECT 1793.0000 856.7200 1796.0000 857.2000 ;
        RECT 1781.4600 845.8400 1783.0600 846.3200 ;
        RECT 1781.4600 851.2800 1783.0600 851.7600 ;
        RECT 1781.4600 856.7200 1783.0600 857.2000 ;
        RECT 1793.0000 834.9600 1796.0000 835.4400 ;
        RECT 1793.0000 840.4000 1796.0000 840.8800 ;
        RECT 1781.4600 834.9600 1783.0600 835.4400 ;
        RECT 1781.4600 840.4000 1783.0600 840.8800 ;
        RECT 1793.0000 818.6400 1796.0000 819.1200 ;
        RECT 1793.0000 824.0800 1796.0000 824.5600 ;
        RECT 1793.0000 829.5200 1796.0000 830.0000 ;
        RECT 1781.4600 818.6400 1783.0600 819.1200 ;
        RECT 1781.4600 824.0800 1783.0600 824.5600 ;
        RECT 1781.4600 829.5200 1783.0600 830.0000 ;
        RECT 1736.4600 862.1600 1738.0600 862.6400 ;
        RECT 1736.4600 867.6000 1738.0600 868.0800 ;
        RECT 1736.4600 845.8400 1738.0600 846.3200 ;
        RECT 1736.4600 851.2800 1738.0600 851.7600 ;
        RECT 1736.4600 856.7200 1738.0600 857.2000 ;
        RECT 1736.4600 834.9600 1738.0600 835.4400 ;
        RECT 1736.4600 840.4000 1738.0600 840.8800 ;
        RECT 1736.4600 818.6400 1738.0600 819.1200 ;
        RECT 1736.4600 824.0800 1738.0600 824.5600 ;
        RECT 1736.4600 829.5200 1738.0600 830.0000 ;
        RECT 1793.0000 807.7600 1796.0000 808.2400 ;
        RECT 1793.0000 813.2000 1796.0000 813.6800 ;
        RECT 1781.4600 807.7600 1783.0600 808.2400 ;
        RECT 1781.4600 813.2000 1783.0600 813.6800 ;
        RECT 1793.0000 791.4400 1796.0000 791.9200 ;
        RECT 1793.0000 796.8800 1796.0000 797.3600 ;
        RECT 1793.0000 802.3200 1796.0000 802.8000 ;
        RECT 1781.4600 791.4400 1783.0600 791.9200 ;
        RECT 1781.4600 796.8800 1783.0600 797.3600 ;
        RECT 1781.4600 802.3200 1783.0600 802.8000 ;
        RECT 1793.0000 780.5600 1796.0000 781.0400 ;
        RECT 1793.0000 786.0000 1796.0000 786.4800 ;
        RECT 1781.4600 780.5600 1783.0600 781.0400 ;
        RECT 1781.4600 786.0000 1783.0600 786.4800 ;
        RECT 1793.0000 775.1200 1796.0000 775.6000 ;
        RECT 1781.4600 775.1200 1783.0600 775.6000 ;
        RECT 1736.4600 807.7600 1738.0600 808.2400 ;
        RECT 1736.4600 813.2000 1738.0600 813.6800 ;
        RECT 1736.4600 791.4400 1738.0600 791.9200 ;
        RECT 1736.4600 796.8800 1738.0600 797.3600 ;
        RECT 1736.4600 802.3200 1738.0600 802.8000 ;
        RECT 1736.4600 780.5600 1738.0600 781.0400 ;
        RECT 1736.4600 786.0000 1738.0600 786.4800 ;
        RECT 1736.4600 775.1200 1738.0600 775.6000 ;
        RECT 1691.4600 862.1600 1693.0600 862.6400 ;
        RECT 1691.4600 867.6000 1693.0600 868.0800 ;
        RECT 1691.4600 845.8400 1693.0600 846.3200 ;
        RECT 1691.4600 851.2800 1693.0600 851.7600 ;
        RECT 1691.4600 856.7200 1693.0600 857.2000 ;
        RECT 1646.4600 862.1600 1648.0600 862.6400 ;
        RECT 1646.4600 867.6000 1648.0600 868.0800 ;
        RECT 1646.4600 845.8400 1648.0600 846.3200 ;
        RECT 1646.4600 851.2800 1648.0600 851.7600 ;
        RECT 1646.4600 856.7200 1648.0600 857.2000 ;
        RECT 1691.4600 834.9600 1693.0600 835.4400 ;
        RECT 1691.4600 840.4000 1693.0600 840.8800 ;
        RECT 1691.4600 818.6400 1693.0600 819.1200 ;
        RECT 1691.4600 824.0800 1693.0600 824.5600 ;
        RECT 1691.4600 829.5200 1693.0600 830.0000 ;
        RECT 1646.4600 834.9600 1648.0600 835.4400 ;
        RECT 1646.4600 840.4000 1648.0600 840.8800 ;
        RECT 1646.4600 818.6400 1648.0600 819.1200 ;
        RECT 1646.4600 824.0800 1648.0600 824.5600 ;
        RECT 1646.4600 829.5200 1648.0600 830.0000 ;
        RECT 1596.9000 862.1600 1599.9000 862.6400 ;
        RECT 1596.9000 867.6000 1599.9000 868.0800 ;
        RECT 1596.9000 851.2800 1599.9000 851.7600 ;
        RECT 1596.9000 845.8400 1599.9000 846.3200 ;
        RECT 1596.9000 856.7200 1599.9000 857.2000 ;
        RECT 1596.9000 834.9600 1599.9000 835.4400 ;
        RECT 1596.9000 840.4000 1599.9000 840.8800 ;
        RECT 1596.9000 824.0800 1599.9000 824.5600 ;
        RECT 1596.9000 818.6400 1599.9000 819.1200 ;
        RECT 1596.9000 829.5200 1599.9000 830.0000 ;
        RECT 1691.4600 807.7600 1693.0600 808.2400 ;
        RECT 1691.4600 813.2000 1693.0600 813.6800 ;
        RECT 1691.4600 791.4400 1693.0600 791.9200 ;
        RECT 1691.4600 796.8800 1693.0600 797.3600 ;
        RECT 1691.4600 802.3200 1693.0600 802.8000 ;
        RECT 1646.4600 807.7600 1648.0600 808.2400 ;
        RECT 1646.4600 813.2000 1648.0600 813.6800 ;
        RECT 1646.4600 791.4400 1648.0600 791.9200 ;
        RECT 1646.4600 796.8800 1648.0600 797.3600 ;
        RECT 1646.4600 802.3200 1648.0600 802.8000 ;
        RECT 1691.4600 786.0000 1693.0600 786.4800 ;
        RECT 1691.4600 780.5600 1693.0600 781.0400 ;
        RECT 1691.4600 775.1200 1693.0600 775.6000 ;
        RECT 1646.4600 786.0000 1648.0600 786.4800 ;
        RECT 1646.4600 780.5600 1648.0600 781.0400 ;
        RECT 1646.4600 775.1200 1648.0600 775.6000 ;
        RECT 1596.9000 807.7600 1599.9000 808.2400 ;
        RECT 1596.9000 813.2000 1599.9000 813.6800 ;
        RECT 1596.9000 796.8800 1599.9000 797.3600 ;
        RECT 1596.9000 791.4400 1599.9000 791.9200 ;
        RECT 1596.9000 802.3200 1599.9000 802.8000 ;
        RECT 1596.9000 780.5600 1599.9000 781.0400 ;
        RECT 1596.9000 786.0000 1599.9000 786.4800 ;
        RECT 1596.9000 775.1200 1599.9000 775.6000 ;
        RECT 1596.9000 973.3100 1796.0000 976.3100 ;
        RECT 1596.9000 768.2100 1796.0000 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1817.1200 2833.6100 1819.1200 2854.5400 ;
        RECT 2014.2200 2833.6100 2016.2200 2854.5400 ;
      LAYER met3 ;
        RECT 2014.2200 2850.0400 2016.2200 2850.5200 ;
        RECT 1817.1200 2850.0400 1819.1200 2850.5200 ;
        RECT 2014.2200 2839.1600 2016.2200 2839.6400 ;
        RECT 1817.1200 2839.1600 1819.1200 2839.6400 ;
        RECT 2014.2200 2844.6000 2016.2200 2845.0800 ;
        RECT 1817.1200 2844.6000 1819.1200 2845.0800 ;
        RECT 1817.1200 2852.5400 2016.2200 2854.5400 ;
        RECT 1817.1200 2833.6100 2016.2200 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1817.1200 79.2900 1819.1200 518.0800 ;
        RECT 2014.2200 79.2900 2016.2200 518.0800 ;
        RECT 1821.6800 79.2900 1823.2800 518.0800 ;
        RECT 1866.6800 79.2900 1868.2800 518.0800 ;
        RECT 1911.6800 79.2900 1913.2800 518.0800 ;
        RECT 1956.6800 79.2900 1958.2800 518.0800 ;
        RECT 2001.6800 79.2900 2003.2800 518.0800 ;
      LAYER met3 ;
        RECT 2014.2200 510.5200 2016.2200 511.0000 ;
        RECT 2014.2200 505.0800 2016.2200 505.5600 ;
        RECT 2014.2200 499.6400 2016.2200 500.1200 ;
        RECT 2014.2200 494.2000 2016.2200 494.6800 ;
        RECT 2014.2200 488.7600 2016.2200 489.2400 ;
        RECT 2014.2200 483.3200 2016.2200 483.8000 ;
        RECT 2014.2200 477.8800 2016.2200 478.3600 ;
        RECT 2014.2200 472.4400 2016.2200 472.9200 ;
        RECT 2014.2200 461.5600 2016.2200 462.0400 ;
        RECT 2014.2200 456.1200 2016.2200 456.6000 ;
        RECT 2014.2200 450.6800 2016.2200 451.1600 ;
        RECT 2014.2200 445.2400 2016.2200 445.7200 ;
        RECT 2014.2200 439.8000 2016.2200 440.2800 ;
        RECT 2014.2200 434.3600 2016.2200 434.8400 ;
        RECT 2014.2200 428.9200 2016.2200 429.4000 ;
        RECT 2014.2200 423.4800 2016.2200 423.9600 ;
        RECT 2014.2200 418.0400 2016.2200 418.5200 ;
        RECT 2014.2200 412.6000 2016.2200 413.0800 ;
        RECT 2014.2200 467.0000 2016.2200 467.4800 ;
        RECT 2014.2200 407.1600 2016.2200 407.6400 ;
        RECT 2014.2200 401.7200 2016.2200 402.2000 ;
        RECT 2014.2200 396.2800 2016.2200 396.7600 ;
        RECT 2014.2200 390.8400 2016.2200 391.3200 ;
        RECT 2014.2200 385.4000 2016.2200 385.8800 ;
        RECT 2014.2200 379.9600 2016.2200 380.4400 ;
        RECT 2014.2200 374.5200 2016.2200 375.0000 ;
        RECT 2014.2200 369.0800 2016.2200 369.5600 ;
        RECT 2014.2200 363.6400 2016.2200 364.1200 ;
        RECT 2014.2200 358.2000 2016.2200 358.6800 ;
        RECT 2014.2200 352.7600 2016.2200 353.2400 ;
        RECT 2014.2200 347.3200 2016.2200 347.8000 ;
        RECT 2014.2200 341.8800 2016.2200 342.3600 ;
        RECT 2014.2200 336.4400 2016.2200 336.9200 ;
        RECT 2014.2200 331.0000 2016.2200 331.4800 ;
        RECT 2014.2200 325.5600 2016.2200 326.0400 ;
        RECT 2014.2200 320.1200 2016.2200 320.6000 ;
        RECT 2014.2200 314.6800 2016.2200 315.1600 ;
        RECT 2014.2200 309.2400 2016.2200 309.7200 ;
        RECT 2014.2200 303.8000 2016.2200 304.2800 ;
        RECT 1817.1200 510.5200 1819.1200 511.0000 ;
        RECT 1817.1200 505.0800 1819.1200 505.5600 ;
        RECT 1817.1200 499.6400 1819.1200 500.1200 ;
        RECT 1817.1200 494.2000 1819.1200 494.6800 ;
        RECT 1817.1200 488.7600 1819.1200 489.2400 ;
        RECT 1817.1200 483.3200 1819.1200 483.8000 ;
        RECT 1817.1200 477.8800 1819.1200 478.3600 ;
        RECT 1817.1200 472.4400 1819.1200 472.9200 ;
        RECT 1817.1200 461.5600 1819.1200 462.0400 ;
        RECT 1817.1200 456.1200 1819.1200 456.6000 ;
        RECT 1817.1200 450.6800 1819.1200 451.1600 ;
        RECT 1817.1200 445.2400 1819.1200 445.7200 ;
        RECT 1817.1200 439.8000 1819.1200 440.2800 ;
        RECT 1817.1200 434.3600 1819.1200 434.8400 ;
        RECT 1817.1200 428.9200 1819.1200 429.4000 ;
        RECT 1817.1200 423.4800 1819.1200 423.9600 ;
        RECT 1817.1200 418.0400 1819.1200 418.5200 ;
        RECT 1817.1200 412.6000 1819.1200 413.0800 ;
        RECT 1817.1200 467.0000 1819.1200 467.4800 ;
        RECT 1817.1200 407.1600 1819.1200 407.6400 ;
        RECT 1817.1200 401.7200 1819.1200 402.2000 ;
        RECT 1817.1200 396.2800 1819.1200 396.7600 ;
        RECT 1817.1200 390.8400 1819.1200 391.3200 ;
        RECT 1817.1200 385.4000 1819.1200 385.8800 ;
        RECT 1817.1200 379.9600 1819.1200 380.4400 ;
        RECT 1817.1200 374.5200 1819.1200 375.0000 ;
        RECT 1817.1200 369.0800 1819.1200 369.5600 ;
        RECT 1817.1200 363.6400 1819.1200 364.1200 ;
        RECT 1817.1200 358.2000 1819.1200 358.6800 ;
        RECT 1817.1200 352.7600 1819.1200 353.2400 ;
        RECT 1817.1200 347.3200 1819.1200 347.8000 ;
        RECT 1817.1200 341.8800 1819.1200 342.3600 ;
        RECT 1817.1200 336.4400 1819.1200 336.9200 ;
        RECT 1817.1200 331.0000 1819.1200 331.4800 ;
        RECT 1817.1200 325.5600 1819.1200 326.0400 ;
        RECT 1817.1200 320.1200 1819.1200 320.6000 ;
        RECT 1817.1200 314.6800 1819.1200 315.1600 ;
        RECT 1817.1200 309.2400 1819.1200 309.7200 ;
        RECT 1817.1200 303.8000 1819.1200 304.2800 ;
        RECT 2014.2200 292.9200 2016.2200 293.4000 ;
        RECT 2014.2200 287.4800 2016.2200 287.9600 ;
        RECT 2014.2200 282.0400 2016.2200 282.5200 ;
        RECT 2014.2200 276.6000 2016.2200 277.0800 ;
        RECT 2014.2200 271.1600 2016.2200 271.6400 ;
        RECT 2014.2200 265.7200 2016.2200 266.2000 ;
        RECT 2014.2200 260.2800 2016.2200 260.7600 ;
        RECT 2014.2200 254.8400 2016.2200 255.3200 ;
        RECT 2014.2200 249.4000 2016.2200 249.8800 ;
        RECT 2014.2200 243.9600 2016.2200 244.4400 ;
        RECT 2014.2200 238.5200 2016.2200 239.0000 ;
        RECT 2014.2200 233.0800 2016.2200 233.5600 ;
        RECT 2014.2200 227.6400 2016.2200 228.1200 ;
        RECT 2014.2200 222.2000 2016.2200 222.6800 ;
        RECT 2014.2200 216.7600 2016.2200 217.2400 ;
        RECT 2014.2200 211.3200 2016.2200 211.8000 ;
        RECT 2014.2200 205.8800 2016.2200 206.3600 ;
        RECT 2014.2200 200.4400 2016.2200 200.9200 ;
        RECT 2014.2200 195.0000 2016.2200 195.4800 ;
        RECT 2014.2200 189.5600 2016.2200 190.0400 ;
        RECT 2014.2200 184.1200 2016.2200 184.6000 ;
        RECT 2014.2200 178.6800 2016.2200 179.1600 ;
        RECT 2014.2200 173.2400 2016.2200 173.7200 ;
        RECT 2014.2200 167.8000 2016.2200 168.2800 ;
        RECT 2014.2200 162.3600 2016.2200 162.8400 ;
        RECT 2014.2200 156.9200 2016.2200 157.4000 ;
        RECT 2014.2200 151.4800 2016.2200 151.9600 ;
        RECT 2014.2200 146.0400 2016.2200 146.5200 ;
        RECT 2014.2200 140.6000 2016.2200 141.0800 ;
        RECT 2014.2200 135.1600 2016.2200 135.6400 ;
        RECT 2014.2200 124.2800 2016.2200 124.7600 ;
        RECT 2014.2200 118.8400 2016.2200 119.3200 ;
        RECT 2014.2200 113.4000 2016.2200 113.8800 ;
        RECT 2014.2200 107.9600 2016.2200 108.4400 ;
        RECT 2014.2200 102.5200 2016.2200 103.0000 ;
        RECT 2014.2200 97.0800 2016.2200 97.5600 ;
        RECT 2014.2200 91.6400 2016.2200 92.1200 ;
        RECT 2014.2200 86.2000 2016.2200 86.6800 ;
        RECT 2014.2200 129.7200 2016.2200 130.2000 ;
        RECT 1817.1200 292.9200 1819.1200 293.4000 ;
        RECT 1817.1200 287.4800 1819.1200 287.9600 ;
        RECT 1817.1200 282.0400 1819.1200 282.5200 ;
        RECT 1817.1200 276.6000 1819.1200 277.0800 ;
        RECT 1817.1200 271.1600 1819.1200 271.6400 ;
        RECT 1817.1200 265.7200 1819.1200 266.2000 ;
        RECT 1817.1200 260.2800 1819.1200 260.7600 ;
        RECT 1817.1200 254.8400 1819.1200 255.3200 ;
        RECT 1817.1200 249.4000 1819.1200 249.8800 ;
        RECT 1817.1200 243.9600 1819.1200 244.4400 ;
        RECT 1817.1200 238.5200 1819.1200 239.0000 ;
        RECT 1817.1200 233.0800 1819.1200 233.5600 ;
        RECT 1817.1200 227.6400 1819.1200 228.1200 ;
        RECT 1817.1200 222.2000 1819.1200 222.6800 ;
        RECT 1817.1200 216.7600 1819.1200 217.2400 ;
        RECT 1817.1200 211.3200 1819.1200 211.8000 ;
        RECT 1817.1200 205.8800 1819.1200 206.3600 ;
        RECT 1817.1200 200.4400 1819.1200 200.9200 ;
        RECT 1817.1200 195.0000 1819.1200 195.4800 ;
        RECT 1817.1200 189.5600 1819.1200 190.0400 ;
        RECT 1817.1200 184.1200 1819.1200 184.6000 ;
        RECT 1817.1200 178.6800 1819.1200 179.1600 ;
        RECT 1817.1200 173.2400 1819.1200 173.7200 ;
        RECT 1817.1200 167.8000 1819.1200 168.2800 ;
        RECT 1817.1200 162.3600 1819.1200 162.8400 ;
        RECT 1817.1200 156.9200 1819.1200 157.4000 ;
        RECT 1817.1200 151.4800 1819.1200 151.9600 ;
        RECT 1817.1200 146.0400 1819.1200 146.5200 ;
        RECT 1817.1200 140.6000 1819.1200 141.0800 ;
        RECT 1817.1200 135.1600 1819.1200 135.6400 ;
        RECT 1817.1200 124.2800 1819.1200 124.7600 ;
        RECT 1817.1200 118.8400 1819.1200 119.3200 ;
        RECT 1817.1200 113.4000 1819.1200 113.8800 ;
        RECT 1817.1200 107.9600 1819.1200 108.4400 ;
        RECT 1817.1200 102.5200 1819.1200 103.0000 ;
        RECT 1817.1200 97.0800 1819.1200 97.5600 ;
        RECT 1817.1200 91.6400 1819.1200 92.1200 ;
        RECT 1817.1200 86.2000 1819.1200 86.6800 ;
        RECT 1817.1200 129.7200 1819.1200 130.2000 ;
        RECT 2014.2200 298.3600 2016.2200 298.8400 ;
        RECT 1817.1200 298.3600 1819.1200 298.8400 ;
        RECT 1817.1200 516.0800 2016.2200 518.0800 ;
        RECT 1817.1200 79.2900 2016.2200 81.2900 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'S_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1817.1200 37.6700 1819.1200 58.6000 ;
        RECT 2014.2200 37.6700 2016.2200 58.6000 ;
      LAYER met3 ;
        RECT 2014.2200 54.1000 2016.2200 54.5800 ;
        RECT 1817.1200 54.1000 1819.1200 54.5800 ;
        RECT 2014.2200 43.2200 2016.2200 43.7000 ;
        RECT 1817.1200 43.2200 1819.1200 43.7000 ;
        RECT 2014.2200 48.6600 2016.2200 49.1400 ;
        RECT 1817.1200 48.6600 1819.1200 49.1400 ;
        RECT 1817.1200 56.6000 2016.2200 58.6000 ;
        RECT 1817.1200 37.6700 2016.2200 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1817.1200 2375.6900 1819.1200 2814.4800 ;
        RECT 2014.2200 2375.6900 2016.2200 2814.4800 ;
        RECT 1821.6800 2375.6900 1823.2800 2814.4800 ;
        RECT 1866.6800 2375.6900 1868.2800 2814.4800 ;
        RECT 1911.6800 2375.6900 1913.2800 2814.4800 ;
        RECT 1956.6800 2375.6900 1958.2800 2814.4800 ;
        RECT 2001.6800 2375.6900 2003.2800 2814.4800 ;
      LAYER met3 ;
        RECT 2014.2200 2806.9200 2016.2200 2807.4000 ;
        RECT 2014.2200 2801.4800 2016.2200 2801.9600 ;
        RECT 2014.2200 2796.0400 2016.2200 2796.5200 ;
        RECT 2014.2200 2790.6000 2016.2200 2791.0800 ;
        RECT 2014.2200 2785.1600 2016.2200 2785.6400 ;
        RECT 2014.2200 2779.7200 2016.2200 2780.2000 ;
        RECT 2014.2200 2774.2800 2016.2200 2774.7600 ;
        RECT 2014.2200 2768.8400 2016.2200 2769.3200 ;
        RECT 2014.2200 2757.9600 2016.2200 2758.4400 ;
        RECT 2014.2200 2752.5200 2016.2200 2753.0000 ;
        RECT 2014.2200 2747.0800 2016.2200 2747.5600 ;
        RECT 2014.2200 2741.6400 2016.2200 2742.1200 ;
        RECT 2014.2200 2736.2000 2016.2200 2736.6800 ;
        RECT 2014.2200 2730.7600 2016.2200 2731.2400 ;
        RECT 2014.2200 2725.3200 2016.2200 2725.8000 ;
        RECT 2014.2200 2719.8800 2016.2200 2720.3600 ;
        RECT 2014.2200 2714.4400 2016.2200 2714.9200 ;
        RECT 2014.2200 2709.0000 2016.2200 2709.4800 ;
        RECT 2014.2200 2763.4000 2016.2200 2763.8800 ;
        RECT 2014.2200 2703.5600 2016.2200 2704.0400 ;
        RECT 2014.2200 2698.1200 2016.2200 2698.6000 ;
        RECT 2014.2200 2692.6800 2016.2200 2693.1600 ;
        RECT 2014.2200 2687.2400 2016.2200 2687.7200 ;
        RECT 2014.2200 2681.8000 2016.2200 2682.2800 ;
        RECT 2014.2200 2676.3600 2016.2200 2676.8400 ;
        RECT 2014.2200 2670.9200 2016.2200 2671.4000 ;
        RECT 2014.2200 2665.4800 2016.2200 2665.9600 ;
        RECT 2014.2200 2660.0400 2016.2200 2660.5200 ;
        RECT 2014.2200 2654.6000 2016.2200 2655.0800 ;
        RECT 2014.2200 2649.1600 2016.2200 2649.6400 ;
        RECT 2014.2200 2643.7200 2016.2200 2644.2000 ;
        RECT 2014.2200 2638.2800 2016.2200 2638.7600 ;
        RECT 2014.2200 2632.8400 2016.2200 2633.3200 ;
        RECT 2014.2200 2627.4000 2016.2200 2627.8800 ;
        RECT 2014.2200 2621.9600 2016.2200 2622.4400 ;
        RECT 2014.2200 2616.5200 2016.2200 2617.0000 ;
        RECT 2014.2200 2611.0800 2016.2200 2611.5600 ;
        RECT 2014.2200 2605.6400 2016.2200 2606.1200 ;
        RECT 2014.2200 2600.2000 2016.2200 2600.6800 ;
        RECT 1817.1200 2806.9200 1819.1200 2807.4000 ;
        RECT 1817.1200 2801.4800 1819.1200 2801.9600 ;
        RECT 1817.1200 2796.0400 1819.1200 2796.5200 ;
        RECT 1817.1200 2790.6000 1819.1200 2791.0800 ;
        RECT 1817.1200 2785.1600 1819.1200 2785.6400 ;
        RECT 1817.1200 2779.7200 1819.1200 2780.2000 ;
        RECT 1817.1200 2774.2800 1819.1200 2774.7600 ;
        RECT 1817.1200 2768.8400 1819.1200 2769.3200 ;
        RECT 1817.1200 2757.9600 1819.1200 2758.4400 ;
        RECT 1817.1200 2752.5200 1819.1200 2753.0000 ;
        RECT 1817.1200 2747.0800 1819.1200 2747.5600 ;
        RECT 1817.1200 2741.6400 1819.1200 2742.1200 ;
        RECT 1817.1200 2736.2000 1819.1200 2736.6800 ;
        RECT 1817.1200 2730.7600 1819.1200 2731.2400 ;
        RECT 1817.1200 2725.3200 1819.1200 2725.8000 ;
        RECT 1817.1200 2719.8800 1819.1200 2720.3600 ;
        RECT 1817.1200 2714.4400 1819.1200 2714.9200 ;
        RECT 1817.1200 2709.0000 1819.1200 2709.4800 ;
        RECT 1817.1200 2763.4000 1819.1200 2763.8800 ;
        RECT 1817.1200 2703.5600 1819.1200 2704.0400 ;
        RECT 1817.1200 2698.1200 1819.1200 2698.6000 ;
        RECT 1817.1200 2692.6800 1819.1200 2693.1600 ;
        RECT 1817.1200 2687.2400 1819.1200 2687.7200 ;
        RECT 1817.1200 2681.8000 1819.1200 2682.2800 ;
        RECT 1817.1200 2676.3600 1819.1200 2676.8400 ;
        RECT 1817.1200 2670.9200 1819.1200 2671.4000 ;
        RECT 1817.1200 2665.4800 1819.1200 2665.9600 ;
        RECT 1817.1200 2660.0400 1819.1200 2660.5200 ;
        RECT 1817.1200 2654.6000 1819.1200 2655.0800 ;
        RECT 1817.1200 2649.1600 1819.1200 2649.6400 ;
        RECT 1817.1200 2643.7200 1819.1200 2644.2000 ;
        RECT 1817.1200 2638.2800 1819.1200 2638.7600 ;
        RECT 1817.1200 2632.8400 1819.1200 2633.3200 ;
        RECT 1817.1200 2627.4000 1819.1200 2627.8800 ;
        RECT 1817.1200 2621.9600 1819.1200 2622.4400 ;
        RECT 1817.1200 2616.5200 1819.1200 2617.0000 ;
        RECT 1817.1200 2611.0800 1819.1200 2611.5600 ;
        RECT 1817.1200 2605.6400 1819.1200 2606.1200 ;
        RECT 1817.1200 2600.2000 1819.1200 2600.6800 ;
        RECT 2014.2200 2589.3200 2016.2200 2589.8000 ;
        RECT 2014.2200 2583.8800 2016.2200 2584.3600 ;
        RECT 2014.2200 2578.4400 2016.2200 2578.9200 ;
        RECT 2014.2200 2573.0000 2016.2200 2573.4800 ;
        RECT 2014.2200 2567.5600 2016.2200 2568.0400 ;
        RECT 2014.2200 2562.1200 2016.2200 2562.6000 ;
        RECT 2014.2200 2556.6800 2016.2200 2557.1600 ;
        RECT 2014.2200 2551.2400 2016.2200 2551.7200 ;
        RECT 2014.2200 2545.8000 2016.2200 2546.2800 ;
        RECT 2014.2200 2540.3600 2016.2200 2540.8400 ;
        RECT 2014.2200 2534.9200 2016.2200 2535.4000 ;
        RECT 2014.2200 2529.4800 2016.2200 2529.9600 ;
        RECT 2014.2200 2524.0400 2016.2200 2524.5200 ;
        RECT 2014.2200 2518.6000 2016.2200 2519.0800 ;
        RECT 2014.2200 2513.1600 2016.2200 2513.6400 ;
        RECT 2014.2200 2507.7200 2016.2200 2508.2000 ;
        RECT 2014.2200 2502.2800 2016.2200 2502.7600 ;
        RECT 2014.2200 2496.8400 2016.2200 2497.3200 ;
        RECT 2014.2200 2491.4000 2016.2200 2491.8800 ;
        RECT 2014.2200 2485.9600 2016.2200 2486.4400 ;
        RECT 2014.2200 2480.5200 2016.2200 2481.0000 ;
        RECT 2014.2200 2475.0800 2016.2200 2475.5600 ;
        RECT 2014.2200 2469.6400 2016.2200 2470.1200 ;
        RECT 2014.2200 2464.2000 2016.2200 2464.6800 ;
        RECT 2014.2200 2458.7600 2016.2200 2459.2400 ;
        RECT 2014.2200 2453.3200 2016.2200 2453.8000 ;
        RECT 2014.2200 2447.8800 2016.2200 2448.3600 ;
        RECT 2014.2200 2442.4400 2016.2200 2442.9200 ;
        RECT 2014.2200 2437.0000 2016.2200 2437.4800 ;
        RECT 2014.2200 2431.5600 2016.2200 2432.0400 ;
        RECT 2014.2200 2420.6800 2016.2200 2421.1600 ;
        RECT 2014.2200 2415.2400 2016.2200 2415.7200 ;
        RECT 2014.2200 2409.8000 2016.2200 2410.2800 ;
        RECT 2014.2200 2404.3600 2016.2200 2404.8400 ;
        RECT 2014.2200 2398.9200 2016.2200 2399.4000 ;
        RECT 2014.2200 2393.4800 2016.2200 2393.9600 ;
        RECT 2014.2200 2388.0400 2016.2200 2388.5200 ;
        RECT 2014.2200 2382.6000 2016.2200 2383.0800 ;
        RECT 2014.2200 2426.1200 2016.2200 2426.6000 ;
        RECT 1817.1200 2589.3200 1819.1200 2589.8000 ;
        RECT 1817.1200 2583.8800 1819.1200 2584.3600 ;
        RECT 1817.1200 2578.4400 1819.1200 2578.9200 ;
        RECT 1817.1200 2573.0000 1819.1200 2573.4800 ;
        RECT 1817.1200 2567.5600 1819.1200 2568.0400 ;
        RECT 1817.1200 2562.1200 1819.1200 2562.6000 ;
        RECT 1817.1200 2556.6800 1819.1200 2557.1600 ;
        RECT 1817.1200 2551.2400 1819.1200 2551.7200 ;
        RECT 1817.1200 2545.8000 1819.1200 2546.2800 ;
        RECT 1817.1200 2540.3600 1819.1200 2540.8400 ;
        RECT 1817.1200 2534.9200 1819.1200 2535.4000 ;
        RECT 1817.1200 2529.4800 1819.1200 2529.9600 ;
        RECT 1817.1200 2524.0400 1819.1200 2524.5200 ;
        RECT 1817.1200 2518.6000 1819.1200 2519.0800 ;
        RECT 1817.1200 2513.1600 1819.1200 2513.6400 ;
        RECT 1817.1200 2507.7200 1819.1200 2508.2000 ;
        RECT 1817.1200 2502.2800 1819.1200 2502.7600 ;
        RECT 1817.1200 2496.8400 1819.1200 2497.3200 ;
        RECT 1817.1200 2491.4000 1819.1200 2491.8800 ;
        RECT 1817.1200 2485.9600 1819.1200 2486.4400 ;
        RECT 1817.1200 2480.5200 1819.1200 2481.0000 ;
        RECT 1817.1200 2475.0800 1819.1200 2475.5600 ;
        RECT 1817.1200 2469.6400 1819.1200 2470.1200 ;
        RECT 1817.1200 2464.2000 1819.1200 2464.6800 ;
        RECT 1817.1200 2458.7600 1819.1200 2459.2400 ;
        RECT 1817.1200 2453.3200 1819.1200 2453.8000 ;
        RECT 1817.1200 2447.8800 1819.1200 2448.3600 ;
        RECT 1817.1200 2442.4400 1819.1200 2442.9200 ;
        RECT 1817.1200 2437.0000 1819.1200 2437.4800 ;
        RECT 1817.1200 2431.5600 1819.1200 2432.0400 ;
        RECT 1817.1200 2420.6800 1819.1200 2421.1600 ;
        RECT 1817.1200 2415.2400 1819.1200 2415.7200 ;
        RECT 1817.1200 2409.8000 1819.1200 2410.2800 ;
        RECT 1817.1200 2404.3600 1819.1200 2404.8400 ;
        RECT 1817.1200 2398.9200 1819.1200 2399.4000 ;
        RECT 1817.1200 2393.4800 1819.1200 2393.9600 ;
        RECT 1817.1200 2388.0400 1819.1200 2388.5200 ;
        RECT 1817.1200 2382.6000 1819.1200 2383.0800 ;
        RECT 1817.1200 2426.1200 1819.1200 2426.6000 ;
        RECT 2014.2200 2594.7600 2016.2200 2595.2400 ;
        RECT 1817.1200 2594.7600 1819.1200 2595.2400 ;
        RECT 1817.1200 2812.4800 2016.2200 2814.4800 ;
        RECT 1817.1200 2375.6900 2016.2200 2377.6900 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1817.1200 1916.4100 1819.1200 2355.2000 ;
        RECT 2014.2200 1916.4100 2016.2200 2355.2000 ;
        RECT 1821.6800 1916.4100 1823.2800 2355.2000 ;
        RECT 1866.6800 1916.4100 1868.2800 2355.2000 ;
        RECT 1911.6800 1916.4100 1913.2800 2355.2000 ;
        RECT 1956.6800 1916.4100 1958.2800 2355.2000 ;
        RECT 2001.6800 1916.4100 2003.2800 2355.2000 ;
      LAYER met3 ;
        RECT 2014.2200 2347.6400 2016.2200 2348.1200 ;
        RECT 2014.2200 2342.2000 2016.2200 2342.6800 ;
        RECT 2014.2200 2336.7600 2016.2200 2337.2400 ;
        RECT 2014.2200 2331.3200 2016.2200 2331.8000 ;
        RECT 2014.2200 2325.8800 2016.2200 2326.3600 ;
        RECT 2014.2200 2320.4400 2016.2200 2320.9200 ;
        RECT 2014.2200 2315.0000 2016.2200 2315.4800 ;
        RECT 2014.2200 2309.5600 2016.2200 2310.0400 ;
        RECT 2014.2200 2298.6800 2016.2200 2299.1600 ;
        RECT 2014.2200 2293.2400 2016.2200 2293.7200 ;
        RECT 2014.2200 2287.8000 2016.2200 2288.2800 ;
        RECT 2014.2200 2282.3600 2016.2200 2282.8400 ;
        RECT 2014.2200 2276.9200 2016.2200 2277.4000 ;
        RECT 2014.2200 2271.4800 2016.2200 2271.9600 ;
        RECT 2014.2200 2266.0400 2016.2200 2266.5200 ;
        RECT 2014.2200 2260.6000 2016.2200 2261.0800 ;
        RECT 2014.2200 2255.1600 2016.2200 2255.6400 ;
        RECT 2014.2200 2249.7200 2016.2200 2250.2000 ;
        RECT 2014.2200 2304.1200 2016.2200 2304.6000 ;
        RECT 2014.2200 2244.2800 2016.2200 2244.7600 ;
        RECT 2014.2200 2238.8400 2016.2200 2239.3200 ;
        RECT 2014.2200 2233.4000 2016.2200 2233.8800 ;
        RECT 2014.2200 2227.9600 2016.2200 2228.4400 ;
        RECT 2014.2200 2222.5200 2016.2200 2223.0000 ;
        RECT 2014.2200 2217.0800 2016.2200 2217.5600 ;
        RECT 2014.2200 2211.6400 2016.2200 2212.1200 ;
        RECT 2014.2200 2206.2000 2016.2200 2206.6800 ;
        RECT 2014.2200 2200.7600 2016.2200 2201.2400 ;
        RECT 2014.2200 2195.3200 2016.2200 2195.8000 ;
        RECT 2014.2200 2189.8800 2016.2200 2190.3600 ;
        RECT 2014.2200 2184.4400 2016.2200 2184.9200 ;
        RECT 2014.2200 2179.0000 2016.2200 2179.4800 ;
        RECT 2014.2200 2173.5600 2016.2200 2174.0400 ;
        RECT 2014.2200 2168.1200 2016.2200 2168.6000 ;
        RECT 2014.2200 2162.6800 2016.2200 2163.1600 ;
        RECT 2014.2200 2157.2400 2016.2200 2157.7200 ;
        RECT 2014.2200 2151.8000 2016.2200 2152.2800 ;
        RECT 2014.2200 2146.3600 2016.2200 2146.8400 ;
        RECT 2014.2200 2140.9200 2016.2200 2141.4000 ;
        RECT 1817.1200 2347.6400 1819.1200 2348.1200 ;
        RECT 1817.1200 2342.2000 1819.1200 2342.6800 ;
        RECT 1817.1200 2336.7600 1819.1200 2337.2400 ;
        RECT 1817.1200 2331.3200 1819.1200 2331.8000 ;
        RECT 1817.1200 2325.8800 1819.1200 2326.3600 ;
        RECT 1817.1200 2320.4400 1819.1200 2320.9200 ;
        RECT 1817.1200 2315.0000 1819.1200 2315.4800 ;
        RECT 1817.1200 2309.5600 1819.1200 2310.0400 ;
        RECT 1817.1200 2298.6800 1819.1200 2299.1600 ;
        RECT 1817.1200 2293.2400 1819.1200 2293.7200 ;
        RECT 1817.1200 2287.8000 1819.1200 2288.2800 ;
        RECT 1817.1200 2282.3600 1819.1200 2282.8400 ;
        RECT 1817.1200 2276.9200 1819.1200 2277.4000 ;
        RECT 1817.1200 2271.4800 1819.1200 2271.9600 ;
        RECT 1817.1200 2266.0400 1819.1200 2266.5200 ;
        RECT 1817.1200 2260.6000 1819.1200 2261.0800 ;
        RECT 1817.1200 2255.1600 1819.1200 2255.6400 ;
        RECT 1817.1200 2249.7200 1819.1200 2250.2000 ;
        RECT 1817.1200 2304.1200 1819.1200 2304.6000 ;
        RECT 1817.1200 2244.2800 1819.1200 2244.7600 ;
        RECT 1817.1200 2238.8400 1819.1200 2239.3200 ;
        RECT 1817.1200 2233.4000 1819.1200 2233.8800 ;
        RECT 1817.1200 2227.9600 1819.1200 2228.4400 ;
        RECT 1817.1200 2222.5200 1819.1200 2223.0000 ;
        RECT 1817.1200 2217.0800 1819.1200 2217.5600 ;
        RECT 1817.1200 2211.6400 1819.1200 2212.1200 ;
        RECT 1817.1200 2206.2000 1819.1200 2206.6800 ;
        RECT 1817.1200 2200.7600 1819.1200 2201.2400 ;
        RECT 1817.1200 2195.3200 1819.1200 2195.8000 ;
        RECT 1817.1200 2189.8800 1819.1200 2190.3600 ;
        RECT 1817.1200 2184.4400 1819.1200 2184.9200 ;
        RECT 1817.1200 2179.0000 1819.1200 2179.4800 ;
        RECT 1817.1200 2173.5600 1819.1200 2174.0400 ;
        RECT 1817.1200 2168.1200 1819.1200 2168.6000 ;
        RECT 1817.1200 2162.6800 1819.1200 2163.1600 ;
        RECT 1817.1200 2157.2400 1819.1200 2157.7200 ;
        RECT 1817.1200 2151.8000 1819.1200 2152.2800 ;
        RECT 1817.1200 2146.3600 1819.1200 2146.8400 ;
        RECT 1817.1200 2140.9200 1819.1200 2141.4000 ;
        RECT 2014.2200 2130.0400 2016.2200 2130.5200 ;
        RECT 2014.2200 2124.6000 2016.2200 2125.0800 ;
        RECT 2014.2200 2119.1600 2016.2200 2119.6400 ;
        RECT 2014.2200 2113.7200 2016.2200 2114.2000 ;
        RECT 2014.2200 2108.2800 2016.2200 2108.7600 ;
        RECT 2014.2200 2102.8400 2016.2200 2103.3200 ;
        RECT 2014.2200 2097.4000 2016.2200 2097.8800 ;
        RECT 2014.2200 2091.9600 2016.2200 2092.4400 ;
        RECT 2014.2200 2086.5200 2016.2200 2087.0000 ;
        RECT 2014.2200 2081.0800 2016.2200 2081.5600 ;
        RECT 2014.2200 2075.6400 2016.2200 2076.1200 ;
        RECT 2014.2200 2070.2000 2016.2200 2070.6800 ;
        RECT 2014.2200 2064.7600 2016.2200 2065.2400 ;
        RECT 2014.2200 2059.3200 2016.2200 2059.8000 ;
        RECT 2014.2200 2053.8800 2016.2200 2054.3600 ;
        RECT 2014.2200 2048.4400 2016.2200 2048.9200 ;
        RECT 2014.2200 2043.0000 2016.2200 2043.4800 ;
        RECT 2014.2200 2037.5600 2016.2200 2038.0400 ;
        RECT 2014.2200 2032.1200 2016.2200 2032.6000 ;
        RECT 2014.2200 2026.6800 2016.2200 2027.1600 ;
        RECT 2014.2200 2021.2400 2016.2200 2021.7200 ;
        RECT 2014.2200 2015.8000 2016.2200 2016.2800 ;
        RECT 2014.2200 2010.3600 2016.2200 2010.8400 ;
        RECT 2014.2200 2004.9200 2016.2200 2005.4000 ;
        RECT 2014.2200 1999.4800 2016.2200 1999.9600 ;
        RECT 2014.2200 1994.0400 2016.2200 1994.5200 ;
        RECT 2014.2200 1988.6000 2016.2200 1989.0800 ;
        RECT 2014.2200 1983.1600 2016.2200 1983.6400 ;
        RECT 2014.2200 1977.7200 2016.2200 1978.2000 ;
        RECT 2014.2200 1972.2800 2016.2200 1972.7600 ;
        RECT 2014.2200 1961.4000 2016.2200 1961.8800 ;
        RECT 2014.2200 1955.9600 2016.2200 1956.4400 ;
        RECT 2014.2200 1950.5200 2016.2200 1951.0000 ;
        RECT 2014.2200 1945.0800 2016.2200 1945.5600 ;
        RECT 2014.2200 1939.6400 2016.2200 1940.1200 ;
        RECT 2014.2200 1934.2000 2016.2200 1934.6800 ;
        RECT 2014.2200 1928.7600 2016.2200 1929.2400 ;
        RECT 2014.2200 1923.3200 2016.2200 1923.8000 ;
        RECT 2014.2200 1966.8400 2016.2200 1967.3200 ;
        RECT 1817.1200 2130.0400 1819.1200 2130.5200 ;
        RECT 1817.1200 2124.6000 1819.1200 2125.0800 ;
        RECT 1817.1200 2119.1600 1819.1200 2119.6400 ;
        RECT 1817.1200 2113.7200 1819.1200 2114.2000 ;
        RECT 1817.1200 2108.2800 1819.1200 2108.7600 ;
        RECT 1817.1200 2102.8400 1819.1200 2103.3200 ;
        RECT 1817.1200 2097.4000 1819.1200 2097.8800 ;
        RECT 1817.1200 2091.9600 1819.1200 2092.4400 ;
        RECT 1817.1200 2086.5200 1819.1200 2087.0000 ;
        RECT 1817.1200 2081.0800 1819.1200 2081.5600 ;
        RECT 1817.1200 2075.6400 1819.1200 2076.1200 ;
        RECT 1817.1200 2070.2000 1819.1200 2070.6800 ;
        RECT 1817.1200 2064.7600 1819.1200 2065.2400 ;
        RECT 1817.1200 2059.3200 1819.1200 2059.8000 ;
        RECT 1817.1200 2053.8800 1819.1200 2054.3600 ;
        RECT 1817.1200 2048.4400 1819.1200 2048.9200 ;
        RECT 1817.1200 2043.0000 1819.1200 2043.4800 ;
        RECT 1817.1200 2037.5600 1819.1200 2038.0400 ;
        RECT 1817.1200 2032.1200 1819.1200 2032.6000 ;
        RECT 1817.1200 2026.6800 1819.1200 2027.1600 ;
        RECT 1817.1200 2021.2400 1819.1200 2021.7200 ;
        RECT 1817.1200 2015.8000 1819.1200 2016.2800 ;
        RECT 1817.1200 2010.3600 1819.1200 2010.8400 ;
        RECT 1817.1200 2004.9200 1819.1200 2005.4000 ;
        RECT 1817.1200 1999.4800 1819.1200 1999.9600 ;
        RECT 1817.1200 1994.0400 1819.1200 1994.5200 ;
        RECT 1817.1200 1988.6000 1819.1200 1989.0800 ;
        RECT 1817.1200 1983.1600 1819.1200 1983.6400 ;
        RECT 1817.1200 1977.7200 1819.1200 1978.2000 ;
        RECT 1817.1200 1972.2800 1819.1200 1972.7600 ;
        RECT 1817.1200 1961.4000 1819.1200 1961.8800 ;
        RECT 1817.1200 1955.9600 1819.1200 1956.4400 ;
        RECT 1817.1200 1950.5200 1819.1200 1951.0000 ;
        RECT 1817.1200 1945.0800 1819.1200 1945.5600 ;
        RECT 1817.1200 1939.6400 1819.1200 1940.1200 ;
        RECT 1817.1200 1934.2000 1819.1200 1934.6800 ;
        RECT 1817.1200 1928.7600 1819.1200 1929.2400 ;
        RECT 1817.1200 1923.3200 1819.1200 1923.8000 ;
        RECT 1817.1200 1966.8400 1819.1200 1967.3200 ;
        RECT 2014.2200 2135.4800 2016.2200 2135.9600 ;
        RECT 1817.1200 2135.4800 1819.1200 2135.9600 ;
        RECT 1817.1200 2353.2000 2016.2200 2355.2000 ;
        RECT 1817.1200 1916.4100 2016.2200 1918.4100 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1817.1200 1457.1300 1819.1200 1895.9200 ;
        RECT 2014.2200 1457.1300 2016.2200 1895.9200 ;
        RECT 1821.6800 1457.1300 1823.2800 1895.9200 ;
        RECT 1866.6800 1457.1300 1868.2800 1895.9200 ;
        RECT 1911.6800 1457.1300 1913.2800 1895.9200 ;
        RECT 1956.6800 1457.1300 1958.2800 1895.9200 ;
        RECT 2001.6800 1457.1300 2003.2800 1895.9200 ;
      LAYER met3 ;
        RECT 2014.2200 1888.3600 2016.2200 1888.8400 ;
        RECT 2014.2200 1882.9200 2016.2200 1883.4000 ;
        RECT 2014.2200 1877.4800 2016.2200 1877.9600 ;
        RECT 2014.2200 1872.0400 2016.2200 1872.5200 ;
        RECT 2014.2200 1866.6000 2016.2200 1867.0800 ;
        RECT 2014.2200 1861.1600 2016.2200 1861.6400 ;
        RECT 2014.2200 1855.7200 2016.2200 1856.2000 ;
        RECT 2014.2200 1850.2800 2016.2200 1850.7600 ;
        RECT 2014.2200 1839.4000 2016.2200 1839.8800 ;
        RECT 2014.2200 1833.9600 2016.2200 1834.4400 ;
        RECT 2014.2200 1828.5200 2016.2200 1829.0000 ;
        RECT 2014.2200 1823.0800 2016.2200 1823.5600 ;
        RECT 2014.2200 1817.6400 2016.2200 1818.1200 ;
        RECT 2014.2200 1812.2000 2016.2200 1812.6800 ;
        RECT 2014.2200 1806.7600 2016.2200 1807.2400 ;
        RECT 2014.2200 1801.3200 2016.2200 1801.8000 ;
        RECT 2014.2200 1795.8800 2016.2200 1796.3600 ;
        RECT 2014.2200 1790.4400 2016.2200 1790.9200 ;
        RECT 2014.2200 1844.8400 2016.2200 1845.3200 ;
        RECT 2014.2200 1785.0000 2016.2200 1785.4800 ;
        RECT 2014.2200 1779.5600 2016.2200 1780.0400 ;
        RECT 2014.2200 1774.1200 2016.2200 1774.6000 ;
        RECT 2014.2200 1768.6800 2016.2200 1769.1600 ;
        RECT 2014.2200 1763.2400 2016.2200 1763.7200 ;
        RECT 2014.2200 1757.8000 2016.2200 1758.2800 ;
        RECT 2014.2200 1752.3600 2016.2200 1752.8400 ;
        RECT 2014.2200 1746.9200 2016.2200 1747.4000 ;
        RECT 2014.2200 1741.4800 2016.2200 1741.9600 ;
        RECT 2014.2200 1736.0400 2016.2200 1736.5200 ;
        RECT 2014.2200 1730.6000 2016.2200 1731.0800 ;
        RECT 2014.2200 1725.1600 2016.2200 1725.6400 ;
        RECT 2014.2200 1719.7200 2016.2200 1720.2000 ;
        RECT 2014.2200 1714.2800 2016.2200 1714.7600 ;
        RECT 2014.2200 1708.8400 2016.2200 1709.3200 ;
        RECT 2014.2200 1703.4000 2016.2200 1703.8800 ;
        RECT 2014.2200 1697.9600 2016.2200 1698.4400 ;
        RECT 2014.2200 1692.5200 2016.2200 1693.0000 ;
        RECT 2014.2200 1687.0800 2016.2200 1687.5600 ;
        RECT 2014.2200 1681.6400 2016.2200 1682.1200 ;
        RECT 1817.1200 1888.3600 1819.1200 1888.8400 ;
        RECT 1817.1200 1882.9200 1819.1200 1883.4000 ;
        RECT 1817.1200 1877.4800 1819.1200 1877.9600 ;
        RECT 1817.1200 1872.0400 1819.1200 1872.5200 ;
        RECT 1817.1200 1866.6000 1819.1200 1867.0800 ;
        RECT 1817.1200 1861.1600 1819.1200 1861.6400 ;
        RECT 1817.1200 1855.7200 1819.1200 1856.2000 ;
        RECT 1817.1200 1850.2800 1819.1200 1850.7600 ;
        RECT 1817.1200 1839.4000 1819.1200 1839.8800 ;
        RECT 1817.1200 1833.9600 1819.1200 1834.4400 ;
        RECT 1817.1200 1828.5200 1819.1200 1829.0000 ;
        RECT 1817.1200 1823.0800 1819.1200 1823.5600 ;
        RECT 1817.1200 1817.6400 1819.1200 1818.1200 ;
        RECT 1817.1200 1812.2000 1819.1200 1812.6800 ;
        RECT 1817.1200 1806.7600 1819.1200 1807.2400 ;
        RECT 1817.1200 1801.3200 1819.1200 1801.8000 ;
        RECT 1817.1200 1795.8800 1819.1200 1796.3600 ;
        RECT 1817.1200 1790.4400 1819.1200 1790.9200 ;
        RECT 1817.1200 1844.8400 1819.1200 1845.3200 ;
        RECT 1817.1200 1785.0000 1819.1200 1785.4800 ;
        RECT 1817.1200 1779.5600 1819.1200 1780.0400 ;
        RECT 1817.1200 1774.1200 1819.1200 1774.6000 ;
        RECT 1817.1200 1768.6800 1819.1200 1769.1600 ;
        RECT 1817.1200 1763.2400 1819.1200 1763.7200 ;
        RECT 1817.1200 1757.8000 1819.1200 1758.2800 ;
        RECT 1817.1200 1752.3600 1819.1200 1752.8400 ;
        RECT 1817.1200 1746.9200 1819.1200 1747.4000 ;
        RECT 1817.1200 1741.4800 1819.1200 1741.9600 ;
        RECT 1817.1200 1736.0400 1819.1200 1736.5200 ;
        RECT 1817.1200 1730.6000 1819.1200 1731.0800 ;
        RECT 1817.1200 1725.1600 1819.1200 1725.6400 ;
        RECT 1817.1200 1719.7200 1819.1200 1720.2000 ;
        RECT 1817.1200 1714.2800 1819.1200 1714.7600 ;
        RECT 1817.1200 1708.8400 1819.1200 1709.3200 ;
        RECT 1817.1200 1703.4000 1819.1200 1703.8800 ;
        RECT 1817.1200 1697.9600 1819.1200 1698.4400 ;
        RECT 1817.1200 1692.5200 1819.1200 1693.0000 ;
        RECT 1817.1200 1687.0800 1819.1200 1687.5600 ;
        RECT 1817.1200 1681.6400 1819.1200 1682.1200 ;
        RECT 2014.2200 1670.7600 2016.2200 1671.2400 ;
        RECT 2014.2200 1665.3200 2016.2200 1665.8000 ;
        RECT 2014.2200 1659.8800 2016.2200 1660.3600 ;
        RECT 2014.2200 1654.4400 2016.2200 1654.9200 ;
        RECT 2014.2200 1649.0000 2016.2200 1649.4800 ;
        RECT 2014.2200 1643.5600 2016.2200 1644.0400 ;
        RECT 2014.2200 1638.1200 2016.2200 1638.6000 ;
        RECT 2014.2200 1632.6800 2016.2200 1633.1600 ;
        RECT 2014.2200 1627.2400 2016.2200 1627.7200 ;
        RECT 2014.2200 1621.8000 2016.2200 1622.2800 ;
        RECT 2014.2200 1616.3600 2016.2200 1616.8400 ;
        RECT 2014.2200 1610.9200 2016.2200 1611.4000 ;
        RECT 2014.2200 1605.4800 2016.2200 1605.9600 ;
        RECT 2014.2200 1600.0400 2016.2200 1600.5200 ;
        RECT 2014.2200 1594.6000 2016.2200 1595.0800 ;
        RECT 2014.2200 1589.1600 2016.2200 1589.6400 ;
        RECT 2014.2200 1583.7200 2016.2200 1584.2000 ;
        RECT 2014.2200 1578.2800 2016.2200 1578.7600 ;
        RECT 2014.2200 1572.8400 2016.2200 1573.3200 ;
        RECT 2014.2200 1567.4000 2016.2200 1567.8800 ;
        RECT 2014.2200 1561.9600 2016.2200 1562.4400 ;
        RECT 2014.2200 1556.5200 2016.2200 1557.0000 ;
        RECT 2014.2200 1551.0800 2016.2200 1551.5600 ;
        RECT 2014.2200 1545.6400 2016.2200 1546.1200 ;
        RECT 2014.2200 1540.2000 2016.2200 1540.6800 ;
        RECT 2014.2200 1534.7600 2016.2200 1535.2400 ;
        RECT 2014.2200 1529.3200 2016.2200 1529.8000 ;
        RECT 2014.2200 1523.8800 2016.2200 1524.3600 ;
        RECT 2014.2200 1518.4400 2016.2200 1518.9200 ;
        RECT 2014.2200 1513.0000 2016.2200 1513.4800 ;
        RECT 2014.2200 1502.1200 2016.2200 1502.6000 ;
        RECT 2014.2200 1496.6800 2016.2200 1497.1600 ;
        RECT 2014.2200 1491.2400 2016.2200 1491.7200 ;
        RECT 2014.2200 1485.8000 2016.2200 1486.2800 ;
        RECT 2014.2200 1480.3600 2016.2200 1480.8400 ;
        RECT 2014.2200 1474.9200 2016.2200 1475.4000 ;
        RECT 2014.2200 1469.4800 2016.2200 1469.9600 ;
        RECT 2014.2200 1464.0400 2016.2200 1464.5200 ;
        RECT 2014.2200 1507.5600 2016.2200 1508.0400 ;
        RECT 1817.1200 1670.7600 1819.1200 1671.2400 ;
        RECT 1817.1200 1665.3200 1819.1200 1665.8000 ;
        RECT 1817.1200 1659.8800 1819.1200 1660.3600 ;
        RECT 1817.1200 1654.4400 1819.1200 1654.9200 ;
        RECT 1817.1200 1649.0000 1819.1200 1649.4800 ;
        RECT 1817.1200 1643.5600 1819.1200 1644.0400 ;
        RECT 1817.1200 1638.1200 1819.1200 1638.6000 ;
        RECT 1817.1200 1632.6800 1819.1200 1633.1600 ;
        RECT 1817.1200 1627.2400 1819.1200 1627.7200 ;
        RECT 1817.1200 1621.8000 1819.1200 1622.2800 ;
        RECT 1817.1200 1616.3600 1819.1200 1616.8400 ;
        RECT 1817.1200 1610.9200 1819.1200 1611.4000 ;
        RECT 1817.1200 1605.4800 1819.1200 1605.9600 ;
        RECT 1817.1200 1600.0400 1819.1200 1600.5200 ;
        RECT 1817.1200 1594.6000 1819.1200 1595.0800 ;
        RECT 1817.1200 1589.1600 1819.1200 1589.6400 ;
        RECT 1817.1200 1583.7200 1819.1200 1584.2000 ;
        RECT 1817.1200 1578.2800 1819.1200 1578.7600 ;
        RECT 1817.1200 1572.8400 1819.1200 1573.3200 ;
        RECT 1817.1200 1567.4000 1819.1200 1567.8800 ;
        RECT 1817.1200 1561.9600 1819.1200 1562.4400 ;
        RECT 1817.1200 1556.5200 1819.1200 1557.0000 ;
        RECT 1817.1200 1551.0800 1819.1200 1551.5600 ;
        RECT 1817.1200 1545.6400 1819.1200 1546.1200 ;
        RECT 1817.1200 1540.2000 1819.1200 1540.6800 ;
        RECT 1817.1200 1534.7600 1819.1200 1535.2400 ;
        RECT 1817.1200 1529.3200 1819.1200 1529.8000 ;
        RECT 1817.1200 1523.8800 1819.1200 1524.3600 ;
        RECT 1817.1200 1518.4400 1819.1200 1518.9200 ;
        RECT 1817.1200 1513.0000 1819.1200 1513.4800 ;
        RECT 1817.1200 1502.1200 1819.1200 1502.6000 ;
        RECT 1817.1200 1496.6800 1819.1200 1497.1600 ;
        RECT 1817.1200 1491.2400 1819.1200 1491.7200 ;
        RECT 1817.1200 1485.8000 1819.1200 1486.2800 ;
        RECT 1817.1200 1480.3600 1819.1200 1480.8400 ;
        RECT 1817.1200 1474.9200 1819.1200 1475.4000 ;
        RECT 1817.1200 1469.4800 1819.1200 1469.9600 ;
        RECT 1817.1200 1464.0400 1819.1200 1464.5200 ;
        RECT 1817.1200 1507.5600 1819.1200 1508.0400 ;
        RECT 2014.2200 1676.2000 2016.2200 1676.6800 ;
        RECT 1817.1200 1676.2000 1819.1200 1676.6800 ;
        RECT 1817.1200 1893.9200 2016.2200 1895.9200 ;
        RECT 1817.1200 1457.1300 2016.2200 1459.1300 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1817.1200 997.8500 1819.1200 1436.6400 ;
        RECT 2014.2200 997.8500 2016.2200 1436.6400 ;
        RECT 1821.6800 997.8500 1823.2800 1436.6400 ;
        RECT 1866.6800 997.8500 1868.2800 1436.6400 ;
        RECT 1911.6800 997.8500 1913.2800 1436.6400 ;
        RECT 1956.6800 997.8500 1958.2800 1436.6400 ;
        RECT 2001.6800 997.8500 2003.2800 1436.6400 ;
      LAYER met3 ;
        RECT 2014.2200 1429.0800 2016.2200 1429.5600 ;
        RECT 2014.2200 1423.6400 2016.2200 1424.1200 ;
        RECT 2014.2200 1418.2000 2016.2200 1418.6800 ;
        RECT 2014.2200 1412.7600 2016.2200 1413.2400 ;
        RECT 2014.2200 1407.3200 2016.2200 1407.8000 ;
        RECT 2014.2200 1401.8800 2016.2200 1402.3600 ;
        RECT 2014.2200 1396.4400 2016.2200 1396.9200 ;
        RECT 2014.2200 1391.0000 2016.2200 1391.4800 ;
        RECT 2014.2200 1380.1200 2016.2200 1380.6000 ;
        RECT 2014.2200 1374.6800 2016.2200 1375.1600 ;
        RECT 2014.2200 1369.2400 2016.2200 1369.7200 ;
        RECT 2014.2200 1363.8000 2016.2200 1364.2800 ;
        RECT 2014.2200 1358.3600 2016.2200 1358.8400 ;
        RECT 2014.2200 1352.9200 2016.2200 1353.4000 ;
        RECT 2014.2200 1347.4800 2016.2200 1347.9600 ;
        RECT 2014.2200 1342.0400 2016.2200 1342.5200 ;
        RECT 2014.2200 1336.6000 2016.2200 1337.0800 ;
        RECT 2014.2200 1331.1600 2016.2200 1331.6400 ;
        RECT 2014.2200 1385.5600 2016.2200 1386.0400 ;
        RECT 2014.2200 1325.7200 2016.2200 1326.2000 ;
        RECT 2014.2200 1320.2800 2016.2200 1320.7600 ;
        RECT 2014.2200 1314.8400 2016.2200 1315.3200 ;
        RECT 2014.2200 1309.4000 2016.2200 1309.8800 ;
        RECT 2014.2200 1303.9600 2016.2200 1304.4400 ;
        RECT 2014.2200 1298.5200 2016.2200 1299.0000 ;
        RECT 2014.2200 1293.0800 2016.2200 1293.5600 ;
        RECT 2014.2200 1287.6400 2016.2200 1288.1200 ;
        RECT 2014.2200 1282.2000 2016.2200 1282.6800 ;
        RECT 2014.2200 1276.7600 2016.2200 1277.2400 ;
        RECT 2014.2200 1271.3200 2016.2200 1271.8000 ;
        RECT 2014.2200 1265.8800 2016.2200 1266.3600 ;
        RECT 2014.2200 1260.4400 2016.2200 1260.9200 ;
        RECT 2014.2200 1255.0000 2016.2200 1255.4800 ;
        RECT 2014.2200 1249.5600 2016.2200 1250.0400 ;
        RECT 2014.2200 1244.1200 2016.2200 1244.6000 ;
        RECT 2014.2200 1238.6800 2016.2200 1239.1600 ;
        RECT 2014.2200 1233.2400 2016.2200 1233.7200 ;
        RECT 2014.2200 1227.8000 2016.2200 1228.2800 ;
        RECT 2014.2200 1222.3600 2016.2200 1222.8400 ;
        RECT 1817.1200 1429.0800 1819.1200 1429.5600 ;
        RECT 1817.1200 1423.6400 1819.1200 1424.1200 ;
        RECT 1817.1200 1418.2000 1819.1200 1418.6800 ;
        RECT 1817.1200 1412.7600 1819.1200 1413.2400 ;
        RECT 1817.1200 1407.3200 1819.1200 1407.8000 ;
        RECT 1817.1200 1401.8800 1819.1200 1402.3600 ;
        RECT 1817.1200 1396.4400 1819.1200 1396.9200 ;
        RECT 1817.1200 1391.0000 1819.1200 1391.4800 ;
        RECT 1817.1200 1380.1200 1819.1200 1380.6000 ;
        RECT 1817.1200 1374.6800 1819.1200 1375.1600 ;
        RECT 1817.1200 1369.2400 1819.1200 1369.7200 ;
        RECT 1817.1200 1363.8000 1819.1200 1364.2800 ;
        RECT 1817.1200 1358.3600 1819.1200 1358.8400 ;
        RECT 1817.1200 1352.9200 1819.1200 1353.4000 ;
        RECT 1817.1200 1347.4800 1819.1200 1347.9600 ;
        RECT 1817.1200 1342.0400 1819.1200 1342.5200 ;
        RECT 1817.1200 1336.6000 1819.1200 1337.0800 ;
        RECT 1817.1200 1331.1600 1819.1200 1331.6400 ;
        RECT 1817.1200 1385.5600 1819.1200 1386.0400 ;
        RECT 1817.1200 1325.7200 1819.1200 1326.2000 ;
        RECT 1817.1200 1320.2800 1819.1200 1320.7600 ;
        RECT 1817.1200 1314.8400 1819.1200 1315.3200 ;
        RECT 1817.1200 1309.4000 1819.1200 1309.8800 ;
        RECT 1817.1200 1303.9600 1819.1200 1304.4400 ;
        RECT 1817.1200 1298.5200 1819.1200 1299.0000 ;
        RECT 1817.1200 1293.0800 1819.1200 1293.5600 ;
        RECT 1817.1200 1287.6400 1819.1200 1288.1200 ;
        RECT 1817.1200 1282.2000 1819.1200 1282.6800 ;
        RECT 1817.1200 1276.7600 1819.1200 1277.2400 ;
        RECT 1817.1200 1271.3200 1819.1200 1271.8000 ;
        RECT 1817.1200 1265.8800 1819.1200 1266.3600 ;
        RECT 1817.1200 1260.4400 1819.1200 1260.9200 ;
        RECT 1817.1200 1255.0000 1819.1200 1255.4800 ;
        RECT 1817.1200 1249.5600 1819.1200 1250.0400 ;
        RECT 1817.1200 1244.1200 1819.1200 1244.6000 ;
        RECT 1817.1200 1238.6800 1819.1200 1239.1600 ;
        RECT 1817.1200 1233.2400 1819.1200 1233.7200 ;
        RECT 1817.1200 1227.8000 1819.1200 1228.2800 ;
        RECT 1817.1200 1222.3600 1819.1200 1222.8400 ;
        RECT 2014.2200 1211.4800 2016.2200 1211.9600 ;
        RECT 2014.2200 1206.0400 2016.2200 1206.5200 ;
        RECT 2014.2200 1200.6000 2016.2200 1201.0800 ;
        RECT 2014.2200 1195.1600 2016.2200 1195.6400 ;
        RECT 2014.2200 1189.7200 2016.2200 1190.2000 ;
        RECT 2014.2200 1184.2800 2016.2200 1184.7600 ;
        RECT 2014.2200 1178.8400 2016.2200 1179.3200 ;
        RECT 2014.2200 1173.4000 2016.2200 1173.8800 ;
        RECT 2014.2200 1167.9600 2016.2200 1168.4400 ;
        RECT 2014.2200 1162.5200 2016.2200 1163.0000 ;
        RECT 2014.2200 1157.0800 2016.2200 1157.5600 ;
        RECT 2014.2200 1151.6400 2016.2200 1152.1200 ;
        RECT 2014.2200 1146.2000 2016.2200 1146.6800 ;
        RECT 2014.2200 1140.7600 2016.2200 1141.2400 ;
        RECT 2014.2200 1135.3200 2016.2200 1135.8000 ;
        RECT 2014.2200 1129.8800 2016.2200 1130.3600 ;
        RECT 2014.2200 1124.4400 2016.2200 1124.9200 ;
        RECT 2014.2200 1119.0000 2016.2200 1119.4800 ;
        RECT 2014.2200 1113.5600 2016.2200 1114.0400 ;
        RECT 2014.2200 1108.1200 2016.2200 1108.6000 ;
        RECT 2014.2200 1102.6800 2016.2200 1103.1600 ;
        RECT 2014.2200 1097.2400 2016.2200 1097.7200 ;
        RECT 2014.2200 1091.8000 2016.2200 1092.2800 ;
        RECT 2014.2200 1086.3600 2016.2200 1086.8400 ;
        RECT 2014.2200 1080.9200 2016.2200 1081.4000 ;
        RECT 2014.2200 1075.4800 2016.2200 1075.9600 ;
        RECT 2014.2200 1070.0400 2016.2200 1070.5200 ;
        RECT 2014.2200 1064.6000 2016.2200 1065.0800 ;
        RECT 2014.2200 1059.1600 2016.2200 1059.6400 ;
        RECT 2014.2200 1053.7200 2016.2200 1054.2000 ;
        RECT 2014.2200 1042.8400 2016.2200 1043.3200 ;
        RECT 2014.2200 1037.4000 2016.2200 1037.8800 ;
        RECT 2014.2200 1031.9600 2016.2200 1032.4400 ;
        RECT 2014.2200 1026.5200 2016.2200 1027.0000 ;
        RECT 2014.2200 1021.0800 2016.2200 1021.5600 ;
        RECT 2014.2200 1015.6400 2016.2200 1016.1200 ;
        RECT 2014.2200 1010.2000 2016.2200 1010.6800 ;
        RECT 2014.2200 1004.7600 2016.2200 1005.2400 ;
        RECT 2014.2200 1048.2800 2016.2200 1048.7600 ;
        RECT 1817.1200 1211.4800 1819.1200 1211.9600 ;
        RECT 1817.1200 1206.0400 1819.1200 1206.5200 ;
        RECT 1817.1200 1200.6000 1819.1200 1201.0800 ;
        RECT 1817.1200 1195.1600 1819.1200 1195.6400 ;
        RECT 1817.1200 1189.7200 1819.1200 1190.2000 ;
        RECT 1817.1200 1184.2800 1819.1200 1184.7600 ;
        RECT 1817.1200 1178.8400 1819.1200 1179.3200 ;
        RECT 1817.1200 1173.4000 1819.1200 1173.8800 ;
        RECT 1817.1200 1167.9600 1819.1200 1168.4400 ;
        RECT 1817.1200 1162.5200 1819.1200 1163.0000 ;
        RECT 1817.1200 1157.0800 1819.1200 1157.5600 ;
        RECT 1817.1200 1151.6400 1819.1200 1152.1200 ;
        RECT 1817.1200 1146.2000 1819.1200 1146.6800 ;
        RECT 1817.1200 1140.7600 1819.1200 1141.2400 ;
        RECT 1817.1200 1135.3200 1819.1200 1135.8000 ;
        RECT 1817.1200 1129.8800 1819.1200 1130.3600 ;
        RECT 1817.1200 1124.4400 1819.1200 1124.9200 ;
        RECT 1817.1200 1119.0000 1819.1200 1119.4800 ;
        RECT 1817.1200 1113.5600 1819.1200 1114.0400 ;
        RECT 1817.1200 1108.1200 1819.1200 1108.6000 ;
        RECT 1817.1200 1102.6800 1819.1200 1103.1600 ;
        RECT 1817.1200 1097.2400 1819.1200 1097.7200 ;
        RECT 1817.1200 1091.8000 1819.1200 1092.2800 ;
        RECT 1817.1200 1086.3600 1819.1200 1086.8400 ;
        RECT 1817.1200 1080.9200 1819.1200 1081.4000 ;
        RECT 1817.1200 1075.4800 1819.1200 1075.9600 ;
        RECT 1817.1200 1070.0400 1819.1200 1070.5200 ;
        RECT 1817.1200 1064.6000 1819.1200 1065.0800 ;
        RECT 1817.1200 1059.1600 1819.1200 1059.6400 ;
        RECT 1817.1200 1053.7200 1819.1200 1054.2000 ;
        RECT 1817.1200 1042.8400 1819.1200 1043.3200 ;
        RECT 1817.1200 1037.4000 1819.1200 1037.8800 ;
        RECT 1817.1200 1031.9600 1819.1200 1032.4400 ;
        RECT 1817.1200 1026.5200 1819.1200 1027.0000 ;
        RECT 1817.1200 1021.0800 1819.1200 1021.5600 ;
        RECT 1817.1200 1015.6400 1819.1200 1016.1200 ;
        RECT 1817.1200 1010.2000 1819.1200 1010.6800 ;
        RECT 1817.1200 1004.7600 1819.1200 1005.2400 ;
        RECT 1817.1200 1048.2800 1819.1200 1048.7600 ;
        RECT 2014.2200 1216.9200 2016.2200 1217.4000 ;
        RECT 1817.1200 1216.9200 1819.1200 1217.4000 ;
        RECT 1817.1200 1434.6400 2016.2200 1436.6400 ;
        RECT 1817.1200 997.8500 2016.2200 999.8500 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1817.1200 538.5700 1819.1200 977.3600 ;
        RECT 2014.2200 538.5700 2016.2200 977.3600 ;
        RECT 1821.6800 538.5700 1823.2800 977.3600 ;
        RECT 1866.6800 538.5700 1868.2800 977.3600 ;
        RECT 1911.6800 538.5700 1913.2800 977.3600 ;
        RECT 1956.6800 538.5700 1958.2800 977.3600 ;
        RECT 2001.6800 538.5700 2003.2800 977.3600 ;
      LAYER met3 ;
        RECT 2014.2200 969.8000 2016.2200 970.2800 ;
        RECT 2014.2200 964.3600 2016.2200 964.8400 ;
        RECT 2014.2200 958.9200 2016.2200 959.4000 ;
        RECT 2014.2200 953.4800 2016.2200 953.9600 ;
        RECT 2014.2200 948.0400 2016.2200 948.5200 ;
        RECT 2014.2200 942.6000 2016.2200 943.0800 ;
        RECT 2014.2200 937.1600 2016.2200 937.6400 ;
        RECT 2014.2200 931.7200 2016.2200 932.2000 ;
        RECT 2014.2200 920.8400 2016.2200 921.3200 ;
        RECT 2014.2200 915.4000 2016.2200 915.8800 ;
        RECT 2014.2200 909.9600 2016.2200 910.4400 ;
        RECT 2014.2200 904.5200 2016.2200 905.0000 ;
        RECT 2014.2200 899.0800 2016.2200 899.5600 ;
        RECT 2014.2200 893.6400 2016.2200 894.1200 ;
        RECT 2014.2200 888.2000 2016.2200 888.6800 ;
        RECT 2014.2200 882.7600 2016.2200 883.2400 ;
        RECT 2014.2200 877.3200 2016.2200 877.8000 ;
        RECT 2014.2200 871.8800 2016.2200 872.3600 ;
        RECT 2014.2200 926.2800 2016.2200 926.7600 ;
        RECT 2014.2200 866.4400 2016.2200 866.9200 ;
        RECT 2014.2200 861.0000 2016.2200 861.4800 ;
        RECT 2014.2200 855.5600 2016.2200 856.0400 ;
        RECT 2014.2200 850.1200 2016.2200 850.6000 ;
        RECT 2014.2200 844.6800 2016.2200 845.1600 ;
        RECT 2014.2200 839.2400 2016.2200 839.7200 ;
        RECT 2014.2200 833.8000 2016.2200 834.2800 ;
        RECT 2014.2200 828.3600 2016.2200 828.8400 ;
        RECT 2014.2200 822.9200 2016.2200 823.4000 ;
        RECT 2014.2200 817.4800 2016.2200 817.9600 ;
        RECT 2014.2200 812.0400 2016.2200 812.5200 ;
        RECT 2014.2200 806.6000 2016.2200 807.0800 ;
        RECT 2014.2200 801.1600 2016.2200 801.6400 ;
        RECT 2014.2200 795.7200 2016.2200 796.2000 ;
        RECT 2014.2200 790.2800 2016.2200 790.7600 ;
        RECT 2014.2200 784.8400 2016.2200 785.3200 ;
        RECT 2014.2200 779.4000 2016.2200 779.8800 ;
        RECT 2014.2200 773.9600 2016.2200 774.4400 ;
        RECT 2014.2200 768.5200 2016.2200 769.0000 ;
        RECT 2014.2200 763.0800 2016.2200 763.5600 ;
        RECT 1817.1200 969.8000 1819.1200 970.2800 ;
        RECT 1817.1200 964.3600 1819.1200 964.8400 ;
        RECT 1817.1200 958.9200 1819.1200 959.4000 ;
        RECT 1817.1200 953.4800 1819.1200 953.9600 ;
        RECT 1817.1200 948.0400 1819.1200 948.5200 ;
        RECT 1817.1200 942.6000 1819.1200 943.0800 ;
        RECT 1817.1200 937.1600 1819.1200 937.6400 ;
        RECT 1817.1200 931.7200 1819.1200 932.2000 ;
        RECT 1817.1200 920.8400 1819.1200 921.3200 ;
        RECT 1817.1200 915.4000 1819.1200 915.8800 ;
        RECT 1817.1200 909.9600 1819.1200 910.4400 ;
        RECT 1817.1200 904.5200 1819.1200 905.0000 ;
        RECT 1817.1200 899.0800 1819.1200 899.5600 ;
        RECT 1817.1200 893.6400 1819.1200 894.1200 ;
        RECT 1817.1200 888.2000 1819.1200 888.6800 ;
        RECT 1817.1200 882.7600 1819.1200 883.2400 ;
        RECT 1817.1200 877.3200 1819.1200 877.8000 ;
        RECT 1817.1200 871.8800 1819.1200 872.3600 ;
        RECT 1817.1200 926.2800 1819.1200 926.7600 ;
        RECT 1817.1200 866.4400 1819.1200 866.9200 ;
        RECT 1817.1200 861.0000 1819.1200 861.4800 ;
        RECT 1817.1200 855.5600 1819.1200 856.0400 ;
        RECT 1817.1200 850.1200 1819.1200 850.6000 ;
        RECT 1817.1200 844.6800 1819.1200 845.1600 ;
        RECT 1817.1200 839.2400 1819.1200 839.7200 ;
        RECT 1817.1200 833.8000 1819.1200 834.2800 ;
        RECT 1817.1200 828.3600 1819.1200 828.8400 ;
        RECT 1817.1200 822.9200 1819.1200 823.4000 ;
        RECT 1817.1200 817.4800 1819.1200 817.9600 ;
        RECT 1817.1200 812.0400 1819.1200 812.5200 ;
        RECT 1817.1200 806.6000 1819.1200 807.0800 ;
        RECT 1817.1200 801.1600 1819.1200 801.6400 ;
        RECT 1817.1200 795.7200 1819.1200 796.2000 ;
        RECT 1817.1200 790.2800 1819.1200 790.7600 ;
        RECT 1817.1200 784.8400 1819.1200 785.3200 ;
        RECT 1817.1200 779.4000 1819.1200 779.8800 ;
        RECT 1817.1200 773.9600 1819.1200 774.4400 ;
        RECT 1817.1200 768.5200 1819.1200 769.0000 ;
        RECT 1817.1200 763.0800 1819.1200 763.5600 ;
        RECT 2014.2200 752.2000 2016.2200 752.6800 ;
        RECT 2014.2200 746.7600 2016.2200 747.2400 ;
        RECT 2014.2200 741.3200 2016.2200 741.8000 ;
        RECT 2014.2200 735.8800 2016.2200 736.3600 ;
        RECT 2014.2200 730.4400 2016.2200 730.9200 ;
        RECT 2014.2200 725.0000 2016.2200 725.4800 ;
        RECT 2014.2200 719.5600 2016.2200 720.0400 ;
        RECT 2014.2200 714.1200 2016.2200 714.6000 ;
        RECT 2014.2200 708.6800 2016.2200 709.1600 ;
        RECT 2014.2200 703.2400 2016.2200 703.7200 ;
        RECT 2014.2200 697.8000 2016.2200 698.2800 ;
        RECT 2014.2200 692.3600 2016.2200 692.8400 ;
        RECT 2014.2200 686.9200 2016.2200 687.4000 ;
        RECT 2014.2200 681.4800 2016.2200 681.9600 ;
        RECT 2014.2200 676.0400 2016.2200 676.5200 ;
        RECT 2014.2200 670.6000 2016.2200 671.0800 ;
        RECT 2014.2200 665.1600 2016.2200 665.6400 ;
        RECT 2014.2200 659.7200 2016.2200 660.2000 ;
        RECT 2014.2200 654.2800 2016.2200 654.7600 ;
        RECT 2014.2200 648.8400 2016.2200 649.3200 ;
        RECT 2014.2200 643.4000 2016.2200 643.8800 ;
        RECT 2014.2200 637.9600 2016.2200 638.4400 ;
        RECT 2014.2200 632.5200 2016.2200 633.0000 ;
        RECT 2014.2200 627.0800 2016.2200 627.5600 ;
        RECT 2014.2200 621.6400 2016.2200 622.1200 ;
        RECT 2014.2200 616.2000 2016.2200 616.6800 ;
        RECT 2014.2200 610.7600 2016.2200 611.2400 ;
        RECT 2014.2200 605.3200 2016.2200 605.8000 ;
        RECT 2014.2200 599.8800 2016.2200 600.3600 ;
        RECT 2014.2200 594.4400 2016.2200 594.9200 ;
        RECT 2014.2200 583.5600 2016.2200 584.0400 ;
        RECT 2014.2200 578.1200 2016.2200 578.6000 ;
        RECT 2014.2200 572.6800 2016.2200 573.1600 ;
        RECT 2014.2200 567.2400 2016.2200 567.7200 ;
        RECT 2014.2200 561.8000 2016.2200 562.2800 ;
        RECT 2014.2200 556.3600 2016.2200 556.8400 ;
        RECT 2014.2200 550.9200 2016.2200 551.4000 ;
        RECT 2014.2200 545.4800 2016.2200 545.9600 ;
        RECT 2014.2200 589.0000 2016.2200 589.4800 ;
        RECT 1817.1200 752.2000 1819.1200 752.6800 ;
        RECT 1817.1200 746.7600 1819.1200 747.2400 ;
        RECT 1817.1200 741.3200 1819.1200 741.8000 ;
        RECT 1817.1200 735.8800 1819.1200 736.3600 ;
        RECT 1817.1200 730.4400 1819.1200 730.9200 ;
        RECT 1817.1200 725.0000 1819.1200 725.4800 ;
        RECT 1817.1200 719.5600 1819.1200 720.0400 ;
        RECT 1817.1200 714.1200 1819.1200 714.6000 ;
        RECT 1817.1200 708.6800 1819.1200 709.1600 ;
        RECT 1817.1200 703.2400 1819.1200 703.7200 ;
        RECT 1817.1200 697.8000 1819.1200 698.2800 ;
        RECT 1817.1200 692.3600 1819.1200 692.8400 ;
        RECT 1817.1200 686.9200 1819.1200 687.4000 ;
        RECT 1817.1200 681.4800 1819.1200 681.9600 ;
        RECT 1817.1200 676.0400 1819.1200 676.5200 ;
        RECT 1817.1200 670.6000 1819.1200 671.0800 ;
        RECT 1817.1200 665.1600 1819.1200 665.6400 ;
        RECT 1817.1200 659.7200 1819.1200 660.2000 ;
        RECT 1817.1200 654.2800 1819.1200 654.7600 ;
        RECT 1817.1200 648.8400 1819.1200 649.3200 ;
        RECT 1817.1200 643.4000 1819.1200 643.8800 ;
        RECT 1817.1200 637.9600 1819.1200 638.4400 ;
        RECT 1817.1200 632.5200 1819.1200 633.0000 ;
        RECT 1817.1200 627.0800 1819.1200 627.5600 ;
        RECT 1817.1200 621.6400 1819.1200 622.1200 ;
        RECT 1817.1200 616.2000 1819.1200 616.6800 ;
        RECT 1817.1200 610.7600 1819.1200 611.2400 ;
        RECT 1817.1200 605.3200 1819.1200 605.8000 ;
        RECT 1817.1200 599.8800 1819.1200 600.3600 ;
        RECT 1817.1200 594.4400 1819.1200 594.9200 ;
        RECT 1817.1200 583.5600 1819.1200 584.0400 ;
        RECT 1817.1200 578.1200 1819.1200 578.6000 ;
        RECT 1817.1200 572.6800 1819.1200 573.1600 ;
        RECT 1817.1200 567.2400 1819.1200 567.7200 ;
        RECT 1817.1200 561.8000 1819.1200 562.2800 ;
        RECT 1817.1200 556.3600 1819.1200 556.8400 ;
        RECT 1817.1200 550.9200 1819.1200 551.4000 ;
        RECT 1817.1200 545.4800 1819.1200 545.9600 ;
        RECT 1817.1200 589.0000 1819.1200 589.4800 ;
        RECT 2014.2200 757.6400 2016.2200 758.1200 ;
        RECT 1817.1200 757.6400 1819.1200 758.1200 ;
        RECT 1817.1200 975.3600 2016.2200 977.3600 ;
        RECT 1817.1200 538.5700 2016.2200 540.5700 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 2037.3400 2833.6100 2039.3400 2854.5400 ;
        RECT 2234.4400 2833.6100 2236.4400 2854.5400 ;
      LAYER met3 ;
        RECT 2234.4400 2850.0400 2236.4400 2850.5200 ;
        RECT 2037.3400 2850.0400 2039.3400 2850.5200 ;
        RECT 2234.4400 2839.1600 2236.4400 2839.6400 ;
        RECT 2037.3400 2839.1600 2039.3400 2839.6400 ;
        RECT 2234.4400 2844.6000 2236.4400 2845.0800 ;
        RECT 2037.3400 2844.6000 2039.3400 2845.0800 ;
        RECT 2037.3400 2852.5400 2236.4400 2854.5400 ;
        RECT 2037.3400 2833.6100 2236.4400 2835.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 538.5700 2223.5000 746.6700 ;
        RECT 2176.9000 538.5700 2178.5000 746.6700 ;
        RECT 2131.9000 538.5700 2133.5000 746.6700 ;
        RECT 2086.9000 538.5700 2088.5000 746.6700 ;
        RECT 2233.4400 538.5700 2236.4400 746.6700 ;
        RECT 2037.3400 538.5700 2040.3400 746.6700 ;
      LAYER met3 ;
        RECT 2233.4400 741.3200 2236.4400 741.8000 ;
        RECT 2221.9000 741.3200 2223.5000 741.8000 ;
        RECT 2233.4400 730.4400 2236.4400 730.9200 ;
        RECT 2233.4400 735.8800 2236.4400 736.3600 ;
        RECT 2221.9000 730.4400 2223.5000 730.9200 ;
        RECT 2221.9000 735.8800 2223.5000 736.3600 ;
        RECT 2233.4400 714.1200 2236.4400 714.6000 ;
        RECT 2233.4400 719.5600 2236.4400 720.0400 ;
        RECT 2221.9000 714.1200 2223.5000 714.6000 ;
        RECT 2221.9000 719.5600 2223.5000 720.0400 ;
        RECT 2233.4400 703.2400 2236.4400 703.7200 ;
        RECT 2233.4400 708.6800 2236.4400 709.1600 ;
        RECT 2221.9000 703.2400 2223.5000 703.7200 ;
        RECT 2221.9000 708.6800 2223.5000 709.1600 ;
        RECT 2233.4400 725.0000 2236.4400 725.4800 ;
        RECT 2221.9000 725.0000 2223.5000 725.4800 ;
        RECT 2176.9000 730.4400 2178.5000 730.9200 ;
        RECT 2176.9000 735.8800 2178.5000 736.3600 ;
        RECT 2176.9000 741.3200 2178.5000 741.8000 ;
        RECT 2176.9000 714.1200 2178.5000 714.6000 ;
        RECT 2176.9000 719.5600 2178.5000 720.0400 ;
        RECT 2176.9000 708.6800 2178.5000 709.1600 ;
        RECT 2176.9000 703.2400 2178.5000 703.7200 ;
        RECT 2176.9000 725.0000 2178.5000 725.4800 ;
        RECT 2233.4400 686.9200 2236.4400 687.4000 ;
        RECT 2233.4400 692.3600 2236.4400 692.8400 ;
        RECT 2221.9000 686.9200 2223.5000 687.4000 ;
        RECT 2221.9000 692.3600 2223.5000 692.8400 ;
        RECT 2233.4400 670.6000 2236.4400 671.0800 ;
        RECT 2233.4400 676.0400 2236.4400 676.5200 ;
        RECT 2233.4400 681.4800 2236.4400 681.9600 ;
        RECT 2221.9000 670.6000 2223.5000 671.0800 ;
        RECT 2221.9000 676.0400 2223.5000 676.5200 ;
        RECT 2221.9000 681.4800 2223.5000 681.9600 ;
        RECT 2233.4400 659.7200 2236.4400 660.2000 ;
        RECT 2233.4400 665.1600 2236.4400 665.6400 ;
        RECT 2221.9000 659.7200 2223.5000 660.2000 ;
        RECT 2221.9000 665.1600 2223.5000 665.6400 ;
        RECT 2233.4400 643.4000 2236.4400 643.8800 ;
        RECT 2233.4400 648.8400 2236.4400 649.3200 ;
        RECT 2233.4400 654.2800 2236.4400 654.7600 ;
        RECT 2221.9000 643.4000 2223.5000 643.8800 ;
        RECT 2221.9000 648.8400 2223.5000 649.3200 ;
        RECT 2221.9000 654.2800 2223.5000 654.7600 ;
        RECT 2176.9000 686.9200 2178.5000 687.4000 ;
        RECT 2176.9000 692.3600 2178.5000 692.8400 ;
        RECT 2176.9000 670.6000 2178.5000 671.0800 ;
        RECT 2176.9000 676.0400 2178.5000 676.5200 ;
        RECT 2176.9000 681.4800 2178.5000 681.9600 ;
        RECT 2176.9000 659.7200 2178.5000 660.2000 ;
        RECT 2176.9000 665.1600 2178.5000 665.6400 ;
        RECT 2176.9000 643.4000 2178.5000 643.8800 ;
        RECT 2176.9000 648.8400 2178.5000 649.3200 ;
        RECT 2176.9000 654.2800 2178.5000 654.7600 ;
        RECT 2233.4400 697.8000 2236.4400 698.2800 ;
        RECT 2176.9000 697.8000 2178.5000 698.2800 ;
        RECT 2221.9000 697.8000 2223.5000 698.2800 ;
        RECT 2131.9000 730.4400 2133.5000 730.9200 ;
        RECT 2131.9000 735.8800 2133.5000 736.3600 ;
        RECT 2131.9000 741.3200 2133.5000 741.8000 ;
        RECT 2086.9000 730.4400 2088.5000 730.9200 ;
        RECT 2086.9000 735.8800 2088.5000 736.3600 ;
        RECT 2086.9000 741.3200 2088.5000 741.8000 ;
        RECT 2131.9000 714.1200 2133.5000 714.6000 ;
        RECT 2131.9000 719.5600 2133.5000 720.0400 ;
        RECT 2131.9000 703.2400 2133.5000 703.7200 ;
        RECT 2131.9000 708.6800 2133.5000 709.1600 ;
        RECT 2086.9000 714.1200 2088.5000 714.6000 ;
        RECT 2086.9000 719.5600 2088.5000 720.0400 ;
        RECT 2086.9000 703.2400 2088.5000 703.7200 ;
        RECT 2086.9000 708.6800 2088.5000 709.1600 ;
        RECT 2086.9000 725.0000 2088.5000 725.4800 ;
        RECT 2131.9000 725.0000 2133.5000 725.4800 ;
        RECT 2037.3400 741.3200 2040.3400 741.8000 ;
        RECT 2037.3400 735.8800 2040.3400 736.3600 ;
        RECT 2037.3400 730.4400 2040.3400 730.9200 ;
        RECT 2037.3400 719.5600 2040.3400 720.0400 ;
        RECT 2037.3400 714.1200 2040.3400 714.6000 ;
        RECT 2037.3400 708.6800 2040.3400 709.1600 ;
        RECT 2037.3400 703.2400 2040.3400 703.7200 ;
        RECT 2037.3400 725.0000 2040.3400 725.4800 ;
        RECT 2131.9000 686.9200 2133.5000 687.4000 ;
        RECT 2131.9000 692.3600 2133.5000 692.8400 ;
        RECT 2131.9000 670.6000 2133.5000 671.0800 ;
        RECT 2131.9000 676.0400 2133.5000 676.5200 ;
        RECT 2131.9000 681.4800 2133.5000 681.9600 ;
        RECT 2086.9000 686.9200 2088.5000 687.4000 ;
        RECT 2086.9000 692.3600 2088.5000 692.8400 ;
        RECT 2086.9000 670.6000 2088.5000 671.0800 ;
        RECT 2086.9000 676.0400 2088.5000 676.5200 ;
        RECT 2086.9000 681.4800 2088.5000 681.9600 ;
        RECT 2131.9000 659.7200 2133.5000 660.2000 ;
        RECT 2131.9000 665.1600 2133.5000 665.6400 ;
        RECT 2131.9000 643.4000 2133.5000 643.8800 ;
        RECT 2131.9000 648.8400 2133.5000 649.3200 ;
        RECT 2131.9000 654.2800 2133.5000 654.7600 ;
        RECT 2086.9000 659.7200 2088.5000 660.2000 ;
        RECT 2086.9000 665.1600 2088.5000 665.6400 ;
        RECT 2086.9000 643.4000 2088.5000 643.8800 ;
        RECT 2086.9000 648.8400 2088.5000 649.3200 ;
        RECT 2086.9000 654.2800 2088.5000 654.7600 ;
        RECT 2037.3400 686.9200 2040.3400 687.4000 ;
        RECT 2037.3400 692.3600 2040.3400 692.8400 ;
        RECT 2037.3400 676.0400 2040.3400 676.5200 ;
        RECT 2037.3400 670.6000 2040.3400 671.0800 ;
        RECT 2037.3400 681.4800 2040.3400 681.9600 ;
        RECT 2037.3400 659.7200 2040.3400 660.2000 ;
        RECT 2037.3400 665.1600 2040.3400 665.6400 ;
        RECT 2037.3400 648.8400 2040.3400 649.3200 ;
        RECT 2037.3400 643.4000 2040.3400 643.8800 ;
        RECT 2037.3400 654.2800 2040.3400 654.7600 ;
        RECT 2037.3400 697.8000 2040.3400 698.2800 ;
        RECT 2086.9000 697.8000 2088.5000 698.2800 ;
        RECT 2131.9000 697.8000 2133.5000 698.2800 ;
        RECT 2233.4400 632.5200 2236.4400 633.0000 ;
        RECT 2233.4400 637.9600 2236.4400 638.4400 ;
        RECT 2221.9000 632.5200 2223.5000 633.0000 ;
        RECT 2221.9000 637.9600 2223.5000 638.4400 ;
        RECT 2233.4400 616.2000 2236.4400 616.6800 ;
        RECT 2233.4400 621.6400 2236.4400 622.1200 ;
        RECT 2233.4400 627.0800 2236.4400 627.5600 ;
        RECT 2221.9000 616.2000 2223.5000 616.6800 ;
        RECT 2221.9000 621.6400 2223.5000 622.1200 ;
        RECT 2221.9000 627.0800 2223.5000 627.5600 ;
        RECT 2233.4400 605.3200 2236.4400 605.8000 ;
        RECT 2233.4400 610.7600 2236.4400 611.2400 ;
        RECT 2221.9000 605.3200 2223.5000 605.8000 ;
        RECT 2221.9000 610.7600 2223.5000 611.2400 ;
        RECT 2233.4400 589.0000 2236.4400 589.4800 ;
        RECT 2233.4400 594.4400 2236.4400 594.9200 ;
        RECT 2233.4400 599.8800 2236.4400 600.3600 ;
        RECT 2221.9000 589.0000 2223.5000 589.4800 ;
        RECT 2221.9000 594.4400 2223.5000 594.9200 ;
        RECT 2221.9000 599.8800 2223.5000 600.3600 ;
        RECT 2176.9000 632.5200 2178.5000 633.0000 ;
        RECT 2176.9000 637.9600 2178.5000 638.4400 ;
        RECT 2176.9000 616.2000 2178.5000 616.6800 ;
        RECT 2176.9000 621.6400 2178.5000 622.1200 ;
        RECT 2176.9000 627.0800 2178.5000 627.5600 ;
        RECT 2176.9000 605.3200 2178.5000 605.8000 ;
        RECT 2176.9000 610.7600 2178.5000 611.2400 ;
        RECT 2176.9000 589.0000 2178.5000 589.4800 ;
        RECT 2176.9000 594.4400 2178.5000 594.9200 ;
        RECT 2176.9000 599.8800 2178.5000 600.3600 ;
        RECT 2233.4400 578.1200 2236.4400 578.6000 ;
        RECT 2233.4400 583.5600 2236.4400 584.0400 ;
        RECT 2221.9000 578.1200 2223.5000 578.6000 ;
        RECT 2221.9000 583.5600 2223.5000 584.0400 ;
        RECT 2233.4400 561.8000 2236.4400 562.2800 ;
        RECT 2233.4400 567.2400 2236.4400 567.7200 ;
        RECT 2233.4400 572.6800 2236.4400 573.1600 ;
        RECT 2221.9000 561.8000 2223.5000 562.2800 ;
        RECT 2221.9000 567.2400 2223.5000 567.7200 ;
        RECT 2221.9000 572.6800 2223.5000 573.1600 ;
        RECT 2233.4400 550.9200 2236.4400 551.4000 ;
        RECT 2233.4400 556.3600 2236.4400 556.8400 ;
        RECT 2221.9000 550.9200 2223.5000 551.4000 ;
        RECT 2221.9000 556.3600 2223.5000 556.8400 ;
        RECT 2233.4400 545.4800 2236.4400 545.9600 ;
        RECT 2221.9000 545.4800 2223.5000 545.9600 ;
        RECT 2176.9000 578.1200 2178.5000 578.6000 ;
        RECT 2176.9000 583.5600 2178.5000 584.0400 ;
        RECT 2176.9000 561.8000 2178.5000 562.2800 ;
        RECT 2176.9000 567.2400 2178.5000 567.7200 ;
        RECT 2176.9000 572.6800 2178.5000 573.1600 ;
        RECT 2176.9000 550.9200 2178.5000 551.4000 ;
        RECT 2176.9000 556.3600 2178.5000 556.8400 ;
        RECT 2176.9000 545.4800 2178.5000 545.9600 ;
        RECT 2131.9000 632.5200 2133.5000 633.0000 ;
        RECT 2131.9000 637.9600 2133.5000 638.4400 ;
        RECT 2131.9000 616.2000 2133.5000 616.6800 ;
        RECT 2131.9000 621.6400 2133.5000 622.1200 ;
        RECT 2131.9000 627.0800 2133.5000 627.5600 ;
        RECT 2086.9000 632.5200 2088.5000 633.0000 ;
        RECT 2086.9000 637.9600 2088.5000 638.4400 ;
        RECT 2086.9000 616.2000 2088.5000 616.6800 ;
        RECT 2086.9000 621.6400 2088.5000 622.1200 ;
        RECT 2086.9000 627.0800 2088.5000 627.5600 ;
        RECT 2131.9000 605.3200 2133.5000 605.8000 ;
        RECT 2131.9000 610.7600 2133.5000 611.2400 ;
        RECT 2131.9000 589.0000 2133.5000 589.4800 ;
        RECT 2131.9000 594.4400 2133.5000 594.9200 ;
        RECT 2131.9000 599.8800 2133.5000 600.3600 ;
        RECT 2086.9000 605.3200 2088.5000 605.8000 ;
        RECT 2086.9000 610.7600 2088.5000 611.2400 ;
        RECT 2086.9000 589.0000 2088.5000 589.4800 ;
        RECT 2086.9000 594.4400 2088.5000 594.9200 ;
        RECT 2086.9000 599.8800 2088.5000 600.3600 ;
        RECT 2037.3400 632.5200 2040.3400 633.0000 ;
        RECT 2037.3400 637.9600 2040.3400 638.4400 ;
        RECT 2037.3400 621.6400 2040.3400 622.1200 ;
        RECT 2037.3400 616.2000 2040.3400 616.6800 ;
        RECT 2037.3400 627.0800 2040.3400 627.5600 ;
        RECT 2037.3400 605.3200 2040.3400 605.8000 ;
        RECT 2037.3400 610.7600 2040.3400 611.2400 ;
        RECT 2037.3400 594.4400 2040.3400 594.9200 ;
        RECT 2037.3400 589.0000 2040.3400 589.4800 ;
        RECT 2037.3400 599.8800 2040.3400 600.3600 ;
        RECT 2131.9000 578.1200 2133.5000 578.6000 ;
        RECT 2131.9000 583.5600 2133.5000 584.0400 ;
        RECT 2131.9000 561.8000 2133.5000 562.2800 ;
        RECT 2131.9000 567.2400 2133.5000 567.7200 ;
        RECT 2131.9000 572.6800 2133.5000 573.1600 ;
        RECT 2086.9000 578.1200 2088.5000 578.6000 ;
        RECT 2086.9000 583.5600 2088.5000 584.0400 ;
        RECT 2086.9000 561.8000 2088.5000 562.2800 ;
        RECT 2086.9000 567.2400 2088.5000 567.7200 ;
        RECT 2086.9000 572.6800 2088.5000 573.1600 ;
        RECT 2131.9000 556.3600 2133.5000 556.8400 ;
        RECT 2131.9000 550.9200 2133.5000 551.4000 ;
        RECT 2131.9000 545.4800 2133.5000 545.9600 ;
        RECT 2086.9000 556.3600 2088.5000 556.8400 ;
        RECT 2086.9000 550.9200 2088.5000 551.4000 ;
        RECT 2086.9000 545.4800 2088.5000 545.9600 ;
        RECT 2037.3400 578.1200 2040.3400 578.6000 ;
        RECT 2037.3400 583.5600 2040.3400 584.0400 ;
        RECT 2037.3400 567.2400 2040.3400 567.7200 ;
        RECT 2037.3400 561.8000 2040.3400 562.2800 ;
        RECT 2037.3400 572.6800 2040.3400 573.1600 ;
        RECT 2037.3400 550.9200 2040.3400 551.4000 ;
        RECT 2037.3400 556.3600 2040.3400 556.8400 ;
        RECT 2037.3400 545.4800 2040.3400 545.9600 ;
        RECT 2037.3400 743.6700 2236.4400 746.6700 ;
        RECT 2037.3400 538.5700 2236.4400 541.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 308.9300 2223.5000 517.0300 ;
        RECT 2176.9000 308.9300 2178.5000 517.0300 ;
        RECT 2131.9000 308.9300 2133.5000 517.0300 ;
        RECT 2086.9000 308.9300 2088.5000 517.0300 ;
        RECT 2233.4400 308.9300 2236.4400 517.0300 ;
        RECT 2037.3400 308.9300 2040.3400 517.0300 ;
      LAYER met3 ;
        RECT 2233.4400 511.6800 2236.4400 512.1600 ;
        RECT 2221.9000 511.6800 2223.5000 512.1600 ;
        RECT 2233.4400 500.8000 2236.4400 501.2800 ;
        RECT 2233.4400 506.2400 2236.4400 506.7200 ;
        RECT 2221.9000 500.8000 2223.5000 501.2800 ;
        RECT 2221.9000 506.2400 2223.5000 506.7200 ;
        RECT 2233.4400 484.4800 2236.4400 484.9600 ;
        RECT 2233.4400 489.9200 2236.4400 490.4000 ;
        RECT 2221.9000 484.4800 2223.5000 484.9600 ;
        RECT 2221.9000 489.9200 2223.5000 490.4000 ;
        RECT 2233.4400 473.6000 2236.4400 474.0800 ;
        RECT 2233.4400 479.0400 2236.4400 479.5200 ;
        RECT 2221.9000 473.6000 2223.5000 474.0800 ;
        RECT 2221.9000 479.0400 2223.5000 479.5200 ;
        RECT 2233.4400 495.3600 2236.4400 495.8400 ;
        RECT 2221.9000 495.3600 2223.5000 495.8400 ;
        RECT 2176.9000 500.8000 2178.5000 501.2800 ;
        RECT 2176.9000 506.2400 2178.5000 506.7200 ;
        RECT 2176.9000 511.6800 2178.5000 512.1600 ;
        RECT 2176.9000 484.4800 2178.5000 484.9600 ;
        RECT 2176.9000 489.9200 2178.5000 490.4000 ;
        RECT 2176.9000 479.0400 2178.5000 479.5200 ;
        RECT 2176.9000 473.6000 2178.5000 474.0800 ;
        RECT 2176.9000 495.3600 2178.5000 495.8400 ;
        RECT 2233.4400 457.2800 2236.4400 457.7600 ;
        RECT 2233.4400 462.7200 2236.4400 463.2000 ;
        RECT 2221.9000 457.2800 2223.5000 457.7600 ;
        RECT 2221.9000 462.7200 2223.5000 463.2000 ;
        RECT 2233.4400 440.9600 2236.4400 441.4400 ;
        RECT 2233.4400 446.4000 2236.4400 446.8800 ;
        RECT 2233.4400 451.8400 2236.4400 452.3200 ;
        RECT 2221.9000 440.9600 2223.5000 441.4400 ;
        RECT 2221.9000 446.4000 2223.5000 446.8800 ;
        RECT 2221.9000 451.8400 2223.5000 452.3200 ;
        RECT 2233.4400 430.0800 2236.4400 430.5600 ;
        RECT 2233.4400 435.5200 2236.4400 436.0000 ;
        RECT 2221.9000 430.0800 2223.5000 430.5600 ;
        RECT 2221.9000 435.5200 2223.5000 436.0000 ;
        RECT 2233.4400 413.7600 2236.4400 414.2400 ;
        RECT 2233.4400 419.2000 2236.4400 419.6800 ;
        RECT 2233.4400 424.6400 2236.4400 425.1200 ;
        RECT 2221.9000 413.7600 2223.5000 414.2400 ;
        RECT 2221.9000 419.2000 2223.5000 419.6800 ;
        RECT 2221.9000 424.6400 2223.5000 425.1200 ;
        RECT 2176.9000 457.2800 2178.5000 457.7600 ;
        RECT 2176.9000 462.7200 2178.5000 463.2000 ;
        RECT 2176.9000 440.9600 2178.5000 441.4400 ;
        RECT 2176.9000 446.4000 2178.5000 446.8800 ;
        RECT 2176.9000 451.8400 2178.5000 452.3200 ;
        RECT 2176.9000 430.0800 2178.5000 430.5600 ;
        RECT 2176.9000 435.5200 2178.5000 436.0000 ;
        RECT 2176.9000 413.7600 2178.5000 414.2400 ;
        RECT 2176.9000 419.2000 2178.5000 419.6800 ;
        RECT 2176.9000 424.6400 2178.5000 425.1200 ;
        RECT 2233.4400 468.1600 2236.4400 468.6400 ;
        RECT 2176.9000 468.1600 2178.5000 468.6400 ;
        RECT 2221.9000 468.1600 2223.5000 468.6400 ;
        RECT 2131.9000 500.8000 2133.5000 501.2800 ;
        RECT 2131.9000 506.2400 2133.5000 506.7200 ;
        RECT 2131.9000 511.6800 2133.5000 512.1600 ;
        RECT 2086.9000 500.8000 2088.5000 501.2800 ;
        RECT 2086.9000 506.2400 2088.5000 506.7200 ;
        RECT 2086.9000 511.6800 2088.5000 512.1600 ;
        RECT 2131.9000 484.4800 2133.5000 484.9600 ;
        RECT 2131.9000 489.9200 2133.5000 490.4000 ;
        RECT 2131.9000 473.6000 2133.5000 474.0800 ;
        RECT 2131.9000 479.0400 2133.5000 479.5200 ;
        RECT 2086.9000 484.4800 2088.5000 484.9600 ;
        RECT 2086.9000 489.9200 2088.5000 490.4000 ;
        RECT 2086.9000 473.6000 2088.5000 474.0800 ;
        RECT 2086.9000 479.0400 2088.5000 479.5200 ;
        RECT 2086.9000 495.3600 2088.5000 495.8400 ;
        RECT 2131.9000 495.3600 2133.5000 495.8400 ;
        RECT 2037.3400 511.6800 2040.3400 512.1600 ;
        RECT 2037.3400 506.2400 2040.3400 506.7200 ;
        RECT 2037.3400 500.8000 2040.3400 501.2800 ;
        RECT 2037.3400 489.9200 2040.3400 490.4000 ;
        RECT 2037.3400 484.4800 2040.3400 484.9600 ;
        RECT 2037.3400 479.0400 2040.3400 479.5200 ;
        RECT 2037.3400 473.6000 2040.3400 474.0800 ;
        RECT 2037.3400 495.3600 2040.3400 495.8400 ;
        RECT 2131.9000 457.2800 2133.5000 457.7600 ;
        RECT 2131.9000 462.7200 2133.5000 463.2000 ;
        RECT 2131.9000 440.9600 2133.5000 441.4400 ;
        RECT 2131.9000 446.4000 2133.5000 446.8800 ;
        RECT 2131.9000 451.8400 2133.5000 452.3200 ;
        RECT 2086.9000 457.2800 2088.5000 457.7600 ;
        RECT 2086.9000 462.7200 2088.5000 463.2000 ;
        RECT 2086.9000 440.9600 2088.5000 441.4400 ;
        RECT 2086.9000 446.4000 2088.5000 446.8800 ;
        RECT 2086.9000 451.8400 2088.5000 452.3200 ;
        RECT 2131.9000 430.0800 2133.5000 430.5600 ;
        RECT 2131.9000 435.5200 2133.5000 436.0000 ;
        RECT 2131.9000 413.7600 2133.5000 414.2400 ;
        RECT 2131.9000 419.2000 2133.5000 419.6800 ;
        RECT 2131.9000 424.6400 2133.5000 425.1200 ;
        RECT 2086.9000 430.0800 2088.5000 430.5600 ;
        RECT 2086.9000 435.5200 2088.5000 436.0000 ;
        RECT 2086.9000 413.7600 2088.5000 414.2400 ;
        RECT 2086.9000 419.2000 2088.5000 419.6800 ;
        RECT 2086.9000 424.6400 2088.5000 425.1200 ;
        RECT 2037.3400 457.2800 2040.3400 457.7600 ;
        RECT 2037.3400 462.7200 2040.3400 463.2000 ;
        RECT 2037.3400 446.4000 2040.3400 446.8800 ;
        RECT 2037.3400 440.9600 2040.3400 441.4400 ;
        RECT 2037.3400 451.8400 2040.3400 452.3200 ;
        RECT 2037.3400 430.0800 2040.3400 430.5600 ;
        RECT 2037.3400 435.5200 2040.3400 436.0000 ;
        RECT 2037.3400 419.2000 2040.3400 419.6800 ;
        RECT 2037.3400 413.7600 2040.3400 414.2400 ;
        RECT 2037.3400 424.6400 2040.3400 425.1200 ;
        RECT 2037.3400 468.1600 2040.3400 468.6400 ;
        RECT 2086.9000 468.1600 2088.5000 468.6400 ;
        RECT 2131.9000 468.1600 2133.5000 468.6400 ;
        RECT 2233.4400 402.8800 2236.4400 403.3600 ;
        RECT 2233.4400 408.3200 2236.4400 408.8000 ;
        RECT 2221.9000 402.8800 2223.5000 403.3600 ;
        RECT 2221.9000 408.3200 2223.5000 408.8000 ;
        RECT 2233.4400 386.5600 2236.4400 387.0400 ;
        RECT 2233.4400 392.0000 2236.4400 392.4800 ;
        RECT 2233.4400 397.4400 2236.4400 397.9200 ;
        RECT 2221.9000 386.5600 2223.5000 387.0400 ;
        RECT 2221.9000 392.0000 2223.5000 392.4800 ;
        RECT 2221.9000 397.4400 2223.5000 397.9200 ;
        RECT 2233.4400 375.6800 2236.4400 376.1600 ;
        RECT 2233.4400 381.1200 2236.4400 381.6000 ;
        RECT 2221.9000 375.6800 2223.5000 376.1600 ;
        RECT 2221.9000 381.1200 2223.5000 381.6000 ;
        RECT 2233.4400 359.3600 2236.4400 359.8400 ;
        RECT 2233.4400 364.8000 2236.4400 365.2800 ;
        RECT 2233.4400 370.2400 2236.4400 370.7200 ;
        RECT 2221.9000 359.3600 2223.5000 359.8400 ;
        RECT 2221.9000 364.8000 2223.5000 365.2800 ;
        RECT 2221.9000 370.2400 2223.5000 370.7200 ;
        RECT 2176.9000 402.8800 2178.5000 403.3600 ;
        RECT 2176.9000 408.3200 2178.5000 408.8000 ;
        RECT 2176.9000 386.5600 2178.5000 387.0400 ;
        RECT 2176.9000 392.0000 2178.5000 392.4800 ;
        RECT 2176.9000 397.4400 2178.5000 397.9200 ;
        RECT 2176.9000 375.6800 2178.5000 376.1600 ;
        RECT 2176.9000 381.1200 2178.5000 381.6000 ;
        RECT 2176.9000 359.3600 2178.5000 359.8400 ;
        RECT 2176.9000 364.8000 2178.5000 365.2800 ;
        RECT 2176.9000 370.2400 2178.5000 370.7200 ;
        RECT 2233.4400 348.4800 2236.4400 348.9600 ;
        RECT 2233.4400 353.9200 2236.4400 354.4000 ;
        RECT 2221.9000 348.4800 2223.5000 348.9600 ;
        RECT 2221.9000 353.9200 2223.5000 354.4000 ;
        RECT 2233.4400 332.1600 2236.4400 332.6400 ;
        RECT 2233.4400 337.6000 2236.4400 338.0800 ;
        RECT 2233.4400 343.0400 2236.4400 343.5200 ;
        RECT 2221.9000 332.1600 2223.5000 332.6400 ;
        RECT 2221.9000 337.6000 2223.5000 338.0800 ;
        RECT 2221.9000 343.0400 2223.5000 343.5200 ;
        RECT 2233.4400 321.2800 2236.4400 321.7600 ;
        RECT 2233.4400 326.7200 2236.4400 327.2000 ;
        RECT 2221.9000 321.2800 2223.5000 321.7600 ;
        RECT 2221.9000 326.7200 2223.5000 327.2000 ;
        RECT 2233.4400 315.8400 2236.4400 316.3200 ;
        RECT 2221.9000 315.8400 2223.5000 316.3200 ;
        RECT 2176.9000 348.4800 2178.5000 348.9600 ;
        RECT 2176.9000 353.9200 2178.5000 354.4000 ;
        RECT 2176.9000 332.1600 2178.5000 332.6400 ;
        RECT 2176.9000 337.6000 2178.5000 338.0800 ;
        RECT 2176.9000 343.0400 2178.5000 343.5200 ;
        RECT 2176.9000 321.2800 2178.5000 321.7600 ;
        RECT 2176.9000 326.7200 2178.5000 327.2000 ;
        RECT 2176.9000 315.8400 2178.5000 316.3200 ;
        RECT 2131.9000 402.8800 2133.5000 403.3600 ;
        RECT 2131.9000 408.3200 2133.5000 408.8000 ;
        RECT 2131.9000 386.5600 2133.5000 387.0400 ;
        RECT 2131.9000 392.0000 2133.5000 392.4800 ;
        RECT 2131.9000 397.4400 2133.5000 397.9200 ;
        RECT 2086.9000 402.8800 2088.5000 403.3600 ;
        RECT 2086.9000 408.3200 2088.5000 408.8000 ;
        RECT 2086.9000 386.5600 2088.5000 387.0400 ;
        RECT 2086.9000 392.0000 2088.5000 392.4800 ;
        RECT 2086.9000 397.4400 2088.5000 397.9200 ;
        RECT 2131.9000 375.6800 2133.5000 376.1600 ;
        RECT 2131.9000 381.1200 2133.5000 381.6000 ;
        RECT 2131.9000 359.3600 2133.5000 359.8400 ;
        RECT 2131.9000 364.8000 2133.5000 365.2800 ;
        RECT 2131.9000 370.2400 2133.5000 370.7200 ;
        RECT 2086.9000 375.6800 2088.5000 376.1600 ;
        RECT 2086.9000 381.1200 2088.5000 381.6000 ;
        RECT 2086.9000 359.3600 2088.5000 359.8400 ;
        RECT 2086.9000 364.8000 2088.5000 365.2800 ;
        RECT 2086.9000 370.2400 2088.5000 370.7200 ;
        RECT 2037.3400 402.8800 2040.3400 403.3600 ;
        RECT 2037.3400 408.3200 2040.3400 408.8000 ;
        RECT 2037.3400 392.0000 2040.3400 392.4800 ;
        RECT 2037.3400 386.5600 2040.3400 387.0400 ;
        RECT 2037.3400 397.4400 2040.3400 397.9200 ;
        RECT 2037.3400 375.6800 2040.3400 376.1600 ;
        RECT 2037.3400 381.1200 2040.3400 381.6000 ;
        RECT 2037.3400 364.8000 2040.3400 365.2800 ;
        RECT 2037.3400 359.3600 2040.3400 359.8400 ;
        RECT 2037.3400 370.2400 2040.3400 370.7200 ;
        RECT 2131.9000 348.4800 2133.5000 348.9600 ;
        RECT 2131.9000 353.9200 2133.5000 354.4000 ;
        RECT 2131.9000 332.1600 2133.5000 332.6400 ;
        RECT 2131.9000 337.6000 2133.5000 338.0800 ;
        RECT 2131.9000 343.0400 2133.5000 343.5200 ;
        RECT 2086.9000 348.4800 2088.5000 348.9600 ;
        RECT 2086.9000 353.9200 2088.5000 354.4000 ;
        RECT 2086.9000 332.1600 2088.5000 332.6400 ;
        RECT 2086.9000 337.6000 2088.5000 338.0800 ;
        RECT 2086.9000 343.0400 2088.5000 343.5200 ;
        RECT 2131.9000 326.7200 2133.5000 327.2000 ;
        RECT 2131.9000 321.2800 2133.5000 321.7600 ;
        RECT 2131.9000 315.8400 2133.5000 316.3200 ;
        RECT 2086.9000 326.7200 2088.5000 327.2000 ;
        RECT 2086.9000 321.2800 2088.5000 321.7600 ;
        RECT 2086.9000 315.8400 2088.5000 316.3200 ;
        RECT 2037.3400 348.4800 2040.3400 348.9600 ;
        RECT 2037.3400 353.9200 2040.3400 354.4000 ;
        RECT 2037.3400 337.6000 2040.3400 338.0800 ;
        RECT 2037.3400 332.1600 2040.3400 332.6400 ;
        RECT 2037.3400 343.0400 2040.3400 343.5200 ;
        RECT 2037.3400 321.2800 2040.3400 321.7600 ;
        RECT 2037.3400 326.7200 2040.3400 327.2000 ;
        RECT 2037.3400 315.8400 2040.3400 316.3200 ;
        RECT 2037.3400 514.0300 2236.4400 517.0300 ;
        RECT 2037.3400 308.9300 2236.4400 311.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 79.2900 2223.5000 287.3900 ;
        RECT 2176.9000 79.2900 2178.5000 287.3900 ;
        RECT 2131.9000 79.2900 2133.5000 287.3900 ;
        RECT 2086.9000 79.2900 2088.5000 287.3900 ;
        RECT 2233.4400 79.2900 2236.4400 287.3900 ;
        RECT 2037.3400 79.2900 2040.3400 287.3900 ;
      LAYER met3 ;
        RECT 2233.4400 282.0400 2236.4400 282.5200 ;
        RECT 2221.9000 282.0400 2223.5000 282.5200 ;
        RECT 2233.4400 271.1600 2236.4400 271.6400 ;
        RECT 2233.4400 276.6000 2236.4400 277.0800 ;
        RECT 2221.9000 271.1600 2223.5000 271.6400 ;
        RECT 2221.9000 276.6000 2223.5000 277.0800 ;
        RECT 2233.4400 254.8400 2236.4400 255.3200 ;
        RECT 2233.4400 260.2800 2236.4400 260.7600 ;
        RECT 2221.9000 254.8400 2223.5000 255.3200 ;
        RECT 2221.9000 260.2800 2223.5000 260.7600 ;
        RECT 2233.4400 243.9600 2236.4400 244.4400 ;
        RECT 2233.4400 249.4000 2236.4400 249.8800 ;
        RECT 2221.9000 243.9600 2223.5000 244.4400 ;
        RECT 2221.9000 249.4000 2223.5000 249.8800 ;
        RECT 2233.4400 265.7200 2236.4400 266.2000 ;
        RECT 2221.9000 265.7200 2223.5000 266.2000 ;
        RECT 2176.9000 271.1600 2178.5000 271.6400 ;
        RECT 2176.9000 276.6000 2178.5000 277.0800 ;
        RECT 2176.9000 282.0400 2178.5000 282.5200 ;
        RECT 2176.9000 254.8400 2178.5000 255.3200 ;
        RECT 2176.9000 260.2800 2178.5000 260.7600 ;
        RECT 2176.9000 249.4000 2178.5000 249.8800 ;
        RECT 2176.9000 243.9600 2178.5000 244.4400 ;
        RECT 2176.9000 265.7200 2178.5000 266.2000 ;
        RECT 2233.4400 227.6400 2236.4400 228.1200 ;
        RECT 2233.4400 233.0800 2236.4400 233.5600 ;
        RECT 2221.9000 227.6400 2223.5000 228.1200 ;
        RECT 2221.9000 233.0800 2223.5000 233.5600 ;
        RECT 2233.4400 211.3200 2236.4400 211.8000 ;
        RECT 2233.4400 216.7600 2236.4400 217.2400 ;
        RECT 2233.4400 222.2000 2236.4400 222.6800 ;
        RECT 2221.9000 211.3200 2223.5000 211.8000 ;
        RECT 2221.9000 216.7600 2223.5000 217.2400 ;
        RECT 2221.9000 222.2000 2223.5000 222.6800 ;
        RECT 2233.4400 200.4400 2236.4400 200.9200 ;
        RECT 2233.4400 205.8800 2236.4400 206.3600 ;
        RECT 2221.9000 200.4400 2223.5000 200.9200 ;
        RECT 2221.9000 205.8800 2223.5000 206.3600 ;
        RECT 2233.4400 184.1200 2236.4400 184.6000 ;
        RECT 2233.4400 189.5600 2236.4400 190.0400 ;
        RECT 2233.4400 195.0000 2236.4400 195.4800 ;
        RECT 2221.9000 184.1200 2223.5000 184.6000 ;
        RECT 2221.9000 189.5600 2223.5000 190.0400 ;
        RECT 2221.9000 195.0000 2223.5000 195.4800 ;
        RECT 2176.9000 227.6400 2178.5000 228.1200 ;
        RECT 2176.9000 233.0800 2178.5000 233.5600 ;
        RECT 2176.9000 211.3200 2178.5000 211.8000 ;
        RECT 2176.9000 216.7600 2178.5000 217.2400 ;
        RECT 2176.9000 222.2000 2178.5000 222.6800 ;
        RECT 2176.9000 200.4400 2178.5000 200.9200 ;
        RECT 2176.9000 205.8800 2178.5000 206.3600 ;
        RECT 2176.9000 184.1200 2178.5000 184.6000 ;
        RECT 2176.9000 189.5600 2178.5000 190.0400 ;
        RECT 2176.9000 195.0000 2178.5000 195.4800 ;
        RECT 2233.4400 238.5200 2236.4400 239.0000 ;
        RECT 2176.9000 238.5200 2178.5000 239.0000 ;
        RECT 2221.9000 238.5200 2223.5000 239.0000 ;
        RECT 2131.9000 271.1600 2133.5000 271.6400 ;
        RECT 2131.9000 276.6000 2133.5000 277.0800 ;
        RECT 2131.9000 282.0400 2133.5000 282.5200 ;
        RECT 2086.9000 271.1600 2088.5000 271.6400 ;
        RECT 2086.9000 276.6000 2088.5000 277.0800 ;
        RECT 2086.9000 282.0400 2088.5000 282.5200 ;
        RECT 2131.9000 254.8400 2133.5000 255.3200 ;
        RECT 2131.9000 260.2800 2133.5000 260.7600 ;
        RECT 2131.9000 243.9600 2133.5000 244.4400 ;
        RECT 2131.9000 249.4000 2133.5000 249.8800 ;
        RECT 2086.9000 254.8400 2088.5000 255.3200 ;
        RECT 2086.9000 260.2800 2088.5000 260.7600 ;
        RECT 2086.9000 243.9600 2088.5000 244.4400 ;
        RECT 2086.9000 249.4000 2088.5000 249.8800 ;
        RECT 2086.9000 265.7200 2088.5000 266.2000 ;
        RECT 2131.9000 265.7200 2133.5000 266.2000 ;
        RECT 2037.3400 282.0400 2040.3400 282.5200 ;
        RECT 2037.3400 276.6000 2040.3400 277.0800 ;
        RECT 2037.3400 271.1600 2040.3400 271.6400 ;
        RECT 2037.3400 260.2800 2040.3400 260.7600 ;
        RECT 2037.3400 254.8400 2040.3400 255.3200 ;
        RECT 2037.3400 249.4000 2040.3400 249.8800 ;
        RECT 2037.3400 243.9600 2040.3400 244.4400 ;
        RECT 2037.3400 265.7200 2040.3400 266.2000 ;
        RECT 2131.9000 227.6400 2133.5000 228.1200 ;
        RECT 2131.9000 233.0800 2133.5000 233.5600 ;
        RECT 2131.9000 211.3200 2133.5000 211.8000 ;
        RECT 2131.9000 216.7600 2133.5000 217.2400 ;
        RECT 2131.9000 222.2000 2133.5000 222.6800 ;
        RECT 2086.9000 227.6400 2088.5000 228.1200 ;
        RECT 2086.9000 233.0800 2088.5000 233.5600 ;
        RECT 2086.9000 211.3200 2088.5000 211.8000 ;
        RECT 2086.9000 216.7600 2088.5000 217.2400 ;
        RECT 2086.9000 222.2000 2088.5000 222.6800 ;
        RECT 2131.9000 200.4400 2133.5000 200.9200 ;
        RECT 2131.9000 205.8800 2133.5000 206.3600 ;
        RECT 2131.9000 184.1200 2133.5000 184.6000 ;
        RECT 2131.9000 189.5600 2133.5000 190.0400 ;
        RECT 2131.9000 195.0000 2133.5000 195.4800 ;
        RECT 2086.9000 200.4400 2088.5000 200.9200 ;
        RECT 2086.9000 205.8800 2088.5000 206.3600 ;
        RECT 2086.9000 184.1200 2088.5000 184.6000 ;
        RECT 2086.9000 189.5600 2088.5000 190.0400 ;
        RECT 2086.9000 195.0000 2088.5000 195.4800 ;
        RECT 2037.3400 227.6400 2040.3400 228.1200 ;
        RECT 2037.3400 233.0800 2040.3400 233.5600 ;
        RECT 2037.3400 216.7600 2040.3400 217.2400 ;
        RECT 2037.3400 211.3200 2040.3400 211.8000 ;
        RECT 2037.3400 222.2000 2040.3400 222.6800 ;
        RECT 2037.3400 200.4400 2040.3400 200.9200 ;
        RECT 2037.3400 205.8800 2040.3400 206.3600 ;
        RECT 2037.3400 189.5600 2040.3400 190.0400 ;
        RECT 2037.3400 184.1200 2040.3400 184.6000 ;
        RECT 2037.3400 195.0000 2040.3400 195.4800 ;
        RECT 2037.3400 238.5200 2040.3400 239.0000 ;
        RECT 2086.9000 238.5200 2088.5000 239.0000 ;
        RECT 2131.9000 238.5200 2133.5000 239.0000 ;
        RECT 2233.4400 173.2400 2236.4400 173.7200 ;
        RECT 2233.4400 178.6800 2236.4400 179.1600 ;
        RECT 2221.9000 173.2400 2223.5000 173.7200 ;
        RECT 2221.9000 178.6800 2223.5000 179.1600 ;
        RECT 2233.4400 156.9200 2236.4400 157.4000 ;
        RECT 2233.4400 162.3600 2236.4400 162.8400 ;
        RECT 2233.4400 167.8000 2236.4400 168.2800 ;
        RECT 2221.9000 156.9200 2223.5000 157.4000 ;
        RECT 2221.9000 162.3600 2223.5000 162.8400 ;
        RECT 2221.9000 167.8000 2223.5000 168.2800 ;
        RECT 2233.4400 146.0400 2236.4400 146.5200 ;
        RECT 2233.4400 151.4800 2236.4400 151.9600 ;
        RECT 2221.9000 146.0400 2223.5000 146.5200 ;
        RECT 2221.9000 151.4800 2223.5000 151.9600 ;
        RECT 2233.4400 129.7200 2236.4400 130.2000 ;
        RECT 2233.4400 135.1600 2236.4400 135.6400 ;
        RECT 2233.4400 140.6000 2236.4400 141.0800 ;
        RECT 2221.9000 129.7200 2223.5000 130.2000 ;
        RECT 2221.9000 135.1600 2223.5000 135.6400 ;
        RECT 2221.9000 140.6000 2223.5000 141.0800 ;
        RECT 2176.9000 173.2400 2178.5000 173.7200 ;
        RECT 2176.9000 178.6800 2178.5000 179.1600 ;
        RECT 2176.9000 156.9200 2178.5000 157.4000 ;
        RECT 2176.9000 162.3600 2178.5000 162.8400 ;
        RECT 2176.9000 167.8000 2178.5000 168.2800 ;
        RECT 2176.9000 146.0400 2178.5000 146.5200 ;
        RECT 2176.9000 151.4800 2178.5000 151.9600 ;
        RECT 2176.9000 129.7200 2178.5000 130.2000 ;
        RECT 2176.9000 135.1600 2178.5000 135.6400 ;
        RECT 2176.9000 140.6000 2178.5000 141.0800 ;
        RECT 2233.4400 118.8400 2236.4400 119.3200 ;
        RECT 2233.4400 124.2800 2236.4400 124.7600 ;
        RECT 2221.9000 118.8400 2223.5000 119.3200 ;
        RECT 2221.9000 124.2800 2223.5000 124.7600 ;
        RECT 2233.4400 102.5200 2236.4400 103.0000 ;
        RECT 2233.4400 107.9600 2236.4400 108.4400 ;
        RECT 2233.4400 113.4000 2236.4400 113.8800 ;
        RECT 2221.9000 102.5200 2223.5000 103.0000 ;
        RECT 2221.9000 107.9600 2223.5000 108.4400 ;
        RECT 2221.9000 113.4000 2223.5000 113.8800 ;
        RECT 2233.4400 91.6400 2236.4400 92.1200 ;
        RECT 2233.4400 97.0800 2236.4400 97.5600 ;
        RECT 2221.9000 91.6400 2223.5000 92.1200 ;
        RECT 2221.9000 97.0800 2223.5000 97.5600 ;
        RECT 2233.4400 86.2000 2236.4400 86.6800 ;
        RECT 2221.9000 86.2000 2223.5000 86.6800 ;
        RECT 2176.9000 118.8400 2178.5000 119.3200 ;
        RECT 2176.9000 124.2800 2178.5000 124.7600 ;
        RECT 2176.9000 102.5200 2178.5000 103.0000 ;
        RECT 2176.9000 107.9600 2178.5000 108.4400 ;
        RECT 2176.9000 113.4000 2178.5000 113.8800 ;
        RECT 2176.9000 91.6400 2178.5000 92.1200 ;
        RECT 2176.9000 97.0800 2178.5000 97.5600 ;
        RECT 2176.9000 86.2000 2178.5000 86.6800 ;
        RECT 2131.9000 173.2400 2133.5000 173.7200 ;
        RECT 2131.9000 178.6800 2133.5000 179.1600 ;
        RECT 2131.9000 156.9200 2133.5000 157.4000 ;
        RECT 2131.9000 162.3600 2133.5000 162.8400 ;
        RECT 2131.9000 167.8000 2133.5000 168.2800 ;
        RECT 2086.9000 173.2400 2088.5000 173.7200 ;
        RECT 2086.9000 178.6800 2088.5000 179.1600 ;
        RECT 2086.9000 156.9200 2088.5000 157.4000 ;
        RECT 2086.9000 162.3600 2088.5000 162.8400 ;
        RECT 2086.9000 167.8000 2088.5000 168.2800 ;
        RECT 2131.9000 146.0400 2133.5000 146.5200 ;
        RECT 2131.9000 151.4800 2133.5000 151.9600 ;
        RECT 2131.9000 129.7200 2133.5000 130.2000 ;
        RECT 2131.9000 135.1600 2133.5000 135.6400 ;
        RECT 2131.9000 140.6000 2133.5000 141.0800 ;
        RECT 2086.9000 146.0400 2088.5000 146.5200 ;
        RECT 2086.9000 151.4800 2088.5000 151.9600 ;
        RECT 2086.9000 129.7200 2088.5000 130.2000 ;
        RECT 2086.9000 135.1600 2088.5000 135.6400 ;
        RECT 2086.9000 140.6000 2088.5000 141.0800 ;
        RECT 2037.3400 173.2400 2040.3400 173.7200 ;
        RECT 2037.3400 178.6800 2040.3400 179.1600 ;
        RECT 2037.3400 162.3600 2040.3400 162.8400 ;
        RECT 2037.3400 156.9200 2040.3400 157.4000 ;
        RECT 2037.3400 167.8000 2040.3400 168.2800 ;
        RECT 2037.3400 146.0400 2040.3400 146.5200 ;
        RECT 2037.3400 151.4800 2040.3400 151.9600 ;
        RECT 2037.3400 135.1600 2040.3400 135.6400 ;
        RECT 2037.3400 129.7200 2040.3400 130.2000 ;
        RECT 2037.3400 140.6000 2040.3400 141.0800 ;
        RECT 2131.9000 118.8400 2133.5000 119.3200 ;
        RECT 2131.9000 124.2800 2133.5000 124.7600 ;
        RECT 2131.9000 102.5200 2133.5000 103.0000 ;
        RECT 2131.9000 107.9600 2133.5000 108.4400 ;
        RECT 2131.9000 113.4000 2133.5000 113.8800 ;
        RECT 2086.9000 118.8400 2088.5000 119.3200 ;
        RECT 2086.9000 124.2800 2088.5000 124.7600 ;
        RECT 2086.9000 102.5200 2088.5000 103.0000 ;
        RECT 2086.9000 107.9600 2088.5000 108.4400 ;
        RECT 2086.9000 113.4000 2088.5000 113.8800 ;
        RECT 2131.9000 97.0800 2133.5000 97.5600 ;
        RECT 2131.9000 91.6400 2133.5000 92.1200 ;
        RECT 2131.9000 86.2000 2133.5000 86.6800 ;
        RECT 2086.9000 97.0800 2088.5000 97.5600 ;
        RECT 2086.9000 91.6400 2088.5000 92.1200 ;
        RECT 2086.9000 86.2000 2088.5000 86.6800 ;
        RECT 2037.3400 118.8400 2040.3400 119.3200 ;
        RECT 2037.3400 124.2800 2040.3400 124.7600 ;
        RECT 2037.3400 107.9600 2040.3400 108.4400 ;
        RECT 2037.3400 102.5200 2040.3400 103.0000 ;
        RECT 2037.3400 113.4000 2040.3400 113.8800 ;
        RECT 2037.3400 91.6400 2040.3400 92.1200 ;
        RECT 2037.3400 97.0800 2040.3400 97.5600 ;
        RECT 2037.3400 86.2000 2040.3400 86.6800 ;
        RECT 2037.3400 284.3900 2236.4400 287.3900 ;
        RECT 2037.3400 79.2900 2236.4400 82.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 2037.3400 37.6700 2039.3400 58.6000 ;
        RECT 2234.4400 37.6700 2236.4400 58.6000 ;
      LAYER met3 ;
        RECT 2234.4400 54.1000 2236.4400 54.5800 ;
        RECT 2037.3400 54.1000 2039.3400 54.5800 ;
        RECT 2234.4400 43.2200 2236.4400 43.7000 ;
        RECT 2037.3400 43.2200 2039.3400 43.7000 ;
        RECT 2234.4400 48.6600 2236.4400 49.1400 ;
        RECT 2037.3400 48.6600 2039.3400 49.1400 ;
        RECT 2037.3400 56.6000 2236.4400 58.6000 ;
        RECT 2037.3400 37.6700 2236.4400 39.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 2605.3300 2223.5000 2813.4300 ;
        RECT 2176.9000 2605.3300 2178.5000 2813.4300 ;
        RECT 2131.9000 2605.3300 2133.5000 2813.4300 ;
        RECT 2086.9000 2605.3300 2088.5000 2813.4300 ;
        RECT 2233.4400 2605.3300 2236.4400 2813.4300 ;
        RECT 2037.3400 2605.3300 2040.3400 2813.4300 ;
      LAYER met3 ;
        RECT 2233.4400 2808.0800 2236.4400 2808.5600 ;
        RECT 2221.9000 2808.0800 2223.5000 2808.5600 ;
        RECT 2233.4400 2797.2000 2236.4400 2797.6800 ;
        RECT 2233.4400 2802.6400 2236.4400 2803.1200 ;
        RECT 2221.9000 2797.2000 2223.5000 2797.6800 ;
        RECT 2221.9000 2802.6400 2223.5000 2803.1200 ;
        RECT 2233.4400 2780.8800 2236.4400 2781.3600 ;
        RECT 2233.4400 2786.3200 2236.4400 2786.8000 ;
        RECT 2221.9000 2780.8800 2223.5000 2781.3600 ;
        RECT 2221.9000 2786.3200 2223.5000 2786.8000 ;
        RECT 2233.4400 2770.0000 2236.4400 2770.4800 ;
        RECT 2233.4400 2775.4400 2236.4400 2775.9200 ;
        RECT 2221.9000 2770.0000 2223.5000 2770.4800 ;
        RECT 2221.9000 2775.4400 2223.5000 2775.9200 ;
        RECT 2233.4400 2791.7600 2236.4400 2792.2400 ;
        RECT 2221.9000 2791.7600 2223.5000 2792.2400 ;
        RECT 2176.9000 2797.2000 2178.5000 2797.6800 ;
        RECT 2176.9000 2802.6400 2178.5000 2803.1200 ;
        RECT 2176.9000 2808.0800 2178.5000 2808.5600 ;
        RECT 2176.9000 2780.8800 2178.5000 2781.3600 ;
        RECT 2176.9000 2786.3200 2178.5000 2786.8000 ;
        RECT 2176.9000 2775.4400 2178.5000 2775.9200 ;
        RECT 2176.9000 2770.0000 2178.5000 2770.4800 ;
        RECT 2176.9000 2791.7600 2178.5000 2792.2400 ;
        RECT 2233.4400 2753.6800 2236.4400 2754.1600 ;
        RECT 2233.4400 2759.1200 2236.4400 2759.6000 ;
        RECT 2221.9000 2753.6800 2223.5000 2754.1600 ;
        RECT 2221.9000 2759.1200 2223.5000 2759.6000 ;
        RECT 2233.4400 2737.3600 2236.4400 2737.8400 ;
        RECT 2233.4400 2742.8000 2236.4400 2743.2800 ;
        RECT 2233.4400 2748.2400 2236.4400 2748.7200 ;
        RECT 2221.9000 2737.3600 2223.5000 2737.8400 ;
        RECT 2221.9000 2742.8000 2223.5000 2743.2800 ;
        RECT 2221.9000 2748.2400 2223.5000 2748.7200 ;
        RECT 2233.4400 2726.4800 2236.4400 2726.9600 ;
        RECT 2233.4400 2731.9200 2236.4400 2732.4000 ;
        RECT 2221.9000 2726.4800 2223.5000 2726.9600 ;
        RECT 2221.9000 2731.9200 2223.5000 2732.4000 ;
        RECT 2233.4400 2710.1600 2236.4400 2710.6400 ;
        RECT 2233.4400 2715.6000 2236.4400 2716.0800 ;
        RECT 2233.4400 2721.0400 2236.4400 2721.5200 ;
        RECT 2221.9000 2710.1600 2223.5000 2710.6400 ;
        RECT 2221.9000 2715.6000 2223.5000 2716.0800 ;
        RECT 2221.9000 2721.0400 2223.5000 2721.5200 ;
        RECT 2176.9000 2753.6800 2178.5000 2754.1600 ;
        RECT 2176.9000 2759.1200 2178.5000 2759.6000 ;
        RECT 2176.9000 2737.3600 2178.5000 2737.8400 ;
        RECT 2176.9000 2742.8000 2178.5000 2743.2800 ;
        RECT 2176.9000 2748.2400 2178.5000 2748.7200 ;
        RECT 2176.9000 2726.4800 2178.5000 2726.9600 ;
        RECT 2176.9000 2731.9200 2178.5000 2732.4000 ;
        RECT 2176.9000 2710.1600 2178.5000 2710.6400 ;
        RECT 2176.9000 2715.6000 2178.5000 2716.0800 ;
        RECT 2176.9000 2721.0400 2178.5000 2721.5200 ;
        RECT 2233.4400 2764.5600 2236.4400 2765.0400 ;
        RECT 2176.9000 2764.5600 2178.5000 2765.0400 ;
        RECT 2221.9000 2764.5600 2223.5000 2765.0400 ;
        RECT 2131.9000 2797.2000 2133.5000 2797.6800 ;
        RECT 2131.9000 2802.6400 2133.5000 2803.1200 ;
        RECT 2131.9000 2808.0800 2133.5000 2808.5600 ;
        RECT 2086.9000 2797.2000 2088.5000 2797.6800 ;
        RECT 2086.9000 2802.6400 2088.5000 2803.1200 ;
        RECT 2086.9000 2808.0800 2088.5000 2808.5600 ;
        RECT 2131.9000 2780.8800 2133.5000 2781.3600 ;
        RECT 2131.9000 2786.3200 2133.5000 2786.8000 ;
        RECT 2131.9000 2770.0000 2133.5000 2770.4800 ;
        RECT 2131.9000 2775.4400 2133.5000 2775.9200 ;
        RECT 2086.9000 2780.8800 2088.5000 2781.3600 ;
        RECT 2086.9000 2786.3200 2088.5000 2786.8000 ;
        RECT 2086.9000 2770.0000 2088.5000 2770.4800 ;
        RECT 2086.9000 2775.4400 2088.5000 2775.9200 ;
        RECT 2086.9000 2791.7600 2088.5000 2792.2400 ;
        RECT 2131.9000 2791.7600 2133.5000 2792.2400 ;
        RECT 2037.3400 2808.0800 2040.3400 2808.5600 ;
        RECT 2037.3400 2802.6400 2040.3400 2803.1200 ;
        RECT 2037.3400 2797.2000 2040.3400 2797.6800 ;
        RECT 2037.3400 2786.3200 2040.3400 2786.8000 ;
        RECT 2037.3400 2780.8800 2040.3400 2781.3600 ;
        RECT 2037.3400 2775.4400 2040.3400 2775.9200 ;
        RECT 2037.3400 2770.0000 2040.3400 2770.4800 ;
        RECT 2037.3400 2791.7600 2040.3400 2792.2400 ;
        RECT 2131.9000 2753.6800 2133.5000 2754.1600 ;
        RECT 2131.9000 2759.1200 2133.5000 2759.6000 ;
        RECT 2131.9000 2737.3600 2133.5000 2737.8400 ;
        RECT 2131.9000 2742.8000 2133.5000 2743.2800 ;
        RECT 2131.9000 2748.2400 2133.5000 2748.7200 ;
        RECT 2086.9000 2753.6800 2088.5000 2754.1600 ;
        RECT 2086.9000 2759.1200 2088.5000 2759.6000 ;
        RECT 2086.9000 2737.3600 2088.5000 2737.8400 ;
        RECT 2086.9000 2742.8000 2088.5000 2743.2800 ;
        RECT 2086.9000 2748.2400 2088.5000 2748.7200 ;
        RECT 2131.9000 2726.4800 2133.5000 2726.9600 ;
        RECT 2131.9000 2731.9200 2133.5000 2732.4000 ;
        RECT 2131.9000 2710.1600 2133.5000 2710.6400 ;
        RECT 2131.9000 2715.6000 2133.5000 2716.0800 ;
        RECT 2131.9000 2721.0400 2133.5000 2721.5200 ;
        RECT 2086.9000 2726.4800 2088.5000 2726.9600 ;
        RECT 2086.9000 2731.9200 2088.5000 2732.4000 ;
        RECT 2086.9000 2710.1600 2088.5000 2710.6400 ;
        RECT 2086.9000 2715.6000 2088.5000 2716.0800 ;
        RECT 2086.9000 2721.0400 2088.5000 2721.5200 ;
        RECT 2037.3400 2753.6800 2040.3400 2754.1600 ;
        RECT 2037.3400 2759.1200 2040.3400 2759.6000 ;
        RECT 2037.3400 2742.8000 2040.3400 2743.2800 ;
        RECT 2037.3400 2737.3600 2040.3400 2737.8400 ;
        RECT 2037.3400 2748.2400 2040.3400 2748.7200 ;
        RECT 2037.3400 2726.4800 2040.3400 2726.9600 ;
        RECT 2037.3400 2731.9200 2040.3400 2732.4000 ;
        RECT 2037.3400 2715.6000 2040.3400 2716.0800 ;
        RECT 2037.3400 2710.1600 2040.3400 2710.6400 ;
        RECT 2037.3400 2721.0400 2040.3400 2721.5200 ;
        RECT 2037.3400 2764.5600 2040.3400 2765.0400 ;
        RECT 2086.9000 2764.5600 2088.5000 2765.0400 ;
        RECT 2131.9000 2764.5600 2133.5000 2765.0400 ;
        RECT 2233.4400 2699.2800 2236.4400 2699.7600 ;
        RECT 2233.4400 2704.7200 2236.4400 2705.2000 ;
        RECT 2221.9000 2699.2800 2223.5000 2699.7600 ;
        RECT 2221.9000 2704.7200 2223.5000 2705.2000 ;
        RECT 2233.4400 2682.9600 2236.4400 2683.4400 ;
        RECT 2233.4400 2688.4000 2236.4400 2688.8800 ;
        RECT 2233.4400 2693.8400 2236.4400 2694.3200 ;
        RECT 2221.9000 2682.9600 2223.5000 2683.4400 ;
        RECT 2221.9000 2688.4000 2223.5000 2688.8800 ;
        RECT 2221.9000 2693.8400 2223.5000 2694.3200 ;
        RECT 2233.4400 2672.0800 2236.4400 2672.5600 ;
        RECT 2233.4400 2677.5200 2236.4400 2678.0000 ;
        RECT 2221.9000 2672.0800 2223.5000 2672.5600 ;
        RECT 2221.9000 2677.5200 2223.5000 2678.0000 ;
        RECT 2233.4400 2655.7600 2236.4400 2656.2400 ;
        RECT 2233.4400 2661.2000 2236.4400 2661.6800 ;
        RECT 2233.4400 2666.6400 2236.4400 2667.1200 ;
        RECT 2221.9000 2655.7600 2223.5000 2656.2400 ;
        RECT 2221.9000 2661.2000 2223.5000 2661.6800 ;
        RECT 2221.9000 2666.6400 2223.5000 2667.1200 ;
        RECT 2176.9000 2699.2800 2178.5000 2699.7600 ;
        RECT 2176.9000 2704.7200 2178.5000 2705.2000 ;
        RECT 2176.9000 2682.9600 2178.5000 2683.4400 ;
        RECT 2176.9000 2688.4000 2178.5000 2688.8800 ;
        RECT 2176.9000 2693.8400 2178.5000 2694.3200 ;
        RECT 2176.9000 2672.0800 2178.5000 2672.5600 ;
        RECT 2176.9000 2677.5200 2178.5000 2678.0000 ;
        RECT 2176.9000 2655.7600 2178.5000 2656.2400 ;
        RECT 2176.9000 2661.2000 2178.5000 2661.6800 ;
        RECT 2176.9000 2666.6400 2178.5000 2667.1200 ;
        RECT 2233.4400 2644.8800 2236.4400 2645.3600 ;
        RECT 2233.4400 2650.3200 2236.4400 2650.8000 ;
        RECT 2221.9000 2644.8800 2223.5000 2645.3600 ;
        RECT 2221.9000 2650.3200 2223.5000 2650.8000 ;
        RECT 2233.4400 2628.5600 2236.4400 2629.0400 ;
        RECT 2233.4400 2634.0000 2236.4400 2634.4800 ;
        RECT 2233.4400 2639.4400 2236.4400 2639.9200 ;
        RECT 2221.9000 2628.5600 2223.5000 2629.0400 ;
        RECT 2221.9000 2634.0000 2223.5000 2634.4800 ;
        RECT 2221.9000 2639.4400 2223.5000 2639.9200 ;
        RECT 2233.4400 2617.6800 2236.4400 2618.1600 ;
        RECT 2233.4400 2623.1200 2236.4400 2623.6000 ;
        RECT 2221.9000 2617.6800 2223.5000 2618.1600 ;
        RECT 2221.9000 2623.1200 2223.5000 2623.6000 ;
        RECT 2233.4400 2612.2400 2236.4400 2612.7200 ;
        RECT 2221.9000 2612.2400 2223.5000 2612.7200 ;
        RECT 2176.9000 2644.8800 2178.5000 2645.3600 ;
        RECT 2176.9000 2650.3200 2178.5000 2650.8000 ;
        RECT 2176.9000 2628.5600 2178.5000 2629.0400 ;
        RECT 2176.9000 2634.0000 2178.5000 2634.4800 ;
        RECT 2176.9000 2639.4400 2178.5000 2639.9200 ;
        RECT 2176.9000 2617.6800 2178.5000 2618.1600 ;
        RECT 2176.9000 2623.1200 2178.5000 2623.6000 ;
        RECT 2176.9000 2612.2400 2178.5000 2612.7200 ;
        RECT 2131.9000 2699.2800 2133.5000 2699.7600 ;
        RECT 2131.9000 2704.7200 2133.5000 2705.2000 ;
        RECT 2131.9000 2682.9600 2133.5000 2683.4400 ;
        RECT 2131.9000 2688.4000 2133.5000 2688.8800 ;
        RECT 2131.9000 2693.8400 2133.5000 2694.3200 ;
        RECT 2086.9000 2699.2800 2088.5000 2699.7600 ;
        RECT 2086.9000 2704.7200 2088.5000 2705.2000 ;
        RECT 2086.9000 2682.9600 2088.5000 2683.4400 ;
        RECT 2086.9000 2688.4000 2088.5000 2688.8800 ;
        RECT 2086.9000 2693.8400 2088.5000 2694.3200 ;
        RECT 2131.9000 2672.0800 2133.5000 2672.5600 ;
        RECT 2131.9000 2677.5200 2133.5000 2678.0000 ;
        RECT 2131.9000 2655.7600 2133.5000 2656.2400 ;
        RECT 2131.9000 2661.2000 2133.5000 2661.6800 ;
        RECT 2131.9000 2666.6400 2133.5000 2667.1200 ;
        RECT 2086.9000 2672.0800 2088.5000 2672.5600 ;
        RECT 2086.9000 2677.5200 2088.5000 2678.0000 ;
        RECT 2086.9000 2655.7600 2088.5000 2656.2400 ;
        RECT 2086.9000 2661.2000 2088.5000 2661.6800 ;
        RECT 2086.9000 2666.6400 2088.5000 2667.1200 ;
        RECT 2037.3400 2699.2800 2040.3400 2699.7600 ;
        RECT 2037.3400 2704.7200 2040.3400 2705.2000 ;
        RECT 2037.3400 2688.4000 2040.3400 2688.8800 ;
        RECT 2037.3400 2682.9600 2040.3400 2683.4400 ;
        RECT 2037.3400 2693.8400 2040.3400 2694.3200 ;
        RECT 2037.3400 2672.0800 2040.3400 2672.5600 ;
        RECT 2037.3400 2677.5200 2040.3400 2678.0000 ;
        RECT 2037.3400 2661.2000 2040.3400 2661.6800 ;
        RECT 2037.3400 2655.7600 2040.3400 2656.2400 ;
        RECT 2037.3400 2666.6400 2040.3400 2667.1200 ;
        RECT 2131.9000 2644.8800 2133.5000 2645.3600 ;
        RECT 2131.9000 2650.3200 2133.5000 2650.8000 ;
        RECT 2131.9000 2628.5600 2133.5000 2629.0400 ;
        RECT 2131.9000 2634.0000 2133.5000 2634.4800 ;
        RECT 2131.9000 2639.4400 2133.5000 2639.9200 ;
        RECT 2086.9000 2644.8800 2088.5000 2645.3600 ;
        RECT 2086.9000 2650.3200 2088.5000 2650.8000 ;
        RECT 2086.9000 2628.5600 2088.5000 2629.0400 ;
        RECT 2086.9000 2634.0000 2088.5000 2634.4800 ;
        RECT 2086.9000 2639.4400 2088.5000 2639.9200 ;
        RECT 2131.9000 2623.1200 2133.5000 2623.6000 ;
        RECT 2131.9000 2617.6800 2133.5000 2618.1600 ;
        RECT 2131.9000 2612.2400 2133.5000 2612.7200 ;
        RECT 2086.9000 2623.1200 2088.5000 2623.6000 ;
        RECT 2086.9000 2617.6800 2088.5000 2618.1600 ;
        RECT 2086.9000 2612.2400 2088.5000 2612.7200 ;
        RECT 2037.3400 2644.8800 2040.3400 2645.3600 ;
        RECT 2037.3400 2650.3200 2040.3400 2650.8000 ;
        RECT 2037.3400 2634.0000 2040.3400 2634.4800 ;
        RECT 2037.3400 2628.5600 2040.3400 2629.0400 ;
        RECT 2037.3400 2639.4400 2040.3400 2639.9200 ;
        RECT 2037.3400 2617.6800 2040.3400 2618.1600 ;
        RECT 2037.3400 2623.1200 2040.3400 2623.6000 ;
        RECT 2037.3400 2612.2400 2040.3400 2612.7200 ;
        RECT 2037.3400 2810.4300 2236.4400 2813.4300 ;
        RECT 2037.3400 2605.3300 2236.4400 2608.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 2375.6900 2223.5000 2583.7900 ;
        RECT 2176.9000 2375.6900 2178.5000 2583.7900 ;
        RECT 2131.9000 2375.6900 2133.5000 2583.7900 ;
        RECT 2086.9000 2375.6900 2088.5000 2583.7900 ;
        RECT 2233.4400 2375.6900 2236.4400 2583.7900 ;
        RECT 2037.3400 2375.6900 2040.3400 2583.7900 ;
      LAYER met3 ;
        RECT 2233.4400 2578.4400 2236.4400 2578.9200 ;
        RECT 2221.9000 2578.4400 2223.5000 2578.9200 ;
        RECT 2233.4400 2567.5600 2236.4400 2568.0400 ;
        RECT 2233.4400 2573.0000 2236.4400 2573.4800 ;
        RECT 2221.9000 2567.5600 2223.5000 2568.0400 ;
        RECT 2221.9000 2573.0000 2223.5000 2573.4800 ;
        RECT 2233.4400 2551.2400 2236.4400 2551.7200 ;
        RECT 2233.4400 2556.6800 2236.4400 2557.1600 ;
        RECT 2221.9000 2551.2400 2223.5000 2551.7200 ;
        RECT 2221.9000 2556.6800 2223.5000 2557.1600 ;
        RECT 2233.4400 2540.3600 2236.4400 2540.8400 ;
        RECT 2233.4400 2545.8000 2236.4400 2546.2800 ;
        RECT 2221.9000 2540.3600 2223.5000 2540.8400 ;
        RECT 2221.9000 2545.8000 2223.5000 2546.2800 ;
        RECT 2233.4400 2562.1200 2236.4400 2562.6000 ;
        RECT 2221.9000 2562.1200 2223.5000 2562.6000 ;
        RECT 2176.9000 2567.5600 2178.5000 2568.0400 ;
        RECT 2176.9000 2573.0000 2178.5000 2573.4800 ;
        RECT 2176.9000 2578.4400 2178.5000 2578.9200 ;
        RECT 2176.9000 2551.2400 2178.5000 2551.7200 ;
        RECT 2176.9000 2556.6800 2178.5000 2557.1600 ;
        RECT 2176.9000 2545.8000 2178.5000 2546.2800 ;
        RECT 2176.9000 2540.3600 2178.5000 2540.8400 ;
        RECT 2176.9000 2562.1200 2178.5000 2562.6000 ;
        RECT 2233.4400 2524.0400 2236.4400 2524.5200 ;
        RECT 2233.4400 2529.4800 2236.4400 2529.9600 ;
        RECT 2221.9000 2524.0400 2223.5000 2524.5200 ;
        RECT 2221.9000 2529.4800 2223.5000 2529.9600 ;
        RECT 2233.4400 2507.7200 2236.4400 2508.2000 ;
        RECT 2233.4400 2513.1600 2236.4400 2513.6400 ;
        RECT 2233.4400 2518.6000 2236.4400 2519.0800 ;
        RECT 2221.9000 2507.7200 2223.5000 2508.2000 ;
        RECT 2221.9000 2513.1600 2223.5000 2513.6400 ;
        RECT 2221.9000 2518.6000 2223.5000 2519.0800 ;
        RECT 2233.4400 2496.8400 2236.4400 2497.3200 ;
        RECT 2233.4400 2502.2800 2236.4400 2502.7600 ;
        RECT 2221.9000 2496.8400 2223.5000 2497.3200 ;
        RECT 2221.9000 2502.2800 2223.5000 2502.7600 ;
        RECT 2233.4400 2480.5200 2236.4400 2481.0000 ;
        RECT 2233.4400 2485.9600 2236.4400 2486.4400 ;
        RECT 2233.4400 2491.4000 2236.4400 2491.8800 ;
        RECT 2221.9000 2480.5200 2223.5000 2481.0000 ;
        RECT 2221.9000 2485.9600 2223.5000 2486.4400 ;
        RECT 2221.9000 2491.4000 2223.5000 2491.8800 ;
        RECT 2176.9000 2524.0400 2178.5000 2524.5200 ;
        RECT 2176.9000 2529.4800 2178.5000 2529.9600 ;
        RECT 2176.9000 2507.7200 2178.5000 2508.2000 ;
        RECT 2176.9000 2513.1600 2178.5000 2513.6400 ;
        RECT 2176.9000 2518.6000 2178.5000 2519.0800 ;
        RECT 2176.9000 2496.8400 2178.5000 2497.3200 ;
        RECT 2176.9000 2502.2800 2178.5000 2502.7600 ;
        RECT 2176.9000 2480.5200 2178.5000 2481.0000 ;
        RECT 2176.9000 2485.9600 2178.5000 2486.4400 ;
        RECT 2176.9000 2491.4000 2178.5000 2491.8800 ;
        RECT 2233.4400 2534.9200 2236.4400 2535.4000 ;
        RECT 2176.9000 2534.9200 2178.5000 2535.4000 ;
        RECT 2221.9000 2534.9200 2223.5000 2535.4000 ;
        RECT 2131.9000 2567.5600 2133.5000 2568.0400 ;
        RECT 2131.9000 2573.0000 2133.5000 2573.4800 ;
        RECT 2131.9000 2578.4400 2133.5000 2578.9200 ;
        RECT 2086.9000 2567.5600 2088.5000 2568.0400 ;
        RECT 2086.9000 2573.0000 2088.5000 2573.4800 ;
        RECT 2086.9000 2578.4400 2088.5000 2578.9200 ;
        RECT 2131.9000 2551.2400 2133.5000 2551.7200 ;
        RECT 2131.9000 2556.6800 2133.5000 2557.1600 ;
        RECT 2131.9000 2540.3600 2133.5000 2540.8400 ;
        RECT 2131.9000 2545.8000 2133.5000 2546.2800 ;
        RECT 2086.9000 2551.2400 2088.5000 2551.7200 ;
        RECT 2086.9000 2556.6800 2088.5000 2557.1600 ;
        RECT 2086.9000 2540.3600 2088.5000 2540.8400 ;
        RECT 2086.9000 2545.8000 2088.5000 2546.2800 ;
        RECT 2086.9000 2562.1200 2088.5000 2562.6000 ;
        RECT 2131.9000 2562.1200 2133.5000 2562.6000 ;
        RECT 2037.3400 2578.4400 2040.3400 2578.9200 ;
        RECT 2037.3400 2573.0000 2040.3400 2573.4800 ;
        RECT 2037.3400 2567.5600 2040.3400 2568.0400 ;
        RECT 2037.3400 2556.6800 2040.3400 2557.1600 ;
        RECT 2037.3400 2551.2400 2040.3400 2551.7200 ;
        RECT 2037.3400 2545.8000 2040.3400 2546.2800 ;
        RECT 2037.3400 2540.3600 2040.3400 2540.8400 ;
        RECT 2037.3400 2562.1200 2040.3400 2562.6000 ;
        RECT 2131.9000 2524.0400 2133.5000 2524.5200 ;
        RECT 2131.9000 2529.4800 2133.5000 2529.9600 ;
        RECT 2131.9000 2507.7200 2133.5000 2508.2000 ;
        RECT 2131.9000 2513.1600 2133.5000 2513.6400 ;
        RECT 2131.9000 2518.6000 2133.5000 2519.0800 ;
        RECT 2086.9000 2524.0400 2088.5000 2524.5200 ;
        RECT 2086.9000 2529.4800 2088.5000 2529.9600 ;
        RECT 2086.9000 2507.7200 2088.5000 2508.2000 ;
        RECT 2086.9000 2513.1600 2088.5000 2513.6400 ;
        RECT 2086.9000 2518.6000 2088.5000 2519.0800 ;
        RECT 2131.9000 2496.8400 2133.5000 2497.3200 ;
        RECT 2131.9000 2502.2800 2133.5000 2502.7600 ;
        RECT 2131.9000 2480.5200 2133.5000 2481.0000 ;
        RECT 2131.9000 2485.9600 2133.5000 2486.4400 ;
        RECT 2131.9000 2491.4000 2133.5000 2491.8800 ;
        RECT 2086.9000 2496.8400 2088.5000 2497.3200 ;
        RECT 2086.9000 2502.2800 2088.5000 2502.7600 ;
        RECT 2086.9000 2480.5200 2088.5000 2481.0000 ;
        RECT 2086.9000 2485.9600 2088.5000 2486.4400 ;
        RECT 2086.9000 2491.4000 2088.5000 2491.8800 ;
        RECT 2037.3400 2524.0400 2040.3400 2524.5200 ;
        RECT 2037.3400 2529.4800 2040.3400 2529.9600 ;
        RECT 2037.3400 2513.1600 2040.3400 2513.6400 ;
        RECT 2037.3400 2507.7200 2040.3400 2508.2000 ;
        RECT 2037.3400 2518.6000 2040.3400 2519.0800 ;
        RECT 2037.3400 2496.8400 2040.3400 2497.3200 ;
        RECT 2037.3400 2502.2800 2040.3400 2502.7600 ;
        RECT 2037.3400 2485.9600 2040.3400 2486.4400 ;
        RECT 2037.3400 2480.5200 2040.3400 2481.0000 ;
        RECT 2037.3400 2491.4000 2040.3400 2491.8800 ;
        RECT 2037.3400 2534.9200 2040.3400 2535.4000 ;
        RECT 2086.9000 2534.9200 2088.5000 2535.4000 ;
        RECT 2131.9000 2534.9200 2133.5000 2535.4000 ;
        RECT 2233.4400 2469.6400 2236.4400 2470.1200 ;
        RECT 2233.4400 2475.0800 2236.4400 2475.5600 ;
        RECT 2221.9000 2469.6400 2223.5000 2470.1200 ;
        RECT 2221.9000 2475.0800 2223.5000 2475.5600 ;
        RECT 2233.4400 2453.3200 2236.4400 2453.8000 ;
        RECT 2233.4400 2458.7600 2236.4400 2459.2400 ;
        RECT 2233.4400 2464.2000 2236.4400 2464.6800 ;
        RECT 2221.9000 2453.3200 2223.5000 2453.8000 ;
        RECT 2221.9000 2458.7600 2223.5000 2459.2400 ;
        RECT 2221.9000 2464.2000 2223.5000 2464.6800 ;
        RECT 2233.4400 2442.4400 2236.4400 2442.9200 ;
        RECT 2233.4400 2447.8800 2236.4400 2448.3600 ;
        RECT 2221.9000 2442.4400 2223.5000 2442.9200 ;
        RECT 2221.9000 2447.8800 2223.5000 2448.3600 ;
        RECT 2233.4400 2426.1200 2236.4400 2426.6000 ;
        RECT 2233.4400 2431.5600 2236.4400 2432.0400 ;
        RECT 2233.4400 2437.0000 2236.4400 2437.4800 ;
        RECT 2221.9000 2426.1200 2223.5000 2426.6000 ;
        RECT 2221.9000 2431.5600 2223.5000 2432.0400 ;
        RECT 2221.9000 2437.0000 2223.5000 2437.4800 ;
        RECT 2176.9000 2469.6400 2178.5000 2470.1200 ;
        RECT 2176.9000 2475.0800 2178.5000 2475.5600 ;
        RECT 2176.9000 2453.3200 2178.5000 2453.8000 ;
        RECT 2176.9000 2458.7600 2178.5000 2459.2400 ;
        RECT 2176.9000 2464.2000 2178.5000 2464.6800 ;
        RECT 2176.9000 2442.4400 2178.5000 2442.9200 ;
        RECT 2176.9000 2447.8800 2178.5000 2448.3600 ;
        RECT 2176.9000 2426.1200 2178.5000 2426.6000 ;
        RECT 2176.9000 2431.5600 2178.5000 2432.0400 ;
        RECT 2176.9000 2437.0000 2178.5000 2437.4800 ;
        RECT 2233.4400 2415.2400 2236.4400 2415.7200 ;
        RECT 2233.4400 2420.6800 2236.4400 2421.1600 ;
        RECT 2221.9000 2415.2400 2223.5000 2415.7200 ;
        RECT 2221.9000 2420.6800 2223.5000 2421.1600 ;
        RECT 2233.4400 2398.9200 2236.4400 2399.4000 ;
        RECT 2233.4400 2404.3600 2236.4400 2404.8400 ;
        RECT 2233.4400 2409.8000 2236.4400 2410.2800 ;
        RECT 2221.9000 2398.9200 2223.5000 2399.4000 ;
        RECT 2221.9000 2404.3600 2223.5000 2404.8400 ;
        RECT 2221.9000 2409.8000 2223.5000 2410.2800 ;
        RECT 2233.4400 2388.0400 2236.4400 2388.5200 ;
        RECT 2233.4400 2393.4800 2236.4400 2393.9600 ;
        RECT 2221.9000 2388.0400 2223.5000 2388.5200 ;
        RECT 2221.9000 2393.4800 2223.5000 2393.9600 ;
        RECT 2233.4400 2382.6000 2236.4400 2383.0800 ;
        RECT 2221.9000 2382.6000 2223.5000 2383.0800 ;
        RECT 2176.9000 2415.2400 2178.5000 2415.7200 ;
        RECT 2176.9000 2420.6800 2178.5000 2421.1600 ;
        RECT 2176.9000 2398.9200 2178.5000 2399.4000 ;
        RECT 2176.9000 2404.3600 2178.5000 2404.8400 ;
        RECT 2176.9000 2409.8000 2178.5000 2410.2800 ;
        RECT 2176.9000 2388.0400 2178.5000 2388.5200 ;
        RECT 2176.9000 2393.4800 2178.5000 2393.9600 ;
        RECT 2176.9000 2382.6000 2178.5000 2383.0800 ;
        RECT 2131.9000 2469.6400 2133.5000 2470.1200 ;
        RECT 2131.9000 2475.0800 2133.5000 2475.5600 ;
        RECT 2131.9000 2453.3200 2133.5000 2453.8000 ;
        RECT 2131.9000 2458.7600 2133.5000 2459.2400 ;
        RECT 2131.9000 2464.2000 2133.5000 2464.6800 ;
        RECT 2086.9000 2469.6400 2088.5000 2470.1200 ;
        RECT 2086.9000 2475.0800 2088.5000 2475.5600 ;
        RECT 2086.9000 2453.3200 2088.5000 2453.8000 ;
        RECT 2086.9000 2458.7600 2088.5000 2459.2400 ;
        RECT 2086.9000 2464.2000 2088.5000 2464.6800 ;
        RECT 2131.9000 2442.4400 2133.5000 2442.9200 ;
        RECT 2131.9000 2447.8800 2133.5000 2448.3600 ;
        RECT 2131.9000 2426.1200 2133.5000 2426.6000 ;
        RECT 2131.9000 2431.5600 2133.5000 2432.0400 ;
        RECT 2131.9000 2437.0000 2133.5000 2437.4800 ;
        RECT 2086.9000 2442.4400 2088.5000 2442.9200 ;
        RECT 2086.9000 2447.8800 2088.5000 2448.3600 ;
        RECT 2086.9000 2426.1200 2088.5000 2426.6000 ;
        RECT 2086.9000 2431.5600 2088.5000 2432.0400 ;
        RECT 2086.9000 2437.0000 2088.5000 2437.4800 ;
        RECT 2037.3400 2469.6400 2040.3400 2470.1200 ;
        RECT 2037.3400 2475.0800 2040.3400 2475.5600 ;
        RECT 2037.3400 2458.7600 2040.3400 2459.2400 ;
        RECT 2037.3400 2453.3200 2040.3400 2453.8000 ;
        RECT 2037.3400 2464.2000 2040.3400 2464.6800 ;
        RECT 2037.3400 2442.4400 2040.3400 2442.9200 ;
        RECT 2037.3400 2447.8800 2040.3400 2448.3600 ;
        RECT 2037.3400 2431.5600 2040.3400 2432.0400 ;
        RECT 2037.3400 2426.1200 2040.3400 2426.6000 ;
        RECT 2037.3400 2437.0000 2040.3400 2437.4800 ;
        RECT 2131.9000 2415.2400 2133.5000 2415.7200 ;
        RECT 2131.9000 2420.6800 2133.5000 2421.1600 ;
        RECT 2131.9000 2398.9200 2133.5000 2399.4000 ;
        RECT 2131.9000 2404.3600 2133.5000 2404.8400 ;
        RECT 2131.9000 2409.8000 2133.5000 2410.2800 ;
        RECT 2086.9000 2415.2400 2088.5000 2415.7200 ;
        RECT 2086.9000 2420.6800 2088.5000 2421.1600 ;
        RECT 2086.9000 2398.9200 2088.5000 2399.4000 ;
        RECT 2086.9000 2404.3600 2088.5000 2404.8400 ;
        RECT 2086.9000 2409.8000 2088.5000 2410.2800 ;
        RECT 2131.9000 2393.4800 2133.5000 2393.9600 ;
        RECT 2131.9000 2388.0400 2133.5000 2388.5200 ;
        RECT 2131.9000 2382.6000 2133.5000 2383.0800 ;
        RECT 2086.9000 2393.4800 2088.5000 2393.9600 ;
        RECT 2086.9000 2388.0400 2088.5000 2388.5200 ;
        RECT 2086.9000 2382.6000 2088.5000 2383.0800 ;
        RECT 2037.3400 2415.2400 2040.3400 2415.7200 ;
        RECT 2037.3400 2420.6800 2040.3400 2421.1600 ;
        RECT 2037.3400 2404.3600 2040.3400 2404.8400 ;
        RECT 2037.3400 2398.9200 2040.3400 2399.4000 ;
        RECT 2037.3400 2409.8000 2040.3400 2410.2800 ;
        RECT 2037.3400 2388.0400 2040.3400 2388.5200 ;
        RECT 2037.3400 2393.4800 2040.3400 2393.9600 ;
        RECT 2037.3400 2382.6000 2040.3400 2383.0800 ;
        RECT 2037.3400 2580.7900 2236.4400 2583.7900 ;
        RECT 2037.3400 2375.6900 2236.4400 2378.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 2146.0500 2223.5000 2354.1500 ;
        RECT 2176.9000 2146.0500 2178.5000 2354.1500 ;
        RECT 2131.9000 2146.0500 2133.5000 2354.1500 ;
        RECT 2086.9000 2146.0500 2088.5000 2354.1500 ;
        RECT 2233.4400 2146.0500 2236.4400 2354.1500 ;
        RECT 2037.3400 2146.0500 2040.3400 2354.1500 ;
      LAYER met3 ;
        RECT 2233.4400 2348.8000 2236.4400 2349.2800 ;
        RECT 2221.9000 2348.8000 2223.5000 2349.2800 ;
        RECT 2233.4400 2337.9200 2236.4400 2338.4000 ;
        RECT 2233.4400 2343.3600 2236.4400 2343.8400 ;
        RECT 2221.9000 2337.9200 2223.5000 2338.4000 ;
        RECT 2221.9000 2343.3600 2223.5000 2343.8400 ;
        RECT 2233.4400 2321.6000 2236.4400 2322.0800 ;
        RECT 2233.4400 2327.0400 2236.4400 2327.5200 ;
        RECT 2221.9000 2321.6000 2223.5000 2322.0800 ;
        RECT 2221.9000 2327.0400 2223.5000 2327.5200 ;
        RECT 2233.4400 2310.7200 2236.4400 2311.2000 ;
        RECT 2233.4400 2316.1600 2236.4400 2316.6400 ;
        RECT 2221.9000 2310.7200 2223.5000 2311.2000 ;
        RECT 2221.9000 2316.1600 2223.5000 2316.6400 ;
        RECT 2233.4400 2332.4800 2236.4400 2332.9600 ;
        RECT 2221.9000 2332.4800 2223.5000 2332.9600 ;
        RECT 2176.9000 2337.9200 2178.5000 2338.4000 ;
        RECT 2176.9000 2343.3600 2178.5000 2343.8400 ;
        RECT 2176.9000 2348.8000 2178.5000 2349.2800 ;
        RECT 2176.9000 2321.6000 2178.5000 2322.0800 ;
        RECT 2176.9000 2327.0400 2178.5000 2327.5200 ;
        RECT 2176.9000 2316.1600 2178.5000 2316.6400 ;
        RECT 2176.9000 2310.7200 2178.5000 2311.2000 ;
        RECT 2176.9000 2332.4800 2178.5000 2332.9600 ;
        RECT 2233.4400 2294.4000 2236.4400 2294.8800 ;
        RECT 2233.4400 2299.8400 2236.4400 2300.3200 ;
        RECT 2221.9000 2294.4000 2223.5000 2294.8800 ;
        RECT 2221.9000 2299.8400 2223.5000 2300.3200 ;
        RECT 2233.4400 2278.0800 2236.4400 2278.5600 ;
        RECT 2233.4400 2283.5200 2236.4400 2284.0000 ;
        RECT 2233.4400 2288.9600 2236.4400 2289.4400 ;
        RECT 2221.9000 2278.0800 2223.5000 2278.5600 ;
        RECT 2221.9000 2283.5200 2223.5000 2284.0000 ;
        RECT 2221.9000 2288.9600 2223.5000 2289.4400 ;
        RECT 2233.4400 2267.2000 2236.4400 2267.6800 ;
        RECT 2233.4400 2272.6400 2236.4400 2273.1200 ;
        RECT 2221.9000 2267.2000 2223.5000 2267.6800 ;
        RECT 2221.9000 2272.6400 2223.5000 2273.1200 ;
        RECT 2233.4400 2250.8800 2236.4400 2251.3600 ;
        RECT 2233.4400 2256.3200 2236.4400 2256.8000 ;
        RECT 2233.4400 2261.7600 2236.4400 2262.2400 ;
        RECT 2221.9000 2250.8800 2223.5000 2251.3600 ;
        RECT 2221.9000 2256.3200 2223.5000 2256.8000 ;
        RECT 2221.9000 2261.7600 2223.5000 2262.2400 ;
        RECT 2176.9000 2294.4000 2178.5000 2294.8800 ;
        RECT 2176.9000 2299.8400 2178.5000 2300.3200 ;
        RECT 2176.9000 2278.0800 2178.5000 2278.5600 ;
        RECT 2176.9000 2283.5200 2178.5000 2284.0000 ;
        RECT 2176.9000 2288.9600 2178.5000 2289.4400 ;
        RECT 2176.9000 2267.2000 2178.5000 2267.6800 ;
        RECT 2176.9000 2272.6400 2178.5000 2273.1200 ;
        RECT 2176.9000 2250.8800 2178.5000 2251.3600 ;
        RECT 2176.9000 2256.3200 2178.5000 2256.8000 ;
        RECT 2176.9000 2261.7600 2178.5000 2262.2400 ;
        RECT 2233.4400 2305.2800 2236.4400 2305.7600 ;
        RECT 2176.9000 2305.2800 2178.5000 2305.7600 ;
        RECT 2221.9000 2305.2800 2223.5000 2305.7600 ;
        RECT 2131.9000 2337.9200 2133.5000 2338.4000 ;
        RECT 2131.9000 2343.3600 2133.5000 2343.8400 ;
        RECT 2131.9000 2348.8000 2133.5000 2349.2800 ;
        RECT 2086.9000 2337.9200 2088.5000 2338.4000 ;
        RECT 2086.9000 2343.3600 2088.5000 2343.8400 ;
        RECT 2086.9000 2348.8000 2088.5000 2349.2800 ;
        RECT 2131.9000 2321.6000 2133.5000 2322.0800 ;
        RECT 2131.9000 2327.0400 2133.5000 2327.5200 ;
        RECT 2131.9000 2310.7200 2133.5000 2311.2000 ;
        RECT 2131.9000 2316.1600 2133.5000 2316.6400 ;
        RECT 2086.9000 2321.6000 2088.5000 2322.0800 ;
        RECT 2086.9000 2327.0400 2088.5000 2327.5200 ;
        RECT 2086.9000 2310.7200 2088.5000 2311.2000 ;
        RECT 2086.9000 2316.1600 2088.5000 2316.6400 ;
        RECT 2086.9000 2332.4800 2088.5000 2332.9600 ;
        RECT 2131.9000 2332.4800 2133.5000 2332.9600 ;
        RECT 2037.3400 2348.8000 2040.3400 2349.2800 ;
        RECT 2037.3400 2343.3600 2040.3400 2343.8400 ;
        RECT 2037.3400 2337.9200 2040.3400 2338.4000 ;
        RECT 2037.3400 2327.0400 2040.3400 2327.5200 ;
        RECT 2037.3400 2321.6000 2040.3400 2322.0800 ;
        RECT 2037.3400 2316.1600 2040.3400 2316.6400 ;
        RECT 2037.3400 2310.7200 2040.3400 2311.2000 ;
        RECT 2037.3400 2332.4800 2040.3400 2332.9600 ;
        RECT 2131.9000 2294.4000 2133.5000 2294.8800 ;
        RECT 2131.9000 2299.8400 2133.5000 2300.3200 ;
        RECT 2131.9000 2278.0800 2133.5000 2278.5600 ;
        RECT 2131.9000 2283.5200 2133.5000 2284.0000 ;
        RECT 2131.9000 2288.9600 2133.5000 2289.4400 ;
        RECT 2086.9000 2294.4000 2088.5000 2294.8800 ;
        RECT 2086.9000 2299.8400 2088.5000 2300.3200 ;
        RECT 2086.9000 2278.0800 2088.5000 2278.5600 ;
        RECT 2086.9000 2283.5200 2088.5000 2284.0000 ;
        RECT 2086.9000 2288.9600 2088.5000 2289.4400 ;
        RECT 2131.9000 2267.2000 2133.5000 2267.6800 ;
        RECT 2131.9000 2272.6400 2133.5000 2273.1200 ;
        RECT 2131.9000 2250.8800 2133.5000 2251.3600 ;
        RECT 2131.9000 2256.3200 2133.5000 2256.8000 ;
        RECT 2131.9000 2261.7600 2133.5000 2262.2400 ;
        RECT 2086.9000 2267.2000 2088.5000 2267.6800 ;
        RECT 2086.9000 2272.6400 2088.5000 2273.1200 ;
        RECT 2086.9000 2250.8800 2088.5000 2251.3600 ;
        RECT 2086.9000 2256.3200 2088.5000 2256.8000 ;
        RECT 2086.9000 2261.7600 2088.5000 2262.2400 ;
        RECT 2037.3400 2294.4000 2040.3400 2294.8800 ;
        RECT 2037.3400 2299.8400 2040.3400 2300.3200 ;
        RECT 2037.3400 2283.5200 2040.3400 2284.0000 ;
        RECT 2037.3400 2278.0800 2040.3400 2278.5600 ;
        RECT 2037.3400 2288.9600 2040.3400 2289.4400 ;
        RECT 2037.3400 2267.2000 2040.3400 2267.6800 ;
        RECT 2037.3400 2272.6400 2040.3400 2273.1200 ;
        RECT 2037.3400 2256.3200 2040.3400 2256.8000 ;
        RECT 2037.3400 2250.8800 2040.3400 2251.3600 ;
        RECT 2037.3400 2261.7600 2040.3400 2262.2400 ;
        RECT 2037.3400 2305.2800 2040.3400 2305.7600 ;
        RECT 2086.9000 2305.2800 2088.5000 2305.7600 ;
        RECT 2131.9000 2305.2800 2133.5000 2305.7600 ;
        RECT 2233.4400 2240.0000 2236.4400 2240.4800 ;
        RECT 2233.4400 2245.4400 2236.4400 2245.9200 ;
        RECT 2221.9000 2240.0000 2223.5000 2240.4800 ;
        RECT 2221.9000 2245.4400 2223.5000 2245.9200 ;
        RECT 2233.4400 2223.6800 2236.4400 2224.1600 ;
        RECT 2233.4400 2229.1200 2236.4400 2229.6000 ;
        RECT 2233.4400 2234.5600 2236.4400 2235.0400 ;
        RECT 2221.9000 2223.6800 2223.5000 2224.1600 ;
        RECT 2221.9000 2229.1200 2223.5000 2229.6000 ;
        RECT 2221.9000 2234.5600 2223.5000 2235.0400 ;
        RECT 2233.4400 2212.8000 2236.4400 2213.2800 ;
        RECT 2233.4400 2218.2400 2236.4400 2218.7200 ;
        RECT 2221.9000 2212.8000 2223.5000 2213.2800 ;
        RECT 2221.9000 2218.2400 2223.5000 2218.7200 ;
        RECT 2233.4400 2196.4800 2236.4400 2196.9600 ;
        RECT 2233.4400 2201.9200 2236.4400 2202.4000 ;
        RECT 2233.4400 2207.3600 2236.4400 2207.8400 ;
        RECT 2221.9000 2196.4800 2223.5000 2196.9600 ;
        RECT 2221.9000 2201.9200 2223.5000 2202.4000 ;
        RECT 2221.9000 2207.3600 2223.5000 2207.8400 ;
        RECT 2176.9000 2240.0000 2178.5000 2240.4800 ;
        RECT 2176.9000 2245.4400 2178.5000 2245.9200 ;
        RECT 2176.9000 2223.6800 2178.5000 2224.1600 ;
        RECT 2176.9000 2229.1200 2178.5000 2229.6000 ;
        RECT 2176.9000 2234.5600 2178.5000 2235.0400 ;
        RECT 2176.9000 2212.8000 2178.5000 2213.2800 ;
        RECT 2176.9000 2218.2400 2178.5000 2218.7200 ;
        RECT 2176.9000 2196.4800 2178.5000 2196.9600 ;
        RECT 2176.9000 2201.9200 2178.5000 2202.4000 ;
        RECT 2176.9000 2207.3600 2178.5000 2207.8400 ;
        RECT 2233.4400 2185.6000 2236.4400 2186.0800 ;
        RECT 2233.4400 2191.0400 2236.4400 2191.5200 ;
        RECT 2221.9000 2185.6000 2223.5000 2186.0800 ;
        RECT 2221.9000 2191.0400 2223.5000 2191.5200 ;
        RECT 2233.4400 2169.2800 2236.4400 2169.7600 ;
        RECT 2233.4400 2174.7200 2236.4400 2175.2000 ;
        RECT 2233.4400 2180.1600 2236.4400 2180.6400 ;
        RECT 2221.9000 2169.2800 2223.5000 2169.7600 ;
        RECT 2221.9000 2174.7200 2223.5000 2175.2000 ;
        RECT 2221.9000 2180.1600 2223.5000 2180.6400 ;
        RECT 2233.4400 2158.4000 2236.4400 2158.8800 ;
        RECT 2233.4400 2163.8400 2236.4400 2164.3200 ;
        RECT 2221.9000 2158.4000 2223.5000 2158.8800 ;
        RECT 2221.9000 2163.8400 2223.5000 2164.3200 ;
        RECT 2233.4400 2152.9600 2236.4400 2153.4400 ;
        RECT 2221.9000 2152.9600 2223.5000 2153.4400 ;
        RECT 2176.9000 2185.6000 2178.5000 2186.0800 ;
        RECT 2176.9000 2191.0400 2178.5000 2191.5200 ;
        RECT 2176.9000 2169.2800 2178.5000 2169.7600 ;
        RECT 2176.9000 2174.7200 2178.5000 2175.2000 ;
        RECT 2176.9000 2180.1600 2178.5000 2180.6400 ;
        RECT 2176.9000 2158.4000 2178.5000 2158.8800 ;
        RECT 2176.9000 2163.8400 2178.5000 2164.3200 ;
        RECT 2176.9000 2152.9600 2178.5000 2153.4400 ;
        RECT 2131.9000 2240.0000 2133.5000 2240.4800 ;
        RECT 2131.9000 2245.4400 2133.5000 2245.9200 ;
        RECT 2131.9000 2223.6800 2133.5000 2224.1600 ;
        RECT 2131.9000 2229.1200 2133.5000 2229.6000 ;
        RECT 2131.9000 2234.5600 2133.5000 2235.0400 ;
        RECT 2086.9000 2240.0000 2088.5000 2240.4800 ;
        RECT 2086.9000 2245.4400 2088.5000 2245.9200 ;
        RECT 2086.9000 2223.6800 2088.5000 2224.1600 ;
        RECT 2086.9000 2229.1200 2088.5000 2229.6000 ;
        RECT 2086.9000 2234.5600 2088.5000 2235.0400 ;
        RECT 2131.9000 2212.8000 2133.5000 2213.2800 ;
        RECT 2131.9000 2218.2400 2133.5000 2218.7200 ;
        RECT 2131.9000 2196.4800 2133.5000 2196.9600 ;
        RECT 2131.9000 2201.9200 2133.5000 2202.4000 ;
        RECT 2131.9000 2207.3600 2133.5000 2207.8400 ;
        RECT 2086.9000 2212.8000 2088.5000 2213.2800 ;
        RECT 2086.9000 2218.2400 2088.5000 2218.7200 ;
        RECT 2086.9000 2196.4800 2088.5000 2196.9600 ;
        RECT 2086.9000 2201.9200 2088.5000 2202.4000 ;
        RECT 2086.9000 2207.3600 2088.5000 2207.8400 ;
        RECT 2037.3400 2240.0000 2040.3400 2240.4800 ;
        RECT 2037.3400 2245.4400 2040.3400 2245.9200 ;
        RECT 2037.3400 2229.1200 2040.3400 2229.6000 ;
        RECT 2037.3400 2223.6800 2040.3400 2224.1600 ;
        RECT 2037.3400 2234.5600 2040.3400 2235.0400 ;
        RECT 2037.3400 2212.8000 2040.3400 2213.2800 ;
        RECT 2037.3400 2218.2400 2040.3400 2218.7200 ;
        RECT 2037.3400 2201.9200 2040.3400 2202.4000 ;
        RECT 2037.3400 2196.4800 2040.3400 2196.9600 ;
        RECT 2037.3400 2207.3600 2040.3400 2207.8400 ;
        RECT 2131.9000 2185.6000 2133.5000 2186.0800 ;
        RECT 2131.9000 2191.0400 2133.5000 2191.5200 ;
        RECT 2131.9000 2169.2800 2133.5000 2169.7600 ;
        RECT 2131.9000 2174.7200 2133.5000 2175.2000 ;
        RECT 2131.9000 2180.1600 2133.5000 2180.6400 ;
        RECT 2086.9000 2185.6000 2088.5000 2186.0800 ;
        RECT 2086.9000 2191.0400 2088.5000 2191.5200 ;
        RECT 2086.9000 2169.2800 2088.5000 2169.7600 ;
        RECT 2086.9000 2174.7200 2088.5000 2175.2000 ;
        RECT 2086.9000 2180.1600 2088.5000 2180.6400 ;
        RECT 2131.9000 2163.8400 2133.5000 2164.3200 ;
        RECT 2131.9000 2158.4000 2133.5000 2158.8800 ;
        RECT 2131.9000 2152.9600 2133.5000 2153.4400 ;
        RECT 2086.9000 2163.8400 2088.5000 2164.3200 ;
        RECT 2086.9000 2158.4000 2088.5000 2158.8800 ;
        RECT 2086.9000 2152.9600 2088.5000 2153.4400 ;
        RECT 2037.3400 2185.6000 2040.3400 2186.0800 ;
        RECT 2037.3400 2191.0400 2040.3400 2191.5200 ;
        RECT 2037.3400 2174.7200 2040.3400 2175.2000 ;
        RECT 2037.3400 2169.2800 2040.3400 2169.7600 ;
        RECT 2037.3400 2180.1600 2040.3400 2180.6400 ;
        RECT 2037.3400 2158.4000 2040.3400 2158.8800 ;
        RECT 2037.3400 2163.8400 2040.3400 2164.3200 ;
        RECT 2037.3400 2152.9600 2040.3400 2153.4400 ;
        RECT 2037.3400 2351.1500 2236.4400 2354.1500 ;
        RECT 2037.3400 2146.0500 2236.4400 2149.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 1916.4100 2223.5000 2124.5100 ;
        RECT 2176.9000 1916.4100 2178.5000 2124.5100 ;
        RECT 2131.9000 1916.4100 2133.5000 2124.5100 ;
        RECT 2086.9000 1916.4100 2088.5000 2124.5100 ;
        RECT 2233.4400 1916.4100 2236.4400 2124.5100 ;
        RECT 2037.3400 1916.4100 2040.3400 2124.5100 ;
      LAYER met3 ;
        RECT 2233.4400 2119.1600 2236.4400 2119.6400 ;
        RECT 2221.9000 2119.1600 2223.5000 2119.6400 ;
        RECT 2233.4400 2108.2800 2236.4400 2108.7600 ;
        RECT 2233.4400 2113.7200 2236.4400 2114.2000 ;
        RECT 2221.9000 2108.2800 2223.5000 2108.7600 ;
        RECT 2221.9000 2113.7200 2223.5000 2114.2000 ;
        RECT 2233.4400 2091.9600 2236.4400 2092.4400 ;
        RECT 2233.4400 2097.4000 2236.4400 2097.8800 ;
        RECT 2221.9000 2091.9600 2223.5000 2092.4400 ;
        RECT 2221.9000 2097.4000 2223.5000 2097.8800 ;
        RECT 2233.4400 2081.0800 2236.4400 2081.5600 ;
        RECT 2233.4400 2086.5200 2236.4400 2087.0000 ;
        RECT 2221.9000 2081.0800 2223.5000 2081.5600 ;
        RECT 2221.9000 2086.5200 2223.5000 2087.0000 ;
        RECT 2233.4400 2102.8400 2236.4400 2103.3200 ;
        RECT 2221.9000 2102.8400 2223.5000 2103.3200 ;
        RECT 2176.9000 2108.2800 2178.5000 2108.7600 ;
        RECT 2176.9000 2113.7200 2178.5000 2114.2000 ;
        RECT 2176.9000 2119.1600 2178.5000 2119.6400 ;
        RECT 2176.9000 2091.9600 2178.5000 2092.4400 ;
        RECT 2176.9000 2097.4000 2178.5000 2097.8800 ;
        RECT 2176.9000 2086.5200 2178.5000 2087.0000 ;
        RECT 2176.9000 2081.0800 2178.5000 2081.5600 ;
        RECT 2176.9000 2102.8400 2178.5000 2103.3200 ;
        RECT 2233.4400 2064.7600 2236.4400 2065.2400 ;
        RECT 2233.4400 2070.2000 2236.4400 2070.6800 ;
        RECT 2221.9000 2064.7600 2223.5000 2065.2400 ;
        RECT 2221.9000 2070.2000 2223.5000 2070.6800 ;
        RECT 2233.4400 2048.4400 2236.4400 2048.9200 ;
        RECT 2233.4400 2053.8800 2236.4400 2054.3600 ;
        RECT 2233.4400 2059.3200 2236.4400 2059.8000 ;
        RECT 2221.9000 2048.4400 2223.5000 2048.9200 ;
        RECT 2221.9000 2053.8800 2223.5000 2054.3600 ;
        RECT 2221.9000 2059.3200 2223.5000 2059.8000 ;
        RECT 2233.4400 2037.5600 2236.4400 2038.0400 ;
        RECT 2233.4400 2043.0000 2236.4400 2043.4800 ;
        RECT 2221.9000 2037.5600 2223.5000 2038.0400 ;
        RECT 2221.9000 2043.0000 2223.5000 2043.4800 ;
        RECT 2233.4400 2021.2400 2236.4400 2021.7200 ;
        RECT 2233.4400 2026.6800 2236.4400 2027.1600 ;
        RECT 2233.4400 2032.1200 2236.4400 2032.6000 ;
        RECT 2221.9000 2021.2400 2223.5000 2021.7200 ;
        RECT 2221.9000 2026.6800 2223.5000 2027.1600 ;
        RECT 2221.9000 2032.1200 2223.5000 2032.6000 ;
        RECT 2176.9000 2064.7600 2178.5000 2065.2400 ;
        RECT 2176.9000 2070.2000 2178.5000 2070.6800 ;
        RECT 2176.9000 2048.4400 2178.5000 2048.9200 ;
        RECT 2176.9000 2053.8800 2178.5000 2054.3600 ;
        RECT 2176.9000 2059.3200 2178.5000 2059.8000 ;
        RECT 2176.9000 2037.5600 2178.5000 2038.0400 ;
        RECT 2176.9000 2043.0000 2178.5000 2043.4800 ;
        RECT 2176.9000 2021.2400 2178.5000 2021.7200 ;
        RECT 2176.9000 2026.6800 2178.5000 2027.1600 ;
        RECT 2176.9000 2032.1200 2178.5000 2032.6000 ;
        RECT 2233.4400 2075.6400 2236.4400 2076.1200 ;
        RECT 2176.9000 2075.6400 2178.5000 2076.1200 ;
        RECT 2221.9000 2075.6400 2223.5000 2076.1200 ;
        RECT 2131.9000 2108.2800 2133.5000 2108.7600 ;
        RECT 2131.9000 2113.7200 2133.5000 2114.2000 ;
        RECT 2131.9000 2119.1600 2133.5000 2119.6400 ;
        RECT 2086.9000 2108.2800 2088.5000 2108.7600 ;
        RECT 2086.9000 2113.7200 2088.5000 2114.2000 ;
        RECT 2086.9000 2119.1600 2088.5000 2119.6400 ;
        RECT 2131.9000 2091.9600 2133.5000 2092.4400 ;
        RECT 2131.9000 2097.4000 2133.5000 2097.8800 ;
        RECT 2131.9000 2081.0800 2133.5000 2081.5600 ;
        RECT 2131.9000 2086.5200 2133.5000 2087.0000 ;
        RECT 2086.9000 2091.9600 2088.5000 2092.4400 ;
        RECT 2086.9000 2097.4000 2088.5000 2097.8800 ;
        RECT 2086.9000 2081.0800 2088.5000 2081.5600 ;
        RECT 2086.9000 2086.5200 2088.5000 2087.0000 ;
        RECT 2086.9000 2102.8400 2088.5000 2103.3200 ;
        RECT 2131.9000 2102.8400 2133.5000 2103.3200 ;
        RECT 2037.3400 2119.1600 2040.3400 2119.6400 ;
        RECT 2037.3400 2113.7200 2040.3400 2114.2000 ;
        RECT 2037.3400 2108.2800 2040.3400 2108.7600 ;
        RECT 2037.3400 2097.4000 2040.3400 2097.8800 ;
        RECT 2037.3400 2091.9600 2040.3400 2092.4400 ;
        RECT 2037.3400 2086.5200 2040.3400 2087.0000 ;
        RECT 2037.3400 2081.0800 2040.3400 2081.5600 ;
        RECT 2037.3400 2102.8400 2040.3400 2103.3200 ;
        RECT 2131.9000 2064.7600 2133.5000 2065.2400 ;
        RECT 2131.9000 2070.2000 2133.5000 2070.6800 ;
        RECT 2131.9000 2048.4400 2133.5000 2048.9200 ;
        RECT 2131.9000 2053.8800 2133.5000 2054.3600 ;
        RECT 2131.9000 2059.3200 2133.5000 2059.8000 ;
        RECT 2086.9000 2064.7600 2088.5000 2065.2400 ;
        RECT 2086.9000 2070.2000 2088.5000 2070.6800 ;
        RECT 2086.9000 2048.4400 2088.5000 2048.9200 ;
        RECT 2086.9000 2053.8800 2088.5000 2054.3600 ;
        RECT 2086.9000 2059.3200 2088.5000 2059.8000 ;
        RECT 2131.9000 2037.5600 2133.5000 2038.0400 ;
        RECT 2131.9000 2043.0000 2133.5000 2043.4800 ;
        RECT 2131.9000 2021.2400 2133.5000 2021.7200 ;
        RECT 2131.9000 2026.6800 2133.5000 2027.1600 ;
        RECT 2131.9000 2032.1200 2133.5000 2032.6000 ;
        RECT 2086.9000 2037.5600 2088.5000 2038.0400 ;
        RECT 2086.9000 2043.0000 2088.5000 2043.4800 ;
        RECT 2086.9000 2021.2400 2088.5000 2021.7200 ;
        RECT 2086.9000 2026.6800 2088.5000 2027.1600 ;
        RECT 2086.9000 2032.1200 2088.5000 2032.6000 ;
        RECT 2037.3400 2064.7600 2040.3400 2065.2400 ;
        RECT 2037.3400 2070.2000 2040.3400 2070.6800 ;
        RECT 2037.3400 2053.8800 2040.3400 2054.3600 ;
        RECT 2037.3400 2048.4400 2040.3400 2048.9200 ;
        RECT 2037.3400 2059.3200 2040.3400 2059.8000 ;
        RECT 2037.3400 2037.5600 2040.3400 2038.0400 ;
        RECT 2037.3400 2043.0000 2040.3400 2043.4800 ;
        RECT 2037.3400 2026.6800 2040.3400 2027.1600 ;
        RECT 2037.3400 2021.2400 2040.3400 2021.7200 ;
        RECT 2037.3400 2032.1200 2040.3400 2032.6000 ;
        RECT 2037.3400 2075.6400 2040.3400 2076.1200 ;
        RECT 2086.9000 2075.6400 2088.5000 2076.1200 ;
        RECT 2131.9000 2075.6400 2133.5000 2076.1200 ;
        RECT 2233.4400 2010.3600 2236.4400 2010.8400 ;
        RECT 2233.4400 2015.8000 2236.4400 2016.2800 ;
        RECT 2221.9000 2010.3600 2223.5000 2010.8400 ;
        RECT 2221.9000 2015.8000 2223.5000 2016.2800 ;
        RECT 2233.4400 1994.0400 2236.4400 1994.5200 ;
        RECT 2233.4400 1999.4800 2236.4400 1999.9600 ;
        RECT 2233.4400 2004.9200 2236.4400 2005.4000 ;
        RECT 2221.9000 1994.0400 2223.5000 1994.5200 ;
        RECT 2221.9000 1999.4800 2223.5000 1999.9600 ;
        RECT 2221.9000 2004.9200 2223.5000 2005.4000 ;
        RECT 2233.4400 1983.1600 2236.4400 1983.6400 ;
        RECT 2233.4400 1988.6000 2236.4400 1989.0800 ;
        RECT 2221.9000 1983.1600 2223.5000 1983.6400 ;
        RECT 2221.9000 1988.6000 2223.5000 1989.0800 ;
        RECT 2233.4400 1966.8400 2236.4400 1967.3200 ;
        RECT 2233.4400 1972.2800 2236.4400 1972.7600 ;
        RECT 2233.4400 1977.7200 2236.4400 1978.2000 ;
        RECT 2221.9000 1966.8400 2223.5000 1967.3200 ;
        RECT 2221.9000 1972.2800 2223.5000 1972.7600 ;
        RECT 2221.9000 1977.7200 2223.5000 1978.2000 ;
        RECT 2176.9000 2010.3600 2178.5000 2010.8400 ;
        RECT 2176.9000 2015.8000 2178.5000 2016.2800 ;
        RECT 2176.9000 1994.0400 2178.5000 1994.5200 ;
        RECT 2176.9000 1999.4800 2178.5000 1999.9600 ;
        RECT 2176.9000 2004.9200 2178.5000 2005.4000 ;
        RECT 2176.9000 1983.1600 2178.5000 1983.6400 ;
        RECT 2176.9000 1988.6000 2178.5000 1989.0800 ;
        RECT 2176.9000 1966.8400 2178.5000 1967.3200 ;
        RECT 2176.9000 1972.2800 2178.5000 1972.7600 ;
        RECT 2176.9000 1977.7200 2178.5000 1978.2000 ;
        RECT 2233.4400 1955.9600 2236.4400 1956.4400 ;
        RECT 2233.4400 1961.4000 2236.4400 1961.8800 ;
        RECT 2221.9000 1955.9600 2223.5000 1956.4400 ;
        RECT 2221.9000 1961.4000 2223.5000 1961.8800 ;
        RECT 2233.4400 1939.6400 2236.4400 1940.1200 ;
        RECT 2233.4400 1945.0800 2236.4400 1945.5600 ;
        RECT 2233.4400 1950.5200 2236.4400 1951.0000 ;
        RECT 2221.9000 1939.6400 2223.5000 1940.1200 ;
        RECT 2221.9000 1945.0800 2223.5000 1945.5600 ;
        RECT 2221.9000 1950.5200 2223.5000 1951.0000 ;
        RECT 2233.4400 1928.7600 2236.4400 1929.2400 ;
        RECT 2233.4400 1934.2000 2236.4400 1934.6800 ;
        RECT 2221.9000 1928.7600 2223.5000 1929.2400 ;
        RECT 2221.9000 1934.2000 2223.5000 1934.6800 ;
        RECT 2233.4400 1923.3200 2236.4400 1923.8000 ;
        RECT 2221.9000 1923.3200 2223.5000 1923.8000 ;
        RECT 2176.9000 1955.9600 2178.5000 1956.4400 ;
        RECT 2176.9000 1961.4000 2178.5000 1961.8800 ;
        RECT 2176.9000 1939.6400 2178.5000 1940.1200 ;
        RECT 2176.9000 1945.0800 2178.5000 1945.5600 ;
        RECT 2176.9000 1950.5200 2178.5000 1951.0000 ;
        RECT 2176.9000 1928.7600 2178.5000 1929.2400 ;
        RECT 2176.9000 1934.2000 2178.5000 1934.6800 ;
        RECT 2176.9000 1923.3200 2178.5000 1923.8000 ;
        RECT 2131.9000 2010.3600 2133.5000 2010.8400 ;
        RECT 2131.9000 2015.8000 2133.5000 2016.2800 ;
        RECT 2131.9000 1994.0400 2133.5000 1994.5200 ;
        RECT 2131.9000 1999.4800 2133.5000 1999.9600 ;
        RECT 2131.9000 2004.9200 2133.5000 2005.4000 ;
        RECT 2086.9000 2010.3600 2088.5000 2010.8400 ;
        RECT 2086.9000 2015.8000 2088.5000 2016.2800 ;
        RECT 2086.9000 1994.0400 2088.5000 1994.5200 ;
        RECT 2086.9000 1999.4800 2088.5000 1999.9600 ;
        RECT 2086.9000 2004.9200 2088.5000 2005.4000 ;
        RECT 2131.9000 1983.1600 2133.5000 1983.6400 ;
        RECT 2131.9000 1988.6000 2133.5000 1989.0800 ;
        RECT 2131.9000 1966.8400 2133.5000 1967.3200 ;
        RECT 2131.9000 1972.2800 2133.5000 1972.7600 ;
        RECT 2131.9000 1977.7200 2133.5000 1978.2000 ;
        RECT 2086.9000 1983.1600 2088.5000 1983.6400 ;
        RECT 2086.9000 1988.6000 2088.5000 1989.0800 ;
        RECT 2086.9000 1966.8400 2088.5000 1967.3200 ;
        RECT 2086.9000 1972.2800 2088.5000 1972.7600 ;
        RECT 2086.9000 1977.7200 2088.5000 1978.2000 ;
        RECT 2037.3400 2010.3600 2040.3400 2010.8400 ;
        RECT 2037.3400 2015.8000 2040.3400 2016.2800 ;
        RECT 2037.3400 1999.4800 2040.3400 1999.9600 ;
        RECT 2037.3400 1994.0400 2040.3400 1994.5200 ;
        RECT 2037.3400 2004.9200 2040.3400 2005.4000 ;
        RECT 2037.3400 1983.1600 2040.3400 1983.6400 ;
        RECT 2037.3400 1988.6000 2040.3400 1989.0800 ;
        RECT 2037.3400 1972.2800 2040.3400 1972.7600 ;
        RECT 2037.3400 1966.8400 2040.3400 1967.3200 ;
        RECT 2037.3400 1977.7200 2040.3400 1978.2000 ;
        RECT 2131.9000 1955.9600 2133.5000 1956.4400 ;
        RECT 2131.9000 1961.4000 2133.5000 1961.8800 ;
        RECT 2131.9000 1939.6400 2133.5000 1940.1200 ;
        RECT 2131.9000 1945.0800 2133.5000 1945.5600 ;
        RECT 2131.9000 1950.5200 2133.5000 1951.0000 ;
        RECT 2086.9000 1955.9600 2088.5000 1956.4400 ;
        RECT 2086.9000 1961.4000 2088.5000 1961.8800 ;
        RECT 2086.9000 1939.6400 2088.5000 1940.1200 ;
        RECT 2086.9000 1945.0800 2088.5000 1945.5600 ;
        RECT 2086.9000 1950.5200 2088.5000 1951.0000 ;
        RECT 2131.9000 1934.2000 2133.5000 1934.6800 ;
        RECT 2131.9000 1928.7600 2133.5000 1929.2400 ;
        RECT 2131.9000 1923.3200 2133.5000 1923.8000 ;
        RECT 2086.9000 1934.2000 2088.5000 1934.6800 ;
        RECT 2086.9000 1928.7600 2088.5000 1929.2400 ;
        RECT 2086.9000 1923.3200 2088.5000 1923.8000 ;
        RECT 2037.3400 1955.9600 2040.3400 1956.4400 ;
        RECT 2037.3400 1961.4000 2040.3400 1961.8800 ;
        RECT 2037.3400 1945.0800 2040.3400 1945.5600 ;
        RECT 2037.3400 1939.6400 2040.3400 1940.1200 ;
        RECT 2037.3400 1950.5200 2040.3400 1951.0000 ;
        RECT 2037.3400 1928.7600 2040.3400 1929.2400 ;
        RECT 2037.3400 1934.2000 2040.3400 1934.6800 ;
        RECT 2037.3400 1923.3200 2040.3400 1923.8000 ;
        RECT 2037.3400 2121.5100 2236.4400 2124.5100 ;
        RECT 2037.3400 1916.4100 2236.4400 1919.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 1686.7700 2223.5000 1894.8700 ;
        RECT 2176.9000 1686.7700 2178.5000 1894.8700 ;
        RECT 2131.9000 1686.7700 2133.5000 1894.8700 ;
        RECT 2086.9000 1686.7700 2088.5000 1894.8700 ;
        RECT 2233.4400 1686.7700 2236.4400 1894.8700 ;
        RECT 2037.3400 1686.7700 2040.3400 1894.8700 ;
      LAYER met3 ;
        RECT 2233.4400 1889.5200 2236.4400 1890.0000 ;
        RECT 2221.9000 1889.5200 2223.5000 1890.0000 ;
        RECT 2233.4400 1878.6400 2236.4400 1879.1200 ;
        RECT 2233.4400 1884.0800 2236.4400 1884.5600 ;
        RECT 2221.9000 1878.6400 2223.5000 1879.1200 ;
        RECT 2221.9000 1884.0800 2223.5000 1884.5600 ;
        RECT 2233.4400 1862.3200 2236.4400 1862.8000 ;
        RECT 2233.4400 1867.7600 2236.4400 1868.2400 ;
        RECT 2221.9000 1862.3200 2223.5000 1862.8000 ;
        RECT 2221.9000 1867.7600 2223.5000 1868.2400 ;
        RECT 2233.4400 1851.4400 2236.4400 1851.9200 ;
        RECT 2233.4400 1856.8800 2236.4400 1857.3600 ;
        RECT 2221.9000 1851.4400 2223.5000 1851.9200 ;
        RECT 2221.9000 1856.8800 2223.5000 1857.3600 ;
        RECT 2233.4400 1873.2000 2236.4400 1873.6800 ;
        RECT 2221.9000 1873.2000 2223.5000 1873.6800 ;
        RECT 2176.9000 1878.6400 2178.5000 1879.1200 ;
        RECT 2176.9000 1884.0800 2178.5000 1884.5600 ;
        RECT 2176.9000 1889.5200 2178.5000 1890.0000 ;
        RECT 2176.9000 1862.3200 2178.5000 1862.8000 ;
        RECT 2176.9000 1867.7600 2178.5000 1868.2400 ;
        RECT 2176.9000 1856.8800 2178.5000 1857.3600 ;
        RECT 2176.9000 1851.4400 2178.5000 1851.9200 ;
        RECT 2176.9000 1873.2000 2178.5000 1873.6800 ;
        RECT 2233.4400 1835.1200 2236.4400 1835.6000 ;
        RECT 2233.4400 1840.5600 2236.4400 1841.0400 ;
        RECT 2221.9000 1835.1200 2223.5000 1835.6000 ;
        RECT 2221.9000 1840.5600 2223.5000 1841.0400 ;
        RECT 2233.4400 1818.8000 2236.4400 1819.2800 ;
        RECT 2233.4400 1824.2400 2236.4400 1824.7200 ;
        RECT 2233.4400 1829.6800 2236.4400 1830.1600 ;
        RECT 2221.9000 1818.8000 2223.5000 1819.2800 ;
        RECT 2221.9000 1824.2400 2223.5000 1824.7200 ;
        RECT 2221.9000 1829.6800 2223.5000 1830.1600 ;
        RECT 2233.4400 1807.9200 2236.4400 1808.4000 ;
        RECT 2233.4400 1813.3600 2236.4400 1813.8400 ;
        RECT 2221.9000 1807.9200 2223.5000 1808.4000 ;
        RECT 2221.9000 1813.3600 2223.5000 1813.8400 ;
        RECT 2233.4400 1791.6000 2236.4400 1792.0800 ;
        RECT 2233.4400 1797.0400 2236.4400 1797.5200 ;
        RECT 2233.4400 1802.4800 2236.4400 1802.9600 ;
        RECT 2221.9000 1791.6000 2223.5000 1792.0800 ;
        RECT 2221.9000 1797.0400 2223.5000 1797.5200 ;
        RECT 2221.9000 1802.4800 2223.5000 1802.9600 ;
        RECT 2176.9000 1835.1200 2178.5000 1835.6000 ;
        RECT 2176.9000 1840.5600 2178.5000 1841.0400 ;
        RECT 2176.9000 1818.8000 2178.5000 1819.2800 ;
        RECT 2176.9000 1824.2400 2178.5000 1824.7200 ;
        RECT 2176.9000 1829.6800 2178.5000 1830.1600 ;
        RECT 2176.9000 1807.9200 2178.5000 1808.4000 ;
        RECT 2176.9000 1813.3600 2178.5000 1813.8400 ;
        RECT 2176.9000 1791.6000 2178.5000 1792.0800 ;
        RECT 2176.9000 1797.0400 2178.5000 1797.5200 ;
        RECT 2176.9000 1802.4800 2178.5000 1802.9600 ;
        RECT 2233.4400 1846.0000 2236.4400 1846.4800 ;
        RECT 2176.9000 1846.0000 2178.5000 1846.4800 ;
        RECT 2221.9000 1846.0000 2223.5000 1846.4800 ;
        RECT 2131.9000 1878.6400 2133.5000 1879.1200 ;
        RECT 2131.9000 1884.0800 2133.5000 1884.5600 ;
        RECT 2131.9000 1889.5200 2133.5000 1890.0000 ;
        RECT 2086.9000 1878.6400 2088.5000 1879.1200 ;
        RECT 2086.9000 1884.0800 2088.5000 1884.5600 ;
        RECT 2086.9000 1889.5200 2088.5000 1890.0000 ;
        RECT 2131.9000 1862.3200 2133.5000 1862.8000 ;
        RECT 2131.9000 1867.7600 2133.5000 1868.2400 ;
        RECT 2131.9000 1851.4400 2133.5000 1851.9200 ;
        RECT 2131.9000 1856.8800 2133.5000 1857.3600 ;
        RECT 2086.9000 1862.3200 2088.5000 1862.8000 ;
        RECT 2086.9000 1867.7600 2088.5000 1868.2400 ;
        RECT 2086.9000 1851.4400 2088.5000 1851.9200 ;
        RECT 2086.9000 1856.8800 2088.5000 1857.3600 ;
        RECT 2086.9000 1873.2000 2088.5000 1873.6800 ;
        RECT 2131.9000 1873.2000 2133.5000 1873.6800 ;
        RECT 2037.3400 1889.5200 2040.3400 1890.0000 ;
        RECT 2037.3400 1884.0800 2040.3400 1884.5600 ;
        RECT 2037.3400 1878.6400 2040.3400 1879.1200 ;
        RECT 2037.3400 1867.7600 2040.3400 1868.2400 ;
        RECT 2037.3400 1862.3200 2040.3400 1862.8000 ;
        RECT 2037.3400 1856.8800 2040.3400 1857.3600 ;
        RECT 2037.3400 1851.4400 2040.3400 1851.9200 ;
        RECT 2037.3400 1873.2000 2040.3400 1873.6800 ;
        RECT 2131.9000 1835.1200 2133.5000 1835.6000 ;
        RECT 2131.9000 1840.5600 2133.5000 1841.0400 ;
        RECT 2131.9000 1818.8000 2133.5000 1819.2800 ;
        RECT 2131.9000 1824.2400 2133.5000 1824.7200 ;
        RECT 2131.9000 1829.6800 2133.5000 1830.1600 ;
        RECT 2086.9000 1835.1200 2088.5000 1835.6000 ;
        RECT 2086.9000 1840.5600 2088.5000 1841.0400 ;
        RECT 2086.9000 1818.8000 2088.5000 1819.2800 ;
        RECT 2086.9000 1824.2400 2088.5000 1824.7200 ;
        RECT 2086.9000 1829.6800 2088.5000 1830.1600 ;
        RECT 2131.9000 1807.9200 2133.5000 1808.4000 ;
        RECT 2131.9000 1813.3600 2133.5000 1813.8400 ;
        RECT 2131.9000 1791.6000 2133.5000 1792.0800 ;
        RECT 2131.9000 1797.0400 2133.5000 1797.5200 ;
        RECT 2131.9000 1802.4800 2133.5000 1802.9600 ;
        RECT 2086.9000 1807.9200 2088.5000 1808.4000 ;
        RECT 2086.9000 1813.3600 2088.5000 1813.8400 ;
        RECT 2086.9000 1791.6000 2088.5000 1792.0800 ;
        RECT 2086.9000 1797.0400 2088.5000 1797.5200 ;
        RECT 2086.9000 1802.4800 2088.5000 1802.9600 ;
        RECT 2037.3400 1835.1200 2040.3400 1835.6000 ;
        RECT 2037.3400 1840.5600 2040.3400 1841.0400 ;
        RECT 2037.3400 1824.2400 2040.3400 1824.7200 ;
        RECT 2037.3400 1818.8000 2040.3400 1819.2800 ;
        RECT 2037.3400 1829.6800 2040.3400 1830.1600 ;
        RECT 2037.3400 1807.9200 2040.3400 1808.4000 ;
        RECT 2037.3400 1813.3600 2040.3400 1813.8400 ;
        RECT 2037.3400 1797.0400 2040.3400 1797.5200 ;
        RECT 2037.3400 1791.6000 2040.3400 1792.0800 ;
        RECT 2037.3400 1802.4800 2040.3400 1802.9600 ;
        RECT 2037.3400 1846.0000 2040.3400 1846.4800 ;
        RECT 2086.9000 1846.0000 2088.5000 1846.4800 ;
        RECT 2131.9000 1846.0000 2133.5000 1846.4800 ;
        RECT 2233.4400 1780.7200 2236.4400 1781.2000 ;
        RECT 2233.4400 1786.1600 2236.4400 1786.6400 ;
        RECT 2221.9000 1780.7200 2223.5000 1781.2000 ;
        RECT 2221.9000 1786.1600 2223.5000 1786.6400 ;
        RECT 2233.4400 1764.4000 2236.4400 1764.8800 ;
        RECT 2233.4400 1769.8400 2236.4400 1770.3200 ;
        RECT 2233.4400 1775.2800 2236.4400 1775.7600 ;
        RECT 2221.9000 1764.4000 2223.5000 1764.8800 ;
        RECT 2221.9000 1769.8400 2223.5000 1770.3200 ;
        RECT 2221.9000 1775.2800 2223.5000 1775.7600 ;
        RECT 2233.4400 1753.5200 2236.4400 1754.0000 ;
        RECT 2233.4400 1758.9600 2236.4400 1759.4400 ;
        RECT 2221.9000 1753.5200 2223.5000 1754.0000 ;
        RECT 2221.9000 1758.9600 2223.5000 1759.4400 ;
        RECT 2233.4400 1737.2000 2236.4400 1737.6800 ;
        RECT 2233.4400 1742.6400 2236.4400 1743.1200 ;
        RECT 2233.4400 1748.0800 2236.4400 1748.5600 ;
        RECT 2221.9000 1737.2000 2223.5000 1737.6800 ;
        RECT 2221.9000 1742.6400 2223.5000 1743.1200 ;
        RECT 2221.9000 1748.0800 2223.5000 1748.5600 ;
        RECT 2176.9000 1780.7200 2178.5000 1781.2000 ;
        RECT 2176.9000 1786.1600 2178.5000 1786.6400 ;
        RECT 2176.9000 1764.4000 2178.5000 1764.8800 ;
        RECT 2176.9000 1769.8400 2178.5000 1770.3200 ;
        RECT 2176.9000 1775.2800 2178.5000 1775.7600 ;
        RECT 2176.9000 1753.5200 2178.5000 1754.0000 ;
        RECT 2176.9000 1758.9600 2178.5000 1759.4400 ;
        RECT 2176.9000 1737.2000 2178.5000 1737.6800 ;
        RECT 2176.9000 1742.6400 2178.5000 1743.1200 ;
        RECT 2176.9000 1748.0800 2178.5000 1748.5600 ;
        RECT 2233.4400 1726.3200 2236.4400 1726.8000 ;
        RECT 2233.4400 1731.7600 2236.4400 1732.2400 ;
        RECT 2221.9000 1726.3200 2223.5000 1726.8000 ;
        RECT 2221.9000 1731.7600 2223.5000 1732.2400 ;
        RECT 2233.4400 1710.0000 2236.4400 1710.4800 ;
        RECT 2233.4400 1715.4400 2236.4400 1715.9200 ;
        RECT 2233.4400 1720.8800 2236.4400 1721.3600 ;
        RECT 2221.9000 1710.0000 2223.5000 1710.4800 ;
        RECT 2221.9000 1715.4400 2223.5000 1715.9200 ;
        RECT 2221.9000 1720.8800 2223.5000 1721.3600 ;
        RECT 2233.4400 1699.1200 2236.4400 1699.6000 ;
        RECT 2233.4400 1704.5600 2236.4400 1705.0400 ;
        RECT 2221.9000 1699.1200 2223.5000 1699.6000 ;
        RECT 2221.9000 1704.5600 2223.5000 1705.0400 ;
        RECT 2233.4400 1693.6800 2236.4400 1694.1600 ;
        RECT 2221.9000 1693.6800 2223.5000 1694.1600 ;
        RECT 2176.9000 1726.3200 2178.5000 1726.8000 ;
        RECT 2176.9000 1731.7600 2178.5000 1732.2400 ;
        RECT 2176.9000 1710.0000 2178.5000 1710.4800 ;
        RECT 2176.9000 1715.4400 2178.5000 1715.9200 ;
        RECT 2176.9000 1720.8800 2178.5000 1721.3600 ;
        RECT 2176.9000 1699.1200 2178.5000 1699.6000 ;
        RECT 2176.9000 1704.5600 2178.5000 1705.0400 ;
        RECT 2176.9000 1693.6800 2178.5000 1694.1600 ;
        RECT 2131.9000 1780.7200 2133.5000 1781.2000 ;
        RECT 2131.9000 1786.1600 2133.5000 1786.6400 ;
        RECT 2131.9000 1764.4000 2133.5000 1764.8800 ;
        RECT 2131.9000 1769.8400 2133.5000 1770.3200 ;
        RECT 2131.9000 1775.2800 2133.5000 1775.7600 ;
        RECT 2086.9000 1780.7200 2088.5000 1781.2000 ;
        RECT 2086.9000 1786.1600 2088.5000 1786.6400 ;
        RECT 2086.9000 1764.4000 2088.5000 1764.8800 ;
        RECT 2086.9000 1769.8400 2088.5000 1770.3200 ;
        RECT 2086.9000 1775.2800 2088.5000 1775.7600 ;
        RECT 2131.9000 1753.5200 2133.5000 1754.0000 ;
        RECT 2131.9000 1758.9600 2133.5000 1759.4400 ;
        RECT 2131.9000 1737.2000 2133.5000 1737.6800 ;
        RECT 2131.9000 1742.6400 2133.5000 1743.1200 ;
        RECT 2131.9000 1748.0800 2133.5000 1748.5600 ;
        RECT 2086.9000 1753.5200 2088.5000 1754.0000 ;
        RECT 2086.9000 1758.9600 2088.5000 1759.4400 ;
        RECT 2086.9000 1737.2000 2088.5000 1737.6800 ;
        RECT 2086.9000 1742.6400 2088.5000 1743.1200 ;
        RECT 2086.9000 1748.0800 2088.5000 1748.5600 ;
        RECT 2037.3400 1780.7200 2040.3400 1781.2000 ;
        RECT 2037.3400 1786.1600 2040.3400 1786.6400 ;
        RECT 2037.3400 1769.8400 2040.3400 1770.3200 ;
        RECT 2037.3400 1764.4000 2040.3400 1764.8800 ;
        RECT 2037.3400 1775.2800 2040.3400 1775.7600 ;
        RECT 2037.3400 1753.5200 2040.3400 1754.0000 ;
        RECT 2037.3400 1758.9600 2040.3400 1759.4400 ;
        RECT 2037.3400 1742.6400 2040.3400 1743.1200 ;
        RECT 2037.3400 1737.2000 2040.3400 1737.6800 ;
        RECT 2037.3400 1748.0800 2040.3400 1748.5600 ;
        RECT 2131.9000 1726.3200 2133.5000 1726.8000 ;
        RECT 2131.9000 1731.7600 2133.5000 1732.2400 ;
        RECT 2131.9000 1710.0000 2133.5000 1710.4800 ;
        RECT 2131.9000 1715.4400 2133.5000 1715.9200 ;
        RECT 2131.9000 1720.8800 2133.5000 1721.3600 ;
        RECT 2086.9000 1726.3200 2088.5000 1726.8000 ;
        RECT 2086.9000 1731.7600 2088.5000 1732.2400 ;
        RECT 2086.9000 1710.0000 2088.5000 1710.4800 ;
        RECT 2086.9000 1715.4400 2088.5000 1715.9200 ;
        RECT 2086.9000 1720.8800 2088.5000 1721.3600 ;
        RECT 2131.9000 1704.5600 2133.5000 1705.0400 ;
        RECT 2131.9000 1699.1200 2133.5000 1699.6000 ;
        RECT 2131.9000 1693.6800 2133.5000 1694.1600 ;
        RECT 2086.9000 1704.5600 2088.5000 1705.0400 ;
        RECT 2086.9000 1699.1200 2088.5000 1699.6000 ;
        RECT 2086.9000 1693.6800 2088.5000 1694.1600 ;
        RECT 2037.3400 1726.3200 2040.3400 1726.8000 ;
        RECT 2037.3400 1731.7600 2040.3400 1732.2400 ;
        RECT 2037.3400 1715.4400 2040.3400 1715.9200 ;
        RECT 2037.3400 1710.0000 2040.3400 1710.4800 ;
        RECT 2037.3400 1720.8800 2040.3400 1721.3600 ;
        RECT 2037.3400 1699.1200 2040.3400 1699.6000 ;
        RECT 2037.3400 1704.5600 2040.3400 1705.0400 ;
        RECT 2037.3400 1693.6800 2040.3400 1694.1600 ;
        RECT 2037.3400 1891.8700 2236.4400 1894.8700 ;
        RECT 2037.3400 1686.7700 2236.4400 1689.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 1457.1300 2223.5000 1665.2300 ;
        RECT 2176.9000 1457.1300 2178.5000 1665.2300 ;
        RECT 2131.9000 1457.1300 2133.5000 1665.2300 ;
        RECT 2086.9000 1457.1300 2088.5000 1665.2300 ;
        RECT 2233.4400 1457.1300 2236.4400 1665.2300 ;
        RECT 2037.3400 1457.1300 2040.3400 1665.2300 ;
      LAYER met3 ;
        RECT 2233.4400 1659.8800 2236.4400 1660.3600 ;
        RECT 2221.9000 1659.8800 2223.5000 1660.3600 ;
        RECT 2233.4400 1649.0000 2236.4400 1649.4800 ;
        RECT 2233.4400 1654.4400 2236.4400 1654.9200 ;
        RECT 2221.9000 1649.0000 2223.5000 1649.4800 ;
        RECT 2221.9000 1654.4400 2223.5000 1654.9200 ;
        RECT 2233.4400 1632.6800 2236.4400 1633.1600 ;
        RECT 2233.4400 1638.1200 2236.4400 1638.6000 ;
        RECT 2221.9000 1632.6800 2223.5000 1633.1600 ;
        RECT 2221.9000 1638.1200 2223.5000 1638.6000 ;
        RECT 2233.4400 1621.8000 2236.4400 1622.2800 ;
        RECT 2233.4400 1627.2400 2236.4400 1627.7200 ;
        RECT 2221.9000 1621.8000 2223.5000 1622.2800 ;
        RECT 2221.9000 1627.2400 2223.5000 1627.7200 ;
        RECT 2233.4400 1643.5600 2236.4400 1644.0400 ;
        RECT 2221.9000 1643.5600 2223.5000 1644.0400 ;
        RECT 2176.9000 1649.0000 2178.5000 1649.4800 ;
        RECT 2176.9000 1654.4400 2178.5000 1654.9200 ;
        RECT 2176.9000 1659.8800 2178.5000 1660.3600 ;
        RECT 2176.9000 1632.6800 2178.5000 1633.1600 ;
        RECT 2176.9000 1638.1200 2178.5000 1638.6000 ;
        RECT 2176.9000 1627.2400 2178.5000 1627.7200 ;
        RECT 2176.9000 1621.8000 2178.5000 1622.2800 ;
        RECT 2176.9000 1643.5600 2178.5000 1644.0400 ;
        RECT 2233.4400 1605.4800 2236.4400 1605.9600 ;
        RECT 2233.4400 1610.9200 2236.4400 1611.4000 ;
        RECT 2221.9000 1605.4800 2223.5000 1605.9600 ;
        RECT 2221.9000 1610.9200 2223.5000 1611.4000 ;
        RECT 2233.4400 1589.1600 2236.4400 1589.6400 ;
        RECT 2233.4400 1594.6000 2236.4400 1595.0800 ;
        RECT 2233.4400 1600.0400 2236.4400 1600.5200 ;
        RECT 2221.9000 1589.1600 2223.5000 1589.6400 ;
        RECT 2221.9000 1594.6000 2223.5000 1595.0800 ;
        RECT 2221.9000 1600.0400 2223.5000 1600.5200 ;
        RECT 2233.4400 1578.2800 2236.4400 1578.7600 ;
        RECT 2233.4400 1583.7200 2236.4400 1584.2000 ;
        RECT 2221.9000 1578.2800 2223.5000 1578.7600 ;
        RECT 2221.9000 1583.7200 2223.5000 1584.2000 ;
        RECT 2233.4400 1561.9600 2236.4400 1562.4400 ;
        RECT 2233.4400 1567.4000 2236.4400 1567.8800 ;
        RECT 2233.4400 1572.8400 2236.4400 1573.3200 ;
        RECT 2221.9000 1561.9600 2223.5000 1562.4400 ;
        RECT 2221.9000 1567.4000 2223.5000 1567.8800 ;
        RECT 2221.9000 1572.8400 2223.5000 1573.3200 ;
        RECT 2176.9000 1605.4800 2178.5000 1605.9600 ;
        RECT 2176.9000 1610.9200 2178.5000 1611.4000 ;
        RECT 2176.9000 1589.1600 2178.5000 1589.6400 ;
        RECT 2176.9000 1594.6000 2178.5000 1595.0800 ;
        RECT 2176.9000 1600.0400 2178.5000 1600.5200 ;
        RECT 2176.9000 1578.2800 2178.5000 1578.7600 ;
        RECT 2176.9000 1583.7200 2178.5000 1584.2000 ;
        RECT 2176.9000 1561.9600 2178.5000 1562.4400 ;
        RECT 2176.9000 1567.4000 2178.5000 1567.8800 ;
        RECT 2176.9000 1572.8400 2178.5000 1573.3200 ;
        RECT 2233.4400 1616.3600 2236.4400 1616.8400 ;
        RECT 2176.9000 1616.3600 2178.5000 1616.8400 ;
        RECT 2221.9000 1616.3600 2223.5000 1616.8400 ;
        RECT 2131.9000 1649.0000 2133.5000 1649.4800 ;
        RECT 2131.9000 1654.4400 2133.5000 1654.9200 ;
        RECT 2131.9000 1659.8800 2133.5000 1660.3600 ;
        RECT 2086.9000 1649.0000 2088.5000 1649.4800 ;
        RECT 2086.9000 1654.4400 2088.5000 1654.9200 ;
        RECT 2086.9000 1659.8800 2088.5000 1660.3600 ;
        RECT 2131.9000 1632.6800 2133.5000 1633.1600 ;
        RECT 2131.9000 1638.1200 2133.5000 1638.6000 ;
        RECT 2131.9000 1621.8000 2133.5000 1622.2800 ;
        RECT 2131.9000 1627.2400 2133.5000 1627.7200 ;
        RECT 2086.9000 1632.6800 2088.5000 1633.1600 ;
        RECT 2086.9000 1638.1200 2088.5000 1638.6000 ;
        RECT 2086.9000 1621.8000 2088.5000 1622.2800 ;
        RECT 2086.9000 1627.2400 2088.5000 1627.7200 ;
        RECT 2086.9000 1643.5600 2088.5000 1644.0400 ;
        RECT 2131.9000 1643.5600 2133.5000 1644.0400 ;
        RECT 2037.3400 1659.8800 2040.3400 1660.3600 ;
        RECT 2037.3400 1654.4400 2040.3400 1654.9200 ;
        RECT 2037.3400 1649.0000 2040.3400 1649.4800 ;
        RECT 2037.3400 1638.1200 2040.3400 1638.6000 ;
        RECT 2037.3400 1632.6800 2040.3400 1633.1600 ;
        RECT 2037.3400 1627.2400 2040.3400 1627.7200 ;
        RECT 2037.3400 1621.8000 2040.3400 1622.2800 ;
        RECT 2037.3400 1643.5600 2040.3400 1644.0400 ;
        RECT 2131.9000 1605.4800 2133.5000 1605.9600 ;
        RECT 2131.9000 1610.9200 2133.5000 1611.4000 ;
        RECT 2131.9000 1589.1600 2133.5000 1589.6400 ;
        RECT 2131.9000 1594.6000 2133.5000 1595.0800 ;
        RECT 2131.9000 1600.0400 2133.5000 1600.5200 ;
        RECT 2086.9000 1605.4800 2088.5000 1605.9600 ;
        RECT 2086.9000 1610.9200 2088.5000 1611.4000 ;
        RECT 2086.9000 1589.1600 2088.5000 1589.6400 ;
        RECT 2086.9000 1594.6000 2088.5000 1595.0800 ;
        RECT 2086.9000 1600.0400 2088.5000 1600.5200 ;
        RECT 2131.9000 1578.2800 2133.5000 1578.7600 ;
        RECT 2131.9000 1583.7200 2133.5000 1584.2000 ;
        RECT 2131.9000 1561.9600 2133.5000 1562.4400 ;
        RECT 2131.9000 1567.4000 2133.5000 1567.8800 ;
        RECT 2131.9000 1572.8400 2133.5000 1573.3200 ;
        RECT 2086.9000 1578.2800 2088.5000 1578.7600 ;
        RECT 2086.9000 1583.7200 2088.5000 1584.2000 ;
        RECT 2086.9000 1561.9600 2088.5000 1562.4400 ;
        RECT 2086.9000 1567.4000 2088.5000 1567.8800 ;
        RECT 2086.9000 1572.8400 2088.5000 1573.3200 ;
        RECT 2037.3400 1605.4800 2040.3400 1605.9600 ;
        RECT 2037.3400 1610.9200 2040.3400 1611.4000 ;
        RECT 2037.3400 1594.6000 2040.3400 1595.0800 ;
        RECT 2037.3400 1589.1600 2040.3400 1589.6400 ;
        RECT 2037.3400 1600.0400 2040.3400 1600.5200 ;
        RECT 2037.3400 1578.2800 2040.3400 1578.7600 ;
        RECT 2037.3400 1583.7200 2040.3400 1584.2000 ;
        RECT 2037.3400 1567.4000 2040.3400 1567.8800 ;
        RECT 2037.3400 1561.9600 2040.3400 1562.4400 ;
        RECT 2037.3400 1572.8400 2040.3400 1573.3200 ;
        RECT 2037.3400 1616.3600 2040.3400 1616.8400 ;
        RECT 2086.9000 1616.3600 2088.5000 1616.8400 ;
        RECT 2131.9000 1616.3600 2133.5000 1616.8400 ;
        RECT 2233.4400 1551.0800 2236.4400 1551.5600 ;
        RECT 2233.4400 1556.5200 2236.4400 1557.0000 ;
        RECT 2221.9000 1551.0800 2223.5000 1551.5600 ;
        RECT 2221.9000 1556.5200 2223.5000 1557.0000 ;
        RECT 2233.4400 1534.7600 2236.4400 1535.2400 ;
        RECT 2233.4400 1540.2000 2236.4400 1540.6800 ;
        RECT 2233.4400 1545.6400 2236.4400 1546.1200 ;
        RECT 2221.9000 1534.7600 2223.5000 1535.2400 ;
        RECT 2221.9000 1540.2000 2223.5000 1540.6800 ;
        RECT 2221.9000 1545.6400 2223.5000 1546.1200 ;
        RECT 2233.4400 1523.8800 2236.4400 1524.3600 ;
        RECT 2233.4400 1529.3200 2236.4400 1529.8000 ;
        RECT 2221.9000 1523.8800 2223.5000 1524.3600 ;
        RECT 2221.9000 1529.3200 2223.5000 1529.8000 ;
        RECT 2233.4400 1507.5600 2236.4400 1508.0400 ;
        RECT 2233.4400 1513.0000 2236.4400 1513.4800 ;
        RECT 2233.4400 1518.4400 2236.4400 1518.9200 ;
        RECT 2221.9000 1507.5600 2223.5000 1508.0400 ;
        RECT 2221.9000 1513.0000 2223.5000 1513.4800 ;
        RECT 2221.9000 1518.4400 2223.5000 1518.9200 ;
        RECT 2176.9000 1551.0800 2178.5000 1551.5600 ;
        RECT 2176.9000 1556.5200 2178.5000 1557.0000 ;
        RECT 2176.9000 1534.7600 2178.5000 1535.2400 ;
        RECT 2176.9000 1540.2000 2178.5000 1540.6800 ;
        RECT 2176.9000 1545.6400 2178.5000 1546.1200 ;
        RECT 2176.9000 1523.8800 2178.5000 1524.3600 ;
        RECT 2176.9000 1529.3200 2178.5000 1529.8000 ;
        RECT 2176.9000 1507.5600 2178.5000 1508.0400 ;
        RECT 2176.9000 1513.0000 2178.5000 1513.4800 ;
        RECT 2176.9000 1518.4400 2178.5000 1518.9200 ;
        RECT 2233.4400 1496.6800 2236.4400 1497.1600 ;
        RECT 2233.4400 1502.1200 2236.4400 1502.6000 ;
        RECT 2221.9000 1496.6800 2223.5000 1497.1600 ;
        RECT 2221.9000 1502.1200 2223.5000 1502.6000 ;
        RECT 2233.4400 1480.3600 2236.4400 1480.8400 ;
        RECT 2233.4400 1485.8000 2236.4400 1486.2800 ;
        RECT 2233.4400 1491.2400 2236.4400 1491.7200 ;
        RECT 2221.9000 1480.3600 2223.5000 1480.8400 ;
        RECT 2221.9000 1485.8000 2223.5000 1486.2800 ;
        RECT 2221.9000 1491.2400 2223.5000 1491.7200 ;
        RECT 2233.4400 1469.4800 2236.4400 1469.9600 ;
        RECT 2233.4400 1474.9200 2236.4400 1475.4000 ;
        RECT 2221.9000 1469.4800 2223.5000 1469.9600 ;
        RECT 2221.9000 1474.9200 2223.5000 1475.4000 ;
        RECT 2233.4400 1464.0400 2236.4400 1464.5200 ;
        RECT 2221.9000 1464.0400 2223.5000 1464.5200 ;
        RECT 2176.9000 1496.6800 2178.5000 1497.1600 ;
        RECT 2176.9000 1502.1200 2178.5000 1502.6000 ;
        RECT 2176.9000 1480.3600 2178.5000 1480.8400 ;
        RECT 2176.9000 1485.8000 2178.5000 1486.2800 ;
        RECT 2176.9000 1491.2400 2178.5000 1491.7200 ;
        RECT 2176.9000 1469.4800 2178.5000 1469.9600 ;
        RECT 2176.9000 1474.9200 2178.5000 1475.4000 ;
        RECT 2176.9000 1464.0400 2178.5000 1464.5200 ;
        RECT 2131.9000 1551.0800 2133.5000 1551.5600 ;
        RECT 2131.9000 1556.5200 2133.5000 1557.0000 ;
        RECT 2131.9000 1534.7600 2133.5000 1535.2400 ;
        RECT 2131.9000 1540.2000 2133.5000 1540.6800 ;
        RECT 2131.9000 1545.6400 2133.5000 1546.1200 ;
        RECT 2086.9000 1551.0800 2088.5000 1551.5600 ;
        RECT 2086.9000 1556.5200 2088.5000 1557.0000 ;
        RECT 2086.9000 1534.7600 2088.5000 1535.2400 ;
        RECT 2086.9000 1540.2000 2088.5000 1540.6800 ;
        RECT 2086.9000 1545.6400 2088.5000 1546.1200 ;
        RECT 2131.9000 1523.8800 2133.5000 1524.3600 ;
        RECT 2131.9000 1529.3200 2133.5000 1529.8000 ;
        RECT 2131.9000 1507.5600 2133.5000 1508.0400 ;
        RECT 2131.9000 1513.0000 2133.5000 1513.4800 ;
        RECT 2131.9000 1518.4400 2133.5000 1518.9200 ;
        RECT 2086.9000 1523.8800 2088.5000 1524.3600 ;
        RECT 2086.9000 1529.3200 2088.5000 1529.8000 ;
        RECT 2086.9000 1507.5600 2088.5000 1508.0400 ;
        RECT 2086.9000 1513.0000 2088.5000 1513.4800 ;
        RECT 2086.9000 1518.4400 2088.5000 1518.9200 ;
        RECT 2037.3400 1551.0800 2040.3400 1551.5600 ;
        RECT 2037.3400 1556.5200 2040.3400 1557.0000 ;
        RECT 2037.3400 1540.2000 2040.3400 1540.6800 ;
        RECT 2037.3400 1534.7600 2040.3400 1535.2400 ;
        RECT 2037.3400 1545.6400 2040.3400 1546.1200 ;
        RECT 2037.3400 1523.8800 2040.3400 1524.3600 ;
        RECT 2037.3400 1529.3200 2040.3400 1529.8000 ;
        RECT 2037.3400 1513.0000 2040.3400 1513.4800 ;
        RECT 2037.3400 1507.5600 2040.3400 1508.0400 ;
        RECT 2037.3400 1518.4400 2040.3400 1518.9200 ;
        RECT 2131.9000 1496.6800 2133.5000 1497.1600 ;
        RECT 2131.9000 1502.1200 2133.5000 1502.6000 ;
        RECT 2131.9000 1480.3600 2133.5000 1480.8400 ;
        RECT 2131.9000 1485.8000 2133.5000 1486.2800 ;
        RECT 2131.9000 1491.2400 2133.5000 1491.7200 ;
        RECT 2086.9000 1496.6800 2088.5000 1497.1600 ;
        RECT 2086.9000 1502.1200 2088.5000 1502.6000 ;
        RECT 2086.9000 1480.3600 2088.5000 1480.8400 ;
        RECT 2086.9000 1485.8000 2088.5000 1486.2800 ;
        RECT 2086.9000 1491.2400 2088.5000 1491.7200 ;
        RECT 2131.9000 1474.9200 2133.5000 1475.4000 ;
        RECT 2131.9000 1469.4800 2133.5000 1469.9600 ;
        RECT 2131.9000 1464.0400 2133.5000 1464.5200 ;
        RECT 2086.9000 1474.9200 2088.5000 1475.4000 ;
        RECT 2086.9000 1469.4800 2088.5000 1469.9600 ;
        RECT 2086.9000 1464.0400 2088.5000 1464.5200 ;
        RECT 2037.3400 1496.6800 2040.3400 1497.1600 ;
        RECT 2037.3400 1502.1200 2040.3400 1502.6000 ;
        RECT 2037.3400 1485.8000 2040.3400 1486.2800 ;
        RECT 2037.3400 1480.3600 2040.3400 1480.8400 ;
        RECT 2037.3400 1491.2400 2040.3400 1491.7200 ;
        RECT 2037.3400 1469.4800 2040.3400 1469.9600 ;
        RECT 2037.3400 1474.9200 2040.3400 1475.4000 ;
        RECT 2037.3400 1464.0400 2040.3400 1464.5200 ;
        RECT 2037.3400 1662.2300 2236.4400 1665.2300 ;
        RECT 2037.3400 1457.1300 2236.4400 1460.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 1227.4900 2223.5000 1435.5900 ;
        RECT 2176.9000 1227.4900 2178.5000 1435.5900 ;
        RECT 2131.9000 1227.4900 2133.5000 1435.5900 ;
        RECT 2086.9000 1227.4900 2088.5000 1435.5900 ;
        RECT 2233.4400 1227.4900 2236.4400 1435.5900 ;
        RECT 2037.3400 1227.4900 2040.3400 1435.5900 ;
      LAYER met3 ;
        RECT 2233.4400 1430.2400 2236.4400 1430.7200 ;
        RECT 2221.9000 1430.2400 2223.5000 1430.7200 ;
        RECT 2233.4400 1419.3600 2236.4400 1419.8400 ;
        RECT 2233.4400 1424.8000 2236.4400 1425.2800 ;
        RECT 2221.9000 1419.3600 2223.5000 1419.8400 ;
        RECT 2221.9000 1424.8000 2223.5000 1425.2800 ;
        RECT 2233.4400 1403.0400 2236.4400 1403.5200 ;
        RECT 2233.4400 1408.4800 2236.4400 1408.9600 ;
        RECT 2221.9000 1403.0400 2223.5000 1403.5200 ;
        RECT 2221.9000 1408.4800 2223.5000 1408.9600 ;
        RECT 2233.4400 1392.1600 2236.4400 1392.6400 ;
        RECT 2233.4400 1397.6000 2236.4400 1398.0800 ;
        RECT 2221.9000 1392.1600 2223.5000 1392.6400 ;
        RECT 2221.9000 1397.6000 2223.5000 1398.0800 ;
        RECT 2233.4400 1413.9200 2236.4400 1414.4000 ;
        RECT 2221.9000 1413.9200 2223.5000 1414.4000 ;
        RECT 2176.9000 1419.3600 2178.5000 1419.8400 ;
        RECT 2176.9000 1424.8000 2178.5000 1425.2800 ;
        RECT 2176.9000 1430.2400 2178.5000 1430.7200 ;
        RECT 2176.9000 1403.0400 2178.5000 1403.5200 ;
        RECT 2176.9000 1408.4800 2178.5000 1408.9600 ;
        RECT 2176.9000 1397.6000 2178.5000 1398.0800 ;
        RECT 2176.9000 1392.1600 2178.5000 1392.6400 ;
        RECT 2176.9000 1413.9200 2178.5000 1414.4000 ;
        RECT 2233.4400 1375.8400 2236.4400 1376.3200 ;
        RECT 2233.4400 1381.2800 2236.4400 1381.7600 ;
        RECT 2221.9000 1375.8400 2223.5000 1376.3200 ;
        RECT 2221.9000 1381.2800 2223.5000 1381.7600 ;
        RECT 2233.4400 1359.5200 2236.4400 1360.0000 ;
        RECT 2233.4400 1364.9600 2236.4400 1365.4400 ;
        RECT 2233.4400 1370.4000 2236.4400 1370.8800 ;
        RECT 2221.9000 1359.5200 2223.5000 1360.0000 ;
        RECT 2221.9000 1364.9600 2223.5000 1365.4400 ;
        RECT 2221.9000 1370.4000 2223.5000 1370.8800 ;
        RECT 2233.4400 1348.6400 2236.4400 1349.1200 ;
        RECT 2233.4400 1354.0800 2236.4400 1354.5600 ;
        RECT 2221.9000 1348.6400 2223.5000 1349.1200 ;
        RECT 2221.9000 1354.0800 2223.5000 1354.5600 ;
        RECT 2233.4400 1332.3200 2236.4400 1332.8000 ;
        RECT 2233.4400 1337.7600 2236.4400 1338.2400 ;
        RECT 2233.4400 1343.2000 2236.4400 1343.6800 ;
        RECT 2221.9000 1332.3200 2223.5000 1332.8000 ;
        RECT 2221.9000 1337.7600 2223.5000 1338.2400 ;
        RECT 2221.9000 1343.2000 2223.5000 1343.6800 ;
        RECT 2176.9000 1375.8400 2178.5000 1376.3200 ;
        RECT 2176.9000 1381.2800 2178.5000 1381.7600 ;
        RECT 2176.9000 1359.5200 2178.5000 1360.0000 ;
        RECT 2176.9000 1364.9600 2178.5000 1365.4400 ;
        RECT 2176.9000 1370.4000 2178.5000 1370.8800 ;
        RECT 2176.9000 1348.6400 2178.5000 1349.1200 ;
        RECT 2176.9000 1354.0800 2178.5000 1354.5600 ;
        RECT 2176.9000 1332.3200 2178.5000 1332.8000 ;
        RECT 2176.9000 1337.7600 2178.5000 1338.2400 ;
        RECT 2176.9000 1343.2000 2178.5000 1343.6800 ;
        RECT 2233.4400 1386.7200 2236.4400 1387.2000 ;
        RECT 2176.9000 1386.7200 2178.5000 1387.2000 ;
        RECT 2221.9000 1386.7200 2223.5000 1387.2000 ;
        RECT 2131.9000 1419.3600 2133.5000 1419.8400 ;
        RECT 2131.9000 1424.8000 2133.5000 1425.2800 ;
        RECT 2131.9000 1430.2400 2133.5000 1430.7200 ;
        RECT 2086.9000 1419.3600 2088.5000 1419.8400 ;
        RECT 2086.9000 1424.8000 2088.5000 1425.2800 ;
        RECT 2086.9000 1430.2400 2088.5000 1430.7200 ;
        RECT 2131.9000 1403.0400 2133.5000 1403.5200 ;
        RECT 2131.9000 1408.4800 2133.5000 1408.9600 ;
        RECT 2131.9000 1392.1600 2133.5000 1392.6400 ;
        RECT 2131.9000 1397.6000 2133.5000 1398.0800 ;
        RECT 2086.9000 1403.0400 2088.5000 1403.5200 ;
        RECT 2086.9000 1408.4800 2088.5000 1408.9600 ;
        RECT 2086.9000 1392.1600 2088.5000 1392.6400 ;
        RECT 2086.9000 1397.6000 2088.5000 1398.0800 ;
        RECT 2086.9000 1413.9200 2088.5000 1414.4000 ;
        RECT 2131.9000 1413.9200 2133.5000 1414.4000 ;
        RECT 2037.3400 1430.2400 2040.3400 1430.7200 ;
        RECT 2037.3400 1424.8000 2040.3400 1425.2800 ;
        RECT 2037.3400 1419.3600 2040.3400 1419.8400 ;
        RECT 2037.3400 1408.4800 2040.3400 1408.9600 ;
        RECT 2037.3400 1403.0400 2040.3400 1403.5200 ;
        RECT 2037.3400 1397.6000 2040.3400 1398.0800 ;
        RECT 2037.3400 1392.1600 2040.3400 1392.6400 ;
        RECT 2037.3400 1413.9200 2040.3400 1414.4000 ;
        RECT 2131.9000 1375.8400 2133.5000 1376.3200 ;
        RECT 2131.9000 1381.2800 2133.5000 1381.7600 ;
        RECT 2131.9000 1359.5200 2133.5000 1360.0000 ;
        RECT 2131.9000 1364.9600 2133.5000 1365.4400 ;
        RECT 2131.9000 1370.4000 2133.5000 1370.8800 ;
        RECT 2086.9000 1375.8400 2088.5000 1376.3200 ;
        RECT 2086.9000 1381.2800 2088.5000 1381.7600 ;
        RECT 2086.9000 1359.5200 2088.5000 1360.0000 ;
        RECT 2086.9000 1364.9600 2088.5000 1365.4400 ;
        RECT 2086.9000 1370.4000 2088.5000 1370.8800 ;
        RECT 2131.9000 1348.6400 2133.5000 1349.1200 ;
        RECT 2131.9000 1354.0800 2133.5000 1354.5600 ;
        RECT 2131.9000 1332.3200 2133.5000 1332.8000 ;
        RECT 2131.9000 1337.7600 2133.5000 1338.2400 ;
        RECT 2131.9000 1343.2000 2133.5000 1343.6800 ;
        RECT 2086.9000 1348.6400 2088.5000 1349.1200 ;
        RECT 2086.9000 1354.0800 2088.5000 1354.5600 ;
        RECT 2086.9000 1332.3200 2088.5000 1332.8000 ;
        RECT 2086.9000 1337.7600 2088.5000 1338.2400 ;
        RECT 2086.9000 1343.2000 2088.5000 1343.6800 ;
        RECT 2037.3400 1375.8400 2040.3400 1376.3200 ;
        RECT 2037.3400 1381.2800 2040.3400 1381.7600 ;
        RECT 2037.3400 1364.9600 2040.3400 1365.4400 ;
        RECT 2037.3400 1359.5200 2040.3400 1360.0000 ;
        RECT 2037.3400 1370.4000 2040.3400 1370.8800 ;
        RECT 2037.3400 1348.6400 2040.3400 1349.1200 ;
        RECT 2037.3400 1354.0800 2040.3400 1354.5600 ;
        RECT 2037.3400 1337.7600 2040.3400 1338.2400 ;
        RECT 2037.3400 1332.3200 2040.3400 1332.8000 ;
        RECT 2037.3400 1343.2000 2040.3400 1343.6800 ;
        RECT 2037.3400 1386.7200 2040.3400 1387.2000 ;
        RECT 2086.9000 1386.7200 2088.5000 1387.2000 ;
        RECT 2131.9000 1386.7200 2133.5000 1387.2000 ;
        RECT 2233.4400 1321.4400 2236.4400 1321.9200 ;
        RECT 2233.4400 1326.8800 2236.4400 1327.3600 ;
        RECT 2221.9000 1321.4400 2223.5000 1321.9200 ;
        RECT 2221.9000 1326.8800 2223.5000 1327.3600 ;
        RECT 2233.4400 1305.1200 2236.4400 1305.6000 ;
        RECT 2233.4400 1310.5600 2236.4400 1311.0400 ;
        RECT 2233.4400 1316.0000 2236.4400 1316.4800 ;
        RECT 2221.9000 1305.1200 2223.5000 1305.6000 ;
        RECT 2221.9000 1310.5600 2223.5000 1311.0400 ;
        RECT 2221.9000 1316.0000 2223.5000 1316.4800 ;
        RECT 2233.4400 1294.2400 2236.4400 1294.7200 ;
        RECT 2233.4400 1299.6800 2236.4400 1300.1600 ;
        RECT 2221.9000 1294.2400 2223.5000 1294.7200 ;
        RECT 2221.9000 1299.6800 2223.5000 1300.1600 ;
        RECT 2233.4400 1277.9200 2236.4400 1278.4000 ;
        RECT 2233.4400 1283.3600 2236.4400 1283.8400 ;
        RECT 2233.4400 1288.8000 2236.4400 1289.2800 ;
        RECT 2221.9000 1277.9200 2223.5000 1278.4000 ;
        RECT 2221.9000 1283.3600 2223.5000 1283.8400 ;
        RECT 2221.9000 1288.8000 2223.5000 1289.2800 ;
        RECT 2176.9000 1321.4400 2178.5000 1321.9200 ;
        RECT 2176.9000 1326.8800 2178.5000 1327.3600 ;
        RECT 2176.9000 1305.1200 2178.5000 1305.6000 ;
        RECT 2176.9000 1310.5600 2178.5000 1311.0400 ;
        RECT 2176.9000 1316.0000 2178.5000 1316.4800 ;
        RECT 2176.9000 1294.2400 2178.5000 1294.7200 ;
        RECT 2176.9000 1299.6800 2178.5000 1300.1600 ;
        RECT 2176.9000 1277.9200 2178.5000 1278.4000 ;
        RECT 2176.9000 1283.3600 2178.5000 1283.8400 ;
        RECT 2176.9000 1288.8000 2178.5000 1289.2800 ;
        RECT 2233.4400 1267.0400 2236.4400 1267.5200 ;
        RECT 2233.4400 1272.4800 2236.4400 1272.9600 ;
        RECT 2221.9000 1267.0400 2223.5000 1267.5200 ;
        RECT 2221.9000 1272.4800 2223.5000 1272.9600 ;
        RECT 2233.4400 1250.7200 2236.4400 1251.2000 ;
        RECT 2233.4400 1256.1600 2236.4400 1256.6400 ;
        RECT 2233.4400 1261.6000 2236.4400 1262.0800 ;
        RECT 2221.9000 1250.7200 2223.5000 1251.2000 ;
        RECT 2221.9000 1256.1600 2223.5000 1256.6400 ;
        RECT 2221.9000 1261.6000 2223.5000 1262.0800 ;
        RECT 2233.4400 1239.8400 2236.4400 1240.3200 ;
        RECT 2233.4400 1245.2800 2236.4400 1245.7600 ;
        RECT 2221.9000 1239.8400 2223.5000 1240.3200 ;
        RECT 2221.9000 1245.2800 2223.5000 1245.7600 ;
        RECT 2233.4400 1234.4000 2236.4400 1234.8800 ;
        RECT 2221.9000 1234.4000 2223.5000 1234.8800 ;
        RECT 2176.9000 1267.0400 2178.5000 1267.5200 ;
        RECT 2176.9000 1272.4800 2178.5000 1272.9600 ;
        RECT 2176.9000 1250.7200 2178.5000 1251.2000 ;
        RECT 2176.9000 1256.1600 2178.5000 1256.6400 ;
        RECT 2176.9000 1261.6000 2178.5000 1262.0800 ;
        RECT 2176.9000 1239.8400 2178.5000 1240.3200 ;
        RECT 2176.9000 1245.2800 2178.5000 1245.7600 ;
        RECT 2176.9000 1234.4000 2178.5000 1234.8800 ;
        RECT 2131.9000 1321.4400 2133.5000 1321.9200 ;
        RECT 2131.9000 1326.8800 2133.5000 1327.3600 ;
        RECT 2131.9000 1305.1200 2133.5000 1305.6000 ;
        RECT 2131.9000 1310.5600 2133.5000 1311.0400 ;
        RECT 2131.9000 1316.0000 2133.5000 1316.4800 ;
        RECT 2086.9000 1321.4400 2088.5000 1321.9200 ;
        RECT 2086.9000 1326.8800 2088.5000 1327.3600 ;
        RECT 2086.9000 1305.1200 2088.5000 1305.6000 ;
        RECT 2086.9000 1310.5600 2088.5000 1311.0400 ;
        RECT 2086.9000 1316.0000 2088.5000 1316.4800 ;
        RECT 2131.9000 1294.2400 2133.5000 1294.7200 ;
        RECT 2131.9000 1299.6800 2133.5000 1300.1600 ;
        RECT 2131.9000 1277.9200 2133.5000 1278.4000 ;
        RECT 2131.9000 1283.3600 2133.5000 1283.8400 ;
        RECT 2131.9000 1288.8000 2133.5000 1289.2800 ;
        RECT 2086.9000 1294.2400 2088.5000 1294.7200 ;
        RECT 2086.9000 1299.6800 2088.5000 1300.1600 ;
        RECT 2086.9000 1277.9200 2088.5000 1278.4000 ;
        RECT 2086.9000 1283.3600 2088.5000 1283.8400 ;
        RECT 2086.9000 1288.8000 2088.5000 1289.2800 ;
        RECT 2037.3400 1321.4400 2040.3400 1321.9200 ;
        RECT 2037.3400 1326.8800 2040.3400 1327.3600 ;
        RECT 2037.3400 1310.5600 2040.3400 1311.0400 ;
        RECT 2037.3400 1305.1200 2040.3400 1305.6000 ;
        RECT 2037.3400 1316.0000 2040.3400 1316.4800 ;
        RECT 2037.3400 1294.2400 2040.3400 1294.7200 ;
        RECT 2037.3400 1299.6800 2040.3400 1300.1600 ;
        RECT 2037.3400 1283.3600 2040.3400 1283.8400 ;
        RECT 2037.3400 1277.9200 2040.3400 1278.4000 ;
        RECT 2037.3400 1288.8000 2040.3400 1289.2800 ;
        RECT 2131.9000 1267.0400 2133.5000 1267.5200 ;
        RECT 2131.9000 1272.4800 2133.5000 1272.9600 ;
        RECT 2131.9000 1250.7200 2133.5000 1251.2000 ;
        RECT 2131.9000 1256.1600 2133.5000 1256.6400 ;
        RECT 2131.9000 1261.6000 2133.5000 1262.0800 ;
        RECT 2086.9000 1267.0400 2088.5000 1267.5200 ;
        RECT 2086.9000 1272.4800 2088.5000 1272.9600 ;
        RECT 2086.9000 1250.7200 2088.5000 1251.2000 ;
        RECT 2086.9000 1256.1600 2088.5000 1256.6400 ;
        RECT 2086.9000 1261.6000 2088.5000 1262.0800 ;
        RECT 2131.9000 1245.2800 2133.5000 1245.7600 ;
        RECT 2131.9000 1239.8400 2133.5000 1240.3200 ;
        RECT 2131.9000 1234.4000 2133.5000 1234.8800 ;
        RECT 2086.9000 1245.2800 2088.5000 1245.7600 ;
        RECT 2086.9000 1239.8400 2088.5000 1240.3200 ;
        RECT 2086.9000 1234.4000 2088.5000 1234.8800 ;
        RECT 2037.3400 1267.0400 2040.3400 1267.5200 ;
        RECT 2037.3400 1272.4800 2040.3400 1272.9600 ;
        RECT 2037.3400 1256.1600 2040.3400 1256.6400 ;
        RECT 2037.3400 1250.7200 2040.3400 1251.2000 ;
        RECT 2037.3400 1261.6000 2040.3400 1262.0800 ;
        RECT 2037.3400 1239.8400 2040.3400 1240.3200 ;
        RECT 2037.3400 1245.2800 2040.3400 1245.7600 ;
        RECT 2037.3400 1234.4000 2040.3400 1234.8800 ;
        RECT 2037.3400 1432.5900 2236.4400 1435.5900 ;
        RECT 2037.3400 1227.4900 2236.4400 1230.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 997.8500 2223.5000 1205.9500 ;
        RECT 2176.9000 997.8500 2178.5000 1205.9500 ;
        RECT 2131.9000 997.8500 2133.5000 1205.9500 ;
        RECT 2086.9000 997.8500 2088.5000 1205.9500 ;
        RECT 2233.4400 997.8500 2236.4400 1205.9500 ;
        RECT 2037.3400 997.8500 2040.3400 1205.9500 ;
      LAYER met3 ;
        RECT 2233.4400 1200.6000 2236.4400 1201.0800 ;
        RECT 2221.9000 1200.6000 2223.5000 1201.0800 ;
        RECT 2233.4400 1189.7200 2236.4400 1190.2000 ;
        RECT 2233.4400 1195.1600 2236.4400 1195.6400 ;
        RECT 2221.9000 1189.7200 2223.5000 1190.2000 ;
        RECT 2221.9000 1195.1600 2223.5000 1195.6400 ;
        RECT 2233.4400 1173.4000 2236.4400 1173.8800 ;
        RECT 2233.4400 1178.8400 2236.4400 1179.3200 ;
        RECT 2221.9000 1173.4000 2223.5000 1173.8800 ;
        RECT 2221.9000 1178.8400 2223.5000 1179.3200 ;
        RECT 2233.4400 1162.5200 2236.4400 1163.0000 ;
        RECT 2233.4400 1167.9600 2236.4400 1168.4400 ;
        RECT 2221.9000 1162.5200 2223.5000 1163.0000 ;
        RECT 2221.9000 1167.9600 2223.5000 1168.4400 ;
        RECT 2233.4400 1184.2800 2236.4400 1184.7600 ;
        RECT 2221.9000 1184.2800 2223.5000 1184.7600 ;
        RECT 2176.9000 1189.7200 2178.5000 1190.2000 ;
        RECT 2176.9000 1195.1600 2178.5000 1195.6400 ;
        RECT 2176.9000 1200.6000 2178.5000 1201.0800 ;
        RECT 2176.9000 1173.4000 2178.5000 1173.8800 ;
        RECT 2176.9000 1178.8400 2178.5000 1179.3200 ;
        RECT 2176.9000 1167.9600 2178.5000 1168.4400 ;
        RECT 2176.9000 1162.5200 2178.5000 1163.0000 ;
        RECT 2176.9000 1184.2800 2178.5000 1184.7600 ;
        RECT 2233.4400 1146.2000 2236.4400 1146.6800 ;
        RECT 2233.4400 1151.6400 2236.4400 1152.1200 ;
        RECT 2221.9000 1146.2000 2223.5000 1146.6800 ;
        RECT 2221.9000 1151.6400 2223.5000 1152.1200 ;
        RECT 2233.4400 1129.8800 2236.4400 1130.3600 ;
        RECT 2233.4400 1135.3200 2236.4400 1135.8000 ;
        RECT 2233.4400 1140.7600 2236.4400 1141.2400 ;
        RECT 2221.9000 1129.8800 2223.5000 1130.3600 ;
        RECT 2221.9000 1135.3200 2223.5000 1135.8000 ;
        RECT 2221.9000 1140.7600 2223.5000 1141.2400 ;
        RECT 2233.4400 1119.0000 2236.4400 1119.4800 ;
        RECT 2233.4400 1124.4400 2236.4400 1124.9200 ;
        RECT 2221.9000 1119.0000 2223.5000 1119.4800 ;
        RECT 2221.9000 1124.4400 2223.5000 1124.9200 ;
        RECT 2233.4400 1102.6800 2236.4400 1103.1600 ;
        RECT 2233.4400 1108.1200 2236.4400 1108.6000 ;
        RECT 2233.4400 1113.5600 2236.4400 1114.0400 ;
        RECT 2221.9000 1102.6800 2223.5000 1103.1600 ;
        RECT 2221.9000 1108.1200 2223.5000 1108.6000 ;
        RECT 2221.9000 1113.5600 2223.5000 1114.0400 ;
        RECT 2176.9000 1146.2000 2178.5000 1146.6800 ;
        RECT 2176.9000 1151.6400 2178.5000 1152.1200 ;
        RECT 2176.9000 1129.8800 2178.5000 1130.3600 ;
        RECT 2176.9000 1135.3200 2178.5000 1135.8000 ;
        RECT 2176.9000 1140.7600 2178.5000 1141.2400 ;
        RECT 2176.9000 1119.0000 2178.5000 1119.4800 ;
        RECT 2176.9000 1124.4400 2178.5000 1124.9200 ;
        RECT 2176.9000 1102.6800 2178.5000 1103.1600 ;
        RECT 2176.9000 1108.1200 2178.5000 1108.6000 ;
        RECT 2176.9000 1113.5600 2178.5000 1114.0400 ;
        RECT 2233.4400 1157.0800 2236.4400 1157.5600 ;
        RECT 2176.9000 1157.0800 2178.5000 1157.5600 ;
        RECT 2221.9000 1157.0800 2223.5000 1157.5600 ;
        RECT 2131.9000 1189.7200 2133.5000 1190.2000 ;
        RECT 2131.9000 1195.1600 2133.5000 1195.6400 ;
        RECT 2131.9000 1200.6000 2133.5000 1201.0800 ;
        RECT 2086.9000 1189.7200 2088.5000 1190.2000 ;
        RECT 2086.9000 1195.1600 2088.5000 1195.6400 ;
        RECT 2086.9000 1200.6000 2088.5000 1201.0800 ;
        RECT 2131.9000 1173.4000 2133.5000 1173.8800 ;
        RECT 2131.9000 1178.8400 2133.5000 1179.3200 ;
        RECT 2131.9000 1162.5200 2133.5000 1163.0000 ;
        RECT 2131.9000 1167.9600 2133.5000 1168.4400 ;
        RECT 2086.9000 1173.4000 2088.5000 1173.8800 ;
        RECT 2086.9000 1178.8400 2088.5000 1179.3200 ;
        RECT 2086.9000 1162.5200 2088.5000 1163.0000 ;
        RECT 2086.9000 1167.9600 2088.5000 1168.4400 ;
        RECT 2086.9000 1184.2800 2088.5000 1184.7600 ;
        RECT 2131.9000 1184.2800 2133.5000 1184.7600 ;
        RECT 2037.3400 1200.6000 2040.3400 1201.0800 ;
        RECT 2037.3400 1195.1600 2040.3400 1195.6400 ;
        RECT 2037.3400 1189.7200 2040.3400 1190.2000 ;
        RECT 2037.3400 1178.8400 2040.3400 1179.3200 ;
        RECT 2037.3400 1173.4000 2040.3400 1173.8800 ;
        RECT 2037.3400 1167.9600 2040.3400 1168.4400 ;
        RECT 2037.3400 1162.5200 2040.3400 1163.0000 ;
        RECT 2037.3400 1184.2800 2040.3400 1184.7600 ;
        RECT 2131.9000 1146.2000 2133.5000 1146.6800 ;
        RECT 2131.9000 1151.6400 2133.5000 1152.1200 ;
        RECT 2131.9000 1129.8800 2133.5000 1130.3600 ;
        RECT 2131.9000 1135.3200 2133.5000 1135.8000 ;
        RECT 2131.9000 1140.7600 2133.5000 1141.2400 ;
        RECT 2086.9000 1146.2000 2088.5000 1146.6800 ;
        RECT 2086.9000 1151.6400 2088.5000 1152.1200 ;
        RECT 2086.9000 1129.8800 2088.5000 1130.3600 ;
        RECT 2086.9000 1135.3200 2088.5000 1135.8000 ;
        RECT 2086.9000 1140.7600 2088.5000 1141.2400 ;
        RECT 2131.9000 1119.0000 2133.5000 1119.4800 ;
        RECT 2131.9000 1124.4400 2133.5000 1124.9200 ;
        RECT 2131.9000 1102.6800 2133.5000 1103.1600 ;
        RECT 2131.9000 1108.1200 2133.5000 1108.6000 ;
        RECT 2131.9000 1113.5600 2133.5000 1114.0400 ;
        RECT 2086.9000 1119.0000 2088.5000 1119.4800 ;
        RECT 2086.9000 1124.4400 2088.5000 1124.9200 ;
        RECT 2086.9000 1102.6800 2088.5000 1103.1600 ;
        RECT 2086.9000 1108.1200 2088.5000 1108.6000 ;
        RECT 2086.9000 1113.5600 2088.5000 1114.0400 ;
        RECT 2037.3400 1146.2000 2040.3400 1146.6800 ;
        RECT 2037.3400 1151.6400 2040.3400 1152.1200 ;
        RECT 2037.3400 1135.3200 2040.3400 1135.8000 ;
        RECT 2037.3400 1129.8800 2040.3400 1130.3600 ;
        RECT 2037.3400 1140.7600 2040.3400 1141.2400 ;
        RECT 2037.3400 1119.0000 2040.3400 1119.4800 ;
        RECT 2037.3400 1124.4400 2040.3400 1124.9200 ;
        RECT 2037.3400 1108.1200 2040.3400 1108.6000 ;
        RECT 2037.3400 1102.6800 2040.3400 1103.1600 ;
        RECT 2037.3400 1113.5600 2040.3400 1114.0400 ;
        RECT 2037.3400 1157.0800 2040.3400 1157.5600 ;
        RECT 2086.9000 1157.0800 2088.5000 1157.5600 ;
        RECT 2131.9000 1157.0800 2133.5000 1157.5600 ;
        RECT 2233.4400 1091.8000 2236.4400 1092.2800 ;
        RECT 2233.4400 1097.2400 2236.4400 1097.7200 ;
        RECT 2221.9000 1091.8000 2223.5000 1092.2800 ;
        RECT 2221.9000 1097.2400 2223.5000 1097.7200 ;
        RECT 2233.4400 1075.4800 2236.4400 1075.9600 ;
        RECT 2233.4400 1080.9200 2236.4400 1081.4000 ;
        RECT 2233.4400 1086.3600 2236.4400 1086.8400 ;
        RECT 2221.9000 1075.4800 2223.5000 1075.9600 ;
        RECT 2221.9000 1080.9200 2223.5000 1081.4000 ;
        RECT 2221.9000 1086.3600 2223.5000 1086.8400 ;
        RECT 2233.4400 1064.6000 2236.4400 1065.0800 ;
        RECT 2233.4400 1070.0400 2236.4400 1070.5200 ;
        RECT 2221.9000 1064.6000 2223.5000 1065.0800 ;
        RECT 2221.9000 1070.0400 2223.5000 1070.5200 ;
        RECT 2233.4400 1048.2800 2236.4400 1048.7600 ;
        RECT 2233.4400 1053.7200 2236.4400 1054.2000 ;
        RECT 2233.4400 1059.1600 2236.4400 1059.6400 ;
        RECT 2221.9000 1048.2800 2223.5000 1048.7600 ;
        RECT 2221.9000 1053.7200 2223.5000 1054.2000 ;
        RECT 2221.9000 1059.1600 2223.5000 1059.6400 ;
        RECT 2176.9000 1091.8000 2178.5000 1092.2800 ;
        RECT 2176.9000 1097.2400 2178.5000 1097.7200 ;
        RECT 2176.9000 1075.4800 2178.5000 1075.9600 ;
        RECT 2176.9000 1080.9200 2178.5000 1081.4000 ;
        RECT 2176.9000 1086.3600 2178.5000 1086.8400 ;
        RECT 2176.9000 1064.6000 2178.5000 1065.0800 ;
        RECT 2176.9000 1070.0400 2178.5000 1070.5200 ;
        RECT 2176.9000 1048.2800 2178.5000 1048.7600 ;
        RECT 2176.9000 1053.7200 2178.5000 1054.2000 ;
        RECT 2176.9000 1059.1600 2178.5000 1059.6400 ;
        RECT 2233.4400 1037.4000 2236.4400 1037.8800 ;
        RECT 2233.4400 1042.8400 2236.4400 1043.3200 ;
        RECT 2221.9000 1037.4000 2223.5000 1037.8800 ;
        RECT 2221.9000 1042.8400 2223.5000 1043.3200 ;
        RECT 2233.4400 1021.0800 2236.4400 1021.5600 ;
        RECT 2233.4400 1026.5200 2236.4400 1027.0000 ;
        RECT 2233.4400 1031.9600 2236.4400 1032.4400 ;
        RECT 2221.9000 1021.0800 2223.5000 1021.5600 ;
        RECT 2221.9000 1026.5200 2223.5000 1027.0000 ;
        RECT 2221.9000 1031.9600 2223.5000 1032.4400 ;
        RECT 2233.4400 1010.2000 2236.4400 1010.6800 ;
        RECT 2233.4400 1015.6400 2236.4400 1016.1200 ;
        RECT 2221.9000 1010.2000 2223.5000 1010.6800 ;
        RECT 2221.9000 1015.6400 2223.5000 1016.1200 ;
        RECT 2233.4400 1004.7600 2236.4400 1005.2400 ;
        RECT 2221.9000 1004.7600 2223.5000 1005.2400 ;
        RECT 2176.9000 1037.4000 2178.5000 1037.8800 ;
        RECT 2176.9000 1042.8400 2178.5000 1043.3200 ;
        RECT 2176.9000 1021.0800 2178.5000 1021.5600 ;
        RECT 2176.9000 1026.5200 2178.5000 1027.0000 ;
        RECT 2176.9000 1031.9600 2178.5000 1032.4400 ;
        RECT 2176.9000 1010.2000 2178.5000 1010.6800 ;
        RECT 2176.9000 1015.6400 2178.5000 1016.1200 ;
        RECT 2176.9000 1004.7600 2178.5000 1005.2400 ;
        RECT 2131.9000 1091.8000 2133.5000 1092.2800 ;
        RECT 2131.9000 1097.2400 2133.5000 1097.7200 ;
        RECT 2131.9000 1075.4800 2133.5000 1075.9600 ;
        RECT 2131.9000 1080.9200 2133.5000 1081.4000 ;
        RECT 2131.9000 1086.3600 2133.5000 1086.8400 ;
        RECT 2086.9000 1091.8000 2088.5000 1092.2800 ;
        RECT 2086.9000 1097.2400 2088.5000 1097.7200 ;
        RECT 2086.9000 1075.4800 2088.5000 1075.9600 ;
        RECT 2086.9000 1080.9200 2088.5000 1081.4000 ;
        RECT 2086.9000 1086.3600 2088.5000 1086.8400 ;
        RECT 2131.9000 1064.6000 2133.5000 1065.0800 ;
        RECT 2131.9000 1070.0400 2133.5000 1070.5200 ;
        RECT 2131.9000 1048.2800 2133.5000 1048.7600 ;
        RECT 2131.9000 1053.7200 2133.5000 1054.2000 ;
        RECT 2131.9000 1059.1600 2133.5000 1059.6400 ;
        RECT 2086.9000 1064.6000 2088.5000 1065.0800 ;
        RECT 2086.9000 1070.0400 2088.5000 1070.5200 ;
        RECT 2086.9000 1048.2800 2088.5000 1048.7600 ;
        RECT 2086.9000 1053.7200 2088.5000 1054.2000 ;
        RECT 2086.9000 1059.1600 2088.5000 1059.6400 ;
        RECT 2037.3400 1091.8000 2040.3400 1092.2800 ;
        RECT 2037.3400 1097.2400 2040.3400 1097.7200 ;
        RECT 2037.3400 1080.9200 2040.3400 1081.4000 ;
        RECT 2037.3400 1075.4800 2040.3400 1075.9600 ;
        RECT 2037.3400 1086.3600 2040.3400 1086.8400 ;
        RECT 2037.3400 1064.6000 2040.3400 1065.0800 ;
        RECT 2037.3400 1070.0400 2040.3400 1070.5200 ;
        RECT 2037.3400 1053.7200 2040.3400 1054.2000 ;
        RECT 2037.3400 1048.2800 2040.3400 1048.7600 ;
        RECT 2037.3400 1059.1600 2040.3400 1059.6400 ;
        RECT 2131.9000 1037.4000 2133.5000 1037.8800 ;
        RECT 2131.9000 1042.8400 2133.5000 1043.3200 ;
        RECT 2131.9000 1021.0800 2133.5000 1021.5600 ;
        RECT 2131.9000 1026.5200 2133.5000 1027.0000 ;
        RECT 2131.9000 1031.9600 2133.5000 1032.4400 ;
        RECT 2086.9000 1037.4000 2088.5000 1037.8800 ;
        RECT 2086.9000 1042.8400 2088.5000 1043.3200 ;
        RECT 2086.9000 1021.0800 2088.5000 1021.5600 ;
        RECT 2086.9000 1026.5200 2088.5000 1027.0000 ;
        RECT 2086.9000 1031.9600 2088.5000 1032.4400 ;
        RECT 2131.9000 1015.6400 2133.5000 1016.1200 ;
        RECT 2131.9000 1010.2000 2133.5000 1010.6800 ;
        RECT 2131.9000 1004.7600 2133.5000 1005.2400 ;
        RECT 2086.9000 1015.6400 2088.5000 1016.1200 ;
        RECT 2086.9000 1010.2000 2088.5000 1010.6800 ;
        RECT 2086.9000 1004.7600 2088.5000 1005.2400 ;
        RECT 2037.3400 1037.4000 2040.3400 1037.8800 ;
        RECT 2037.3400 1042.8400 2040.3400 1043.3200 ;
        RECT 2037.3400 1026.5200 2040.3400 1027.0000 ;
        RECT 2037.3400 1021.0800 2040.3400 1021.5600 ;
        RECT 2037.3400 1031.9600 2040.3400 1032.4400 ;
        RECT 2037.3400 1010.2000 2040.3400 1010.6800 ;
        RECT 2037.3400 1015.6400 2040.3400 1016.1200 ;
        RECT 2037.3400 1004.7600 2040.3400 1005.2400 ;
        RECT 2037.3400 1202.9500 2236.4400 1205.9500 ;
        RECT 2037.3400 997.8500 2236.4400 1000.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2221.9000 768.2100 2223.5000 976.3100 ;
        RECT 2176.9000 768.2100 2178.5000 976.3100 ;
        RECT 2131.9000 768.2100 2133.5000 976.3100 ;
        RECT 2086.9000 768.2100 2088.5000 976.3100 ;
        RECT 2233.4400 768.2100 2236.4400 976.3100 ;
        RECT 2037.3400 768.2100 2040.3400 976.3100 ;
      LAYER met3 ;
        RECT 2233.4400 970.9600 2236.4400 971.4400 ;
        RECT 2221.9000 970.9600 2223.5000 971.4400 ;
        RECT 2233.4400 960.0800 2236.4400 960.5600 ;
        RECT 2233.4400 965.5200 2236.4400 966.0000 ;
        RECT 2221.9000 960.0800 2223.5000 960.5600 ;
        RECT 2221.9000 965.5200 2223.5000 966.0000 ;
        RECT 2233.4400 943.7600 2236.4400 944.2400 ;
        RECT 2233.4400 949.2000 2236.4400 949.6800 ;
        RECT 2221.9000 943.7600 2223.5000 944.2400 ;
        RECT 2221.9000 949.2000 2223.5000 949.6800 ;
        RECT 2233.4400 932.8800 2236.4400 933.3600 ;
        RECT 2233.4400 938.3200 2236.4400 938.8000 ;
        RECT 2221.9000 932.8800 2223.5000 933.3600 ;
        RECT 2221.9000 938.3200 2223.5000 938.8000 ;
        RECT 2233.4400 954.6400 2236.4400 955.1200 ;
        RECT 2221.9000 954.6400 2223.5000 955.1200 ;
        RECT 2176.9000 960.0800 2178.5000 960.5600 ;
        RECT 2176.9000 965.5200 2178.5000 966.0000 ;
        RECT 2176.9000 970.9600 2178.5000 971.4400 ;
        RECT 2176.9000 943.7600 2178.5000 944.2400 ;
        RECT 2176.9000 949.2000 2178.5000 949.6800 ;
        RECT 2176.9000 938.3200 2178.5000 938.8000 ;
        RECT 2176.9000 932.8800 2178.5000 933.3600 ;
        RECT 2176.9000 954.6400 2178.5000 955.1200 ;
        RECT 2233.4400 916.5600 2236.4400 917.0400 ;
        RECT 2233.4400 922.0000 2236.4400 922.4800 ;
        RECT 2221.9000 916.5600 2223.5000 917.0400 ;
        RECT 2221.9000 922.0000 2223.5000 922.4800 ;
        RECT 2233.4400 900.2400 2236.4400 900.7200 ;
        RECT 2233.4400 905.6800 2236.4400 906.1600 ;
        RECT 2233.4400 911.1200 2236.4400 911.6000 ;
        RECT 2221.9000 900.2400 2223.5000 900.7200 ;
        RECT 2221.9000 905.6800 2223.5000 906.1600 ;
        RECT 2221.9000 911.1200 2223.5000 911.6000 ;
        RECT 2233.4400 889.3600 2236.4400 889.8400 ;
        RECT 2233.4400 894.8000 2236.4400 895.2800 ;
        RECT 2221.9000 889.3600 2223.5000 889.8400 ;
        RECT 2221.9000 894.8000 2223.5000 895.2800 ;
        RECT 2233.4400 873.0400 2236.4400 873.5200 ;
        RECT 2233.4400 878.4800 2236.4400 878.9600 ;
        RECT 2233.4400 883.9200 2236.4400 884.4000 ;
        RECT 2221.9000 873.0400 2223.5000 873.5200 ;
        RECT 2221.9000 878.4800 2223.5000 878.9600 ;
        RECT 2221.9000 883.9200 2223.5000 884.4000 ;
        RECT 2176.9000 916.5600 2178.5000 917.0400 ;
        RECT 2176.9000 922.0000 2178.5000 922.4800 ;
        RECT 2176.9000 900.2400 2178.5000 900.7200 ;
        RECT 2176.9000 905.6800 2178.5000 906.1600 ;
        RECT 2176.9000 911.1200 2178.5000 911.6000 ;
        RECT 2176.9000 889.3600 2178.5000 889.8400 ;
        RECT 2176.9000 894.8000 2178.5000 895.2800 ;
        RECT 2176.9000 873.0400 2178.5000 873.5200 ;
        RECT 2176.9000 878.4800 2178.5000 878.9600 ;
        RECT 2176.9000 883.9200 2178.5000 884.4000 ;
        RECT 2233.4400 927.4400 2236.4400 927.9200 ;
        RECT 2176.9000 927.4400 2178.5000 927.9200 ;
        RECT 2221.9000 927.4400 2223.5000 927.9200 ;
        RECT 2131.9000 960.0800 2133.5000 960.5600 ;
        RECT 2131.9000 965.5200 2133.5000 966.0000 ;
        RECT 2131.9000 970.9600 2133.5000 971.4400 ;
        RECT 2086.9000 960.0800 2088.5000 960.5600 ;
        RECT 2086.9000 965.5200 2088.5000 966.0000 ;
        RECT 2086.9000 970.9600 2088.5000 971.4400 ;
        RECT 2131.9000 943.7600 2133.5000 944.2400 ;
        RECT 2131.9000 949.2000 2133.5000 949.6800 ;
        RECT 2131.9000 932.8800 2133.5000 933.3600 ;
        RECT 2131.9000 938.3200 2133.5000 938.8000 ;
        RECT 2086.9000 943.7600 2088.5000 944.2400 ;
        RECT 2086.9000 949.2000 2088.5000 949.6800 ;
        RECT 2086.9000 932.8800 2088.5000 933.3600 ;
        RECT 2086.9000 938.3200 2088.5000 938.8000 ;
        RECT 2086.9000 954.6400 2088.5000 955.1200 ;
        RECT 2131.9000 954.6400 2133.5000 955.1200 ;
        RECT 2037.3400 970.9600 2040.3400 971.4400 ;
        RECT 2037.3400 965.5200 2040.3400 966.0000 ;
        RECT 2037.3400 960.0800 2040.3400 960.5600 ;
        RECT 2037.3400 949.2000 2040.3400 949.6800 ;
        RECT 2037.3400 943.7600 2040.3400 944.2400 ;
        RECT 2037.3400 938.3200 2040.3400 938.8000 ;
        RECT 2037.3400 932.8800 2040.3400 933.3600 ;
        RECT 2037.3400 954.6400 2040.3400 955.1200 ;
        RECT 2131.9000 916.5600 2133.5000 917.0400 ;
        RECT 2131.9000 922.0000 2133.5000 922.4800 ;
        RECT 2131.9000 900.2400 2133.5000 900.7200 ;
        RECT 2131.9000 905.6800 2133.5000 906.1600 ;
        RECT 2131.9000 911.1200 2133.5000 911.6000 ;
        RECT 2086.9000 916.5600 2088.5000 917.0400 ;
        RECT 2086.9000 922.0000 2088.5000 922.4800 ;
        RECT 2086.9000 900.2400 2088.5000 900.7200 ;
        RECT 2086.9000 905.6800 2088.5000 906.1600 ;
        RECT 2086.9000 911.1200 2088.5000 911.6000 ;
        RECT 2131.9000 889.3600 2133.5000 889.8400 ;
        RECT 2131.9000 894.8000 2133.5000 895.2800 ;
        RECT 2131.9000 873.0400 2133.5000 873.5200 ;
        RECT 2131.9000 878.4800 2133.5000 878.9600 ;
        RECT 2131.9000 883.9200 2133.5000 884.4000 ;
        RECT 2086.9000 889.3600 2088.5000 889.8400 ;
        RECT 2086.9000 894.8000 2088.5000 895.2800 ;
        RECT 2086.9000 873.0400 2088.5000 873.5200 ;
        RECT 2086.9000 878.4800 2088.5000 878.9600 ;
        RECT 2086.9000 883.9200 2088.5000 884.4000 ;
        RECT 2037.3400 916.5600 2040.3400 917.0400 ;
        RECT 2037.3400 922.0000 2040.3400 922.4800 ;
        RECT 2037.3400 905.6800 2040.3400 906.1600 ;
        RECT 2037.3400 900.2400 2040.3400 900.7200 ;
        RECT 2037.3400 911.1200 2040.3400 911.6000 ;
        RECT 2037.3400 889.3600 2040.3400 889.8400 ;
        RECT 2037.3400 894.8000 2040.3400 895.2800 ;
        RECT 2037.3400 878.4800 2040.3400 878.9600 ;
        RECT 2037.3400 873.0400 2040.3400 873.5200 ;
        RECT 2037.3400 883.9200 2040.3400 884.4000 ;
        RECT 2037.3400 927.4400 2040.3400 927.9200 ;
        RECT 2086.9000 927.4400 2088.5000 927.9200 ;
        RECT 2131.9000 927.4400 2133.5000 927.9200 ;
        RECT 2233.4400 862.1600 2236.4400 862.6400 ;
        RECT 2233.4400 867.6000 2236.4400 868.0800 ;
        RECT 2221.9000 862.1600 2223.5000 862.6400 ;
        RECT 2221.9000 867.6000 2223.5000 868.0800 ;
        RECT 2233.4400 845.8400 2236.4400 846.3200 ;
        RECT 2233.4400 851.2800 2236.4400 851.7600 ;
        RECT 2233.4400 856.7200 2236.4400 857.2000 ;
        RECT 2221.9000 845.8400 2223.5000 846.3200 ;
        RECT 2221.9000 851.2800 2223.5000 851.7600 ;
        RECT 2221.9000 856.7200 2223.5000 857.2000 ;
        RECT 2233.4400 834.9600 2236.4400 835.4400 ;
        RECT 2233.4400 840.4000 2236.4400 840.8800 ;
        RECT 2221.9000 834.9600 2223.5000 835.4400 ;
        RECT 2221.9000 840.4000 2223.5000 840.8800 ;
        RECT 2233.4400 818.6400 2236.4400 819.1200 ;
        RECT 2233.4400 824.0800 2236.4400 824.5600 ;
        RECT 2233.4400 829.5200 2236.4400 830.0000 ;
        RECT 2221.9000 818.6400 2223.5000 819.1200 ;
        RECT 2221.9000 824.0800 2223.5000 824.5600 ;
        RECT 2221.9000 829.5200 2223.5000 830.0000 ;
        RECT 2176.9000 862.1600 2178.5000 862.6400 ;
        RECT 2176.9000 867.6000 2178.5000 868.0800 ;
        RECT 2176.9000 845.8400 2178.5000 846.3200 ;
        RECT 2176.9000 851.2800 2178.5000 851.7600 ;
        RECT 2176.9000 856.7200 2178.5000 857.2000 ;
        RECT 2176.9000 834.9600 2178.5000 835.4400 ;
        RECT 2176.9000 840.4000 2178.5000 840.8800 ;
        RECT 2176.9000 818.6400 2178.5000 819.1200 ;
        RECT 2176.9000 824.0800 2178.5000 824.5600 ;
        RECT 2176.9000 829.5200 2178.5000 830.0000 ;
        RECT 2233.4400 807.7600 2236.4400 808.2400 ;
        RECT 2233.4400 813.2000 2236.4400 813.6800 ;
        RECT 2221.9000 807.7600 2223.5000 808.2400 ;
        RECT 2221.9000 813.2000 2223.5000 813.6800 ;
        RECT 2233.4400 791.4400 2236.4400 791.9200 ;
        RECT 2233.4400 796.8800 2236.4400 797.3600 ;
        RECT 2233.4400 802.3200 2236.4400 802.8000 ;
        RECT 2221.9000 791.4400 2223.5000 791.9200 ;
        RECT 2221.9000 796.8800 2223.5000 797.3600 ;
        RECT 2221.9000 802.3200 2223.5000 802.8000 ;
        RECT 2233.4400 780.5600 2236.4400 781.0400 ;
        RECT 2233.4400 786.0000 2236.4400 786.4800 ;
        RECT 2221.9000 780.5600 2223.5000 781.0400 ;
        RECT 2221.9000 786.0000 2223.5000 786.4800 ;
        RECT 2233.4400 775.1200 2236.4400 775.6000 ;
        RECT 2221.9000 775.1200 2223.5000 775.6000 ;
        RECT 2176.9000 807.7600 2178.5000 808.2400 ;
        RECT 2176.9000 813.2000 2178.5000 813.6800 ;
        RECT 2176.9000 791.4400 2178.5000 791.9200 ;
        RECT 2176.9000 796.8800 2178.5000 797.3600 ;
        RECT 2176.9000 802.3200 2178.5000 802.8000 ;
        RECT 2176.9000 780.5600 2178.5000 781.0400 ;
        RECT 2176.9000 786.0000 2178.5000 786.4800 ;
        RECT 2176.9000 775.1200 2178.5000 775.6000 ;
        RECT 2131.9000 862.1600 2133.5000 862.6400 ;
        RECT 2131.9000 867.6000 2133.5000 868.0800 ;
        RECT 2131.9000 845.8400 2133.5000 846.3200 ;
        RECT 2131.9000 851.2800 2133.5000 851.7600 ;
        RECT 2131.9000 856.7200 2133.5000 857.2000 ;
        RECT 2086.9000 862.1600 2088.5000 862.6400 ;
        RECT 2086.9000 867.6000 2088.5000 868.0800 ;
        RECT 2086.9000 845.8400 2088.5000 846.3200 ;
        RECT 2086.9000 851.2800 2088.5000 851.7600 ;
        RECT 2086.9000 856.7200 2088.5000 857.2000 ;
        RECT 2131.9000 834.9600 2133.5000 835.4400 ;
        RECT 2131.9000 840.4000 2133.5000 840.8800 ;
        RECT 2131.9000 818.6400 2133.5000 819.1200 ;
        RECT 2131.9000 824.0800 2133.5000 824.5600 ;
        RECT 2131.9000 829.5200 2133.5000 830.0000 ;
        RECT 2086.9000 834.9600 2088.5000 835.4400 ;
        RECT 2086.9000 840.4000 2088.5000 840.8800 ;
        RECT 2086.9000 818.6400 2088.5000 819.1200 ;
        RECT 2086.9000 824.0800 2088.5000 824.5600 ;
        RECT 2086.9000 829.5200 2088.5000 830.0000 ;
        RECT 2037.3400 862.1600 2040.3400 862.6400 ;
        RECT 2037.3400 867.6000 2040.3400 868.0800 ;
        RECT 2037.3400 851.2800 2040.3400 851.7600 ;
        RECT 2037.3400 845.8400 2040.3400 846.3200 ;
        RECT 2037.3400 856.7200 2040.3400 857.2000 ;
        RECT 2037.3400 834.9600 2040.3400 835.4400 ;
        RECT 2037.3400 840.4000 2040.3400 840.8800 ;
        RECT 2037.3400 824.0800 2040.3400 824.5600 ;
        RECT 2037.3400 818.6400 2040.3400 819.1200 ;
        RECT 2037.3400 829.5200 2040.3400 830.0000 ;
        RECT 2131.9000 807.7600 2133.5000 808.2400 ;
        RECT 2131.9000 813.2000 2133.5000 813.6800 ;
        RECT 2131.9000 791.4400 2133.5000 791.9200 ;
        RECT 2131.9000 796.8800 2133.5000 797.3600 ;
        RECT 2131.9000 802.3200 2133.5000 802.8000 ;
        RECT 2086.9000 807.7600 2088.5000 808.2400 ;
        RECT 2086.9000 813.2000 2088.5000 813.6800 ;
        RECT 2086.9000 791.4400 2088.5000 791.9200 ;
        RECT 2086.9000 796.8800 2088.5000 797.3600 ;
        RECT 2086.9000 802.3200 2088.5000 802.8000 ;
        RECT 2131.9000 786.0000 2133.5000 786.4800 ;
        RECT 2131.9000 780.5600 2133.5000 781.0400 ;
        RECT 2131.9000 775.1200 2133.5000 775.6000 ;
        RECT 2086.9000 786.0000 2088.5000 786.4800 ;
        RECT 2086.9000 780.5600 2088.5000 781.0400 ;
        RECT 2086.9000 775.1200 2088.5000 775.6000 ;
        RECT 2037.3400 807.7600 2040.3400 808.2400 ;
        RECT 2037.3400 813.2000 2040.3400 813.6800 ;
        RECT 2037.3400 796.8800 2040.3400 797.3600 ;
        RECT 2037.3400 791.4400 2040.3400 791.9200 ;
        RECT 2037.3400 802.3200 2040.3400 802.8000 ;
        RECT 2037.3400 780.5600 2040.3400 781.0400 ;
        RECT 2037.3400 786.0000 2040.3400 786.4800 ;
        RECT 2037.3400 775.1200 2040.3400 775.6000 ;
        RECT 2037.3400 973.3100 2236.4400 976.3100 ;
        RECT 2037.3400 768.2100 2236.4400 771.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 6.0000 6.0000 3384.2000 9.0000 ;
        RECT 6.0000 2880.6600 3384.2000 2883.6600 ;
        RECT 6.0000 597.1400 9.0000 597.6200 ;
        RECT 6.0000 9.6200 9.0000 10.1000 ;
        RECT 6.0000 25.9400 9.0000 26.4200 ;
        RECT 6.0000 20.5000 9.0000 20.9800 ;
        RECT 6.0000 15.0600 9.0000 15.5400 ;
        RECT 6.0000 36.8200 9.0000 37.3000 ;
        RECT 6.0000 31.3800 9.0000 31.8600 ;
        RECT 6.0000 53.1400 9.0000 53.6200 ;
        RECT 6.0000 47.7000 9.0000 48.1800 ;
        RECT 6.0000 42.2600 9.0000 42.7400 ;
        RECT 6.0000 64.0200 9.0000 64.5000 ;
        RECT 6.0000 58.5800 9.0000 59.0600 ;
        RECT 6.0000 80.3400 9.0000 80.8200 ;
        RECT 6.0000 74.9000 9.0000 75.3800 ;
        RECT 6.0000 69.4600 9.0000 69.9400 ;
        RECT 6.0000 91.2200 9.0000 91.7000 ;
        RECT 6.0000 85.7800 9.0000 86.2600 ;
        RECT 6.0000 102.1000 9.0000 102.5800 ;
        RECT 6.0000 96.6600 9.0000 97.1400 ;
        RECT 6.0000 118.4200 9.0000 118.9000 ;
        RECT 6.0000 112.9800 9.0000 113.4600 ;
        RECT 6.0000 107.5400 9.0000 108.0200 ;
        RECT 6.0000 129.3000 9.0000 129.7800 ;
        RECT 6.0000 123.8600 9.0000 124.3400 ;
        RECT 6.0000 145.6200 9.0000 146.1000 ;
        RECT 6.0000 140.1800 9.0000 140.6600 ;
        RECT 6.0000 134.7400 9.0000 135.2200 ;
        RECT 6.0000 156.5000 9.0000 156.9800 ;
        RECT 6.0000 151.0600 9.0000 151.5400 ;
        RECT 6.0000 172.8200 9.0000 173.3000 ;
        RECT 6.0000 167.3800 9.0000 167.8600 ;
        RECT 6.0000 161.9400 9.0000 162.4200 ;
        RECT 6.0000 384.9800 9.0000 385.4600 ;
        RECT 6.0000 183.7000 9.0000 184.1800 ;
        RECT 6.0000 178.2600 9.0000 178.7400 ;
        RECT 6.0000 194.5800 9.0000 195.0600 ;
        RECT 6.0000 189.1400 9.0000 189.6200 ;
        RECT 6.0000 210.9000 9.0000 211.3800 ;
        RECT 6.0000 205.4600 9.0000 205.9400 ;
        RECT 6.0000 200.0200 9.0000 200.5000 ;
        RECT 6.0000 221.7800 9.0000 222.2600 ;
        RECT 6.0000 216.3400 9.0000 216.8200 ;
        RECT 6.0000 238.1000 9.0000 238.5800 ;
        RECT 6.0000 232.6600 9.0000 233.1400 ;
        RECT 6.0000 227.2200 9.0000 227.7000 ;
        RECT 6.0000 248.9800 9.0000 249.4600 ;
        RECT 6.0000 243.5400 9.0000 244.0200 ;
        RECT 6.0000 265.3000 9.0000 265.7800 ;
        RECT 6.0000 259.8600 9.0000 260.3400 ;
        RECT 6.0000 254.4200 9.0000 254.9000 ;
        RECT 6.0000 276.1800 9.0000 276.6600 ;
        RECT 6.0000 270.7400 9.0000 271.2200 ;
        RECT 6.0000 292.5000 9.0000 292.9800 ;
        RECT 6.0000 287.0600 9.0000 287.5400 ;
        RECT 6.0000 281.6200 9.0000 282.1000 ;
        RECT 6.0000 303.3800 9.0000 303.8600 ;
        RECT 6.0000 297.9400 9.0000 298.4200 ;
        RECT 6.0000 314.2600 9.0000 314.7400 ;
        RECT 6.0000 308.8200 9.0000 309.3000 ;
        RECT 6.0000 330.5800 9.0000 331.0600 ;
        RECT 6.0000 325.1400 9.0000 325.6200 ;
        RECT 6.0000 319.7000 9.0000 320.1800 ;
        RECT 6.0000 341.4600 9.0000 341.9400 ;
        RECT 6.0000 336.0200 9.0000 336.5000 ;
        RECT 6.0000 357.7800 9.0000 358.2600 ;
        RECT 6.0000 352.3400 9.0000 352.8200 ;
        RECT 6.0000 346.9000 9.0000 347.3800 ;
        RECT 6.0000 368.6600 9.0000 369.1400 ;
        RECT 6.0000 363.2200 9.0000 363.7000 ;
        RECT 6.0000 379.5400 9.0000 380.0200 ;
        RECT 6.0000 374.1000 9.0000 374.5800 ;
        RECT 6.0000 395.8600 9.0000 396.3400 ;
        RECT 6.0000 390.4200 9.0000 390.9000 ;
        RECT 6.0000 406.7400 9.0000 407.2200 ;
        RECT 6.0000 401.3000 9.0000 401.7800 ;
        RECT 6.0000 423.0600 9.0000 423.5400 ;
        RECT 6.0000 417.6200 9.0000 418.1000 ;
        RECT 6.0000 412.1800 9.0000 412.6600 ;
        RECT 6.0000 433.9400 9.0000 434.4200 ;
        RECT 6.0000 428.5000 9.0000 428.9800 ;
        RECT 6.0000 450.2600 9.0000 450.7400 ;
        RECT 6.0000 444.8200 9.0000 445.3000 ;
        RECT 6.0000 439.3800 9.0000 439.8600 ;
        RECT 6.0000 461.1400 9.0000 461.6200 ;
        RECT 6.0000 455.7000 9.0000 456.1800 ;
        RECT 6.0000 477.4600 9.0000 477.9400 ;
        RECT 6.0000 472.0200 9.0000 472.5000 ;
        RECT 6.0000 466.5800 9.0000 467.0600 ;
        RECT 6.0000 488.3400 9.0000 488.8200 ;
        RECT 6.0000 482.9000 9.0000 483.3800 ;
        RECT 6.0000 499.2200 9.0000 499.7000 ;
        RECT 6.0000 493.7800 9.0000 494.2600 ;
        RECT 6.0000 515.5400 9.0000 516.0200 ;
        RECT 6.0000 510.1000 9.0000 510.5800 ;
        RECT 6.0000 504.6600 9.0000 505.1400 ;
        RECT 6.0000 526.4200 9.0000 526.9000 ;
        RECT 6.0000 520.9800 9.0000 521.4600 ;
        RECT 6.0000 542.7400 9.0000 543.2200 ;
        RECT 6.0000 537.3000 9.0000 537.7800 ;
        RECT 6.0000 531.8600 9.0000 532.3400 ;
        RECT 6.0000 553.6200 9.0000 554.1000 ;
        RECT 6.0000 548.1800 9.0000 548.6600 ;
        RECT 6.0000 569.9400 9.0000 570.4200 ;
        RECT 6.0000 564.5000 9.0000 564.9800 ;
        RECT 6.0000 559.0600 9.0000 559.5400 ;
        RECT 6.0000 580.8200 9.0000 581.3000 ;
        RECT 6.0000 575.3800 9.0000 575.8600 ;
        RECT 6.0000 591.7000 9.0000 592.1800 ;
        RECT 6.0000 586.2600 9.0000 586.7400 ;
        RECT 6.0000 608.0200 9.0000 608.5000 ;
        RECT 6.0000 602.5800 9.0000 603.0600 ;
        RECT 6.0000 618.9000 9.0000 619.3800 ;
        RECT 6.0000 613.4600 9.0000 613.9400 ;
        RECT 6.0000 635.2200 9.0000 635.7000 ;
        RECT 6.0000 629.7800 9.0000 630.2600 ;
        RECT 6.0000 624.3400 9.0000 624.8200 ;
        RECT 6.0000 646.1000 9.0000 646.5800 ;
        RECT 6.0000 640.6600 9.0000 641.1400 ;
        RECT 6.0000 662.4200 9.0000 662.9000 ;
        RECT 6.0000 656.9800 9.0000 657.4600 ;
        RECT 6.0000 651.5400 9.0000 652.0200 ;
        RECT 6.0000 673.3000 9.0000 673.7800 ;
        RECT 6.0000 667.8600 9.0000 668.3400 ;
        RECT 6.0000 689.6200 9.0000 690.1000 ;
        RECT 6.0000 684.1800 9.0000 684.6600 ;
        RECT 6.0000 678.7400 9.0000 679.2200 ;
        RECT 6.0000 700.5000 9.0000 700.9800 ;
        RECT 6.0000 695.0600 9.0000 695.5400 ;
        RECT 6.0000 711.3800 9.0000 711.8600 ;
        RECT 6.0000 705.9400 9.0000 706.4200 ;
        RECT 6.0000 727.7000 9.0000 728.1800 ;
        RECT 6.0000 722.2600 9.0000 722.7400 ;
        RECT 6.0000 716.8200 9.0000 717.3000 ;
        RECT 6.0000 738.5800 9.0000 739.0600 ;
        RECT 6.0000 733.1400 9.0000 733.6200 ;
        RECT 6.0000 754.9000 9.0000 755.3800 ;
        RECT 6.0000 749.4600 9.0000 749.9400 ;
        RECT 6.0000 744.0200 9.0000 744.5000 ;
        RECT 6.0000 765.7800 9.0000 766.2600 ;
        RECT 6.0000 760.3400 9.0000 760.8200 ;
        RECT 6.0000 782.1000 9.0000 782.5800 ;
        RECT 6.0000 776.6600 9.0000 777.1400 ;
        RECT 6.0000 771.2200 9.0000 771.7000 ;
        RECT 6.0000 792.9800 9.0000 793.4600 ;
        RECT 6.0000 787.5400 9.0000 788.0200 ;
        RECT 6.0000 803.8600 9.0000 804.3400 ;
        RECT 6.0000 798.4200 9.0000 798.9000 ;
        RECT 6.0000 820.1800 9.0000 820.6600 ;
        RECT 6.0000 814.7400 9.0000 815.2200 ;
        RECT 6.0000 809.3000 9.0000 809.7800 ;
        RECT 6.0000 831.0600 9.0000 831.5400 ;
        RECT 6.0000 825.6200 9.0000 826.1000 ;
        RECT 6.0000 847.3800 9.0000 847.8600 ;
        RECT 6.0000 841.9400 9.0000 842.4200 ;
        RECT 6.0000 836.5000 9.0000 836.9800 ;
        RECT 6.0000 858.2600 9.0000 858.7400 ;
        RECT 6.0000 852.8200 9.0000 853.3000 ;
        RECT 6.0000 874.5800 9.0000 875.0600 ;
        RECT 6.0000 869.1400 9.0000 869.6200 ;
        RECT 6.0000 863.7000 9.0000 864.1800 ;
        RECT 6.0000 885.4600 9.0000 885.9400 ;
        RECT 6.0000 880.0200 9.0000 880.5000 ;
        RECT 6.0000 901.7800 9.0000 902.2600 ;
        RECT 6.0000 896.3400 9.0000 896.8200 ;
        RECT 6.0000 890.9000 9.0000 891.3800 ;
        RECT 6.0000 912.6600 9.0000 913.1400 ;
        RECT 6.0000 907.2200 9.0000 907.7000 ;
        RECT 6.0000 923.5400 9.0000 924.0200 ;
        RECT 6.0000 918.1000 9.0000 918.5800 ;
        RECT 6.0000 939.8600 9.0000 940.3400 ;
        RECT 6.0000 934.4200 9.0000 934.9000 ;
        RECT 6.0000 928.9800 9.0000 929.4600 ;
        RECT 6.0000 950.7400 9.0000 951.2200 ;
        RECT 6.0000 945.3000 9.0000 945.7800 ;
        RECT 6.0000 967.0600 9.0000 967.5400 ;
        RECT 6.0000 961.6200 9.0000 962.1000 ;
        RECT 6.0000 956.1800 9.0000 956.6600 ;
        RECT 6.0000 994.2600 9.0000 994.7400 ;
        RECT 6.0000 977.9400 9.0000 978.4200 ;
        RECT 6.0000 972.5000 9.0000 972.9800 ;
        RECT 6.0000 988.8200 9.0000 989.3000 ;
        RECT 6.0000 983.3800 9.0000 983.8600 ;
        RECT 6.0000 1005.1400 9.0000 1005.6200 ;
        RECT 6.0000 999.7000 9.0000 1000.1800 ;
        RECT 6.0000 1016.0200 9.0000 1016.5000 ;
        RECT 6.0000 1010.5800 9.0000 1011.0600 ;
        RECT 6.0000 1032.3400 9.0000 1032.8200 ;
        RECT 6.0000 1026.9000 9.0000 1027.3800 ;
        RECT 6.0000 1021.4600 9.0000 1021.9400 ;
        RECT 6.0000 1043.2200 9.0000 1043.7000 ;
        RECT 6.0000 1037.7800 9.0000 1038.2600 ;
        RECT 6.0000 1059.5400 9.0000 1060.0200 ;
        RECT 6.0000 1054.1000 9.0000 1054.5800 ;
        RECT 6.0000 1048.6600 9.0000 1049.1400 ;
        RECT 6.0000 1070.4200 9.0000 1070.9000 ;
        RECT 6.0000 1064.9800 9.0000 1065.4600 ;
        RECT 6.0000 1086.7400 9.0000 1087.2200 ;
        RECT 6.0000 1081.3000 9.0000 1081.7800 ;
        RECT 6.0000 1075.8600 9.0000 1076.3400 ;
        RECT 6.0000 1097.6200 9.0000 1098.1000 ;
        RECT 6.0000 1092.1800 9.0000 1092.6600 ;
        RECT 6.0000 1108.5000 9.0000 1108.9800 ;
        RECT 6.0000 1103.0600 9.0000 1103.5400 ;
        RECT 6.0000 1124.8200 9.0000 1125.3000 ;
        RECT 6.0000 1119.3800 9.0000 1119.8600 ;
        RECT 6.0000 1113.9400 9.0000 1114.4200 ;
        RECT 6.0000 1135.7000 9.0000 1136.1800 ;
        RECT 6.0000 1130.2600 9.0000 1130.7400 ;
        RECT 6.0000 1152.0200 9.0000 1152.5000 ;
        RECT 6.0000 1146.5800 9.0000 1147.0600 ;
        RECT 6.0000 1141.1400 9.0000 1141.6200 ;
        RECT 6.0000 1162.9000 9.0000 1163.3800 ;
        RECT 6.0000 1157.4600 9.0000 1157.9400 ;
        RECT 6.0000 1179.2200 9.0000 1179.7000 ;
        RECT 6.0000 1173.7800 9.0000 1174.2600 ;
        RECT 6.0000 1168.3400 9.0000 1168.8200 ;
        RECT 6.0000 1206.4200 9.0000 1206.9000 ;
        RECT 6.0000 1190.1000 9.0000 1190.5800 ;
        RECT 6.0000 1184.6600 9.0000 1185.1400 ;
        RECT 6.0000 1200.9800 9.0000 1201.4600 ;
        RECT 6.0000 1195.5400 9.0000 1196.0200 ;
        RECT 6.0000 1217.3000 9.0000 1217.7800 ;
        RECT 6.0000 1211.8600 9.0000 1212.3400 ;
        RECT 6.0000 1228.1800 9.0000 1228.6600 ;
        RECT 6.0000 1222.7400 9.0000 1223.2200 ;
        RECT 6.0000 1244.5000 9.0000 1244.9800 ;
        RECT 6.0000 1239.0600 9.0000 1239.5400 ;
        RECT 6.0000 1233.6200 9.0000 1234.1000 ;
        RECT 6.0000 1255.3800 9.0000 1255.8600 ;
        RECT 6.0000 1249.9400 9.0000 1250.4200 ;
        RECT 6.0000 1271.7000 9.0000 1272.1800 ;
        RECT 6.0000 1266.2600 9.0000 1266.7400 ;
        RECT 6.0000 1260.8200 9.0000 1261.3000 ;
        RECT 6.0000 1282.5800 9.0000 1283.0600 ;
        RECT 6.0000 1277.1400 9.0000 1277.6200 ;
        RECT 6.0000 1298.9000 9.0000 1299.3800 ;
        RECT 6.0000 1293.4600 9.0000 1293.9400 ;
        RECT 6.0000 1288.0200 9.0000 1288.5000 ;
        RECT 6.0000 1309.7800 9.0000 1310.2600 ;
        RECT 6.0000 1304.3400 9.0000 1304.8200 ;
        RECT 6.0000 1320.6600 9.0000 1321.1400 ;
        RECT 6.0000 1315.2200 9.0000 1315.7000 ;
        RECT 6.0000 1336.9800 9.0000 1337.4600 ;
        RECT 6.0000 1331.5400 9.0000 1332.0200 ;
        RECT 6.0000 1326.1000 9.0000 1326.5800 ;
        RECT 6.0000 1391.3800 9.0000 1391.8600 ;
        RECT 6.0000 1347.8600 9.0000 1348.3400 ;
        RECT 6.0000 1342.4200 9.0000 1342.9000 ;
        RECT 6.0000 1364.1800 9.0000 1364.6600 ;
        RECT 6.0000 1358.7400 9.0000 1359.2200 ;
        RECT 6.0000 1353.3000 9.0000 1353.7800 ;
        RECT 6.0000 1375.0600 9.0000 1375.5400 ;
        RECT 6.0000 1369.6200 9.0000 1370.1000 ;
        RECT 6.0000 1385.9400 9.0000 1386.4200 ;
        RECT 6.0000 1380.5000 9.0000 1380.9800 ;
        RECT 6.0000 1402.2600 9.0000 1402.7400 ;
        RECT 6.0000 1396.8200 9.0000 1397.3000 ;
        RECT 6.0000 1413.1400 9.0000 1413.6200 ;
        RECT 6.0000 1407.7000 9.0000 1408.1800 ;
        RECT 6.0000 1429.4600 9.0000 1429.9400 ;
        RECT 6.0000 1424.0200 9.0000 1424.5000 ;
        RECT 6.0000 1418.5800 9.0000 1419.0600 ;
        RECT 6.0000 1440.3400 9.0000 1440.8200 ;
        RECT 6.0000 1434.9000 9.0000 1435.3800 ;
        RECT 3381.2000 597.1400 3384.2000 597.6200 ;
        RECT 3381.2000 9.6200 3384.2000 10.1000 ;
        RECT 3381.2000 25.9400 3384.2000 26.4200 ;
        RECT 3381.2000 20.5000 3384.2000 20.9800 ;
        RECT 3381.2000 15.0600 3384.2000 15.5400 ;
        RECT 3381.2000 36.8200 3384.2000 37.3000 ;
        RECT 3381.2000 31.3800 3384.2000 31.8600 ;
        RECT 3381.2000 53.1400 3384.2000 53.6200 ;
        RECT 3381.2000 47.7000 3384.2000 48.1800 ;
        RECT 3381.2000 42.2600 3384.2000 42.7400 ;
        RECT 3381.2000 64.0200 3384.2000 64.5000 ;
        RECT 3381.2000 58.5800 3384.2000 59.0600 ;
        RECT 3381.2000 80.3400 3384.2000 80.8200 ;
        RECT 3381.2000 74.9000 3384.2000 75.3800 ;
        RECT 3381.2000 69.4600 3384.2000 69.9400 ;
        RECT 3381.2000 91.2200 3384.2000 91.7000 ;
        RECT 3381.2000 85.7800 3384.2000 86.2600 ;
        RECT 3381.2000 102.1000 3384.2000 102.5800 ;
        RECT 3381.2000 96.6600 3384.2000 97.1400 ;
        RECT 3381.2000 118.4200 3384.2000 118.9000 ;
        RECT 3381.2000 112.9800 3384.2000 113.4600 ;
        RECT 3381.2000 107.5400 3384.2000 108.0200 ;
        RECT 3381.2000 129.3000 3384.2000 129.7800 ;
        RECT 3381.2000 123.8600 3384.2000 124.3400 ;
        RECT 3381.2000 145.6200 3384.2000 146.1000 ;
        RECT 3381.2000 140.1800 3384.2000 140.6600 ;
        RECT 3381.2000 134.7400 3384.2000 135.2200 ;
        RECT 3381.2000 156.5000 3384.2000 156.9800 ;
        RECT 3381.2000 151.0600 3384.2000 151.5400 ;
        RECT 3381.2000 172.8200 3384.2000 173.3000 ;
        RECT 3381.2000 167.3800 3384.2000 167.8600 ;
        RECT 3381.2000 161.9400 3384.2000 162.4200 ;
        RECT 3381.2000 384.9800 3384.2000 385.4600 ;
        RECT 3381.2000 183.7000 3384.2000 184.1800 ;
        RECT 3381.2000 178.2600 3384.2000 178.7400 ;
        RECT 3381.2000 194.5800 3384.2000 195.0600 ;
        RECT 3381.2000 189.1400 3384.2000 189.6200 ;
        RECT 3381.2000 210.9000 3384.2000 211.3800 ;
        RECT 3381.2000 205.4600 3384.2000 205.9400 ;
        RECT 3381.2000 200.0200 3384.2000 200.5000 ;
        RECT 3381.2000 221.7800 3384.2000 222.2600 ;
        RECT 3381.2000 216.3400 3384.2000 216.8200 ;
        RECT 3381.2000 238.1000 3384.2000 238.5800 ;
        RECT 3381.2000 232.6600 3384.2000 233.1400 ;
        RECT 3381.2000 227.2200 3384.2000 227.7000 ;
        RECT 3381.2000 248.9800 3384.2000 249.4600 ;
        RECT 3381.2000 243.5400 3384.2000 244.0200 ;
        RECT 3381.2000 265.3000 3384.2000 265.7800 ;
        RECT 3381.2000 259.8600 3384.2000 260.3400 ;
        RECT 3381.2000 254.4200 3384.2000 254.9000 ;
        RECT 3381.2000 276.1800 3384.2000 276.6600 ;
        RECT 3381.2000 270.7400 3384.2000 271.2200 ;
        RECT 3381.2000 292.5000 3384.2000 292.9800 ;
        RECT 3381.2000 287.0600 3384.2000 287.5400 ;
        RECT 3381.2000 281.6200 3384.2000 282.1000 ;
        RECT 3381.2000 303.3800 3384.2000 303.8600 ;
        RECT 3381.2000 297.9400 3384.2000 298.4200 ;
        RECT 3381.2000 314.2600 3384.2000 314.7400 ;
        RECT 3381.2000 308.8200 3384.2000 309.3000 ;
        RECT 3381.2000 330.5800 3384.2000 331.0600 ;
        RECT 3381.2000 325.1400 3384.2000 325.6200 ;
        RECT 3381.2000 319.7000 3384.2000 320.1800 ;
        RECT 3381.2000 341.4600 3384.2000 341.9400 ;
        RECT 3381.2000 336.0200 3384.2000 336.5000 ;
        RECT 3381.2000 357.7800 3384.2000 358.2600 ;
        RECT 3381.2000 352.3400 3384.2000 352.8200 ;
        RECT 3381.2000 346.9000 3384.2000 347.3800 ;
        RECT 3381.2000 368.6600 3384.2000 369.1400 ;
        RECT 3381.2000 363.2200 3384.2000 363.7000 ;
        RECT 3381.2000 379.5400 3384.2000 380.0200 ;
        RECT 3381.2000 374.1000 3384.2000 374.5800 ;
        RECT 3381.2000 395.8600 3384.2000 396.3400 ;
        RECT 3381.2000 390.4200 3384.2000 390.9000 ;
        RECT 3381.2000 406.7400 3384.2000 407.2200 ;
        RECT 3381.2000 401.3000 3384.2000 401.7800 ;
        RECT 3381.2000 423.0600 3384.2000 423.5400 ;
        RECT 3381.2000 417.6200 3384.2000 418.1000 ;
        RECT 3381.2000 412.1800 3384.2000 412.6600 ;
        RECT 3381.2000 433.9400 3384.2000 434.4200 ;
        RECT 3381.2000 428.5000 3384.2000 428.9800 ;
        RECT 3381.2000 450.2600 3384.2000 450.7400 ;
        RECT 3381.2000 444.8200 3384.2000 445.3000 ;
        RECT 3381.2000 439.3800 3384.2000 439.8600 ;
        RECT 3381.2000 461.1400 3384.2000 461.6200 ;
        RECT 3381.2000 455.7000 3384.2000 456.1800 ;
        RECT 3381.2000 477.4600 3384.2000 477.9400 ;
        RECT 3381.2000 472.0200 3384.2000 472.5000 ;
        RECT 3381.2000 466.5800 3384.2000 467.0600 ;
        RECT 3381.2000 488.3400 3384.2000 488.8200 ;
        RECT 3381.2000 482.9000 3384.2000 483.3800 ;
        RECT 3381.2000 499.2200 3384.2000 499.7000 ;
        RECT 3381.2000 493.7800 3384.2000 494.2600 ;
        RECT 3381.2000 515.5400 3384.2000 516.0200 ;
        RECT 3381.2000 510.1000 3384.2000 510.5800 ;
        RECT 3381.2000 504.6600 3384.2000 505.1400 ;
        RECT 3381.2000 526.4200 3384.2000 526.9000 ;
        RECT 3381.2000 520.9800 3384.2000 521.4600 ;
        RECT 3381.2000 542.7400 3384.2000 543.2200 ;
        RECT 3381.2000 537.3000 3384.2000 537.7800 ;
        RECT 3381.2000 531.8600 3384.2000 532.3400 ;
        RECT 3381.2000 553.6200 3384.2000 554.1000 ;
        RECT 3381.2000 548.1800 3384.2000 548.6600 ;
        RECT 3381.2000 569.9400 3384.2000 570.4200 ;
        RECT 3381.2000 564.5000 3384.2000 564.9800 ;
        RECT 3381.2000 559.0600 3384.2000 559.5400 ;
        RECT 3381.2000 580.8200 3384.2000 581.3000 ;
        RECT 3381.2000 575.3800 3384.2000 575.8600 ;
        RECT 3381.2000 591.7000 3384.2000 592.1800 ;
        RECT 3381.2000 586.2600 3384.2000 586.7400 ;
        RECT 3381.2000 608.0200 3384.2000 608.5000 ;
        RECT 3381.2000 602.5800 3384.2000 603.0600 ;
        RECT 3381.2000 618.9000 3384.2000 619.3800 ;
        RECT 3381.2000 613.4600 3384.2000 613.9400 ;
        RECT 3381.2000 635.2200 3384.2000 635.7000 ;
        RECT 3381.2000 629.7800 3384.2000 630.2600 ;
        RECT 3381.2000 624.3400 3384.2000 624.8200 ;
        RECT 3381.2000 646.1000 3384.2000 646.5800 ;
        RECT 3381.2000 640.6600 3384.2000 641.1400 ;
        RECT 3381.2000 662.4200 3384.2000 662.9000 ;
        RECT 3381.2000 656.9800 3384.2000 657.4600 ;
        RECT 3381.2000 651.5400 3384.2000 652.0200 ;
        RECT 3381.2000 673.3000 3384.2000 673.7800 ;
        RECT 3381.2000 667.8600 3384.2000 668.3400 ;
        RECT 3381.2000 689.6200 3384.2000 690.1000 ;
        RECT 3381.2000 684.1800 3384.2000 684.6600 ;
        RECT 3381.2000 678.7400 3384.2000 679.2200 ;
        RECT 3381.2000 700.5000 3384.2000 700.9800 ;
        RECT 3381.2000 695.0600 3384.2000 695.5400 ;
        RECT 3381.2000 711.3800 3384.2000 711.8600 ;
        RECT 3381.2000 705.9400 3384.2000 706.4200 ;
        RECT 3381.2000 727.7000 3384.2000 728.1800 ;
        RECT 3381.2000 722.2600 3384.2000 722.7400 ;
        RECT 3381.2000 716.8200 3384.2000 717.3000 ;
        RECT 3381.2000 738.5800 3384.2000 739.0600 ;
        RECT 3381.2000 733.1400 3384.2000 733.6200 ;
        RECT 3381.2000 754.9000 3384.2000 755.3800 ;
        RECT 3381.2000 749.4600 3384.2000 749.9400 ;
        RECT 3381.2000 744.0200 3384.2000 744.5000 ;
        RECT 3381.2000 765.7800 3384.2000 766.2600 ;
        RECT 3381.2000 760.3400 3384.2000 760.8200 ;
        RECT 3381.2000 782.1000 3384.2000 782.5800 ;
        RECT 3381.2000 776.6600 3384.2000 777.1400 ;
        RECT 3381.2000 771.2200 3384.2000 771.7000 ;
        RECT 3381.2000 792.9800 3384.2000 793.4600 ;
        RECT 3381.2000 787.5400 3384.2000 788.0200 ;
        RECT 3381.2000 803.8600 3384.2000 804.3400 ;
        RECT 3381.2000 798.4200 3384.2000 798.9000 ;
        RECT 3381.2000 820.1800 3384.2000 820.6600 ;
        RECT 3381.2000 814.7400 3384.2000 815.2200 ;
        RECT 3381.2000 809.3000 3384.2000 809.7800 ;
        RECT 3381.2000 831.0600 3384.2000 831.5400 ;
        RECT 3381.2000 825.6200 3384.2000 826.1000 ;
        RECT 3381.2000 847.3800 3384.2000 847.8600 ;
        RECT 3381.2000 841.9400 3384.2000 842.4200 ;
        RECT 3381.2000 836.5000 3384.2000 836.9800 ;
        RECT 3381.2000 858.2600 3384.2000 858.7400 ;
        RECT 3381.2000 852.8200 3384.2000 853.3000 ;
        RECT 3381.2000 874.5800 3384.2000 875.0600 ;
        RECT 3381.2000 869.1400 3384.2000 869.6200 ;
        RECT 3381.2000 863.7000 3384.2000 864.1800 ;
        RECT 3381.2000 885.4600 3384.2000 885.9400 ;
        RECT 3381.2000 880.0200 3384.2000 880.5000 ;
        RECT 3381.2000 901.7800 3384.2000 902.2600 ;
        RECT 3381.2000 896.3400 3384.2000 896.8200 ;
        RECT 3381.2000 890.9000 3384.2000 891.3800 ;
        RECT 3381.2000 912.6600 3384.2000 913.1400 ;
        RECT 3381.2000 907.2200 3384.2000 907.7000 ;
        RECT 3381.2000 923.5400 3384.2000 924.0200 ;
        RECT 3381.2000 918.1000 3384.2000 918.5800 ;
        RECT 3381.2000 939.8600 3384.2000 940.3400 ;
        RECT 3381.2000 934.4200 3384.2000 934.9000 ;
        RECT 3381.2000 928.9800 3384.2000 929.4600 ;
        RECT 3381.2000 950.7400 3384.2000 951.2200 ;
        RECT 3381.2000 945.3000 3384.2000 945.7800 ;
        RECT 3381.2000 967.0600 3384.2000 967.5400 ;
        RECT 3381.2000 961.6200 3384.2000 962.1000 ;
        RECT 3381.2000 956.1800 3384.2000 956.6600 ;
        RECT 3381.2000 994.2600 3384.2000 994.7400 ;
        RECT 3381.2000 977.9400 3384.2000 978.4200 ;
        RECT 3381.2000 972.5000 3384.2000 972.9800 ;
        RECT 3381.2000 988.8200 3384.2000 989.3000 ;
        RECT 3381.2000 983.3800 3384.2000 983.8600 ;
        RECT 3381.2000 1005.1400 3384.2000 1005.6200 ;
        RECT 3381.2000 999.7000 3384.2000 1000.1800 ;
        RECT 3381.2000 1016.0200 3384.2000 1016.5000 ;
        RECT 3381.2000 1010.5800 3384.2000 1011.0600 ;
        RECT 3381.2000 1032.3400 3384.2000 1032.8200 ;
        RECT 3381.2000 1026.9000 3384.2000 1027.3800 ;
        RECT 3381.2000 1021.4600 3384.2000 1021.9400 ;
        RECT 3381.2000 1043.2200 3384.2000 1043.7000 ;
        RECT 3381.2000 1037.7800 3384.2000 1038.2600 ;
        RECT 3381.2000 1059.5400 3384.2000 1060.0200 ;
        RECT 3381.2000 1054.1000 3384.2000 1054.5800 ;
        RECT 3381.2000 1048.6600 3384.2000 1049.1400 ;
        RECT 3381.2000 1070.4200 3384.2000 1070.9000 ;
        RECT 3381.2000 1064.9800 3384.2000 1065.4600 ;
        RECT 3381.2000 1086.7400 3384.2000 1087.2200 ;
        RECT 3381.2000 1081.3000 3384.2000 1081.7800 ;
        RECT 3381.2000 1075.8600 3384.2000 1076.3400 ;
        RECT 3381.2000 1097.6200 3384.2000 1098.1000 ;
        RECT 3381.2000 1092.1800 3384.2000 1092.6600 ;
        RECT 3381.2000 1108.5000 3384.2000 1108.9800 ;
        RECT 3381.2000 1103.0600 3384.2000 1103.5400 ;
        RECT 3381.2000 1124.8200 3384.2000 1125.3000 ;
        RECT 3381.2000 1119.3800 3384.2000 1119.8600 ;
        RECT 3381.2000 1113.9400 3384.2000 1114.4200 ;
        RECT 3381.2000 1135.7000 3384.2000 1136.1800 ;
        RECT 3381.2000 1130.2600 3384.2000 1130.7400 ;
        RECT 3381.2000 1152.0200 3384.2000 1152.5000 ;
        RECT 3381.2000 1146.5800 3384.2000 1147.0600 ;
        RECT 3381.2000 1141.1400 3384.2000 1141.6200 ;
        RECT 3381.2000 1162.9000 3384.2000 1163.3800 ;
        RECT 3381.2000 1157.4600 3384.2000 1157.9400 ;
        RECT 3381.2000 1179.2200 3384.2000 1179.7000 ;
        RECT 3381.2000 1173.7800 3384.2000 1174.2600 ;
        RECT 3381.2000 1168.3400 3384.2000 1168.8200 ;
        RECT 3381.2000 1206.4200 3384.2000 1206.9000 ;
        RECT 3381.2000 1190.1000 3384.2000 1190.5800 ;
        RECT 3381.2000 1184.6600 3384.2000 1185.1400 ;
        RECT 3381.2000 1200.9800 3384.2000 1201.4600 ;
        RECT 3381.2000 1195.5400 3384.2000 1196.0200 ;
        RECT 3381.2000 1217.3000 3384.2000 1217.7800 ;
        RECT 3381.2000 1211.8600 3384.2000 1212.3400 ;
        RECT 3381.2000 1228.1800 3384.2000 1228.6600 ;
        RECT 3381.2000 1222.7400 3384.2000 1223.2200 ;
        RECT 3381.2000 1244.5000 3384.2000 1244.9800 ;
        RECT 3381.2000 1239.0600 3384.2000 1239.5400 ;
        RECT 3381.2000 1233.6200 3384.2000 1234.1000 ;
        RECT 3381.2000 1255.3800 3384.2000 1255.8600 ;
        RECT 3381.2000 1249.9400 3384.2000 1250.4200 ;
        RECT 3381.2000 1271.7000 3384.2000 1272.1800 ;
        RECT 3381.2000 1266.2600 3384.2000 1266.7400 ;
        RECT 3381.2000 1260.8200 3384.2000 1261.3000 ;
        RECT 3381.2000 1282.5800 3384.2000 1283.0600 ;
        RECT 3381.2000 1277.1400 3384.2000 1277.6200 ;
        RECT 3381.2000 1298.9000 3384.2000 1299.3800 ;
        RECT 3381.2000 1293.4600 3384.2000 1293.9400 ;
        RECT 3381.2000 1288.0200 3384.2000 1288.5000 ;
        RECT 3381.2000 1309.7800 3384.2000 1310.2600 ;
        RECT 3381.2000 1304.3400 3384.2000 1304.8200 ;
        RECT 3381.2000 1320.6600 3384.2000 1321.1400 ;
        RECT 3381.2000 1315.2200 3384.2000 1315.7000 ;
        RECT 3381.2000 1336.9800 3384.2000 1337.4600 ;
        RECT 3381.2000 1331.5400 3384.2000 1332.0200 ;
        RECT 3381.2000 1326.1000 3384.2000 1326.5800 ;
        RECT 3381.2000 1391.3800 3384.2000 1391.8600 ;
        RECT 3381.2000 1347.8600 3384.2000 1348.3400 ;
        RECT 3381.2000 1342.4200 3384.2000 1342.9000 ;
        RECT 3381.2000 1364.1800 3384.2000 1364.6600 ;
        RECT 3381.2000 1358.7400 3384.2000 1359.2200 ;
        RECT 3381.2000 1353.3000 3384.2000 1353.7800 ;
        RECT 3381.2000 1375.0600 3384.2000 1375.5400 ;
        RECT 3381.2000 1369.6200 3384.2000 1370.1000 ;
        RECT 3381.2000 1385.9400 3384.2000 1386.4200 ;
        RECT 3381.2000 1380.5000 3384.2000 1380.9800 ;
        RECT 3381.2000 1402.2600 3384.2000 1402.7400 ;
        RECT 3381.2000 1396.8200 3384.2000 1397.3000 ;
        RECT 3381.2000 1413.1400 3384.2000 1413.6200 ;
        RECT 3381.2000 1407.7000 3384.2000 1408.1800 ;
        RECT 3381.2000 1429.4600 3384.2000 1429.9400 ;
        RECT 3381.2000 1424.0200 3384.2000 1424.5000 ;
        RECT 3381.2000 1418.5800 3384.2000 1419.0600 ;
        RECT 3381.2000 1440.3400 3384.2000 1440.8200 ;
        RECT 3381.2000 1434.9000 3384.2000 1435.3800 ;
        RECT 6.0000 1456.6600 9.0000 1457.1400 ;
        RECT 6.0000 1451.2200 9.0000 1451.7000 ;
        RECT 6.0000 1445.7800 9.0000 1446.2600 ;
        RECT 6.0000 1467.5400 9.0000 1468.0200 ;
        RECT 6.0000 1462.1000 9.0000 1462.5800 ;
        RECT 6.0000 1483.8600 9.0000 1484.3400 ;
        RECT 6.0000 1478.4200 9.0000 1478.9000 ;
        RECT 6.0000 1472.9800 9.0000 1473.4600 ;
        RECT 6.0000 1494.7400 9.0000 1495.2200 ;
        RECT 6.0000 1489.3000 9.0000 1489.7800 ;
        RECT 6.0000 1505.6200 9.0000 1506.1000 ;
        RECT 6.0000 1500.1800 9.0000 1500.6600 ;
        RECT 6.0000 1521.9400 9.0000 1522.4200 ;
        RECT 6.0000 1516.5000 9.0000 1516.9800 ;
        RECT 6.0000 1511.0600 9.0000 1511.5400 ;
        RECT 6.0000 1532.8200 9.0000 1533.3000 ;
        RECT 6.0000 1527.3800 9.0000 1527.8600 ;
        RECT 6.0000 1549.1400 9.0000 1549.6200 ;
        RECT 6.0000 1543.7000 9.0000 1544.1800 ;
        RECT 6.0000 1538.2600 9.0000 1538.7400 ;
        RECT 6.0000 1603.5400 9.0000 1604.0200 ;
        RECT 6.0000 1560.0200 9.0000 1560.5000 ;
        RECT 6.0000 1554.5800 9.0000 1555.0600 ;
        RECT 6.0000 1576.3400 9.0000 1576.8200 ;
        RECT 6.0000 1570.9000 9.0000 1571.3800 ;
        RECT 6.0000 1565.4600 9.0000 1565.9400 ;
        RECT 6.0000 1587.2200 9.0000 1587.7000 ;
        RECT 6.0000 1581.7800 9.0000 1582.2600 ;
        RECT 6.0000 1598.1000 9.0000 1598.5800 ;
        RECT 6.0000 1592.6600 9.0000 1593.1400 ;
        RECT 6.0000 1614.4200 9.0000 1614.9000 ;
        RECT 6.0000 1608.9800 9.0000 1609.4600 ;
        RECT 6.0000 1625.3000 9.0000 1625.7800 ;
        RECT 6.0000 1619.8600 9.0000 1620.3400 ;
        RECT 6.0000 1641.6200 9.0000 1642.1000 ;
        RECT 6.0000 1636.1800 9.0000 1636.6600 ;
        RECT 6.0000 1630.7400 9.0000 1631.2200 ;
        RECT 6.0000 1652.5000 9.0000 1652.9800 ;
        RECT 6.0000 1647.0600 9.0000 1647.5400 ;
        RECT 6.0000 1668.8200 9.0000 1669.3000 ;
        RECT 6.0000 1663.3800 9.0000 1663.8600 ;
        RECT 6.0000 1657.9400 9.0000 1658.4200 ;
        RECT 6.0000 1679.7000 9.0000 1680.1800 ;
        RECT 6.0000 1674.2600 9.0000 1674.7400 ;
        RECT 6.0000 1696.0200 9.0000 1696.5000 ;
        RECT 6.0000 1690.5800 9.0000 1691.0600 ;
        RECT 6.0000 1685.1400 9.0000 1685.6200 ;
        RECT 6.0000 1706.9000 9.0000 1707.3800 ;
        RECT 6.0000 1701.4600 9.0000 1701.9400 ;
        RECT 6.0000 1717.7800 9.0000 1718.2600 ;
        RECT 6.0000 1712.3400 9.0000 1712.8200 ;
        RECT 6.0000 1734.1000 9.0000 1734.5800 ;
        RECT 6.0000 1728.6600 9.0000 1729.1400 ;
        RECT 6.0000 1723.2200 9.0000 1723.7000 ;
        RECT 6.0000 1744.9800 9.0000 1745.4600 ;
        RECT 6.0000 1739.5400 9.0000 1740.0200 ;
        RECT 6.0000 1761.3000 9.0000 1761.7800 ;
        RECT 6.0000 1755.8600 9.0000 1756.3400 ;
        RECT 6.0000 1750.4200 9.0000 1750.9000 ;
        RECT 6.0000 1772.1800 9.0000 1772.6600 ;
        RECT 6.0000 1766.7400 9.0000 1767.2200 ;
        RECT 6.0000 1788.5000 9.0000 1788.9800 ;
        RECT 6.0000 1783.0600 9.0000 1783.5400 ;
        RECT 6.0000 1777.6200 9.0000 1778.1000 ;
        RECT 6.0000 1799.3800 9.0000 1799.8600 ;
        RECT 6.0000 1793.9400 9.0000 1794.4200 ;
        RECT 6.0000 1810.2600 9.0000 1810.7400 ;
        RECT 6.0000 1804.8200 9.0000 1805.3000 ;
        RECT 6.0000 1826.5800 9.0000 1827.0600 ;
        RECT 6.0000 1821.1400 9.0000 1821.6200 ;
        RECT 6.0000 1815.7000 9.0000 1816.1800 ;
        RECT 6.0000 1837.4600 9.0000 1837.9400 ;
        RECT 6.0000 1832.0200 9.0000 1832.5000 ;
        RECT 6.0000 1853.7800 9.0000 1854.2600 ;
        RECT 6.0000 1848.3400 9.0000 1848.8200 ;
        RECT 6.0000 1842.9000 9.0000 1843.3800 ;
        RECT 6.0000 1864.6600 9.0000 1865.1400 ;
        RECT 6.0000 1859.2200 9.0000 1859.7000 ;
        RECT 6.0000 1880.9800 9.0000 1881.4600 ;
        RECT 6.0000 1875.5400 9.0000 1876.0200 ;
        RECT 6.0000 1870.1000 9.0000 1870.5800 ;
        RECT 6.0000 1891.8600 9.0000 1892.3400 ;
        RECT 6.0000 1886.4200 9.0000 1886.9000 ;
        RECT 6.0000 1908.1800 9.0000 1908.6600 ;
        RECT 6.0000 1902.7400 9.0000 1903.2200 ;
        RECT 6.0000 1897.3000 9.0000 1897.7800 ;
        RECT 6.0000 1919.0600 9.0000 1919.5400 ;
        RECT 6.0000 1913.6200 9.0000 1914.1000 ;
        RECT 6.0000 1929.9400 9.0000 1930.4200 ;
        RECT 6.0000 1924.5000 9.0000 1924.9800 ;
        RECT 6.0000 1946.2600 9.0000 1946.7400 ;
        RECT 6.0000 1940.8200 9.0000 1941.3000 ;
        RECT 6.0000 1935.3800 9.0000 1935.8600 ;
        RECT 6.0000 1957.1400 9.0000 1957.6200 ;
        RECT 6.0000 1951.7000 9.0000 1952.1800 ;
        RECT 6.0000 1973.4600 9.0000 1973.9400 ;
        RECT 6.0000 1968.0200 9.0000 1968.5000 ;
        RECT 6.0000 1962.5800 9.0000 1963.0600 ;
        RECT 6.0000 2000.6600 9.0000 2001.1400 ;
        RECT 6.0000 1984.3400 9.0000 1984.8200 ;
        RECT 6.0000 1978.9000 9.0000 1979.3800 ;
        RECT 6.0000 1995.2200 9.0000 1995.7000 ;
        RECT 6.0000 1989.7800 9.0000 1990.2600 ;
        RECT 6.0000 2011.5400 9.0000 2012.0200 ;
        RECT 6.0000 2006.1000 9.0000 2006.5800 ;
        RECT 6.0000 2022.4200 9.0000 2022.9000 ;
        RECT 6.0000 2016.9800 9.0000 2017.4600 ;
        RECT 6.0000 2038.7400 9.0000 2039.2200 ;
        RECT 6.0000 2033.3000 9.0000 2033.7800 ;
        RECT 6.0000 2027.8600 9.0000 2028.3400 ;
        RECT 6.0000 2049.6200 9.0000 2050.1000 ;
        RECT 6.0000 2044.1800 9.0000 2044.6600 ;
        RECT 6.0000 2065.9400 9.0000 2066.4200 ;
        RECT 6.0000 2060.5000 9.0000 2060.9800 ;
        RECT 6.0000 2055.0600 9.0000 2055.5400 ;
        RECT 6.0000 2076.8200 9.0000 2077.3000 ;
        RECT 6.0000 2071.3800 9.0000 2071.8600 ;
        RECT 6.0000 2093.1400 9.0000 2093.6200 ;
        RECT 6.0000 2087.7000 9.0000 2088.1800 ;
        RECT 6.0000 2082.2600 9.0000 2082.7400 ;
        RECT 6.0000 2104.0200 9.0000 2104.5000 ;
        RECT 6.0000 2098.5800 9.0000 2099.0600 ;
        RECT 6.0000 2114.9000 9.0000 2115.3800 ;
        RECT 6.0000 2109.4600 9.0000 2109.9400 ;
        RECT 6.0000 2131.2200 9.0000 2131.7000 ;
        RECT 6.0000 2125.7800 9.0000 2126.2600 ;
        RECT 6.0000 2120.3400 9.0000 2120.8200 ;
        RECT 6.0000 2142.1000 9.0000 2142.5800 ;
        RECT 6.0000 2136.6600 9.0000 2137.1400 ;
        RECT 6.0000 2158.4200 9.0000 2158.9000 ;
        RECT 6.0000 2152.9800 9.0000 2153.4600 ;
        RECT 6.0000 2147.5400 9.0000 2148.0200 ;
        RECT 6.0000 2169.3000 9.0000 2169.7800 ;
        RECT 6.0000 2163.8600 9.0000 2164.3400 ;
        RECT 6.0000 2185.6200 9.0000 2186.1000 ;
        RECT 6.0000 2180.1800 9.0000 2180.6600 ;
        RECT 6.0000 2174.7400 9.0000 2175.2200 ;
        RECT 6.0000 2212.8200 9.0000 2213.3000 ;
        RECT 6.0000 2196.5000 9.0000 2196.9800 ;
        RECT 6.0000 2191.0600 9.0000 2191.5400 ;
        RECT 6.0000 2207.3800 9.0000 2207.8600 ;
        RECT 6.0000 2201.9400 9.0000 2202.4200 ;
        RECT 6.0000 2223.7000 9.0000 2224.1800 ;
        RECT 6.0000 2218.2600 9.0000 2218.7400 ;
        RECT 6.0000 2234.5800 9.0000 2235.0600 ;
        RECT 6.0000 2229.1400 9.0000 2229.6200 ;
        RECT 6.0000 2250.9000 9.0000 2251.3800 ;
        RECT 6.0000 2245.4600 9.0000 2245.9400 ;
        RECT 6.0000 2240.0200 9.0000 2240.5000 ;
        RECT 6.0000 2261.7800 9.0000 2262.2600 ;
        RECT 6.0000 2256.3400 9.0000 2256.8200 ;
        RECT 6.0000 2278.1000 9.0000 2278.5800 ;
        RECT 6.0000 2272.6600 9.0000 2273.1400 ;
        RECT 6.0000 2267.2200 9.0000 2267.7000 ;
        RECT 6.0000 2288.9800 9.0000 2289.4600 ;
        RECT 6.0000 2283.5400 9.0000 2284.0200 ;
        RECT 6.0000 2305.3000 9.0000 2305.7800 ;
        RECT 6.0000 2299.8600 9.0000 2300.3400 ;
        RECT 6.0000 2294.4200 9.0000 2294.9000 ;
        RECT 6.0000 2316.1800 9.0000 2316.6600 ;
        RECT 6.0000 2310.7400 9.0000 2311.2200 ;
        RECT 6.0000 2327.0600 9.0000 2327.5400 ;
        RECT 6.0000 2321.6200 9.0000 2322.1000 ;
        RECT 6.0000 2343.3800 9.0000 2343.8600 ;
        RECT 6.0000 2337.9400 9.0000 2338.4200 ;
        RECT 6.0000 2332.5000 9.0000 2332.9800 ;
        RECT 6.0000 2354.2600 9.0000 2354.7400 ;
        RECT 6.0000 2348.8200 9.0000 2349.3000 ;
        RECT 6.0000 2370.5800 9.0000 2371.0600 ;
        RECT 6.0000 2365.1400 9.0000 2365.6200 ;
        RECT 6.0000 2359.7000 9.0000 2360.1800 ;
        RECT 6.0000 2381.4600 9.0000 2381.9400 ;
        RECT 6.0000 2376.0200 9.0000 2376.5000 ;
        RECT 6.0000 2397.7800 9.0000 2398.2600 ;
        RECT 6.0000 2392.3400 9.0000 2392.8200 ;
        RECT 6.0000 2386.9000 9.0000 2387.3800 ;
        RECT 6.0000 2408.6600 9.0000 2409.1400 ;
        RECT 6.0000 2403.2200 9.0000 2403.7000 ;
        RECT 6.0000 2419.5400 9.0000 2420.0200 ;
        RECT 6.0000 2414.1000 9.0000 2414.5800 ;
        RECT 6.0000 2435.8600 9.0000 2436.3400 ;
        RECT 6.0000 2430.4200 9.0000 2430.9000 ;
        RECT 6.0000 2424.9800 9.0000 2425.4600 ;
        RECT 6.0000 2446.7400 9.0000 2447.2200 ;
        RECT 6.0000 2441.3000 9.0000 2441.7800 ;
        RECT 6.0000 2463.0600 9.0000 2463.5400 ;
        RECT 6.0000 2457.6200 9.0000 2458.1000 ;
        RECT 6.0000 2452.1800 9.0000 2452.6600 ;
        RECT 6.0000 2473.9400 9.0000 2474.4200 ;
        RECT 6.0000 2468.5000 9.0000 2468.9800 ;
        RECT 6.0000 2490.2600 9.0000 2490.7400 ;
        RECT 6.0000 2484.8200 9.0000 2485.3000 ;
        RECT 6.0000 2479.3800 9.0000 2479.8600 ;
        RECT 6.0000 2501.1400 9.0000 2501.6200 ;
        RECT 6.0000 2495.7000 9.0000 2496.1800 ;
        RECT 6.0000 2609.9400 9.0000 2610.4200 ;
        RECT 6.0000 2517.4600 9.0000 2517.9400 ;
        RECT 6.0000 2512.0200 9.0000 2512.5000 ;
        RECT 6.0000 2506.5800 9.0000 2507.0600 ;
        RECT 6.0000 2528.3400 9.0000 2528.8200 ;
        RECT 6.0000 2522.9000 9.0000 2523.3800 ;
        RECT 6.0000 2539.2200 9.0000 2539.7000 ;
        RECT 6.0000 2533.7800 9.0000 2534.2600 ;
        RECT 6.0000 2555.5400 9.0000 2556.0200 ;
        RECT 6.0000 2550.1000 9.0000 2550.5800 ;
        RECT 6.0000 2544.6600 9.0000 2545.1400 ;
        RECT 6.0000 2566.4200 9.0000 2566.9000 ;
        RECT 6.0000 2560.9800 9.0000 2561.4600 ;
        RECT 6.0000 2582.7400 9.0000 2583.2200 ;
        RECT 6.0000 2577.3000 9.0000 2577.7800 ;
        RECT 6.0000 2571.8600 9.0000 2572.3400 ;
        RECT 6.0000 2593.6200 9.0000 2594.1000 ;
        RECT 6.0000 2588.1800 9.0000 2588.6600 ;
        RECT 6.0000 2604.5000 9.0000 2604.9800 ;
        RECT 6.0000 2599.0600 9.0000 2599.5400 ;
        RECT 6.0000 2620.8200 9.0000 2621.3000 ;
        RECT 6.0000 2615.3800 9.0000 2615.8600 ;
        RECT 6.0000 2631.7000 9.0000 2632.1800 ;
        RECT 6.0000 2626.2600 9.0000 2626.7400 ;
        RECT 6.0000 2648.0200 9.0000 2648.5000 ;
        RECT 6.0000 2642.5800 9.0000 2643.0600 ;
        RECT 6.0000 2637.1400 9.0000 2637.6200 ;
        RECT 6.0000 2658.9000 9.0000 2659.3800 ;
        RECT 6.0000 2653.4600 9.0000 2653.9400 ;
        RECT 6.0000 2675.2200 9.0000 2675.7000 ;
        RECT 6.0000 2669.7800 9.0000 2670.2600 ;
        RECT 6.0000 2664.3400 9.0000 2664.8200 ;
        RECT 6.0000 2686.1000 9.0000 2686.5800 ;
        RECT 6.0000 2680.6600 9.0000 2681.1400 ;
        RECT 6.0000 2702.4200 9.0000 2702.9000 ;
        RECT 6.0000 2696.9800 9.0000 2697.4600 ;
        RECT 6.0000 2691.5400 9.0000 2692.0200 ;
        RECT 6.0000 2713.3000 9.0000 2713.7800 ;
        RECT 6.0000 2707.8600 9.0000 2708.3400 ;
        RECT 6.0000 2724.1800 9.0000 2724.6600 ;
        RECT 6.0000 2718.7400 9.0000 2719.2200 ;
        RECT 6.0000 2740.5000 9.0000 2740.9800 ;
        RECT 6.0000 2735.0600 9.0000 2735.5400 ;
        RECT 6.0000 2729.6200 9.0000 2730.1000 ;
        RECT 6.0000 2751.3800 9.0000 2751.8600 ;
        RECT 6.0000 2745.9400 9.0000 2746.4200 ;
        RECT 6.0000 2767.7000 9.0000 2768.1800 ;
        RECT 6.0000 2762.2600 9.0000 2762.7400 ;
        RECT 6.0000 2756.8200 9.0000 2757.3000 ;
        RECT 6.0000 2778.5800 9.0000 2779.0600 ;
        RECT 6.0000 2773.1400 9.0000 2773.6200 ;
        RECT 6.0000 2794.9000 9.0000 2795.3800 ;
        RECT 6.0000 2789.4600 9.0000 2789.9400 ;
        RECT 6.0000 2784.0200 9.0000 2784.5000 ;
        RECT 6.0000 2805.7800 9.0000 2806.2600 ;
        RECT 6.0000 2800.3400 9.0000 2800.8200 ;
        RECT 6.0000 2816.6600 9.0000 2817.1400 ;
        RECT 6.0000 2811.2200 9.0000 2811.7000 ;
        RECT 6.0000 2832.9800 9.0000 2833.4600 ;
        RECT 6.0000 2827.5400 9.0000 2828.0200 ;
        RECT 6.0000 2822.1000 9.0000 2822.5800 ;
        RECT 6.0000 2843.8600 9.0000 2844.3400 ;
        RECT 6.0000 2838.4200 9.0000 2838.9000 ;
        RECT 6.0000 2860.1800 9.0000 2860.6600 ;
        RECT 6.0000 2854.7400 9.0000 2855.2200 ;
        RECT 6.0000 2849.3000 9.0000 2849.7800 ;
        RECT 6.0000 2871.0600 9.0000 2871.5400 ;
        RECT 6.0000 2865.6200 9.0000 2866.1000 ;
        RECT 6.0000 2876.5000 9.0000 2876.9800 ;
        RECT 3381.2000 1456.6600 3384.2000 1457.1400 ;
        RECT 3381.2000 1451.2200 3384.2000 1451.7000 ;
        RECT 3381.2000 1445.7800 3384.2000 1446.2600 ;
        RECT 3381.2000 1467.5400 3384.2000 1468.0200 ;
        RECT 3381.2000 1462.1000 3384.2000 1462.5800 ;
        RECT 3381.2000 1483.8600 3384.2000 1484.3400 ;
        RECT 3381.2000 1478.4200 3384.2000 1478.9000 ;
        RECT 3381.2000 1472.9800 3384.2000 1473.4600 ;
        RECT 3381.2000 1494.7400 3384.2000 1495.2200 ;
        RECT 3381.2000 1489.3000 3384.2000 1489.7800 ;
        RECT 3381.2000 1505.6200 3384.2000 1506.1000 ;
        RECT 3381.2000 1500.1800 3384.2000 1500.6600 ;
        RECT 3381.2000 1521.9400 3384.2000 1522.4200 ;
        RECT 3381.2000 1516.5000 3384.2000 1516.9800 ;
        RECT 3381.2000 1511.0600 3384.2000 1511.5400 ;
        RECT 3381.2000 1532.8200 3384.2000 1533.3000 ;
        RECT 3381.2000 1527.3800 3384.2000 1527.8600 ;
        RECT 3381.2000 1549.1400 3384.2000 1549.6200 ;
        RECT 3381.2000 1543.7000 3384.2000 1544.1800 ;
        RECT 3381.2000 1538.2600 3384.2000 1538.7400 ;
        RECT 3381.2000 1603.5400 3384.2000 1604.0200 ;
        RECT 3381.2000 1560.0200 3384.2000 1560.5000 ;
        RECT 3381.2000 1554.5800 3384.2000 1555.0600 ;
        RECT 3381.2000 1576.3400 3384.2000 1576.8200 ;
        RECT 3381.2000 1570.9000 3384.2000 1571.3800 ;
        RECT 3381.2000 1565.4600 3384.2000 1565.9400 ;
        RECT 3381.2000 1587.2200 3384.2000 1587.7000 ;
        RECT 3381.2000 1581.7800 3384.2000 1582.2600 ;
        RECT 3381.2000 1598.1000 3384.2000 1598.5800 ;
        RECT 3381.2000 1592.6600 3384.2000 1593.1400 ;
        RECT 3381.2000 1614.4200 3384.2000 1614.9000 ;
        RECT 3381.2000 1608.9800 3384.2000 1609.4600 ;
        RECT 3381.2000 1625.3000 3384.2000 1625.7800 ;
        RECT 3381.2000 1619.8600 3384.2000 1620.3400 ;
        RECT 3381.2000 1641.6200 3384.2000 1642.1000 ;
        RECT 3381.2000 1636.1800 3384.2000 1636.6600 ;
        RECT 3381.2000 1630.7400 3384.2000 1631.2200 ;
        RECT 3381.2000 1652.5000 3384.2000 1652.9800 ;
        RECT 3381.2000 1647.0600 3384.2000 1647.5400 ;
        RECT 3381.2000 1668.8200 3384.2000 1669.3000 ;
        RECT 3381.2000 1663.3800 3384.2000 1663.8600 ;
        RECT 3381.2000 1657.9400 3384.2000 1658.4200 ;
        RECT 3381.2000 1679.7000 3384.2000 1680.1800 ;
        RECT 3381.2000 1674.2600 3384.2000 1674.7400 ;
        RECT 3381.2000 1696.0200 3384.2000 1696.5000 ;
        RECT 3381.2000 1690.5800 3384.2000 1691.0600 ;
        RECT 3381.2000 1685.1400 3384.2000 1685.6200 ;
        RECT 3381.2000 1706.9000 3384.2000 1707.3800 ;
        RECT 3381.2000 1701.4600 3384.2000 1701.9400 ;
        RECT 3381.2000 1717.7800 3384.2000 1718.2600 ;
        RECT 3381.2000 1712.3400 3384.2000 1712.8200 ;
        RECT 3381.2000 1734.1000 3384.2000 1734.5800 ;
        RECT 3381.2000 1728.6600 3384.2000 1729.1400 ;
        RECT 3381.2000 1723.2200 3384.2000 1723.7000 ;
        RECT 3381.2000 1744.9800 3384.2000 1745.4600 ;
        RECT 3381.2000 1739.5400 3384.2000 1740.0200 ;
        RECT 3381.2000 1761.3000 3384.2000 1761.7800 ;
        RECT 3381.2000 1755.8600 3384.2000 1756.3400 ;
        RECT 3381.2000 1750.4200 3384.2000 1750.9000 ;
        RECT 3381.2000 1772.1800 3384.2000 1772.6600 ;
        RECT 3381.2000 1766.7400 3384.2000 1767.2200 ;
        RECT 3381.2000 1788.5000 3384.2000 1788.9800 ;
        RECT 3381.2000 1783.0600 3384.2000 1783.5400 ;
        RECT 3381.2000 1777.6200 3384.2000 1778.1000 ;
        RECT 3381.2000 1799.3800 3384.2000 1799.8600 ;
        RECT 3381.2000 1793.9400 3384.2000 1794.4200 ;
        RECT 3381.2000 1810.2600 3384.2000 1810.7400 ;
        RECT 3381.2000 1804.8200 3384.2000 1805.3000 ;
        RECT 3381.2000 1826.5800 3384.2000 1827.0600 ;
        RECT 3381.2000 1821.1400 3384.2000 1821.6200 ;
        RECT 3381.2000 1815.7000 3384.2000 1816.1800 ;
        RECT 3381.2000 1837.4600 3384.2000 1837.9400 ;
        RECT 3381.2000 1832.0200 3384.2000 1832.5000 ;
        RECT 3381.2000 1853.7800 3384.2000 1854.2600 ;
        RECT 3381.2000 1848.3400 3384.2000 1848.8200 ;
        RECT 3381.2000 1842.9000 3384.2000 1843.3800 ;
        RECT 3381.2000 1864.6600 3384.2000 1865.1400 ;
        RECT 3381.2000 1859.2200 3384.2000 1859.7000 ;
        RECT 3381.2000 1880.9800 3384.2000 1881.4600 ;
        RECT 3381.2000 1875.5400 3384.2000 1876.0200 ;
        RECT 3381.2000 1870.1000 3384.2000 1870.5800 ;
        RECT 3381.2000 1891.8600 3384.2000 1892.3400 ;
        RECT 3381.2000 1886.4200 3384.2000 1886.9000 ;
        RECT 3381.2000 1908.1800 3384.2000 1908.6600 ;
        RECT 3381.2000 1902.7400 3384.2000 1903.2200 ;
        RECT 3381.2000 1897.3000 3384.2000 1897.7800 ;
        RECT 3381.2000 1919.0600 3384.2000 1919.5400 ;
        RECT 3381.2000 1913.6200 3384.2000 1914.1000 ;
        RECT 3381.2000 1929.9400 3384.2000 1930.4200 ;
        RECT 3381.2000 1924.5000 3384.2000 1924.9800 ;
        RECT 3381.2000 1946.2600 3384.2000 1946.7400 ;
        RECT 3381.2000 1940.8200 3384.2000 1941.3000 ;
        RECT 3381.2000 1935.3800 3384.2000 1935.8600 ;
        RECT 3381.2000 1957.1400 3384.2000 1957.6200 ;
        RECT 3381.2000 1951.7000 3384.2000 1952.1800 ;
        RECT 3381.2000 1973.4600 3384.2000 1973.9400 ;
        RECT 3381.2000 1968.0200 3384.2000 1968.5000 ;
        RECT 3381.2000 1962.5800 3384.2000 1963.0600 ;
        RECT 3381.2000 2000.6600 3384.2000 2001.1400 ;
        RECT 3381.2000 1984.3400 3384.2000 1984.8200 ;
        RECT 3381.2000 1978.9000 3384.2000 1979.3800 ;
        RECT 3381.2000 1995.2200 3384.2000 1995.7000 ;
        RECT 3381.2000 1989.7800 3384.2000 1990.2600 ;
        RECT 3381.2000 2011.5400 3384.2000 2012.0200 ;
        RECT 3381.2000 2006.1000 3384.2000 2006.5800 ;
        RECT 3381.2000 2022.4200 3384.2000 2022.9000 ;
        RECT 3381.2000 2016.9800 3384.2000 2017.4600 ;
        RECT 3381.2000 2038.7400 3384.2000 2039.2200 ;
        RECT 3381.2000 2033.3000 3384.2000 2033.7800 ;
        RECT 3381.2000 2027.8600 3384.2000 2028.3400 ;
        RECT 3381.2000 2049.6200 3384.2000 2050.1000 ;
        RECT 3381.2000 2044.1800 3384.2000 2044.6600 ;
        RECT 3381.2000 2065.9400 3384.2000 2066.4200 ;
        RECT 3381.2000 2060.5000 3384.2000 2060.9800 ;
        RECT 3381.2000 2055.0600 3384.2000 2055.5400 ;
        RECT 3381.2000 2076.8200 3384.2000 2077.3000 ;
        RECT 3381.2000 2071.3800 3384.2000 2071.8600 ;
        RECT 3381.2000 2093.1400 3384.2000 2093.6200 ;
        RECT 3381.2000 2087.7000 3384.2000 2088.1800 ;
        RECT 3381.2000 2082.2600 3384.2000 2082.7400 ;
        RECT 3381.2000 2104.0200 3384.2000 2104.5000 ;
        RECT 3381.2000 2098.5800 3384.2000 2099.0600 ;
        RECT 3381.2000 2114.9000 3384.2000 2115.3800 ;
        RECT 3381.2000 2109.4600 3384.2000 2109.9400 ;
        RECT 3381.2000 2131.2200 3384.2000 2131.7000 ;
        RECT 3381.2000 2125.7800 3384.2000 2126.2600 ;
        RECT 3381.2000 2120.3400 3384.2000 2120.8200 ;
        RECT 3381.2000 2142.1000 3384.2000 2142.5800 ;
        RECT 3381.2000 2136.6600 3384.2000 2137.1400 ;
        RECT 3381.2000 2158.4200 3384.2000 2158.9000 ;
        RECT 3381.2000 2152.9800 3384.2000 2153.4600 ;
        RECT 3381.2000 2147.5400 3384.2000 2148.0200 ;
        RECT 3381.2000 2169.3000 3384.2000 2169.7800 ;
        RECT 3381.2000 2163.8600 3384.2000 2164.3400 ;
        RECT 3381.2000 2185.6200 3384.2000 2186.1000 ;
        RECT 3381.2000 2180.1800 3384.2000 2180.6600 ;
        RECT 3381.2000 2174.7400 3384.2000 2175.2200 ;
        RECT 3381.2000 2212.8200 3384.2000 2213.3000 ;
        RECT 3381.2000 2196.5000 3384.2000 2196.9800 ;
        RECT 3381.2000 2191.0600 3384.2000 2191.5400 ;
        RECT 3381.2000 2207.3800 3384.2000 2207.8600 ;
        RECT 3381.2000 2201.9400 3384.2000 2202.4200 ;
        RECT 3381.2000 2223.7000 3384.2000 2224.1800 ;
        RECT 3381.2000 2218.2600 3384.2000 2218.7400 ;
        RECT 3381.2000 2234.5800 3384.2000 2235.0600 ;
        RECT 3381.2000 2229.1400 3384.2000 2229.6200 ;
        RECT 3381.2000 2250.9000 3384.2000 2251.3800 ;
        RECT 3381.2000 2245.4600 3384.2000 2245.9400 ;
        RECT 3381.2000 2240.0200 3384.2000 2240.5000 ;
        RECT 3381.2000 2261.7800 3384.2000 2262.2600 ;
        RECT 3381.2000 2256.3400 3384.2000 2256.8200 ;
        RECT 3381.2000 2278.1000 3384.2000 2278.5800 ;
        RECT 3381.2000 2272.6600 3384.2000 2273.1400 ;
        RECT 3381.2000 2267.2200 3384.2000 2267.7000 ;
        RECT 3381.2000 2288.9800 3384.2000 2289.4600 ;
        RECT 3381.2000 2283.5400 3384.2000 2284.0200 ;
        RECT 3381.2000 2305.3000 3384.2000 2305.7800 ;
        RECT 3381.2000 2299.8600 3384.2000 2300.3400 ;
        RECT 3381.2000 2294.4200 3384.2000 2294.9000 ;
        RECT 3381.2000 2316.1800 3384.2000 2316.6600 ;
        RECT 3381.2000 2310.7400 3384.2000 2311.2200 ;
        RECT 3381.2000 2327.0600 3384.2000 2327.5400 ;
        RECT 3381.2000 2321.6200 3384.2000 2322.1000 ;
        RECT 3381.2000 2343.3800 3384.2000 2343.8600 ;
        RECT 3381.2000 2337.9400 3384.2000 2338.4200 ;
        RECT 3381.2000 2332.5000 3384.2000 2332.9800 ;
        RECT 3381.2000 2354.2600 3384.2000 2354.7400 ;
        RECT 3381.2000 2348.8200 3384.2000 2349.3000 ;
        RECT 3381.2000 2370.5800 3384.2000 2371.0600 ;
        RECT 3381.2000 2365.1400 3384.2000 2365.6200 ;
        RECT 3381.2000 2359.7000 3384.2000 2360.1800 ;
        RECT 3381.2000 2381.4600 3384.2000 2381.9400 ;
        RECT 3381.2000 2376.0200 3384.2000 2376.5000 ;
        RECT 3381.2000 2397.7800 3384.2000 2398.2600 ;
        RECT 3381.2000 2392.3400 3384.2000 2392.8200 ;
        RECT 3381.2000 2386.9000 3384.2000 2387.3800 ;
        RECT 3381.2000 2408.6600 3384.2000 2409.1400 ;
        RECT 3381.2000 2403.2200 3384.2000 2403.7000 ;
        RECT 3381.2000 2419.5400 3384.2000 2420.0200 ;
        RECT 3381.2000 2414.1000 3384.2000 2414.5800 ;
        RECT 3381.2000 2435.8600 3384.2000 2436.3400 ;
        RECT 3381.2000 2430.4200 3384.2000 2430.9000 ;
        RECT 3381.2000 2424.9800 3384.2000 2425.4600 ;
        RECT 3381.2000 2446.7400 3384.2000 2447.2200 ;
        RECT 3381.2000 2441.3000 3384.2000 2441.7800 ;
        RECT 3381.2000 2463.0600 3384.2000 2463.5400 ;
        RECT 3381.2000 2457.6200 3384.2000 2458.1000 ;
        RECT 3381.2000 2452.1800 3384.2000 2452.6600 ;
        RECT 3381.2000 2473.9400 3384.2000 2474.4200 ;
        RECT 3381.2000 2468.5000 3384.2000 2468.9800 ;
        RECT 3381.2000 2490.2600 3384.2000 2490.7400 ;
        RECT 3381.2000 2484.8200 3384.2000 2485.3000 ;
        RECT 3381.2000 2479.3800 3384.2000 2479.8600 ;
        RECT 3381.2000 2501.1400 3384.2000 2501.6200 ;
        RECT 3381.2000 2495.7000 3384.2000 2496.1800 ;
        RECT 3381.2000 2609.9400 3384.2000 2610.4200 ;
        RECT 3381.2000 2517.4600 3384.2000 2517.9400 ;
        RECT 3381.2000 2512.0200 3384.2000 2512.5000 ;
        RECT 3381.2000 2506.5800 3384.2000 2507.0600 ;
        RECT 3381.2000 2528.3400 3384.2000 2528.8200 ;
        RECT 3381.2000 2522.9000 3384.2000 2523.3800 ;
        RECT 3381.2000 2539.2200 3384.2000 2539.7000 ;
        RECT 3381.2000 2533.7800 3384.2000 2534.2600 ;
        RECT 3381.2000 2555.5400 3384.2000 2556.0200 ;
        RECT 3381.2000 2550.1000 3384.2000 2550.5800 ;
        RECT 3381.2000 2544.6600 3384.2000 2545.1400 ;
        RECT 3381.2000 2566.4200 3384.2000 2566.9000 ;
        RECT 3381.2000 2560.9800 3384.2000 2561.4600 ;
        RECT 3381.2000 2582.7400 3384.2000 2583.2200 ;
        RECT 3381.2000 2577.3000 3384.2000 2577.7800 ;
        RECT 3381.2000 2571.8600 3384.2000 2572.3400 ;
        RECT 3381.2000 2593.6200 3384.2000 2594.1000 ;
        RECT 3381.2000 2588.1800 3384.2000 2588.6600 ;
        RECT 3381.2000 2604.5000 3384.2000 2604.9800 ;
        RECT 3381.2000 2599.0600 3384.2000 2599.5400 ;
        RECT 3381.2000 2620.8200 3384.2000 2621.3000 ;
        RECT 3381.2000 2615.3800 3384.2000 2615.8600 ;
        RECT 3381.2000 2631.7000 3384.2000 2632.1800 ;
        RECT 3381.2000 2626.2600 3384.2000 2626.7400 ;
        RECT 3381.2000 2648.0200 3384.2000 2648.5000 ;
        RECT 3381.2000 2642.5800 3384.2000 2643.0600 ;
        RECT 3381.2000 2637.1400 3384.2000 2637.6200 ;
        RECT 3381.2000 2658.9000 3384.2000 2659.3800 ;
        RECT 3381.2000 2653.4600 3384.2000 2653.9400 ;
        RECT 3381.2000 2675.2200 3384.2000 2675.7000 ;
        RECT 3381.2000 2669.7800 3384.2000 2670.2600 ;
        RECT 3381.2000 2664.3400 3384.2000 2664.8200 ;
        RECT 3381.2000 2686.1000 3384.2000 2686.5800 ;
        RECT 3381.2000 2680.6600 3384.2000 2681.1400 ;
        RECT 3381.2000 2702.4200 3384.2000 2702.9000 ;
        RECT 3381.2000 2696.9800 3384.2000 2697.4600 ;
        RECT 3381.2000 2691.5400 3384.2000 2692.0200 ;
        RECT 3381.2000 2713.3000 3384.2000 2713.7800 ;
        RECT 3381.2000 2707.8600 3384.2000 2708.3400 ;
        RECT 3381.2000 2724.1800 3384.2000 2724.6600 ;
        RECT 3381.2000 2718.7400 3384.2000 2719.2200 ;
        RECT 3381.2000 2740.5000 3384.2000 2740.9800 ;
        RECT 3381.2000 2735.0600 3384.2000 2735.5400 ;
        RECT 3381.2000 2729.6200 3384.2000 2730.1000 ;
        RECT 3381.2000 2751.3800 3384.2000 2751.8600 ;
        RECT 3381.2000 2745.9400 3384.2000 2746.4200 ;
        RECT 3381.2000 2767.7000 3384.2000 2768.1800 ;
        RECT 3381.2000 2762.2600 3384.2000 2762.7400 ;
        RECT 3381.2000 2756.8200 3384.2000 2757.3000 ;
        RECT 3381.2000 2778.5800 3384.2000 2779.0600 ;
        RECT 3381.2000 2773.1400 3384.2000 2773.6200 ;
        RECT 3381.2000 2794.9000 3384.2000 2795.3800 ;
        RECT 3381.2000 2789.4600 3384.2000 2789.9400 ;
        RECT 3381.2000 2784.0200 3384.2000 2784.5000 ;
        RECT 3381.2000 2805.7800 3384.2000 2806.2600 ;
        RECT 3381.2000 2800.3400 3384.2000 2800.8200 ;
        RECT 3381.2000 2816.6600 3384.2000 2817.1400 ;
        RECT 3381.2000 2811.2200 3384.2000 2811.7000 ;
        RECT 3381.2000 2832.9800 3384.2000 2833.4600 ;
        RECT 3381.2000 2827.5400 3384.2000 2828.0200 ;
        RECT 3381.2000 2822.1000 3384.2000 2822.5800 ;
        RECT 3381.2000 2843.8600 3384.2000 2844.3400 ;
        RECT 3381.2000 2838.4200 3384.2000 2838.9000 ;
        RECT 3381.2000 2860.1800 3384.2000 2860.6600 ;
        RECT 3381.2000 2854.7400 3384.2000 2855.2200 ;
        RECT 3381.2000 2849.3000 3384.2000 2849.7800 ;
        RECT 3381.2000 2871.0600 3384.2000 2871.5400 ;
        RECT 3381.2000 2865.6200 3384.2000 2866.1000 ;
        RECT 3381.2000 2876.5000 3384.2000 2876.9800 ;
      LAYER met4 ;
        RECT 3381.2000 6.0000 3384.2000 2883.6600 ;
        RECT 6.0000 6.0000 9.0000 2883.6600 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2808.2800 79.2900 2809.7800 518.0800 ;
        RECT 3305.8000 79.2900 3307.3000 518.0800 ;
      LAYER met3 ;
        RECT 3305.8000 105.2400 3307.3000 105.7200 ;
        RECT 3305.8000 99.8000 3307.3000 100.2800 ;
        RECT 3305.8000 94.3600 3307.3000 94.8400 ;
        RECT 3305.8000 88.9200 3307.3000 89.4000 ;
        RECT 3305.8000 83.4800 3307.3000 83.9600 ;
        RECT 2808.2800 105.2400 2809.7800 105.7200 ;
        RECT 2808.2800 99.8000 2809.7800 100.2800 ;
        RECT 2808.2800 94.3600 2809.7800 94.8400 ;
        RECT 2808.2800 88.9200 2809.7800 89.4000 ;
        RECT 2808.2800 83.4800 2809.7800 83.9600 ;
        RECT 2808.2800 516.5800 3307.3000 518.0800 ;
        RECT 2808.2800 79.2900 3307.3000 80.7900 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2808.2800 538.5700 2809.7800 977.3600 ;
        RECT 3305.8000 538.5700 3307.3000 977.3600 ;
      LAYER met3 ;
        RECT 3305.8000 564.5200 3307.3000 565.0000 ;
        RECT 3305.8000 559.0800 3307.3000 559.5600 ;
        RECT 3305.8000 553.6400 3307.3000 554.1200 ;
        RECT 3305.8000 548.2000 3307.3000 548.6800 ;
        RECT 3305.8000 542.7600 3307.3000 543.2400 ;
        RECT 2808.2800 564.5200 2809.7800 565.0000 ;
        RECT 2808.2800 559.0800 2809.7800 559.5600 ;
        RECT 2808.2800 553.6400 2809.7800 554.1200 ;
        RECT 2808.2800 548.2000 2809.7800 548.6800 ;
        RECT 2808.2800 542.7600 2809.7800 543.2400 ;
        RECT 2808.2800 975.8600 3307.3000 977.3600 ;
        RECT 2808.2800 538.5700 3307.3000 540.0700 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2808.2800 997.8500 2809.7800 1436.6400 ;
        RECT 3305.8000 997.8500 3307.3000 1436.6400 ;
      LAYER met3 ;
        RECT 3305.8000 1023.8000 3307.3000 1024.2800 ;
        RECT 3305.8000 1018.3600 3307.3000 1018.8400 ;
        RECT 3305.8000 1012.9200 3307.3000 1013.4000 ;
        RECT 3305.8000 1007.4800 3307.3000 1007.9600 ;
        RECT 3305.8000 1002.0400 3307.3000 1002.5200 ;
        RECT 2808.2800 1023.8000 2809.7800 1024.2800 ;
        RECT 2808.2800 1018.3600 2809.7800 1018.8400 ;
        RECT 2808.2800 1012.9200 2809.7800 1013.4000 ;
        RECT 2808.2800 1007.4800 2809.7800 1007.9600 ;
        RECT 2808.2800 1002.0400 2809.7800 1002.5200 ;
        RECT 2808.2800 1435.1400 3307.3000 1436.6400 ;
        RECT 2808.2800 997.8500 3307.3000 999.3500 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2808.2800 1457.1300 2809.7800 1895.9200 ;
        RECT 3305.8000 1457.1300 3307.3000 1895.9200 ;
      LAYER met3 ;
        RECT 3305.8000 1483.0800 3307.3000 1483.5600 ;
        RECT 3305.8000 1477.6400 3307.3000 1478.1200 ;
        RECT 3305.8000 1472.2000 3307.3000 1472.6800 ;
        RECT 3305.8000 1466.7600 3307.3000 1467.2400 ;
        RECT 3305.8000 1461.3200 3307.3000 1461.8000 ;
        RECT 2808.2800 1483.0800 2809.7800 1483.5600 ;
        RECT 2808.2800 1477.6400 2809.7800 1478.1200 ;
        RECT 2808.2800 1472.2000 2809.7800 1472.6800 ;
        RECT 2808.2800 1466.7600 2809.7800 1467.2400 ;
        RECT 2808.2800 1461.3200 2809.7800 1461.8000 ;
        RECT 2808.2800 1894.4200 3307.3000 1895.9200 ;
        RECT 2808.2800 1457.1300 3307.3000 1458.6300 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2808.2800 1916.4100 2809.7800 2355.2000 ;
        RECT 3305.8000 1916.4100 3307.3000 2355.2000 ;
      LAYER met3 ;
        RECT 3305.8000 1942.3600 3307.3000 1942.8400 ;
        RECT 3305.8000 1936.9200 3307.3000 1937.4000 ;
        RECT 3305.8000 1931.4800 3307.3000 1931.9600 ;
        RECT 3305.8000 1926.0400 3307.3000 1926.5200 ;
        RECT 3305.8000 1920.6000 3307.3000 1921.0800 ;
        RECT 2808.2800 1942.3600 2809.7800 1942.8400 ;
        RECT 2808.2800 1936.9200 2809.7800 1937.4000 ;
        RECT 2808.2800 1931.4800 2809.7800 1931.9600 ;
        RECT 2808.2800 1926.0400 2809.7800 1926.5200 ;
        RECT 2808.2800 1920.6000 2809.7800 1921.0800 ;
        RECT 2808.2800 2353.7000 3307.3000 2355.2000 ;
        RECT 2808.2800 1916.4100 3307.3000 1917.9100 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'BlockRAM_1KB'
    PORT
      LAYER met4 ;
        RECT 2808.2800 2375.6900 2809.7800 2814.4800 ;
        RECT 3305.8000 2375.6900 3307.3000 2814.4800 ;
      LAYER met3 ;
        RECT 3305.8000 2401.6400 3307.3000 2402.1200 ;
        RECT 3305.8000 2396.2000 3307.3000 2396.6800 ;
        RECT 3305.8000 2390.7600 3307.3000 2391.2400 ;
        RECT 3305.8000 2385.3200 3307.3000 2385.8000 ;
        RECT 3305.8000 2379.8800 3307.3000 2380.3600 ;
        RECT 2808.2800 2401.6400 2809.7800 2402.1200 ;
        RECT 2808.2800 2396.2000 2809.7800 2396.6800 ;
        RECT 2808.2800 2390.7600 2809.7800 2391.2400 ;
        RECT 2808.2800 2385.3200 2809.7800 2385.8000 ;
        RECT 2808.2800 2379.8800 2809.7800 2380.3600 ;
        RECT 2808.2800 2812.9800 3307.3000 2814.4800 ;
        RECT 2808.2800 2375.6900 3307.3000 2377.1900 ;
    END
# end of P/G pin shape extracted from block 'BlockRAM_1KB'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 536.9300 228.4500 748.8300 ;
        RECT 161.7100 536.9300 162.7100 748.8300 ;
      LAYER met3 ;
        RECT 227.4500 727.9800 228.4500 728.4600 ;
        RECT 227.4500 733.4200 228.4500 733.9000 ;
        RECT 227.4500 738.8600 228.4500 739.3400 ;
        RECT 227.4500 717.1000 228.4500 717.5800 ;
        RECT 227.4500 722.5400 228.4500 723.0200 ;
        RECT 227.4500 700.7800 228.4500 701.2600 ;
        RECT 227.4500 706.2200 228.4500 706.7000 ;
        RECT 227.4500 711.6600 228.4500 712.1400 ;
        RECT 227.4500 684.4600 228.4500 684.9400 ;
        RECT 227.4500 689.9000 228.4500 690.3800 ;
        RECT 227.4500 695.3400 228.4500 695.8200 ;
        RECT 227.4500 673.5800 228.4500 674.0600 ;
        RECT 227.4500 679.0200 228.4500 679.5000 ;
        RECT 227.4500 657.2600 228.4500 657.7400 ;
        RECT 227.4500 662.7000 228.4500 663.1800 ;
        RECT 227.4500 668.1400 228.4500 668.6200 ;
        RECT 227.4500 646.3800 228.4500 646.8600 ;
        RECT 227.4500 651.8200 228.4500 652.3000 ;
        RECT 161.7100 727.9800 162.7100 728.4600 ;
        RECT 161.7100 733.4200 162.7100 733.9000 ;
        RECT 161.7100 738.8600 162.7100 739.3400 ;
        RECT 161.7100 717.1000 162.7100 717.5800 ;
        RECT 161.7100 722.5400 162.7100 723.0200 ;
        RECT 161.7100 700.7800 162.7100 701.2600 ;
        RECT 161.7100 706.2200 162.7100 706.7000 ;
        RECT 161.7100 711.6600 162.7100 712.1400 ;
        RECT 161.7100 684.4600 162.7100 684.9400 ;
        RECT 161.7100 689.9000 162.7100 690.3800 ;
        RECT 161.7100 695.3400 162.7100 695.8200 ;
        RECT 161.7100 673.5800 162.7100 674.0600 ;
        RECT 161.7100 679.0200 162.7100 679.5000 ;
        RECT 161.7100 657.2600 162.7100 657.7400 ;
        RECT 161.7100 662.7000 162.7100 663.1800 ;
        RECT 161.7100 668.1400 162.7100 668.6200 ;
        RECT 161.7100 646.3800 162.7100 646.8600 ;
        RECT 161.7100 651.8200 162.7100 652.3000 ;
        RECT 227.4500 630.0600 228.4500 630.5400 ;
        RECT 227.4500 635.5000 228.4500 635.9800 ;
        RECT 227.4500 640.9400 228.4500 641.4200 ;
        RECT 227.4500 619.1800 228.4500 619.6600 ;
        RECT 227.4500 624.6200 228.4500 625.1000 ;
        RECT 227.4500 602.8600 228.4500 603.3400 ;
        RECT 227.4500 608.3000 228.4500 608.7800 ;
        RECT 227.4500 613.7400 228.4500 614.2200 ;
        RECT 227.4500 591.9800 228.4500 592.4600 ;
        RECT 227.4500 597.4200 228.4500 597.9000 ;
        RECT 227.4500 575.6600 228.4500 576.1400 ;
        RECT 227.4500 581.1000 228.4500 581.5800 ;
        RECT 227.4500 586.5400 228.4500 587.0200 ;
        RECT 227.4500 564.7800 228.4500 565.2600 ;
        RECT 227.4500 570.2200 228.4500 570.7000 ;
        RECT 227.4500 548.4600 228.4500 548.9400 ;
        RECT 227.4500 553.9000 228.4500 554.3800 ;
        RECT 227.4500 559.3400 228.4500 559.8200 ;
        RECT 227.4500 543.0200 228.4500 543.5000 ;
        RECT 161.7100 630.0600 162.7100 630.5400 ;
        RECT 161.7100 635.5000 162.7100 635.9800 ;
        RECT 161.7100 640.9400 162.7100 641.4200 ;
        RECT 161.7100 619.1800 162.7100 619.6600 ;
        RECT 161.7100 624.6200 162.7100 625.1000 ;
        RECT 161.7100 602.8600 162.7100 603.3400 ;
        RECT 161.7100 608.3000 162.7100 608.7800 ;
        RECT 161.7100 613.7400 162.7100 614.2200 ;
        RECT 161.7100 591.9800 162.7100 592.4600 ;
        RECT 161.7100 597.4200 162.7100 597.9000 ;
        RECT 161.7100 575.6600 162.7100 576.1400 ;
        RECT 161.7100 581.1000 162.7100 581.5800 ;
        RECT 161.7100 586.5400 162.7100 587.0200 ;
        RECT 161.7100 564.7800 162.7100 565.2600 ;
        RECT 161.7100 570.2200 162.7100 570.7000 ;
        RECT 161.7100 548.4600 162.7100 548.9400 ;
        RECT 161.7100 553.9000 162.7100 554.3800 ;
        RECT 161.7100 559.3400 162.7100 559.8200 ;
        RECT 161.7100 543.0200 162.7100 543.5000 ;
        RECT 161.7100 747.8300 228.4500 748.8300 ;
        RECT 161.7100 536.9300 228.4500 537.9300 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 307.2900 228.4500 519.1900 ;
        RECT 161.7100 307.2900 162.7100 519.1900 ;
      LAYER met3 ;
        RECT 227.4500 498.3400 228.4500 498.8200 ;
        RECT 227.4500 503.7800 228.4500 504.2600 ;
        RECT 227.4500 509.2200 228.4500 509.7000 ;
        RECT 227.4500 487.4600 228.4500 487.9400 ;
        RECT 227.4500 492.9000 228.4500 493.3800 ;
        RECT 227.4500 471.1400 228.4500 471.6200 ;
        RECT 227.4500 476.5800 228.4500 477.0600 ;
        RECT 227.4500 482.0200 228.4500 482.5000 ;
        RECT 227.4500 454.8200 228.4500 455.3000 ;
        RECT 227.4500 460.2600 228.4500 460.7400 ;
        RECT 227.4500 465.7000 228.4500 466.1800 ;
        RECT 227.4500 443.9400 228.4500 444.4200 ;
        RECT 227.4500 449.3800 228.4500 449.8600 ;
        RECT 227.4500 427.6200 228.4500 428.1000 ;
        RECT 227.4500 433.0600 228.4500 433.5400 ;
        RECT 227.4500 438.5000 228.4500 438.9800 ;
        RECT 227.4500 416.7400 228.4500 417.2200 ;
        RECT 227.4500 422.1800 228.4500 422.6600 ;
        RECT 161.7100 498.3400 162.7100 498.8200 ;
        RECT 161.7100 503.7800 162.7100 504.2600 ;
        RECT 161.7100 509.2200 162.7100 509.7000 ;
        RECT 161.7100 487.4600 162.7100 487.9400 ;
        RECT 161.7100 492.9000 162.7100 493.3800 ;
        RECT 161.7100 471.1400 162.7100 471.6200 ;
        RECT 161.7100 476.5800 162.7100 477.0600 ;
        RECT 161.7100 482.0200 162.7100 482.5000 ;
        RECT 161.7100 454.8200 162.7100 455.3000 ;
        RECT 161.7100 460.2600 162.7100 460.7400 ;
        RECT 161.7100 465.7000 162.7100 466.1800 ;
        RECT 161.7100 443.9400 162.7100 444.4200 ;
        RECT 161.7100 449.3800 162.7100 449.8600 ;
        RECT 161.7100 427.6200 162.7100 428.1000 ;
        RECT 161.7100 433.0600 162.7100 433.5400 ;
        RECT 161.7100 438.5000 162.7100 438.9800 ;
        RECT 161.7100 416.7400 162.7100 417.2200 ;
        RECT 161.7100 422.1800 162.7100 422.6600 ;
        RECT 227.4500 400.4200 228.4500 400.9000 ;
        RECT 227.4500 405.8600 228.4500 406.3400 ;
        RECT 227.4500 411.3000 228.4500 411.7800 ;
        RECT 227.4500 389.5400 228.4500 390.0200 ;
        RECT 227.4500 394.9800 228.4500 395.4600 ;
        RECT 227.4500 373.2200 228.4500 373.7000 ;
        RECT 227.4500 378.6600 228.4500 379.1400 ;
        RECT 227.4500 384.1000 228.4500 384.5800 ;
        RECT 227.4500 362.3400 228.4500 362.8200 ;
        RECT 227.4500 367.7800 228.4500 368.2600 ;
        RECT 227.4500 346.0200 228.4500 346.5000 ;
        RECT 227.4500 351.4600 228.4500 351.9400 ;
        RECT 227.4500 356.9000 228.4500 357.3800 ;
        RECT 227.4500 335.1400 228.4500 335.6200 ;
        RECT 227.4500 340.5800 228.4500 341.0600 ;
        RECT 227.4500 318.8200 228.4500 319.3000 ;
        RECT 227.4500 324.2600 228.4500 324.7400 ;
        RECT 227.4500 329.7000 228.4500 330.1800 ;
        RECT 227.4500 313.3800 228.4500 313.8600 ;
        RECT 161.7100 400.4200 162.7100 400.9000 ;
        RECT 161.7100 405.8600 162.7100 406.3400 ;
        RECT 161.7100 411.3000 162.7100 411.7800 ;
        RECT 161.7100 389.5400 162.7100 390.0200 ;
        RECT 161.7100 394.9800 162.7100 395.4600 ;
        RECT 161.7100 373.2200 162.7100 373.7000 ;
        RECT 161.7100 378.6600 162.7100 379.1400 ;
        RECT 161.7100 384.1000 162.7100 384.5800 ;
        RECT 161.7100 362.3400 162.7100 362.8200 ;
        RECT 161.7100 367.7800 162.7100 368.2600 ;
        RECT 161.7100 346.0200 162.7100 346.5000 ;
        RECT 161.7100 351.4600 162.7100 351.9400 ;
        RECT 161.7100 356.9000 162.7100 357.3800 ;
        RECT 161.7100 335.1400 162.7100 335.6200 ;
        RECT 161.7100 340.5800 162.7100 341.0600 ;
        RECT 161.7100 318.8200 162.7100 319.3000 ;
        RECT 161.7100 324.2600 162.7100 324.7400 ;
        RECT 161.7100 329.7000 162.7100 330.1800 ;
        RECT 161.7100 313.3800 162.7100 313.8600 ;
        RECT 161.7100 518.1900 228.4500 519.1900 ;
        RECT 161.7100 307.2900 228.4500 308.2900 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 77.6500 228.4500 289.5500 ;
        RECT 161.7100 77.6500 162.7100 289.5500 ;
      LAYER met3 ;
        RECT 227.4500 268.7000 228.4500 269.1800 ;
        RECT 227.4500 274.1400 228.4500 274.6200 ;
        RECT 227.4500 279.5800 228.4500 280.0600 ;
        RECT 227.4500 257.8200 228.4500 258.3000 ;
        RECT 227.4500 263.2600 228.4500 263.7400 ;
        RECT 227.4500 241.5000 228.4500 241.9800 ;
        RECT 227.4500 246.9400 228.4500 247.4200 ;
        RECT 227.4500 252.3800 228.4500 252.8600 ;
        RECT 227.4500 225.1800 228.4500 225.6600 ;
        RECT 227.4500 230.6200 228.4500 231.1000 ;
        RECT 227.4500 236.0600 228.4500 236.5400 ;
        RECT 227.4500 214.3000 228.4500 214.7800 ;
        RECT 227.4500 219.7400 228.4500 220.2200 ;
        RECT 227.4500 197.9800 228.4500 198.4600 ;
        RECT 227.4500 203.4200 228.4500 203.9000 ;
        RECT 227.4500 208.8600 228.4500 209.3400 ;
        RECT 227.4500 187.1000 228.4500 187.5800 ;
        RECT 227.4500 192.5400 228.4500 193.0200 ;
        RECT 161.7100 268.7000 162.7100 269.1800 ;
        RECT 161.7100 274.1400 162.7100 274.6200 ;
        RECT 161.7100 279.5800 162.7100 280.0600 ;
        RECT 161.7100 257.8200 162.7100 258.3000 ;
        RECT 161.7100 263.2600 162.7100 263.7400 ;
        RECT 161.7100 241.5000 162.7100 241.9800 ;
        RECT 161.7100 246.9400 162.7100 247.4200 ;
        RECT 161.7100 252.3800 162.7100 252.8600 ;
        RECT 161.7100 225.1800 162.7100 225.6600 ;
        RECT 161.7100 230.6200 162.7100 231.1000 ;
        RECT 161.7100 236.0600 162.7100 236.5400 ;
        RECT 161.7100 214.3000 162.7100 214.7800 ;
        RECT 161.7100 219.7400 162.7100 220.2200 ;
        RECT 161.7100 197.9800 162.7100 198.4600 ;
        RECT 161.7100 203.4200 162.7100 203.9000 ;
        RECT 161.7100 208.8600 162.7100 209.3400 ;
        RECT 161.7100 187.1000 162.7100 187.5800 ;
        RECT 161.7100 192.5400 162.7100 193.0200 ;
        RECT 227.4500 170.7800 228.4500 171.2600 ;
        RECT 227.4500 176.2200 228.4500 176.7000 ;
        RECT 227.4500 181.6600 228.4500 182.1400 ;
        RECT 227.4500 159.9000 228.4500 160.3800 ;
        RECT 227.4500 165.3400 228.4500 165.8200 ;
        RECT 227.4500 143.5800 228.4500 144.0600 ;
        RECT 227.4500 149.0200 228.4500 149.5000 ;
        RECT 227.4500 154.4600 228.4500 154.9400 ;
        RECT 227.4500 132.7000 228.4500 133.1800 ;
        RECT 227.4500 138.1400 228.4500 138.6200 ;
        RECT 227.4500 116.3800 228.4500 116.8600 ;
        RECT 227.4500 121.8200 228.4500 122.3000 ;
        RECT 227.4500 127.2600 228.4500 127.7400 ;
        RECT 227.4500 105.5000 228.4500 105.9800 ;
        RECT 227.4500 110.9400 228.4500 111.4200 ;
        RECT 227.4500 89.1800 228.4500 89.6600 ;
        RECT 227.4500 94.6200 228.4500 95.1000 ;
        RECT 227.4500 100.0600 228.4500 100.5400 ;
        RECT 227.4500 83.7400 228.4500 84.2200 ;
        RECT 161.7100 170.7800 162.7100 171.2600 ;
        RECT 161.7100 176.2200 162.7100 176.7000 ;
        RECT 161.7100 181.6600 162.7100 182.1400 ;
        RECT 161.7100 159.9000 162.7100 160.3800 ;
        RECT 161.7100 165.3400 162.7100 165.8200 ;
        RECT 161.7100 143.5800 162.7100 144.0600 ;
        RECT 161.7100 149.0200 162.7100 149.5000 ;
        RECT 161.7100 154.4600 162.7100 154.9400 ;
        RECT 161.7100 132.7000 162.7100 133.1800 ;
        RECT 161.7100 138.1400 162.7100 138.6200 ;
        RECT 161.7100 116.3800 162.7100 116.8600 ;
        RECT 161.7100 121.8200 162.7100 122.3000 ;
        RECT 161.7100 127.2600 162.7100 127.7400 ;
        RECT 161.7100 105.5000 162.7100 105.9800 ;
        RECT 161.7100 110.9400 162.7100 111.4200 ;
        RECT 161.7100 89.1800 162.7100 89.6600 ;
        RECT 161.7100 94.6200 162.7100 95.1000 ;
        RECT 161.7100 100.0600 162.7100 100.5400 ;
        RECT 161.7100 83.7400 162.7100 84.2200 ;
        RECT 161.7100 288.5500 228.4500 289.5500 ;
        RECT 161.7100 77.6500 228.4500 78.6500 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 2603.6900 228.4500 2815.5900 ;
        RECT 161.7100 2603.6900 162.7100 2815.5900 ;
      LAYER met3 ;
        RECT 227.4500 2794.7400 228.4500 2795.2200 ;
        RECT 227.4500 2800.1800 228.4500 2800.6600 ;
        RECT 227.4500 2805.6200 228.4500 2806.1000 ;
        RECT 227.4500 2783.8600 228.4500 2784.3400 ;
        RECT 227.4500 2789.3000 228.4500 2789.7800 ;
        RECT 227.4500 2767.5400 228.4500 2768.0200 ;
        RECT 227.4500 2772.9800 228.4500 2773.4600 ;
        RECT 227.4500 2778.4200 228.4500 2778.9000 ;
        RECT 227.4500 2751.2200 228.4500 2751.7000 ;
        RECT 227.4500 2756.6600 228.4500 2757.1400 ;
        RECT 227.4500 2762.1000 228.4500 2762.5800 ;
        RECT 227.4500 2740.3400 228.4500 2740.8200 ;
        RECT 227.4500 2745.7800 228.4500 2746.2600 ;
        RECT 227.4500 2724.0200 228.4500 2724.5000 ;
        RECT 227.4500 2729.4600 228.4500 2729.9400 ;
        RECT 227.4500 2734.9000 228.4500 2735.3800 ;
        RECT 227.4500 2713.1400 228.4500 2713.6200 ;
        RECT 227.4500 2718.5800 228.4500 2719.0600 ;
        RECT 161.7100 2794.7400 162.7100 2795.2200 ;
        RECT 161.7100 2800.1800 162.7100 2800.6600 ;
        RECT 161.7100 2805.6200 162.7100 2806.1000 ;
        RECT 161.7100 2783.8600 162.7100 2784.3400 ;
        RECT 161.7100 2789.3000 162.7100 2789.7800 ;
        RECT 161.7100 2767.5400 162.7100 2768.0200 ;
        RECT 161.7100 2772.9800 162.7100 2773.4600 ;
        RECT 161.7100 2778.4200 162.7100 2778.9000 ;
        RECT 161.7100 2751.2200 162.7100 2751.7000 ;
        RECT 161.7100 2756.6600 162.7100 2757.1400 ;
        RECT 161.7100 2762.1000 162.7100 2762.5800 ;
        RECT 161.7100 2740.3400 162.7100 2740.8200 ;
        RECT 161.7100 2745.7800 162.7100 2746.2600 ;
        RECT 161.7100 2724.0200 162.7100 2724.5000 ;
        RECT 161.7100 2729.4600 162.7100 2729.9400 ;
        RECT 161.7100 2734.9000 162.7100 2735.3800 ;
        RECT 161.7100 2713.1400 162.7100 2713.6200 ;
        RECT 161.7100 2718.5800 162.7100 2719.0600 ;
        RECT 227.4500 2696.8200 228.4500 2697.3000 ;
        RECT 227.4500 2702.2600 228.4500 2702.7400 ;
        RECT 227.4500 2707.7000 228.4500 2708.1800 ;
        RECT 227.4500 2685.9400 228.4500 2686.4200 ;
        RECT 227.4500 2691.3800 228.4500 2691.8600 ;
        RECT 227.4500 2669.6200 228.4500 2670.1000 ;
        RECT 227.4500 2675.0600 228.4500 2675.5400 ;
        RECT 227.4500 2680.5000 228.4500 2680.9800 ;
        RECT 227.4500 2658.7400 228.4500 2659.2200 ;
        RECT 227.4500 2664.1800 228.4500 2664.6600 ;
        RECT 227.4500 2642.4200 228.4500 2642.9000 ;
        RECT 227.4500 2647.8600 228.4500 2648.3400 ;
        RECT 227.4500 2653.3000 228.4500 2653.7800 ;
        RECT 227.4500 2631.5400 228.4500 2632.0200 ;
        RECT 227.4500 2636.9800 228.4500 2637.4600 ;
        RECT 227.4500 2615.2200 228.4500 2615.7000 ;
        RECT 227.4500 2620.6600 228.4500 2621.1400 ;
        RECT 227.4500 2626.1000 228.4500 2626.5800 ;
        RECT 227.4500 2609.7800 228.4500 2610.2600 ;
        RECT 161.7100 2696.8200 162.7100 2697.3000 ;
        RECT 161.7100 2702.2600 162.7100 2702.7400 ;
        RECT 161.7100 2707.7000 162.7100 2708.1800 ;
        RECT 161.7100 2685.9400 162.7100 2686.4200 ;
        RECT 161.7100 2691.3800 162.7100 2691.8600 ;
        RECT 161.7100 2669.6200 162.7100 2670.1000 ;
        RECT 161.7100 2675.0600 162.7100 2675.5400 ;
        RECT 161.7100 2680.5000 162.7100 2680.9800 ;
        RECT 161.7100 2658.7400 162.7100 2659.2200 ;
        RECT 161.7100 2664.1800 162.7100 2664.6600 ;
        RECT 161.7100 2642.4200 162.7100 2642.9000 ;
        RECT 161.7100 2647.8600 162.7100 2648.3400 ;
        RECT 161.7100 2653.3000 162.7100 2653.7800 ;
        RECT 161.7100 2631.5400 162.7100 2632.0200 ;
        RECT 161.7100 2636.9800 162.7100 2637.4600 ;
        RECT 161.7100 2615.2200 162.7100 2615.7000 ;
        RECT 161.7100 2620.6600 162.7100 2621.1400 ;
        RECT 161.7100 2626.1000 162.7100 2626.5800 ;
        RECT 161.7100 2609.7800 162.7100 2610.2600 ;
        RECT 161.7100 2814.5900 228.4500 2815.5900 ;
        RECT 161.7100 2603.6900 228.4500 2604.6900 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 2374.0500 228.4500 2585.9500 ;
        RECT 161.7100 2374.0500 162.7100 2585.9500 ;
      LAYER met3 ;
        RECT 227.4500 2565.1000 228.4500 2565.5800 ;
        RECT 227.4500 2570.5400 228.4500 2571.0200 ;
        RECT 227.4500 2575.9800 228.4500 2576.4600 ;
        RECT 227.4500 2554.2200 228.4500 2554.7000 ;
        RECT 227.4500 2559.6600 228.4500 2560.1400 ;
        RECT 227.4500 2537.9000 228.4500 2538.3800 ;
        RECT 227.4500 2543.3400 228.4500 2543.8200 ;
        RECT 227.4500 2548.7800 228.4500 2549.2600 ;
        RECT 227.4500 2521.5800 228.4500 2522.0600 ;
        RECT 227.4500 2527.0200 228.4500 2527.5000 ;
        RECT 227.4500 2532.4600 228.4500 2532.9400 ;
        RECT 227.4500 2510.7000 228.4500 2511.1800 ;
        RECT 227.4500 2516.1400 228.4500 2516.6200 ;
        RECT 227.4500 2494.3800 228.4500 2494.8600 ;
        RECT 227.4500 2499.8200 228.4500 2500.3000 ;
        RECT 227.4500 2505.2600 228.4500 2505.7400 ;
        RECT 227.4500 2483.5000 228.4500 2483.9800 ;
        RECT 227.4500 2488.9400 228.4500 2489.4200 ;
        RECT 161.7100 2565.1000 162.7100 2565.5800 ;
        RECT 161.7100 2570.5400 162.7100 2571.0200 ;
        RECT 161.7100 2575.9800 162.7100 2576.4600 ;
        RECT 161.7100 2554.2200 162.7100 2554.7000 ;
        RECT 161.7100 2559.6600 162.7100 2560.1400 ;
        RECT 161.7100 2537.9000 162.7100 2538.3800 ;
        RECT 161.7100 2543.3400 162.7100 2543.8200 ;
        RECT 161.7100 2548.7800 162.7100 2549.2600 ;
        RECT 161.7100 2521.5800 162.7100 2522.0600 ;
        RECT 161.7100 2527.0200 162.7100 2527.5000 ;
        RECT 161.7100 2532.4600 162.7100 2532.9400 ;
        RECT 161.7100 2510.7000 162.7100 2511.1800 ;
        RECT 161.7100 2516.1400 162.7100 2516.6200 ;
        RECT 161.7100 2494.3800 162.7100 2494.8600 ;
        RECT 161.7100 2499.8200 162.7100 2500.3000 ;
        RECT 161.7100 2505.2600 162.7100 2505.7400 ;
        RECT 161.7100 2483.5000 162.7100 2483.9800 ;
        RECT 161.7100 2488.9400 162.7100 2489.4200 ;
        RECT 227.4500 2467.1800 228.4500 2467.6600 ;
        RECT 227.4500 2472.6200 228.4500 2473.1000 ;
        RECT 227.4500 2478.0600 228.4500 2478.5400 ;
        RECT 227.4500 2456.3000 228.4500 2456.7800 ;
        RECT 227.4500 2461.7400 228.4500 2462.2200 ;
        RECT 227.4500 2439.9800 228.4500 2440.4600 ;
        RECT 227.4500 2445.4200 228.4500 2445.9000 ;
        RECT 227.4500 2450.8600 228.4500 2451.3400 ;
        RECT 227.4500 2429.1000 228.4500 2429.5800 ;
        RECT 227.4500 2434.5400 228.4500 2435.0200 ;
        RECT 227.4500 2412.7800 228.4500 2413.2600 ;
        RECT 227.4500 2418.2200 228.4500 2418.7000 ;
        RECT 227.4500 2423.6600 228.4500 2424.1400 ;
        RECT 227.4500 2401.9000 228.4500 2402.3800 ;
        RECT 227.4500 2407.3400 228.4500 2407.8200 ;
        RECT 227.4500 2385.5800 228.4500 2386.0600 ;
        RECT 227.4500 2391.0200 228.4500 2391.5000 ;
        RECT 227.4500 2396.4600 228.4500 2396.9400 ;
        RECT 227.4500 2380.1400 228.4500 2380.6200 ;
        RECT 161.7100 2467.1800 162.7100 2467.6600 ;
        RECT 161.7100 2472.6200 162.7100 2473.1000 ;
        RECT 161.7100 2478.0600 162.7100 2478.5400 ;
        RECT 161.7100 2456.3000 162.7100 2456.7800 ;
        RECT 161.7100 2461.7400 162.7100 2462.2200 ;
        RECT 161.7100 2439.9800 162.7100 2440.4600 ;
        RECT 161.7100 2445.4200 162.7100 2445.9000 ;
        RECT 161.7100 2450.8600 162.7100 2451.3400 ;
        RECT 161.7100 2429.1000 162.7100 2429.5800 ;
        RECT 161.7100 2434.5400 162.7100 2435.0200 ;
        RECT 161.7100 2412.7800 162.7100 2413.2600 ;
        RECT 161.7100 2418.2200 162.7100 2418.7000 ;
        RECT 161.7100 2423.6600 162.7100 2424.1400 ;
        RECT 161.7100 2401.9000 162.7100 2402.3800 ;
        RECT 161.7100 2407.3400 162.7100 2407.8200 ;
        RECT 161.7100 2385.5800 162.7100 2386.0600 ;
        RECT 161.7100 2391.0200 162.7100 2391.5000 ;
        RECT 161.7100 2396.4600 162.7100 2396.9400 ;
        RECT 161.7100 2380.1400 162.7100 2380.6200 ;
        RECT 161.7100 2584.9500 228.4500 2585.9500 ;
        RECT 161.7100 2374.0500 228.4500 2375.0500 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 2144.4100 228.4500 2356.3100 ;
        RECT 161.7100 2144.4100 162.7100 2356.3100 ;
      LAYER met3 ;
        RECT 227.4500 2335.4600 228.4500 2335.9400 ;
        RECT 227.4500 2340.9000 228.4500 2341.3800 ;
        RECT 227.4500 2346.3400 228.4500 2346.8200 ;
        RECT 227.4500 2324.5800 228.4500 2325.0600 ;
        RECT 227.4500 2330.0200 228.4500 2330.5000 ;
        RECT 227.4500 2308.2600 228.4500 2308.7400 ;
        RECT 227.4500 2313.7000 228.4500 2314.1800 ;
        RECT 227.4500 2319.1400 228.4500 2319.6200 ;
        RECT 227.4500 2291.9400 228.4500 2292.4200 ;
        RECT 227.4500 2297.3800 228.4500 2297.8600 ;
        RECT 227.4500 2302.8200 228.4500 2303.3000 ;
        RECT 227.4500 2281.0600 228.4500 2281.5400 ;
        RECT 227.4500 2286.5000 228.4500 2286.9800 ;
        RECT 227.4500 2264.7400 228.4500 2265.2200 ;
        RECT 227.4500 2270.1800 228.4500 2270.6600 ;
        RECT 227.4500 2275.6200 228.4500 2276.1000 ;
        RECT 227.4500 2253.8600 228.4500 2254.3400 ;
        RECT 227.4500 2259.3000 228.4500 2259.7800 ;
        RECT 161.7100 2335.4600 162.7100 2335.9400 ;
        RECT 161.7100 2340.9000 162.7100 2341.3800 ;
        RECT 161.7100 2346.3400 162.7100 2346.8200 ;
        RECT 161.7100 2324.5800 162.7100 2325.0600 ;
        RECT 161.7100 2330.0200 162.7100 2330.5000 ;
        RECT 161.7100 2308.2600 162.7100 2308.7400 ;
        RECT 161.7100 2313.7000 162.7100 2314.1800 ;
        RECT 161.7100 2319.1400 162.7100 2319.6200 ;
        RECT 161.7100 2291.9400 162.7100 2292.4200 ;
        RECT 161.7100 2297.3800 162.7100 2297.8600 ;
        RECT 161.7100 2302.8200 162.7100 2303.3000 ;
        RECT 161.7100 2281.0600 162.7100 2281.5400 ;
        RECT 161.7100 2286.5000 162.7100 2286.9800 ;
        RECT 161.7100 2264.7400 162.7100 2265.2200 ;
        RECT 161.7100 2270.1800 162.7100 2270.6600 ;
        RECT 161.7100 2275.6200 162.7100 2276.1000 ;
        RECT 161.7100 2253.8600 162.7100 2254.3400 ;
        RECT 161.7100 2259.3000 162.7100 2259.7800 ;
        RECT 227.4500 2237.5400 228.4500 2238.0200 ;
        RECT 227.4500 2242.9800 228.4500 2243.4600 ;
        RECT 227.4500 2248.4200 228.4500 2248.9000 ;
        RECT 227.4500 2226.6600 228.4500 2227.1400 ;
        RECT 227.4500 2232.1000 228.4500 2232.5800 ;
        RECT 227.4500 2210.3400 228.4500 2210.8200 ;
        RECT 227.4500 2215.7800 228.4500 2216.2600 ;
        RECT 227.4500 2221.2200 228.4500 2221.7000 ;
        RECT 227.4500 2199.4600 228.4500 2199.9400 ;
        RECT 227.4500 2204.9000 228.4500 2205.3800 ;
        RECT 227.4500 2183.1400 228.4500 2183.6200 ;
        RECT 227.4500 2188.5800 228.4500 2189.0600 ;
        RECT 227.4500 2194.0200 228.4500 2194.5000 ;
        RECT 227.4500 2172.2600 228.4500 2172.7400 ;
        RECT 227.4500 2177.7000 228.4500 2178.1800 ;
        RECT 227.4500 2155.9400 228.4500 2156.4200 ;
        RECT 227.4500 2161.3800 228.4500 2161.8600 ;
        RECT 227.4500 2166.8200 228.4500 2167.3000 ;
        RECT 227.4500 2150.5000 228.4500 2150.9800 ;
        RECT 161.7100 2237.5400 162.7100 2238.0200 ;
        RECT 161.7100 2242.9800 162.7100 2243.4600 ;
        RECT 161.7100 2248.4200 162.7100 2248.9000 ;
        RECT 161.7100 2226.6600 162.7100 2227.1400 ;
        RECT 161.7100 2232.1000 162.7100 2232.5800 ;
        RECT 161.7100 2210.3400 162.7100 2210.8200 ;
        RECT 161.7100 2215.7800 162.7100 2216.2600 ;
        RECT 161.7100 2221.2200 162.7100 2221.7000 ;
        RECT 161.7100 2199.4600 162.7100 2199.9400 ;
        RECT 161.7100 2204.9000 162.7100 2205.3800 ;
        RECT 161.7100 2183.1400 162.7100 2183.6200 ;
        RECT 161.7100 2188.5800 162.7100 2189.0600 ;
        RECT 161.7100 2194.0200 162.7100 2194.5000 ;
        RECT 161.7100 2172.2600 162.7100 2172.7400 ;
        RECT 161.7100 2177.7000 162.7100 2178.1800 ;
        RECT 161.7100 2155.9400 162.7100 2156.4200 ;
        RECT 161.7100 2161.3800 162.7100 2161.8600 ;
        RECT 161.7100 2166.8200 162.7100 2167.3000 ;
        RECT 161.7100 2150.5000 162.7100 2150.9800 ;
        RECT 161.7100 2355.3100 228.4500 2356.3100 ;
        RECT 161.7100 2144.4100 228.4500 2145.4100 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 1914.7700 228.4500 2126.6700 ;
        RECT 161.7100 1914.7700 162.7100 2126.6700 ;
      LAYER met3 ;
        RECT 227.4500 2105.8200 228.4500 2106.3000 ;
        RECT 227.4500 2111.2600 228.4500 2111.7400 ;
        RECT 227.4500 2116.7000 228.4500 2117.1800 ;
        RECT 227.4500 2094.9400 228.4500 2095.4200 ;
        RECT 227.4500 2100.3800 228.4500 2100.8600 ;
        RECT 227.4500 2078.6200 228.4500 2079.1000 ;
        RECT 227.4500 2084.0600 228.4500 2084.5400 ;
        RECT 227.4500 2089.5000 228.4500 2089.9800 ;
        RECT 227.4500 2062.3000 228.4500 2062.7800 ;
        RECT 227.4500 2067.7400 228.4500 2068.2200 ;
        RECT 227.4500 2073.1800 228.4500 2073.6600 ;
        RECT 227.4500 2051.4200 228.4500 2051.9000 ;
        RECT 227.4500 2056.8600 228.4500 2057.3400 ;
        RECT 227.4500 2035.1000 228.4500 2035.5800 ;
        RECT 227.4500 2040.5400 228.4500 2041.0200 ;
        RECT 227.4500 2045.9800 228.4500 2046.4600 ;
        RECT 227.4500 2024.2200 228.4500 2024.7000 ;
        RECT 227.4500 2029.6600 228.4500 2030.1400 ;
        RECT 161.7100 2105.8200 162.7100 2106.3000 ;
        RECT 161.7100 2111.2600 162.7100 2111.7400 ;
        RECT 161.7100 2116.7000 162.7100 2117.1800 ;
        RECT 161.7100 2094.9400 162.7100 2095.4200 ;
        RECT 161.7100 2100.3800 162.7100 2100.8600 ;
        RECT 161.7100 2078.6200 162.7100 2079.1000 ;
        RECT 161.7100 2084.0600 162.7100 2084.5400 ;
        RECT 161.7100 2089.5000 162.7100 2089.9800 ;
        RECT 161.7100 2062.3000 162.7100 2062.7800 ;
        RECT 161.7100 2067.7400 162.7100 2068.2200 ;
        RECT 161.7100 2073.1800 162.7100 2073.6600 ;
        RECT 161.7100 2051.4200 162.7100 2051.9000 ;
        RECT 161.7100 2056.8600 162.7100 2057.3400 ;
        RECT 161.7100 2035.1000 162.7100 2035.5800 ;
        RECT 161.7100 2040.5400 162.7100 2041.0200 ;
        RECT 161.7100 2045.9800 162.7100 2046.4600 ;
        RECT 161.7100 2024.2200 162.7100 2024.7000 ;
        RECT 161.7100 2029.6600 162.7100 2030.1400 ;
        RECT 227.4500 2007.9000 228.4500 2008.3800 ;
        RECT 227.4500 2013.3400 228.4500 2013.8200 ;
        RECT 227.4500 2018.7800 228.4500 2019.2600 ;
        RECT 227.4500 1997.0200 228.4500 1997.5000 ;
        RECT 227.4500 2002.4600 228.4500 2002.9400 ;
        RECT 227.4500 1980.7000 228.4500 1981.1800 ;
        RECT 227.4500 1986.1400 228.4500 1986.6200 ;
        RECT 227.4500 1991.5800 228.4500 1992.0600 ;
        RECT 227.4500 1969.8200 228.4500 1970.3000 ;
        RECT 227.4500 1975.2600 228.4500 1975.7400 ;
        RECT 227.4500 1953.5000 228.4500 1953.9800 ;
        RECT 227.4500 1958.9400 228.4500 1959.4200 ;
        RECT 227.4500 1964.3800 228.4500 1964.8600 ;
        RECT 227.4500 1942.6200 228.4500 1943.1000 ;
        RECT 227.4500 1948.0600 228.4500 1948.5400 ;
        RECT 227.4500 1926.3000 228.4500 1926.7800 ;
        RECT 227.4500 1931.7400 228.4500 1932.2200 ;
        RECT 227.4500 1937.1800 228.4500 1937.6600 ;
        RECT 227.4500 1920.8600 228.4500 1921.3400 ;
        RECT 161.7100 2007.9000 162.7100 2008.3800 ;
        RECT 161.7100 2013.3400 162.7100 2013.8200 ;
        RECT 161.7100 2018.7800 162.7100 2019.2600 ;
        RECT 161.7100 1997.0200 162.7100 1997.5000 ;
        RECT 161.7100 2002.4600 162.7100 2002.9400 ;
        RECT 161.7100 1980.7000 162.7100 1981.1800 ;
        RECT 161.7100 1986.1400 162.7100 1986.6200 ;
        RECT 161.7100 1991.5800 162.7100 1992.0600 ;
        RECT 161.7100 1969.8200 162.7100 1970.3000 ;
        RECT 161.7100 1975.2600 162.7100 1975.7400 ;
        RECT 161.7100 1953.5000 162.7100 1953.9800 ;
        RECT 161.7100 1958.9400 162.7100 1959.4200 ;
        RECT 161.7100 1964.3800 162.7100 1964.8600 ;
        RECT 161.7100 1942.6200 162.7100 1943.1000 ;
        RECT 161.7100 1948.0600 162.7100 1948.5400 ;
        RECT 161.7100 1926.3000 162.7100 1926.7800 ;
        RECT 161.7100 1931.7400 162.7100 1932.2200 ;
        RECT 161.7100 1937.1800 162.7100 1937.6600 ;
        RECT 161.7100 1920.8600 162.7100 1921.3400 ;
        RECT 161.7100 2125.6700 228.4500 2126.6700 ;
        RECT 161.7100 1914.7700 228.4500 1915.7700 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 1685.1300 228.4500 1897.0300 ;
        RECT 161.7100 1685.1300 162.7100 1897.0300 ;
      LAYER met3 ;
        RECT 227.4500 1876.1800 228.4500 1876.6600 ;
        RECT 227.4500 1881.6200 228.4500 1882.1000 ;
        RECT 227.4500 1887.0600 228.4500 1887.5400 ;
        RECT 227.4500 1865.3000 228.4500 1865.7800 ;
        RECT 227.4500 1870.7400 228.4500 1871.2200 ;
        RECT 227.4500 1848.9800 228.4500 1849.4600 ;
        RECT 227.4500 1854.4200 228.4500 1854.9000 ;
        RECT 227.4500 1859.8600 228.4500 1860.3400 ;
        RECT 227.4500 1832.6600 228.4500 1833.1400 ;
        RECT 227.4500 1838.1000 228.4500 1838.5800 ;
        RECT 227.4500 1843.5400 228.4500 1844.0200 ;
        RECT 227.4500 1821.7800 228.4500 1822.2600 ;
        RECT 227.4500 1827.2200 228.4500 1827.7000 ;
        RECT 227.4500 1805.4600 228.4500 1805.9400 ;
        RECT 227.4500 1810.9000 228.4500 1811.3800 ;
        RECT 227.4500 1816.3400 228.4500 1816.8200 ;
        RECT 227.4500 1794.5800 228.4500 1795.0600 ;
        RECT 227.4500 1800.0200 228.4500 1800.5000 ;
        RECT 161.7100 1876.1800 162.7100 1876.6600 ;
        RECT 161.7100 1881.6200 162.7100 1882.1000 ;
        RECT 161.7100 1887.0600 162.7100 1887.5400 ;
        RECT 161.7100 1865.3000 162.7100 1865.7800 ;
        RECT 161.7100 1870.7400 162.7100 1871.2200 ;
        RECT 161.7100 1848.9800 162.7100 1849.4600 ;
        RECT 161.7100 1854.4200 162.7100 1854.9000 ;
        RECT 161.7100 1859.8600 162.7100 1860.3400 ;
        RECT 161.7100 1832.6600 162.7100 1833.1400 ;
        RECT 161.7100 1838.1000 162.7100 1838.5800 ;
        RECT 161.7100 1843.5400 162.7100 1844.0200 ;
        RECT 161.7100 1821.7800 162.7100 1822.2600 ;
        RECT 161.7100 1827.2200 162.7100 1827.7000 ;
        RECT 161.7100 1805.4600 162.7100 1805.9400 ;
        RECT 161.7100 1810.9000 162.7100 1811.3800 ;
        RECT 161.7100 1816.3400 162.7100 1816.8200 ;
        RECT 161.7100 1794.5800 162.7100 1795.0600 ;
        RECT 161.7100 1800.0200 162.7100 1800.5000 ;
        RECT 227.4500 1778.2600 228.4500 1778.7400 ;
        RECT 227.4500 1783.7000 228.4500 1784.1800 ;
        RECT 227.4500 1789.1400 228.4500 1789.6200 ;
        RECT 227.4500 1767.3800 228.4500 1767.8600 ;
        RECT 227.4500 1772.8200 228.4500 1773.3000 ;
        RECT 227.4500 1751.0600 228.4500 1751.5400 ;
        RECT 227.4500 1756.5000 228.4500 1756.9800 ;
        RECT 227.4500 1761.9400 228.4500 1762.4200 ;
        RECT 227.4500 1740.1800 228.4500 1740.6600 ;
        RECT 227.4500 1745.6200 228.4500 1746.1000 ;
        RECT 227.4500 1723.8600 228.4500 1724.3400 ;
        RECT 227.4500 1729.3000 228.4500 1729.7800 ;
        RECT 227.4500 1734.7400 228.4500 1735.2200 ;
        RECT 227.4500 1712.9800 228.4500 1713.4600 ;
        RECT 227.4500 1718.4200 228.4500 1718.9000 ;
        RECT 227.4500 1696.6600 228.4500 1697.1400 ;
        RECT 227.4500 1702.1000 228.4500 1702.5800 ;
        RECT 227.4500 1707.5400 228.4500 1708.0200 ;
        RECT 227.4500 1691.2200 228.4500 1691.7000 ;
        RECT 161.7100 1778.2600 162.7100 1778.7400 ;
        RECT 161.7100 1783.7000 162.7100 1784.1800 ;
        RECT 161.7100 1789.1400 162.7100 1789.6200 ;
        RECT 161.7100 1767.3800 162.7100 1767.8600 ;
        RECT 161.7100 1772.8200 162.7100 1773.3000 ;
        RECT 161.7100 1751.0600 162.7100 1751.5400 ;
        RECT 161.7100 1756.5000 162.7100 1756.9800 ;
        RECT 161.7100 1761.9400 162.7100 1762.4200 ;
        RECT 161.7100 1740.1800 162.7100 1740.6600 ;
        RECT 161.7100 1745.6200 162.7100 1746.1000 ;
        RECT 161.7100 1723.8600 162.7100 1724.3400 ;
        RECT 161.7100 1729.3000 162.7100 1729.7800 ;
        RECT 161.7100 1734.7400 162.7100 1735.2200 ;
        RECT 161.7100 1712.9800 162.7100 1713.4600 ;
        RECT 161.7100 1718.4200 162.7100 1718.9000 ;
        RECT 161.7100 1696.6600 162.7100 1697.1400 ;
        RECT 161.7100 1702.1000 162.7100 1702.5800 ;
        RECT 161.7100 1707.5400 162.7100 1708.0200 ;
        RECT 161.7100 1691.2200 162.7100 1691.7000 ;
        RECT 161.7100 1896.0300 228.4500 1897.0300 ;
        RECT 161.7100 1685.1300 228.4500 1686.1300 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 1455.4900 228.4500 1667.3900 ;
        RECT 161.7100 1455.4900 162.7100 1667.3900 ;
      LAYER met3 ;
        RECT 227.4500 1646.5400 228.4500 1647.0200 ;
        RECT 227.4500 1651.9800 228.4500 1652.4600 ;
        RECT 227.4500 1657.4200 228.4500 1657.9000 ;
        RECT 227.4500 1635.6600 228.4500 1636.1400 ;
        RECT 227.4500 1641.1000 228.4500 1641.5800 ;
        RECT 227.4500 1619.3400 228.4500 1619.8200 ;
        RECT 227.4500 1624.7800 228.4500 1625.2600 ;
        RECT 227.4500 1630.2200 228.4500 1630.7000 ;
        RECT 227.4500 1603.0200 228.4500 1603.5000 ;
        RECT 227.4500 1608.4600 228.4500 1608.9400 ;
        RECT 227.4500 1613.9000 228.4500 1614.3800 ;
        RECT 227.4500 1592.1400 228.4500 1592.6200 ;
        RECT 227.4500 1597.5800 228.4500 1598.0600 ;
        RECT 227.4500 1575.8200 228.4500 1576.3000 ;
        RECT 227.4500 1581.2600 228.4500 1581.7400 ;
        RECT 227.4500 1586.7000 228.4500 1587.1800 ;
        RECT 227.4500 1564.9400 228.4500 1565.4200 ;
        RECT 227.4500 1570.3800 228.4500 1570.8600 ;
        RECT 161.7100 1646.5400 162.7100 1647.0200 ;
        RECT 161.7100 1651.9800 162.7100 1652.4600 ;
        RECT 161.7100 1657.4200 162.7100 1657.9000 ;
        RECT 161.7100 1635.6600 162.7100 1636.1400 ;
        RECT 161.7100 1641.1000 162.7100 1641.5800 ;
        RECT 161.7100 1619.3400 162.7100 1619.8200 ;
        RECT 161.7100 1624.7800 162.7100 1625.2600 ;
        RECT 161.7100 1630.2200 162.7100 1630.7000 ;
        RECT 161.7100 1603.0200 162.7100 1603.5000 ;
        RECT 161.7100 1608.4600 162.7100 1608.9400 ;
        RECT 161.7100 1613.9000 162.7100 1614.3800 ;
        RECT 161.7100 1592.1400 162.7100 1592.6200 ;
        RECT 161.7100 1597.5800 162.7100 1598.0600 ;
        RECT 161.7100 1575.8200 162.7100 1576.3000 ;
        RECT 161.7100 1581.2600 162.7100 1581.7400 ;
        RECT 161.7100 1586.7000 162.7100 1587.1800 ;
        RECT 161.7100 1564.9400 162.7100 1565.4200 ;
        RECT 161.7100 1570.3800 162.7100 1570.8600 ;
        RECT 227.4500 1548.6200 228.4500 1549.1000 ;
        RECT 227.4500 1554.0600 228.4500 1554.5400 ;
        RECT 227.4500 1559.5000 228.4500 1559.9800 ;
        RECT 227.4500 1537.7400 228.4500 1538.2200 ;
        RECT 227.4500 1543.1800 228.4500 1543.6600 ;
        RECT 227.4500 1521.4200 228.4500 1521.9000 ;
        RECT 227.4500 1526.8600 228.4500 1527.3400 ;
        RECT 227.4500 1532.3000 228.4500 1532.7800 ;
        RECT 227.4500 1510.5400 228.4500 1511.0200 ;
        RECT 227.4500 1515.9800 228.4500 1516.4600 ;
        RECT 227.4500 1494.2200 228.4500 1494.7000 ;
        RECT 227.4500 1499.6600 228.4500 1500.1400 ;
        RECT 227.4500 1505.1000 228.4500 1505.5800 ;
        RECT 227.4500 1483.3400 228.4500 1483.8200 ;
        RECT 227.4500 1488.7800 228.4500 1489.2600 ;
        RECT 227.4500 1467.0200 228.4500 1467.5000 ;
        RECT 227.4500 1472.4600 228.4500 1472.9400 ;
        RECT 227.4500 1477.9000 228.4500 1478.3800 ;
        RECT 227.4500 1461.5800 228.4500 1462.0600 ;
        RECT 161.7100 1548.6200 162.7100 1549.1000 ;
        RECT 161.7100 1554.0600 162.7100 1554.5400 ;
        RECT 161.7100 1559.5000 162.7100 1559.9800 ;
        RECT 161.7100 1537.7400 162.7100 1538.2200 ;
        RECT 161.7100 1543.1800 162.7100 1543.6600 ;
        RECT 161.7100 1521.4200 162.7100 1521.9000 ;
        RECT 161.7100 1526.8600 162.7100 1527.3400 ;
        RECT 161.7100 1532.3000 162.7100 1532.7800 ;
        RECT 161.7100 1510.5400 162.7100 1511.0200 ;
        RECT 161.7100 1515.9800 162.7100 1516.4600 ;
        RECT 161.7100 1494.2200 162.7100 1494.7000 ;
        RECT 161.7100 1499.6600 162.7100 1500.1400 ;
        RECT 161.7100 1505.1000 162.7100 1505.5800 ;
        RECT 161.7100 1483.3400 162.7100 1483.8200 ;
        RECT 161.7100 1488.7800 162.7100 1489.2600 ;
        RECT 161.7100 1467.0200 162.7100 1467.5000 ;
        RECT 161.7100 1472.4600 162.7100 1472.9400 ;
        RECT 161.7100 1477.9000 162.7100 1478.3800 ;
        RECT 161.7100 1461.5800 162.7100 1462.0600 ;
        RECT 161.7100 1666.3900 228.4500 1667.3900 ;
        RECT 161.7100 1455.4900 228.4500 1456.4900 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 1225.8500 228.4500 1437.7500 ;
        RECT 161.7100 1225.8500 162.7100 1437.7500 ;
      LAYER met3 ;
        RECT 227.4500 1416.9000 228.4500 1417.3800 ;
        RECT 227.4500 1422.3400 228.4500 1422.8200 ;
        RECT 227.4500 1427.7800 228.4500 1428.2600 ;
        RECT 227.4500 1406.0200 228.4500 1406.5000 ;
        RECT 227.4500 1411.4600 228.4500 1411.9400 ;
        RECT 227.4500 1389.7000 228.4500 1390.1800 ;
        RECT 227.4500 1395.1400 228.4500 1395.6200 ;
        RECT 227.4500 1400.5800 228.4500 1401.0600 ;
        RECT 227.4500 1373.3800 228.4500 1373.8600 ;
        RECT 227.4500 1378.8200 228.4500 1379.3000 ;
        RECT 227.4500 1384.2600 228.4500 1384.7400 ;
        RECT 227.4500 1362.5000 228.4500 1362.9800 ;
        RECT 227.4500 1367.9400 228.4500 1368.4200 ;
        RECT 227.4500 1346.1800 228.4500 1346.6600 ;
        RECT 227.4500 1351.6200 228.4500 1352.1000 ;
        RECT 227.4500 1357.0600 228.4500 1357.5400 ;
        RECT 227.4500 1335.3000 228.4500 1335.7800 ;
        RECT 227.4500 1340.7400 228.4500 1341.2200 ;
        RECT 161.7100 1416.9000 162.7100 1417.3800 ;
        RECT 161.7100 1422.3400 162.7100 1422.8200 ;
        RECT 161.7100 1427.7800 162.7100 1428.2600 ;
        RECT 161.7100 1406.0200 162.7100 1406.5000 ;
        RECT 161.7100 1411.4600 162.7100 1411.9400 ;
        RECT 161.7100 1389.7000 162.7100 1390.1800 ;
        RECT 161.7100 1395.1400 162.7100 1395.6200 ;
        RECT 161.7100 1400.5800 162.7100 1401.0600 ;
        RECT 161.7100 1373.3800 162.7100 1373.8600 ;
        RECT 161.7100 1378.8200 162.7100 1379.3000 ;
        RECT 161.7100 1384.2600 162.7100 1384.7400 ;
        RECT 161.7100 1362.5000 162.7100 1362.9800 ;
        RECT 161.7100 1367.9400 162.7100 1368.4200 ;
        RECT 161.7100 1346.1800 162.7100 1346.6600 ;
        RECT 161.7100 1351.6200 162.7100 1352.1000 ;
        RECT 161.7100 1357.0600 162.7100 1357.5400 ;
        RECT 161.7100 1335.3000 162.7100 1335.7800 ;
        RECT 161.7100 1340.7400 162.7100 1341.2200 ;
        RECT 227.4500 1318.9800 228.4500 1319.4600 ;
        RECT 227.4500 1324.4200 228.4500 1324.9000 ;
        RECT 227.4500 1329.8600 228.4500 1330.3400 ;
        RECT 227.4500 1308.1000 228.4500 1308.5800 ;
        RECT 227.4500 1313.5400 228.4500 1314.0200 ;
        RECT 227.4500 1291.7800 228.4500 1292.2600 ;
        RECT 227.4500 1297.2200 228.4500 1297.7000 ;
        RECT 227.4500 1302.6600 228.4500 1303.1400 ;
        RECT 227.4500 1280.9000 228.4500 1281.3800 ;
        RECT 227.4500 1286.3400 228.4500 1286.8200 ;
        RECT 227.4500 1264.5800 228.4500 1265.0600 ;
        RECT 227.4500 1270.0200 228.4500 1270.5000 ;
        RECT 227.4500 1275.4600 228.4500 1275.9400 ;
        RECT 227.4500 1253.7000 228.4500 1254.1800 ;
        RECT 227.4500 1259.1400 228.4500 1259.6200 ;
        RECT 227.4500 1237.3800 228.4500 1237.8600 ;
        RECT 227.4500 1242.8200 228.4500 1243.3000 ;
        RECT 227.4500 1248.2600 228.4500 1248.7400 ;
        RECT 227.4500 1231.9400 228.4500 1232.4200 ;
        RECT 161.7100 1318.9800 162.7100 1319.4600 ;
        RECT 161.7100 1324.4200 162.7100 1324.9000 ;
        RECT 161.7100 1329.8600 162.7100 1330.3400 ;
        RECT 161.7100 1308.1000 162.7100 1308.5800 ;
        RECT 161.7100 1313.5400 162.7100 1314.0200 ;
        RECT 161.7100 1291.7800 162.7100 1292.2600 ;
        RECT 161.7100 1297.2200 162.7100 1297.7000 ;
        RECT 161.7100 1302.6600 162.7100 1303.1400 ;
        RECT 161.7100 1280.9000 162.7100 1281.3800 ;
        RECT 161.7100 1286.3400 162.7100 1286.8200 ;
        RECT 161.7100 1264.5800 162.7100 1265.0600 ;
        RECT 161.7100 1270.0200 162.7100 1270.5000 ;
        RECT 161.7100 1275.4600 162.7100 1275.9400 ;
        RECT 161.7100 1253.7000 162.7100 1254.1800 ;
        RECT 161.7100 1259.1400 162.7100 1259.6200 ;
        RECT 161.7100 1237.3800 162.7100 1237.8600 ;
        RECT 161.7100 1242.8200 162.7100 1243.3000 ;
        RECT 161.7100 1248.2600 162.7100 1248.7400 ;
        RECT 161.7100 1231.9400 162.7100 1232.4200 ;
        RECT 161.7100 1436.7500 228.4500 1437.7500 ;
        RECT 161.7100 1225.8500 228.4500 1226.8500 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 996.2100 228.4500 1208.1100 ;
        RECT 161.7100 996.2100 162.7100 1208.1100 ;
      LAYER met3 ;
        RECT 227.4500 1187.2600 228.4500 1187.7400 ;
        RECT 227.4500 1192.7000 228.4500 1193.1800 ;
        RECT 227.4500 1198.1400 228.4500 1198.6200 ;
        RECT 227.4500 1176.3800 228.4500 1176.8600 ;
        RECT 227.4500 1181.8200 228.4500 1182.3000 ;
        RECT 227.4500 1160.0600 228.4500 1160.5400 ;
        RECT 227.4500 1165.5000 228.4500 1165.9800 ;
        RECT 227.4500 1170.9400 228.4500 1171.4200 ;
        RECT 227.4500 1143.7400 228.4500 1144.2200 ;
        RECT 227.4500 1149.1800 228.4500 1149.6600 ;
        RECT 227.4500 1154.6200 228.4500 1155.1000 ;
        RECT 227.4500 1132.8600 228.4500 1133.3400 ;
        RECT 227.4500 1138.3000 228.4500 1138.7800 ;
        RECT 227.4500 1116.5400 228.4500 1117.0200 ;
        RECT 227.4500 1121.9800 228.4500 1122.4600 ;
        RECT 227.4500 1127.4200 228.4500 1127.9000 ;
        RECT 227.4500 1105.6600 228.4500 1106.1400 ;
        RECT 227.4500 1111.1000 228.4500 1111.5800 ;
        RECT 161.7100 1187.2600 162.7100 1187.7400 ;
        RECT 161.7100 1192.7000 162.7100 1193.1800 ;
        RECT 161.7100 1198.1400 162.7100 1198.6200 ;
        RECT 161.7100 1176.3800 162.7100 1176.8600 ;
        RECT 161.7100 1181.8200 162.7100 1182.3000 ;
        RECT 161.7100 1160.0600 162.7100 1160.5400 ;
        RECT 161.7100 1165.5000 162.7100 1165.9800 ;
        RECT 161.7100 1170.9400 162.7100 1171.4200 ;
        RECT 161.7100 1143.7400 162.7100 1144.2200 ;
        RECT 161.7100 1149.1800 162.7100 1149.6600 ;
        RECT 161.7100 1154.6200 162.7100 1155.1000 ;
        RECT 161.7100 1132.8600 162.7100 1133.3400 ;
        RECT 161.7100 1138.3000 162.7100 1138.7800 ;
        RECT 161.7100 1116.5400 162.7100 1117.0200 ;
        RECT 161.7100 1121.9800 162.7100 1122.4600 ;
        RECT 161.7100 1127.4200 162.7100 1127.9000 ;
        RECT 161.7100 1105.6600 162.7100 1106.1400 ;
        RECT 161.7100 1111.1000 162.7100 1111.5800 ;
        RECT 227.4500 1089.3400 228.4500 1089.8200 ;
        RECT 227.4500 1094.7800 228.4500 1095.2600 ;
        RECT 227.4500 1100.2200 228.4500 1100.7000 ;
        RECT 227.4500 1078.4600 228.4500 1078.9400 ;
        RECT 227.4500 1083.9000 228.4500 1084.3800 ;
        RECT 227.4500 1062.1400 228.4500 1062.6200 ;
        RECT 227.4500 1067.5800 228.4500 1068.0600 ;
        RECT 227.4500 1073.0200 228.4500 1073.5000 ;
        RECT 227.4500 1051.2600 228.4500 1051.7400 ;
        RECT 227.4500 1056.7000 228.4500 1057.1800 ;
        RECT 227.4500 1034.9400 228.4500 1035.4200 ;
        RECT 227.4500 1040.3800 228.4500 1040.8600 ;
        RECT 227.4500 1045.8200 228.4500 1046.3000 ;
        RECT 227.4500 1024.0600 228.4500 1024.5400 ;
        RECT 227.4500 1029.5000 228.4500 1029.9800 ;
        RECT 227.4500 1007.7400 228.4500 1008.2200 ;
        RECT 227.4500 1013.1800 228.4500 1013.6600 ;
        RECT 227.4500 1018.6200 228.4500 1019.1000 ;
        RECT 227.4500 1002.3000 228.4500 1002.7800 ;
        RECT 161.7100 1089.3400 162.7100 1089.8200 ;
        RECT 161.7100 1094.7800 162.7100 1095.2600 ;
        RECT 161.7100 1100.2200 162.7100 1100.7000 ;
        RECT 161.7100 1078.4600 162.7100 1078.9400 ;
        RECT 161.7100 1083.9000 162.7100 1084.3800 ;
        RECT 161.7100 1062.1400 162.7100 1062.6200 ;
        RECT 161.7100 1067.5800 162.7100 1068.0600 ;
        RECT 161.7100 1073.0200 162.7100 1073.5000 ;
        RECT 161.7100 1051.2600 162.7100 1051.7400 ;
        RECT 161.7100 1056.7000 162.7100 1057.1800 ;
        RECT 161.7100 1034.9400 162.7100 1035.4200 ;
        RECT 161.7100 1040.3800 162.7100 1040.8600 ;
        RECT 161.7100 1045.8200 162.7100 1046.3000 ;
        RECT 161.7100 1024.0600 162.7100 1024.5400 ;
        RECT 161.7100 1029.5000 162.7100 1029.9800 ;
        RECT 161.7100 1007.7400 162.7100 1008.2200 ;
        RECT 161.7100 1013.1800 162.7100 1013.6600 ;
        RECT 161.7100 1018.6200 162.7100 1019.1000 ;
        RECT 161.7100 1002.3000 162.7100 1002.7800 ;
        RECT 161.7100 1207.1100 228.4500 1208.1100 ;
        RECT 161.7100 996.2100 228.4500 997.2100 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'W_IO'
    PORT
      LAYER met4 ;
        RECT 227.4500 766.5700 228.4500 978.4700 ;
        RECT 161.7100 766.5700 162.7100 978.4700 ;
      LAYER met3 ;
        RECT 227.4500 957.6200 228.4500 958.1000 ;
        RECT 227.4500 963.0600 228.4500 963.5400 ;
        RECT 227.4500 968.5000 228.4500 968.9800 ;
        RECT 227.4500 946.7400 228.4500 947.2200 ;
        RECT 227.4500 952.1800 228.4500 952.6600 ;
        RECT 227.4500 930.4200 228.4500 930.9000 ;
        RECT 227.4500 935.8600 228.4500 936.3400 ;
        RECT 227.4500 941.3000 228.4500 941.7800 ;
        RECT 227.4500 914.1000 228.4500 914.5800 ;
        RECT 227.4500 919.5400 228.4500 920.0200 ;
        RECT 227.4500 924.9800 228.4500 925.4600 ;
        RECT 227.4500 903.2200 228.4500 903.7000 ;
        RECT 227.4500 908.6600 228.4500 909.1400 ;
        RECT 227.4500 886.9000 228.4500 887.3800 ;
        RECT 227.4500 892.3400 228.4500 892.8200 ;
        RECT 227.4500 897.7800 228.4500 898.2600 ;
        RECT 227.4500 876.0200 228.4500 876.5000 ;
        RECT 227.4500 881.4600 228.4500 881.9400 ;
        RECT 161.7100 957.6200 162.7100 958.1000 ;
        RECT 161.7100 963.0600 162.7100 963.5400 ;
        RECT 161.7100 968.5000 162.7100 968.9800 ;
        RECT 161.7100 946.7400 162.7100 947.2200 ;
        RECT 161.7100 952.1800 162.7100 952.6600 ;
        RECT 161.7100 930.4200 162.7100 930.9000 ;
        RECT 161.7100 935.8600 162.7100 936.3400 ;
        RECT 161.7100 941.3000 162.7100 941.7800 ;
        RECT 161.7100 914.1000 162.7100 914.5800 ;
        RECT 161.7100 919.5400 162.7100 920.0200 ;
        RECT 161.7100 924.9800 162.7100 925.4600 ;
        RECT 161.7100 903.2200 162.7100 903.7000 ;
        RECT 161.7100 908.6600 162.7100 909.1400 ;
        RECT 161.7100 886.9000 162.7100 887.3800 ;
        RECT 161.7100 892.3400 162.7100 892.8200 ;
        RECT 161.7100 897.7800 162.7100 898.2600 ;
        RECT 161.7100 876.0200 162.7100 876.5000 ;
        RECT 161.7100 881.4600 162.7100 881.9400 ;
        RECT 227.4500 859.7000 228.4500 860.1800 ;
        RECT 227.4500 865.1400 228.4500 865.6200 ;
        RECT 227.4500 870.5800 228.4500 871.0600 ;
        RECT 227.4500 848.8200 228.4500 849.3000 ;
        RECT 227.4500 854.2600 228.4500 854.7400 ;
        RECT 227.4500 832.5000 228.4500 832.9800 ;
        RECT 227.4500 837.9400 228.4500 838.4200 ;
        RECT 227.4500 843.3800 228.4500 843.8600 ;
        RECT 227.4500 821.6200 228.4500 822.1000 ;
        RECT 227.4500 827.0600 228.4500 827.5400 ;
        RECT 227.4500 805.3000 228.4500 805.7800 ;
        RECT 227.4500 810.7400 228.4500 811.2200 ;
        RECT 227.4500 816.1800 228.4500 816.6600 ;
        RECT 227.4500 794.4200 228.4500 794.9000 ;
        RECT 227.4500 799.8600 228.4500 800.3400 ;
        RECT 227.4500 778.1000 228.4500 778.5800 ;
        RECT 227.4500 783.5400 228.4500 784.0200 ;
        RECT 227.4500 788.9800 228.4500 789.4600 ;
        RECT 227.4500 772.6600 228.4500 773.1400 ;
        RECT 161.7100 859.7000 162.7100 860.1800 ;
        RECT 161.7100 865.1400 162.7100 865.6200 ;
        RECT 161.7100 870.5800 162.7100 871.0600 ;
        RECT 161.7100 848.8200 162.7100 849.3000 ;
        RECT 161.7100 854.2600 162.7100 854.7400 ;
        RECT 161.7100 832.5000 162.7100 832.9800 ;
        RECT 161.7100 837.9400 162.7100 838.4200 ;
        RECT 161.7100 843.3800 162.7100 843.8600 ;
        RECT 161.7100 821.6200 162.7100 822.1000 ;
        RECT 161.7100 827.0600 162.7100 827.5400 ;
        RECT 161.7100 805.3000 162.7100 805.7800 ;
        RECT 161.7100 810.7400 162.7100 811.2200 ;
        RECT 161.7100 816.1800 162.7100 816.6600 ;
        RECT 161.7100 794.4200 162.7100 794.9000 ;
        RECT 161.7100 799.8600 162.7100 800.3400 ;
        RECT 161.7100 778.1000 162.7100 778.5800 ;
        RECT 161.7100 783.5400 162.7100 784.0200 ;
        RECT 161.7100 788.9800 162.7100 789.4600 ;
        RECT 161.7100 772.6600 162.7100 773.1400 ;
        RECT 161.7100 977.4700 228.4500 978.4700 ;
        RECT 161.7100 766.5700 228.4500 767.5700 ;
    END
# end of P/G pin shape extracted from block 'W_IO'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 2254.5600 2830.6100 2256.5600 2857.5400 ;
        RECT 2457.6600 2830.6100 2459.6600 2857.5400 ;
      LAYER met3 ;
        RECT 2457.6600 2847.3200 2459.6600 2847.8000 ;
        RECT 2254.5600 2847.3200 2256.5600 2847.8000 ;
        RECT 2457.6600 2841.8800 2459.6600 2842.3600 ;
        RECT 2457.6600 2836.4400 2459.6600 2836.9200 ;
        RECT 2254.5600 2841.8800 2256.5600 2842.3600 ;
        RECT 2254.5600 2836.4400 2256.5600 2836.9200 ;
        RECT 2254.5600 2855.5400 2459.6600 2857.5400 ;
        RECT 2254.5600 2830.6100 2459.6600 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 534.5700 2446.9200 750.6700 ;
        RECT 2400.3200 534.5700 2401.9200 750.6700 ;
        RECT 2355.3200 534.5700 2356.9200 750.6700 ;
        RECT 2310.3200 534.5700 2311.9200 750.6700 ;
        RECT 2265.3200 534.5700 2266.9200 750.6700 ;
        RECT 2457.6600 534.5700 2460.6600 750.6700 ;
        RECT 2253.5600 534.5700 2256.5600 750.6700 ;
      LAYER met3 ;
        RECT 2457.6600 727.7200 2460.6600 728.2000 ;
        RECT 2457.6600 733.1600 2460.6600 733.6400 ;
        RECT 2445.3200 727.7200 2446.9200 728.2000 ;
        RECT 2445.3200 733.1600 2446.9200 733.6400 ;
        RECT 2457.6600 738.6000 2460.6600 739.0800 ;
        RECT 2445.3200 738.6000 2446.9200 739.0800 ;
        RECT 2457.6600 716.8400 2460.6600 717.3200 ;
        RECT 2457.6600 722.2800 2460.6600 722.7600 ;
        RECT 2445.3200 716.8400 2446.9200 717.3200 ;
        RECT 2445.3200 722.2800 2446.9200 722.7600 ;
        RECT 2457.6600 700.5200 2460.6600 701.0000 ;
        RECT 2457.6600 705.9600 2460.6600 706.4400 ;
        RECT 2445.3200 700.5200 2446.9200 701.0000 ;
        RECT 2445.3200 705.9600 2446.9200 706.4400 ;
        RECT 2457.6600 711.4000 2460.6600 711.8800 ;
        RECT 2445.3200 711.4000 2446.9200 711.8800 ;
        RECT 2400.3200 727.7200 2401.9200 728.2000 ;
        RECT 2400.3200 733.1600 2401.9200 733.6400 ;
        RECT 2400.3200 738.6000 2401.9200 739.0800 ;
        RECT 2400.3200 716.8400 2401.9200 717.3200 ;
        RECT 2400.3200 722.2800 2401.9200 722.7600 ;
        RECT 2400.3200 700.5200 2401.9200 701.0000 ;
        RECT 2400.3200 705.9600 2401.9200 706.4400 ;
        RECT 2400.3200 711.4000 2401.9200 711.8800 ;
        RECT 2457.6600 684.2000 2460.6600 684.6800 ;
        RECT 2457.6600 689.6400 2460.6600 690.1200 ;
        RECT 2457.6600 695.0800 2460.6600 695.5600 ;
        RECT 2445.3200 684.2000 2446.9200 684.6800 ;
        RECT 2445.3200 689.6400 2446.9200 690.1200 ;
        RECT 2445.3200 695.0800 2446.9200 695.5600 ;
        RECT 2457.6600 673.3200 2460.6600 673.8000 ;
        RECT 2457.6600 678.7600 2460.6600 679.2400 ;
        RECT 2445.3200 673.3200 2446.9200 673.8000 ;
        RECT 2445.3200 678.7600 2446.9200 679.2400 ;
        RECT 2457.6600 657.0000 2460.6600 657.4800 ;
        RECT 2457.6600 662.4400 2460.6600 662.9200 ;
        RECT 2457.6600 667.8800 2460.6600 668.3600 ;
        RECT 2445.3200 657.0000 2446.9200 657.4800 ;
        RECT 2445.3200 662.4400 2446.9200 662.9200 ;
        RECT 2445.3200 667.8800 2446.9200 668.3600 ;
        RECT 2457.6600 646.1200 2460.6600 646.6000 ;
        RECT 2457.6600 651.5600 2460.6600 652.0400 ;
        RECT 2445.3200 646.1200 2446.9200 646.6000 ;
        RECT 2445.3200 651.5600 2446.9200 652.0400 ;
        RECT 2400.3200 684.2000 2401.9200 684.6800 ;
        RECT 2400.3200 689.6400 2401.9200 690.1200 ;
        RECT 2400.3200 695.0800 2401.9200 695.5600 ;
        RECT 2400.3200 673.3200 2401.9200 673.8000 ;
        RECT 2400.3200 678.7600 2401.9200 679.2400 ;
        RECT 2400.3200 657.0000 2401.9200 657.4800 ;
        RECT 2400.3200 662.4400 2401.9200 662.9200 ;
        RECT 2400.3200 667.8800 2401.9200 668.3600 ;
        RECT 2400.3200 646.1200 2401.9200 646.6000 ;
        RECT 2400.3200 651.5600 2401.9200 652.0400 ;
        RECT 2355.3200 727.7200 2356.9200 728.2000 ;
        RECT 2355.3200 733.1600 2356.9200 733.6400 ;
        RECT 2355.3200 738.6000 2356.9200 739.0800 ;
        RECT 2310.3200 727.7200 2311.9200 728.2000 ;
        RECT 2310.3200 733.1600 2311.9200 733.6400 ;
        RECT 2310.3200 738.6000 2311.9200 739.0800 ;
        RECT 2355.3200 716.8400 2356.9200 717.3200 ;
        RECT 2355.3200 722.2800 2356.9200 722.7600 ;
        RECT 2355.3200 700.5200 2356.9200 701.0000 ;
        RECT 2355.3200 705.9600 2356.9200 706.4400 ;
        RECT 2355.3200 711.4000 2356.9200 711.8800 ;
        RECT 2310.3200 716.8400 2311.9200 717.3200 ;
        RECT 2310.3200 722.2800 2311.9200 722.7600 ;
        RECT 2310.3200 700.5200 2311.9200 701.0000 ;
        RECT 2310.3200 705.9600 2311.9200 706.4400 ;
        RECT 2310.3200 711.4000 2311.9200 711.8800 ;
        RECT 2265.3200 727.7200 2266.9200 728.2000 ;
        RECT 2265.3200 733.1600 2266.9200 733.6400 ;
        RECT 2253.5600 733.1600 2256.5600 733.6400 ;
        RECT 2253.5600 727.7200 2256.5600 728.2000 ;
        RECT 2253.5600 738.6000 2256.5600 739.0800 ;
        RECT 2265.3200 738.6000 2266.9200 739.0800 ;
        RECT 2265.3200 716.8400 2266.9200 717.3200 ;
        RECT 2265.3200 722.2800 2266.9200 722.7600 ;
        RECT 2253.5600 722.2800 2256.5600 722.7600 ;
        RECT 2253.5600 716.8400 2256.5600 717.3200 ;
        RECT 2265.3200 700.5200 2266.9200 701.0000 ;
        RECT 2265.3200 705.9600 2266.9200 706.4400 ;
        RECT 2253.5600 705.9600 2256.5600 706.4400 ;
        RECT 2253.5600 700.5200 2256.5600 701.0000 ;
        RECT 2253.5600 711.4000 2256.5600 711.8800 ;
        RECT 2265.3200 711.4000 2266.9200 711.8800 ;
        RECT 2355.3200 684.2000 2356.9200 684.6800 ;
        RECT 2355.3200 689.6400 2356.9200 690.1200 ;
        RECT 2355.3200 695.0800 2356.9200 695.5600 ;
        RECT 2355.3200 673.3200 2356.9200 673.8000 ;
        RECT 2355.3200 678.7600 2356.9200 679.2400 ;
        RECT 2310.3200 684.2000 2311.9200 684.6800 ;
        RECT 2310.3200 689.6400 2311.9200 690.1200 ;
        RECT 2310.3200 695.0800 2311.9200 695.5600 ;
        RECT 2310.3200 673.3200 2311.9200 673.8000 ;
        RECT 2310.3200 678.7600 2311.9200 679.2400 ;
        RECT 2355.3200 657.0000 2356.9200 657.4800 ;
        RECT 2355.3200 662.4400 2356.9200 662.9200 ;
        RECT 2355.3200 667.8800 2356.9200 668.3600 ;
        RECT 2355.3200 646.1200 2356.9200 646.6000 ;
        RECT 2355.3200 651.5600 2356.9200 652.0400 ;
        RECT 2310.3200 657.0000 2311.9200 657.4800 ;
        RECT 2310.3200 662.4400 2311.9200 662.9200 ;
        RECT 2310.3200 667.8800 2311.9200 668.3600 ;
        RECT 2310.3200 646.1200 2311.9200 646.6000 ;
        RECT 2310.3200 651.5600 2311.9200 652.0400 ;
        RECT 2265.3200 684.2000 2266.9200 684.6800 ;
        RECT 2265.3200 689.6400 2266.9200 690.1200 ;
        RECT 2265.3200 695.0800 2266.9200 695.5600 ;
        RECT 2253.5600 684.2000 2256.5600 684.6800 ;
        RECT 2253.5600 689.6400 2256.5600 690.1200 ;
        RECT 2253.5600 695.0800 2256.5600 695.5600 ;
        RECT 2265.3200 673.3200 2266.9200 673.8000 ;
        RECT 2265.3200 678.7600 2266.9200 679.2400 ;
        RECT 2253.5600 673.3200 2256.5600 673.8000 ;
        RECT 2253.5600 678.7600 2256.5600 679.2400 ;
        RECT 2265.3200 657.0000 2266.9200 657.4800 ;
        RECT 2265.3200 662.4400 2266.9200 662.9200 ;
        RECT 2265.3200 667.8800 2266.9200 668.3600 ;
        RECT 2253.5600 657.0000 2256.5600 657.4800 ;
        RECT 2253.5600 662.4400 2256.5600 662.9200 ;
        RECT 2253.5600 667.8800 2256.5600 668.3600 ;
        RECT 2265.3200 646.1200 2266.9200 646.6000 ;
        RECT 2265.3200 651.5600 2266.9200 652.0400 ;
        RECT 2253.5600 646.1200 2256.5600 646.6000 ;
        RECT 2253.5600 651.5600 2256.5600 652.0400 ;
        RECT 2457.6600 629.8000 2460.6600 630.2800 ;
        RECT 2457.6600 635.2400 2460.6600 635.7200 ;
        RECT 2457.6600 640.6800 2460.6600 641.1600 ;
        RECT 2445.3200 629.8000 2446.9200 630.2800 ;
        RECT 2445.3200 635.2400 2446.9200 635.7200 ;
        RECT 2445.3200 640.6800 2446.9200 641.1600 ;
        RECT 2457.6600 618.9200 2460.6600 619.4000 ;
        RECT 2457.6600 624.3600 2460.6600 624.8400 ;
        RECT 2445.3200 618.9200 2446.9200 619.4000 ;
        RECT 2445.3200 624.3600 2446.9200 624.8400 ;
        RECT 2457.6600 602.6000 2460.6600 603.0800 ;
        RECT 2457.6600 608.0400 2460.6600 608.5200 ;
        RECT 2457.6600 613.4800 2460.6600 613.9600 ;
        RECT 2445.3200 602.6000 2446.9200 603.0800 ;
        RECT 2445.3200 608.0400 2446.9200 608.5200 ;
        RECT 2445.3200 613.4800 2446.9200 613.9600 ;
        RECT 2457.6600 591.7200 2460.6600 592.2000 ;
        RECT 2457.6600 597.1600 2460.6600 597.6400 ;
        RECT 2445.3200 591.7200 2446.9200 592.2000 ;
        RECT 2445.3200 597.1600 2446.9200 597.6400 ;
        RECT 2400.3200 629.8000 2401.9200 630.2800 ;
        RECT 2400.3200 635.2400 2401.9200 635.7200 ;
        RECT 2400.3200 640.6800 2401.9200 641.1600 ;
        RECT 2400.3200 618.9200 2401.9200 619.4000 ;
        RECT 2400.3200 624.3600 2401.9200 624.8400 ;
        RECT 2400.3200 602.6000 2401.9200 603.0800 ;
        RECT 2400.3200 608.0400 2401.9200 608.5200 ;
        RECT 2400.3200 613.4800 2401.9200 613.9600 ;
        RECT 2400.3200 591.7200 2401.9200 592.2000 ;
        RECT 2400.3200 597.1600 2401.9200 597.6400 ;
        RECT 2457.6600 575.4000 2460.6600 575.8800 ;
        RECT 2457.6600 580.8400 2460.6600 581.3200 ;
        RECT 2457.6600 586.2800 2460.6600 586.7600 ;
        RECT 2445.3200 575.4000 2446.9200 575.8800 ;
        RECT 2445.3200 580.8400 2446.9200 581.3200 ;
        RECT 2445.3200 586.2800 2446.9200 586.7600 ;
        RECT 2457.6600 564.5200 2460.6600 565.0000 ;
        RECT 2457.6600 569.9600 2460.6600 570.4400 ;
        RECT 2445.3200 564.5200 2446.9200 565.0000 ;
        RECT 2445.3200 569.9600 2446.9200 570.4400 ;
        RECT 2457.6600 548.2000 2460.6600 548.6800 ;
        RECT 2457.6600 553.6400 2460.6600 554.1200 ;
        RECT 2457.6600 559.0800 2460.6600 559.5600 ;
        RECT 2445.3200 548.2000 2446.9200 548.6800 ;
        RECT 2445.3200 553.6400 2446.9200 554.1200 ;
        RECT 2445.3200 559.0800 2446.9200 559.5600 ;
        RECT 2457.6600 542.7600 2460.6600 543.2400 ;
        RECT 2445.3200 542.7600 2446.9200 543.2400 ;
        RECT 2400.3200 575.4000 2401.9200 575.8800 ;
        RECT 2400.3200 580.8400 2401.9200 581.3200 ;
        RECT 2400.3200 586.2800 2401.9200 586.7600 ;
        RECT 2400.3200 564.5200 2401.9200 565.0000 ;
        RECT 2400.3200 569.9600 2401.9200 570.4400 ;
        RECT 2400.3200 548.2000 2401.9200 548.6800 ;
        RECT 2400.3200 553.6400 2401.9200 554.1200 ;
        RECT 2400.3200 559.0800 2401.9200 559.5600 ;
        RECT 2400.3200 542.7600 2401.9200 543.2400 ;
        RECT 2355.3200 629.8000 2356.9200 630.2800 ;
        RECT 2355.3200 635.2400 2356.9200 635.7200 ;
        RECT 2355.3200 640.6800 2356.9200 641.1600 ;
        RECT 2355.3200 618.9200 2356.9200 619.4000 ;
        RECT 2355.3200 624.3600 2356.9200 624.8400 ;
        RECT 2310.3200 629.8000 2311.9200 630.2800 ;
        RECT 2310.3200 635.2400 2311.9200 635.7200 ;
        RECT 2310.3200 640.6800 2311.9200 641.1600 ;
        RECT 2310.3200 618.9200 2311.9200 619.4000 ;
        RECT 2310.3200 624.3600 2311.9200 624.8400 ;
        RECT 2355.3200 602.6000 2356.9200 603.0800 ;
        RECT 2355.3200 608.0400 2356.9200 608.5200 ;
        RECT 2355.3200 613.4800 2356.9200 613.9600 ;
        RECT 2355.3200 591.7200 2356.9200 592.2000 ;
        RECT 2355.3200 597.1600 2356.9200 597.6400 ;
        RECT 2310.3200 602.6000 2311.9200 603.0800 ;
        RECT 2310.3200 608.0400 2311.9200 608.5200 ;
        RECT 2310.3200 613.4800 2311.9200 613.9600 ;
        RECT 2310.3200 591.7200 2311.9200 592.2000 ;
        RECT 2310.3200 597.1600 2311.9200 597.6400 ;
        RECT 2265.3200 629.8000 2266.9200 630.2800 ;
        RECT 2265.3200 635.2400 2266.9200 635.7200 ;
        RECT 2265.3200 640.6800 2266.9200 641.1600 ;
        RECT 2253.5600 629.8000 2256.5600 630.2800 ;
        RECT 2253.5600 635.2400 2256.5600 635.7200 ;
        RECT 2253.5600 640.6800 2256.5600 641.1600 ;
        RECT 2265.3200 618.9200 2266.9200 619.4000 ;
        RECT 2265.3200 624.3600 2266.9200 624.8400 ;
        RECT 2253.5600 618.9200 2256.5600 619.4000 ;
        RECT 2253.5600 624.3600 2256.5600 624.8400 ;
        RECT 2265.3200 602.6000 2266.9200 603.0800 ;
        RECT 2265.3200 608.0400 2266.9200 608.5200 ;
        RECT 2265.3200 613.4800 2266.9200 613.9600 ;
        RECT 2253.5600 602.6000 2256.5600 603.0800 ;
        RECT 2253.5600 608.0400 2256.5600 608.5200 ;
        RECT 2253.5600 613.4800 2256.5600 613.9600 ;
        RECT 2265.3200 591.7200 2266.9200 592.2000 ;
        RECT 2265.3200 597.1600 2266.9200 597.6400 ;
        RECT 2253.5600 591.7200 2256.5600 592.2000 ;
        RECT 2253.5600 597.1600 2256.5600 597.6400 ;
        RECT 2355.3200 575.4000 2356.9200 575.8800 ;
        RECT 2355.3200 580.8400 2356.9200 581.3200 ;
        RECT 2355.3200 586.2800 2356.9200 586.7600 ;
        RECT 2355.3200 564.5200 2356.9200 565.0000 ;
        RECT 2355.3200 569.9600 2356.9200 570.4400 ;
        RECT 2310.3200 575.4000 2311.9200 575.8800 ;
        RECT 2310.3200 580.8400 2311.9200 581.3200 ;
        RECT 2310.3200 586.2800 2311.9200 586.7600 ;
        RECT 2310.3200 564.5200 2311.9200 565.0000 ;
        RECT 2310.3200 569.9600 2311.9200 570.4400 ;
        RECT 2355.3200 548.2000 2356.9200 548.6800 ;
        RECT 2355.3200 553.6400 2356.9200 554.1200 ;
        RECT 2355.3200 559.0800 2356.9200 559.5600 ;
        RECT 2355.3200 542.7600 2356.9200 543.2400 ;
        RECT 2310.3200 548.2000 2311.9200 548.6800 ;
        RECT 2310.3200 553.6400 2311.9200 554.1200 ;
        RECT 2310.3200 559.0800 2311.9200 559.5600 ;
        RECT 2310.3200 542.7600 2311.9200 543.2400 ;
        RECT 2265.3200 575.4000 2266.9200 575.8800 ;
        RECT 2265.3200 580.8400 2266.9200 581.3200 ;
        RECT 2265.3200 586.2800 2266.9200 586.7600 ;
        RECT 2253.5600 575.4000 2256.5600 575.8800 ;
        RECT 2253.5600 580.8400 2256.5600 581.3200 ;
        RECT 2253.5600 586.2800 2256.5600 586.7600 ;
        RECT 2265.3200 564.5200 2266.9200 565.0000 ;
        RECT 2265.3200 569.9600 2266.9200 570.4400 ;
        RECT 2253.5600 564.5200 2256.5600 565.0000 ;
        RECT 2253.5600 569.9600 2256.5600 570.4400 ;
        RECT 2265.3200 548.2000 2266.9200 548.6800 ;
        RECT 2265.3200 553.6400 2266.9200 554.1200 ;
        RECT 2265.3200 559.0800 2266.9200 559.5600 ;
        RECT 2253.5600 548.2000 2256.5600 548.6800 ;
        RECT 2253.5600 553.6400 2256.5600 554.1200 ;
        RECT 2253.5600 559.0800 2256.5600 559.5600 ;
        RECT 2253.5600 542.7600 2256.5600 543.2400 ;
        RECT 2265.3200 542.7600 2266.9200 543.2400 ;
        RECT 2253.5600 747.6700 2460.6600 750.6700 ;
        RECT 2253.5600 534.5700 2460.6600 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 304.9300 2446.9200 521.0300 ;
        RECT 2400.3200 304.9300 2401.9200 521.0300 ;
        RECT 2355.3200 304.9300 2356.9200 521.0300 ;
        RECT 2310.3200 304.9300 2311.9200 521.0300 ;
        RECT 2265.3200 304.9300 2266.9200 521.0300 ;
        RECT 2457.6600 304.9300 2460.6600 521.0300 ;
        RECT 2253.5600 304.9300 2256.5600 521.0300 ;
      LAYER met3 ;
        RECT 2457.6600 498.0800 2460.6600 498.5600 ;
        RECT 2457.6600 503.5200 2460.6600 504.0000 ;
        RECT 2445.3200 498.0800 2446.9200 498.5600 ;
        RECT 2445.3200 503.5200 2446.9200 504.0000 ;
        RECT 2457.6600 508.9600 2460.6600 509.4400 ;
        RECT 2445.3200 508.9600 2446.9200 509.4400 ;
        RECT 2457.6600 487.2000 2460.6600 487.6800 ;
        RECT 2457.6600 492.6400 2460.6600 493.1200 ;
        RECT 2445.3200 487.2000 2446.9200 487.6800 ;
        RECT 2445.3200 492.6400 2446.9200 493.1200 ;
        RECT 2457.6600 470.8800 2460.6600 471.3600 ;
        RECT 2457.6600 476.3200 2460.6600 476.8000 ;
        RECT 2445.3200 470.8800 2446.9200 471.3600 ;
        RECT 2445.3200 476.3200 2446.9200 476.8000 ;
        RECT 2457.6600 481.7600 2460.6600 482.2400 ;
        RECT 2445.3200 481.7600 2446.9200 482.2400 ;
        RECT 2400.3200 498.0800 2401.9200 498.5600 ;
        RECT 2400.3200 503.5200 2401.9200 504.0000 ;
        RECT 2400.3200 508.9600 2401.9200 509.4400 ;
        RECT 2400.3200 487.2000 2401.9200 487.6800 ;
        RECT 2400.3200 492.6400 2401.9200 493.1200 ;
        RECT 2400.3200 470.8800 2401.9200 471.3600 ;
        RECT 2400.3200 476.3200 2401.9200 476.8000 ;
        RECT 2400.3200 481.7600 2401.9200 482.2400 ;
        RECT 2457.6600 454.5600 2460.6600 455.0400 ;
        RECT 2457.6600 460.0000 2460.6600 460.4800 ;
        RECT 2457.6600 465.4400 2460.6600 465.9200 ;
        RECT 2445.3200 454.5600 2446.9200 455.0400 ;
        RECT 2445.3200 460.0000 2446.9200 460.4800 ;
        RECT 2445.3200 465.4400 2446.9200 465.9200 ;
        RECT 2457.6600 443.6800 2460.6600 444.1600 ;
        RECT 2457.6600 449.1200 2460.6600 449.6000 ;
        RECT 2445.3200 443.6800 2446.9200 444.1600 ;
        RECT 2445.3200 449.1200 2446.9200 449.6000 ;
        RECT 2457.6600 427.3600 2460.6600 427.8400 ;
        RECT 2457.6600 432.8000 2460.6600 433.2800 ;
        RECT 2457.6600 438.2400 2460.6600 438.7200 ;
        RECT 2445.3200 427.3600 2446.9200 427.8400 ;
        RECT 2445.3200 432.8000 2446.9200 433.2800 ;
        RECT 2445.3200 438.2400 2446.9200 438.7200 ;
        RECT 2457.6600 416.4800 2460.6600 416.9600 ;
        RECT 2457.6600 421.9200 2460.6600 422.4000 ;
        RECT 2445.3200 416.4800 2446.9200 416.9600 ;
        RECT 2445.3200 421.9200 2446.9200 422.4000 ;
        RECT 2400.3200 454.5600 2401.9200 455.0400 ;
        RECT 2400.3200 460.0000 2401.9200 460.4800 ;
        RECT 2400.3200 465.4400 2401.9200 465.9200 ;
        RECT 2400.3200 443.6800 2401.9200 444.1600 ;
        RECT 2400.3200 449.1200 2401.9200 449.6000 ;
        RECT 2400.3200 427.3600 2401.9200 427.8400 ;
        RECT 2400.3200 432.8000 2401.9200 433.2800 ;
        RECT 2400.3200 438.2400 2401.9200 438.7200 ;
        RECT 2400.3200 416.4800 2401.9200 416.9600 ;
        RECT 2400.3200 421.9200 2401.9200 422.4000 ;
        RECT 2355.3200 498.0800 2356.9200 498.5600 ;
        RECT 2355.3200 503.5200 2356.9200 504.0000 ;
        RECT 2355.3200 508.9600 2356.9200 509.4400 ;
        RECT 2310.3200 498.0800 2311.9200 498.5600 ;
        RECT 2310.3200 503.5200 2311.9200 504.0000 ;
        RECT 2310.3200 508.9600 2311.9200 509.4400 ;
        RECT 2355.3200 487.2000 2356.9200 487.6800 ;
        RECT 2355.3200 492.6400 2356.9200 493.1200 ;
        RECT 2355.3200 470.8800 2356.9200 471.3600 ;
        RECT 2355.3200 476.3200 2356.9200 476.8000 ;
        RECT 2355.3200 481.7600 2356.9200 482.2400 ;
        RECT 2310.3200 487.2000 2311.9200 487.6800 ;
        RECT 2310.3200 492.6400 2311.9200 493.1200 ;
        RECT 2310.3200 470.8800 2311.9200 471.3600 ;
        RECT 2310.3200 476.3200 2311.9200 476.8000 ;
        RECT 2310.3200 481.7600 2311.9200 482.2400 ;
        RECT 2265.3200 498.0800 2266.9200 498.5600 ;
        RECT 2265.3200 503.5200 2266.9200 504.0000 ;
        RECT 2253.5600 503.5200 2256.5600 504.0000 ;
        RECT 2253.5600 498.0800 2256.5600 498.5600 ;
        RECT 2253.5600 508.9600 2256.5600 509.4400 ;
        RECT 2265.3200 508.9600 2266.9200 509.4400 ;
        RECT 2265.3200 487.2000 2266.9200 487.6800 ;
        RECT 2265.3200 492.6400 2266.9200 493.1200 ;
        RECT 2253.5600 492.6400 2256.5600 493.1200 ;
        RECT 2253.5600 487.2000 2256.5600 487.6800 ;
        RECT 2265.3200 470.8800 2266.9200 471.3600 ;
        RECT 2265.3200 476.3200 2266.9200 476.8000 ;
        RECT 2253.5600 476.3200 2256.5600 476.8000 ;
        RECT 2253.5600 470.8800 2256.5600 471.3600 ;
        RECT 2253.5600 481.7600 2256.5600 482.2400 ;
        RECT 2265.3200 481.7600 2266.9200 482.2400 ;
        RECT 2355.3200 454.5600 2356.9200 455.0400 ;
        RECT 2355.3200 460.0000 2356.9200 460.4800 ;
        RECT 2355.3200 465.4400 2356.9200 465.9200 ;
        RECT 2355.3200 443.6800 2356.9200 444.1600 ;
        RECT 2355.3200 449.1200 2356.9200 449.6000 ;
        RECT 2310.3200 454.5600 2311.9200 455.0400 ;
        RECT 2310.3200 460.0000 2311.9200 460.4800 ;
        RECT 2310.3200 465.4400 2311.9200 465.9200 ;
        RECT 2310.3200 443.6800 2311.9200 444.1600 ;
        RECT 2310.3200 449.1200 2311.9200 449.6000 ;
        RECT 2355.3200 427.3600 2356.9200 427.8400 ;
        RECT 2355.3200 432.8000 2356.9200 433.2800 ;
        RECT 2355.3200 438.2400 2356.9200 438.7200 ;
        RECT 2355.3200 416.4800 2356.9200 416.9600 ;
        RECT 2355.3200 421.9200 2356.9200 422.4000 ;
        RECT 2310.3200 427.3600 2311.9200 427.8400 ;
        RECT 2310.3200 432.8000 2311.9200 433.2800 ;
        RECT 2310.3200 438.2400 2311.9200 438.7200 ;
        RECT 2310.3200 416.4800 2311.9200 416.9600 ;
        RECT 2310.3200 421.9200 2311.9200 422.4000 ;
        RECT 2265.3200 454.5600 2266.9200 455.0400 ;
        RECT 2265.3200 460.0000 2266.9200 460.4800 ;
        RECT 2265.3200 465.4400 2266.9200 465.9200 ;
        RECT 2253.5600 454.5600 2256.5600 455.0400 ;
        RECT 2253.5600 460.0000 2256.5600 460.4800 ;
        RECT 2253.5600 465.4400 2256.5600 465.9200 ;
        RECT 2265.3200 443.6800 2266.9200 444.1600 ;
        RECT 2265.3200 449.1200 2266.9200 449.6000 ;
        RECT 2253.5600 443.6800 2256.5600 444.1600 ;
        RECT 2253.5600 449.1200 2256.5600 449.6000 ;
        RECT 2265.3200 427.3600 2266.9200 427.8400 ;
        RECT 2265.3200 432.8000 2266.9200 433.2800 ;
        RECT 2265.3200 438.2400 2266.9200 438.7200 ;
        RECT 2253.5600 427.3600 2256.5600 427.8400 ;
        RECT 2253.5600 432.8000 2256.5600 433.2800 ;
        RECT 2253.5600 438.2400 2256.5600 438.7200 ;
        RECT 2265.3200 416.4800 2266.9200 416.9600 ;
        RECT 2265.3200 421.9200 2266.9200 422.4000 ;
        RECT 2253.5600 416.4800 2256.5600 416.9600 ;
        RECT 2253.5600 421.9200 2256.5600 422.4000 ;
        RECT 2457.6600 400.1600 2460.6600 400.6400 ;
        RECT 2457.6600 405.6000 2460.6600 406.0800 ;
        RECT 2457.6600 411.0400 2460.6600 411.5200 ;
        RECT 2445.3200 400.1600 2446.9200 400.6400 ;
        RECT 2445.3200 405.6000 2446.9200 406.0800 ;
        RECT 2445.3200 411.0400 2446.9200 411.5200 ;
        RECT 2457.6600 389.2800 2460.6600 389.7600 ;
        RECT 2457.6600 394.7200 2460.6600 395.2000 ;
        RECT 2445.3200 389.2800 2446.9200 389.7600 ;
        RECT 2445.3200 394.7200 2446.9200 395.2000 ;
        RECT 2457.6600 372.9600 2460.6600 373.4400 ;
        RECT 2457.6600 378.4000 2460.6600 378.8800 ;
        RECT 2457.6600 383.8400 2460.6600 384.3200 ;
        RECT 2445.3200 372.9600 2446.9200 373.4400 ;
        RECT 2445.3200 378.4000 2446.9200 378.8800 ;
        RECT 2445.3200 383.8400 2446.9200 384.3200 ;
        RECT 2457.6600 362.0800 2460.6600 362.5600 ;
        RECT 2457.6600 367.5200 2460.6600 368.0000 ;
        RECT 2445.3200 362.0800 2446.9200 362.5600 ;
        RECT 2445.3200 367.5200 2446.9200 368.0000 ;
        RECT 2400.3200 400.1600 2401.9200 400.6400 ;
        RECT 2400.3200 405.6000 2401.9200 406.0800 ;
        RECT 2400.3200 411.0400 2401.9200 411.5200 ;
        RECT 2400.3200 389.2800 2401.9200 389.7600 ;
        RECT 2400.3200 394.7200 2401.9200 395.2000 ;
        RECT 2400.3200 372.9600 2401.9200 373.4400 ;
        RECT 2400.3200 378.4000 2401.9200 378.8800 ;
        RECT 2400.3200 383.8400 2401.9200 384.3200 ;
        RECT 2400.3200 362.0800 2401.9200 362.5600 ;
        RECT 2400.3200 367.5200 2401.9200 368.0000 ;
        RECT 2457.6600 345.7600 2460.6600 346.2400 ;
        RECT 2457.6600 351.2000 2460.6600 351.6800 ;
        RECT 2457.6600 356.6400 2460.6600 357.1200 ;
        RECT 2445.3200 345.7600 2446.9200 346.2400 ;
        RECT 2445.3200 351.2000 2446.9200 351.6800 ;
        RECT 2445.3200 356.6400 2446.9200 357.1200 ;
        RECT 2457.6600 334.8800 2460.6600 335.3600 ;
        RECT 2457.6600 340.3200 2460.6600 340.8000 ;
        RECT 2445.3200 334.8800 2446.9200 335.3600 ;
        RECT 2445.3200 340.3200 2446.9200 340.8000 ;
        RECT 2457.6600 318.5600 2460.6600 319.0400 ;
        RECT 2457.6600 324.0000 2460.6600 324.4800 ;
        RECT 2457.6600 329.4400 2460.6600 329.9200 ;
        RECT 2445.3200 318.5600 2446.9200 319.0400 ;
        RECT 2445.3200 324.0000 2446.9200 324.4800 ;
        RECT 2445.3200 329.4400 2446.9200 329.9200 ;
        RECT 2457.6600 313.1200 2460.6600 313.6000 ;
        RECT 2445.3200 313.1200 2446.9200 313.6000 ;
        RECT 2400.3200 345.7600 2401.9200 346.2400 ;
        RECT 2400.3200 351.2000 2401.9200 351.6800 ;
        RECT 2400.3200 356.6400 2401.9200 357.1200 ;
        RECT 2400.3200 334.8800 2401.9200 335.3600 ;
        RECT 2400.3200 340.3200 2401.9200 340.8000 ;
        RECT 2400.3200 318.5600 2401.9200 319.0400 ;
        RECT 2400.3200 324.0000 2401.9200 324.4800 ;
        RECT 2400.3200 329.4400 2401.9200 329.9200 ;
        RECT 2400.3200 313.1200 2401.9200 313.6000 ;
        RECT 2355.3200 400.1600 2356.9200 400.6400 ;
        RECT 2355.3200 405.6000 2356.9200 406.0800 ;
        RECT 2355.3200 411.0400 2356.9200 411.5200 ;
        RECT 2355.3200 389.2800 2356.9200 389.7600 ;
        RECT 2355.3200 394.7200 2356.9200 395.2000 ;
        RECT 2310.3200 400.1600 2311.9200 400.6400 ;
        RECT 2310.3200 405.6000 2311.9200 406.0800 ;
        RECT 2310.3200 411.0400 2311.9200 411.5200 ;
        RECT 2310.3200 389.2800 2311.9200 389.7600 ;
        RECT 2310.3200 394.7200 2311.9200 395.2000 ;
        RECT 2355.3200 372.9600 2356.9200 373.4400 ;
        RECT 2355.3200 378.4000 2356.9200 378.8800 ;
        RECT 2355.3200 383.8400 2356.9200 384.3200 ;
        RECT 2355.3200 362.0800 2356.9200 362.5600 ;
        RECT 2355.3200 367.5200 2356.9200 368.0000 ;
        RECT 2310.3200 372.9600 2311.9200 373.4400 ;
        RECT 2310.3200 378.4000 2311.9200 378.8800 ;
        RECT 2310.3200 383.8400 2311.9200 384.3200 ;
        RECT 2310.3200 362.0800 2311.9200 362.5600 ;
        RECT 2310.3200 367.5200 2311.9200 368.0000 ;
        RECT 2265.3200 400.1600 2266.9200 400.6400 ;
        RECT 2265.3200 405.6000 2266.9200 406.0800 ;
        RECT 2265.3200 411.0400 2266.9200 411.5200 ;
        RECT 2253.5600 400.1600 2256.5600 400.6400 ;
        RECT 2253.5600 405.6000 2256.5600 406.0800 ;
        RECT 2253.5600 411.0400 2256.5600 411.5200 ;
        RECT 2265.3200 389.2800 2266.9200 389.7600 ;
        RECT 2265.3200 394.7200 2266.9200 395.2000 ;
        RECT 2253.5600 389.2800 2256.5600 389.7600 ;
        RECT 2253.5600 394.7200 2256.5600 395.2000 ;
        RECT 2265.3200 372.9600 2266.9200 373.4400 ;
        RECT 2265.3200 378.4000 2266.9200 378.8800 ;
        RECT 2265.3200 383.8400 2266.9200 384.3200 ;
        RECT 2253.5600 372.9600 2256.5600 373.4400 ;
        RECT 2253.5600 378.4000 2256.5600 378.8800 ;
        RECT 2253.5600 383.8400 2256.5600 384.3200 ;
        RECT 2265.3200 362.0800 2266.9200 362.5600 ;
        RECT 2265.3200 367.5200 2266.9200 368.0000 ;
        RECT 2253.5600 362.0800 2256.5600 362.5600 ;
        RECT 2253.5600 367.5200 2256.5600 368.0000 ;
        RECT 2355.3200 345.7600 2356.9200 346.2400 ;
        RECT 2355.3200 351.2000 2356.9200 351.6800 ;
        RECT 2355.3200 356.6400 2356.9200 357.1200 ;
        RECT 2355.3200 334.8800 2356.9200 335.3600 ;
        RECT 2355.3200 340.3200 2356.9200 340.8000 ;
        RECT 2310.3200 345.7600 2311.9200 346.2400 ;
        RECT 2310.3200 351.2000 2311.9200 351.6800 ;
        RECT 2310.3200 356.6400 2311.9200 357.1200 ;
        RECT 2310.3200 334.8800 2311.9200 335.3600 ;
        RECT 2310.3200 340.3200 2311.9200 340.8000 ;
        RECT 2355.3200 318.5600 2356.9200 319.0400 ;
        RECT 2355.3200 324.0000 2356.9200 324.4800 ;
        RECT 2355.3200 329.4400 2356.9200 329.9200 ;
        RECT 2355.3200 313.1200 2356.9200 313.6000 ;
        RECT 2310.3200 318.5600 2311.9200 319.0400 ;
        RECT 2310.3200 324.0000 2311.9200 324.4800 ;
        RECT 2310.3200 329.4400 2311.9200 329.9200 ;
        RECT 2310.3200 313.1200 2311.9200 313.6000 ;
        RECT 2265.3200 345.7600 2266.9200 346.2400 ;
        RECT 2265.3200 351.2000 2266.9200 351.6800 ;
        RECT 2265.3200 356.6400 2266.9200 357.1200 ;
        RECT 2253.5600 345.7600 2256.5600 346.2400 ;
        RECT 2253.5600 351.2000 2256.5600 351.6800 ;
        RECT 2253.5600 356.6400 2256.5600 357.1200 ;
        RECT 2265.3200 334.8800 2266.9200 335.3600 ;
        RECT 2265.3200 340.3200 2266.9200 340.8000 ;
        RECT 2253.5600 334.8800 2256.5600 335.3600 ;
        RECT 2253.5600 340.3200 2256.5600 340.8000 ;
        RECT 2265.3200 318.5600 2266.9200 319.0400 ;
        RECT 2265.3200 324.0000 2266.9200 324.4800 ;
        RECT 2265.3200 329.4400 2266.9200 329.9200 ;
        RECT 2253.5600 318.5600 2256.5600 319.0400 ;
        RECT 2253.5600 324.0000 2256.5600 324.4800 ;
        RECT 2253.5600 329.4400 2256.5600 329.9200 ;
        RECT 2253.5600 313.1200 2256.5600 313.6000 ;
        RECT 2265.3200 313.1200 2266.9200 313.6000 ;
        RECT 2253.5600 518.0300 2460.6600 521.0300 ;
        RECT 2253.5600 304.9300 2460.6600 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 75.2900 2446.9200 291.3900 ;
        RECT 2400.3200 75.2900 2401.9200 291.3900 ;
        RECT 2355.3200 75.2900 2356.9200 291.3900 ;
        RECT 2310.3200 75.2900 2311.9200 291.3900 ;
        RECT 2265.3200 75.2900 2266.9200 291.3900 ;
        RECT 2457.6600 75.2900 2460.6600 291.3900 ;
        RECT 2253.5600 75.2900 2256.5600 291.3900 ;
      LAYER met3 ;
        RECT 2457.6600 268.4400 2460.6600 268.9200 ;
        RECT 2457.6600 273.8800 2460.6600 274.3600 ;
        RECT 2445.3200 268.4400 2446.9200 268.9200 ;
        RECT 2445.3200 273.8800 2446.9200 274.3600 ;
        RECT 2457.6600 279.3200 2460.6600 279.8000 ;
        RECT 2445.3200 279.3200 2446.9200 279.8000 ;
        RECT 2457.6600 257.5600 2460.6600 258.0400 ;
        RECT 2457.6600 263.0000 2460.6600 263.4800 ;
        RECT 2445.3200 257.5600 2446.9200 258.0400 ;
        RECT 2445.3200 263.0000 2446.9200 263.4800 ;
        RECT 2457.6600 241.2400 2460.6600 241.7200 ;
        RECT 2457.6600 246.6800 2460.6600 247.1600 ;
        RECT 2445.3200 241.2400 2446.9200 241.7200 ;
        RECT 2445.3200 246.6800 2446.9200 247.1600 ;
        RECT 2457.6600 252.1200 2460.6600 252.6000 ;
        RECT 2445.3200 252.1200 2446.9200 252.6000 ;
        RECT 2400.3200 268.4400 2401.9200 268.9200 ;
        RECT 2400.3200 273.8800 2401.9200 274.3600 ;
        RECT 2400.3200 279.3200 2401.9200 279.8000 ;
        RECT 2400.3200 257.5600 2401.9200 258.0400 ;
        RECT 2400.3200 263.0000 2401.9200 263.4800 ;
        RECT 2400.3200 241.2400 2401.9200 241.7200 ;
        RECT 2400.3200 246.6800 2401.9200 247.1600 ;
        RECT 2400.3200 252.1200 2401.9200 252.6000 ;
        RECT 2457.6600 224.9200 2460.6600 225.4000 ;
        RECT 2457.6600 230.3600 2460.6600 230.8400 ;
        RECT 2457.6600 235.8000 2460.6600 236.2800 ;
        RECT 2445.3200 224.9200 2446.9200 225.4000 ;
        RECT 2445.3200 230.3600 2446.9200 230.8400 ;
        RECT 2445.3200 235.8000 2446.9200 236.2800 ;
        RECT 2457.6600 214.0400 2460.6600 214.5200 ;
        RECT 2457.6600 219.4800 2460.6600 219.9600 ;
        RECT 2445.3200 214.0400 2446.9200 214.5200 ;
        RECT 2445.3200 219.4800 2446.9200 219.9600 ;
        RECT 2457.6600 197.7200 2460.6600 198.2000 ;
        RECT 2457.6600 203.1600 2460.6600 203.6400 ;
        RECT 2457.6600 208.6000 2460.6600 209.0800 ;
        RECT 2445.3200 197.7200 2446.9200 198.2000 ;
        RECT 2445.3200 203.1600 2446.9200 203.6400 ;
        RECT 2445.3200 208.6000 2446.9200 209.0800 ;
        RECT 2457.6600 186.8400 2460.6600 187.3200 ;
        RECT 2457.6600 192.2800 2460.6600 192.7600 ;
        RECT 2445.3200 186.8400 2446.9200 187.3200 ;
        RECT 2445.3200 192.2800 2446.9200 192.7600 ;
        RECT 2400.3200 224.9200 2401.9200 225.4000 ;
        RECT 2400.3200 230.3600 2401.9200 230.8400 ;
        RECT 2400.3200 235.8000 2401.9200 236.2800 ;
        RECT 2400.3200 214.0400 2401.9200 214.5200 ;
        RECT 2400.3200 219.4800 2401.9200 219.9600 ;
        RECT 2400.3200 197.7200 2401.9200 198.2000 ;
        RECT 2400.3200 203.1600 2401.9200 203.6400 ;
        RECT 2400.3200 208.6000 2401.9200 209.0800 ;
        RECT 2400.3200 186.8400 2401.9200 187.3200 ;
        RECT 2400.3200 192.2800 2401.9200 192.7600 ;
        RECT 2355.3200 268.4400 2356.9200 268.9200 ;
        RECT 2355.3200 273.8800 2356.9200 274.3600 ;
        RECT 2355.3200 279.3200 2356.9200 279.8000 ;
        RECT 2310.3200 268.4400 2311.9200 268.9200 ;
        RECT 2310.3200 273.8800 2311.9200 274.3600 ;
        RECT 2310.3200 279.3200 2311.9200 279.8000 ;
        RECT 2355.3200 257.5600 2356.9200 258.0400 ;
        RECT 2355.3200 263.0000 2356.9200 263.4800 ;
        RECT 2355.3200 241.2400 2356.9200 241.7200 ;
        RECT 2355.3200 246.6800 2356.9200 247.1600 ;
        RECT 2355.3200 252.1200 2356.9200 252.6000 ;
        RECT 2310.3200 257.5600 2311.9200 258.0400 ;
        RECT 2310.3200 263.0000 2311.9200 263.4800 ;
        RECT 2310.3200 241.2400 2311.9200 241.7200 ;
        RECT 2310.3200 246.6800 2311.9200 247.1600 ;
        RECT 2310.3200 252.1200 2311.9200 252.6000 ;
        RECT 2265.3200 268.4400 2266.9200 268.9200 ;
        RECT 2265.3200 273.8800 2266.9200 274.3600 ;
        RECT 2253.5600 273.8800 2256.5600 274.3600 ;
        RECT 2253.5600 268.4400 2256.5600 268.9200 ;
        RECT 2253.5600 279.3200 2256.5600 279.8000 ;
        RECT 2265.3200 279.3200 2266.9200 279.8000 ;
        RECT 2265.3200 257.5600 2266.9200 258.0400 ;
        RECT 2265.3200 263.0000 2266.9200 263.4800 ;
        RECT 2253.5600 263.0000 2256.5600 263.4800 ;
        RECT 2253.5600 257.5600 2256.5600 258.0400 ;
        RECT 2265.3200 241.2400 2266.9200 241.7200 ;
        RECT 2265.3200 246.6800 2266.9200 247.1600 ;
        RECT 2253.5600 246.6800 2256.5600 247.1600 ;
        RECT 2253.5600 241.2400 2256.5600 241.7200 ;
        RECT 2253.5600 252.1200 2256.5600 252.6000 ;
        RECT 2265.3200 252.1200 2266.9200 252.6000 ;
        RECT 2355.3200 224.9200 2356.9200 225.4000 ;
        RECT 2355.3200 230.3600 2356.9200 230.8400 ;
        RECT 2355.3200 235.8000 2356.9200 236.2800 ;
        RECT 2355.3200 214.0400 2356.9200 214.5200 ;
        RECT 2355.3200 219.4800 2356.9200 219.9600 ;
        RECT 2310.3200 224.9200 2311.9200 225.4000 ;
        RECT 2310.3200 230.3600 2311.9200 230.8400 ;
        RECT 2310.3200 235.8000 2311.9200 236.2800 ;
        RECT 2310.3200 214.0400 2311.9200 214.5200 ;
        RECT 2310.3200 219.4800 2311.9200 219.9600 ;
        RECT 2355.3200 197.7200 2356.9200 198.2000 ;
        RECT 2355.3200 203.1600 2356.9200 203.6400 ;
        RECT 2355.3200 208.6000 2356.9200 209.0800 ;
        RECT 2355.3200 186.8400 2356.9200 187.3200 ;
        RECT 2355.3200 192.2800 2356.9200 192.7600 ;
        RECT 2310.3200 197.7200 2311.9200 198.2000 ;
        RECT 2310.3200 203.1600 2311.9200 203.6400 ;
        RECT 2310.3200 208.6000 2311.9200 209.0800 ;
        RECT 2310.3200 186.8400 2311.9200 187.3200 ;
        RECT 2310.3200 192.2800 2311.9200 192.7600 ;
        RECT 2265.3200 224.9200 2266.9200 225.4000 ;
        RECT 2265.3200 230.3600 2266.9200 230.8400 ;
        RECT 2265.3200 235.8000 2266.9200 236.2800 ;
        RECT 2253.5600 224.9200 2256.5600 225.4000 ;
        RECT 2253.5600 230.3600 2256.5600 230.8400 ;
        RECT 2253.5600 235.8000 2256.5600 236.2800 ;
        RECT 2265.3200 214.0400 2266.9200 214.5200 ;
        RECT 2265.3200 219.4800 2266.9200 219.9600 ;
        RECT 2253.5600 214.0400 2256.5600 214.5200 ;
        RECT 2253.5600 219.4800 2256.5600 219.9600 ;
        RECT 2265.3200 197.7200 2266.9200 198.2000 ;
        RECT 2265.3200 203.1600 2266.9200 203.6400 ;
        RECT 2265.3200 208.6000 2266.9200 209.0800 ;
        RECT 2253.5600 197.7200 2256.5600 198.2000 ;
        RECT 2253.5600 203.1600 2256.5600 203.6400 ;
        RECT 2253.5600 208.6000 2256.5600 209.0800 ;
        RECT 2265.3200 186.8400 2266.9200 187.3200 ;
        RECT 2265.3200 192.2800 2266.9200 192.7600 ;
        RECT 2253.5600 186.8400 2256.5600 187.3200 ;
        RECT 2253.5600 192.2800 2256.5600 192.7600 ;
        RECT 2457.6600 170.5200 2460.6600 171.0000 ;
        RECT 2457.6600 175.9600 2460.6600 176.4400 ;
        RECT 2457.6600 181.4000 2460.6600 181.8800 ;
        RECT 2445.3200 170.5200 2446.9200 171.0000 ;
        RECT 2445.3200 175.9600 2446.9200 176.4400 ;
        RECT 2445.3200 181.4000 2446.9200 181.8800 ;
        RECT 2457.6600 159.6400 2460.6600 160.1200 ;
        RECT 2457.6600 165.0800 2460.6600 165.5600 ;
        RECT 2445.3200 159.6400 2446.9200 160.1200 ;
        RECT 2445.3200 165.0800 2446.9200 165.5600 ;
        RECT 2457.6600 143.3200 2460.6600 143.8000 ;
        RECT 2457.6600 148.7600 2460.6600 149.2400 ;
        RECT 2457.6600 154.2000 2460.6600 154.6800 ;
        RECT 2445.3200 143.3200 2446.9200 143.8000 ;
        RECT 2445.3200 148.7600 2446.9200 149.2400 ;
        RECT 2445.3200 154.2000 2446.9200 154.6800 ;
        RECT 2457.6600 132.4400 2460.6600 132.9200 ;
        RECT 2457.6600 137.8800 2460.6600 138.3600 ;
        RECT 2445.3200 132.4400 2446.9200 132.9200 ;
        RECT 2445.3200 137.8800 2446.9200 138.3600 ;
        RECT 2400.3200 170.5200 2401.9200 171.0000 ;
        RECT 2400.3200 175.9600 2401.9200 176.4400 ;
        RECT 2400.3200 181.4000 2401.9200 181.8800 ;
        RECT 2400.3200 159.6400 2401.9200 160.1200 ;
        RECT 2400.3200 165.0800 2401.9200 165.5600 ;
        RECT 2400.3200 143.3200 2401.9200 143.8000 ;
        RECT 2400.3200 148.7600 2401.9200 149.2400 ;
        RECT 2400.3200 154.2000 2401.9200 154.6800 ;
        RECT 2400.3200 132.4400 2401.9200 132.9200 ;
        RECT 2400.3200 137.8800 2401.9200 138.3600 ;
        RECT 2457.6600 116.1200 2460.6600 116.6000 ;
        RECT 2457.6600 121.5600 2460.6600 122.0400 ;
        RECT 2457.6600 127.0000 2460.6600 127.4800 ;
        RECT 2445.3200 116.1200 2446.9200 116.6000 ;
        RECT 2445.3200 121.5600 2446.9200 122.0400 ;
        RECT 2445.3200 127.0000 2446.9200 127.4800 ;
        RECT 2457.6600 105.2400 2460.6600 105.7200 ;
        RECT 2457.6600 110.6800 2460.6600 111.1600 ;
        RECT 2445.3200 105.2400 2446.9200 105.7200 ;
        RECT 2445.3200 110.6800 2446.9200 111.1600 ;
        RECT 2457.6600 88.9200 2460.6600 89.4000 ;
        RECT 2457.6600 94.3600 2460.6600 94.8400 ;
        RECT 2457.6600 99.8000 2460.6600 100.2800 ;
        RECT 2445.3200 88.9200 2446.9200 89.4000 ;
        RECT 2445.3200 94.3600 2446.9200 94.8400 ;
        RECT 2445.3200 99.8000 2446.9200 100.2800 ;
        RECT 2457.6600 83.4800 2460.6600 83.9600 ;
        RECT 2445.3200 83.4800 2446.9200 83.9600 ;
        RECT 2400.3200 116.1200 2401.9200 116.6000 ;
        RECT 2400.3200 121.5600 2401.9200 122.0400 ;
        RECT 2400.3200 127.0000 2401.9200 127.4800 ;
        RECT 2400.3200 105.2400 2401.9200 105.7200 ;
        RECT 2400.3200 110.6800 2401.9200 111.1600 ;
        RECT 2400.3200 88.9200 2401.9200 89.4000 ;
        RECT 2400.3200 94.3600 2401.9200 94.8400 ;
        RECT 2400.3200 99.8000 2401.9200 100.2800 ;
        RECT 2400.3200 83.4800 2401.9200 83.9600 ;
        RECT 2355.3200 170.5200 2356.9200 171.0000 ;
        RECT 2355.3200 175.9600 2356.9200 176.4400 ;
        RECT 2355.3200 181.4000 2356.9200 181.8800 ;
        RECT 2355.3200 159.6400 2356.9200 160.1200 ;
        RECT 2355.3200 165.0800 2356.9200 165.5600 ;
        RECT 2310.3200 170.5200 2311.9200 171.0000 ;
        RECT 2310.3200 175.9600 2311.9200 176.4400 ;
        RECT 2310.3200 181.4000 2311.9200 181.8800 ;
        RECT 2310.3200 159.6400 2311.9200 160.1200 ;
        RECT 2310.3200 165.0800 2311.9200 165.5600 ;
        RECT 2355.3200 143.3200 2356.9200 143.8000 ;
        RECT 2355.3200 148.7600 2356.9200 149.2400 ;
        RECT 2355.3200 154.2000 2356.9200 154.6800 ;
        RECT 2355.3200 132.4400 2356.9200 132.9200 ;
        RECT 2355.3200 137.8800 2356.9200 138.3600 ;
        RECT 2310.3200 143.3200 2311.9200 143.8000 ;
        RECT 2310.3200 148.7600 2311.9200 149.2400 ;
        RECT 2310.3200 154.2000 2311.9200 154.6800 ;
        RECT 2310.3200 132.4400 2311.9200 132.9200 ;
        RECT 2310.3200 137.8800 2311.9200 138.3600 ;
        RECT 2265.3200 170.5200 2266.9200 171.0000 ;
        RECT 2265.3200 175.9600 2266.9200 176.4400 ;
        RECT 2265.3200 181.4000 2266.9200 181.8800 ;
        RECT 2253.5600 170.5200 2256.5600 171.0000 ;
        RECT 2253.5600 175.9600 2256.5600 176.4400 ;
        RECT 2253.5600 181.4000 2256.5600 181.8800 ;
        RECT 2265.3200 159.6400 2266.9200 160.1200 ;
        RECT 2265.3200 165.0800 2266.9200 165.5600 ;
        RECT 2253.5600 159.6400 2256.5600 160.1200 ;
        RECT 2253.5600 165.0800 2256.5600 165.5600 ;
        RECT 2265.3200 143.3200 2266.9200 143.8000 ;
        RECT 2265.3200 148.7600 2266.9200 149.2400 ;
        RECT 2265.3200 154.2000 2266.9200 154.6800 ;
        RECT 2253.5600 143.3200 2256.5600 143.8000 ;
        RECT 2253.5600 148.7600 2256.5600 149.2400 ;
        RECT 2253.5600 154.2000 2256.5600 154.6800 ;
        RECT 2265.3200 132.4400 2266.9200 132.9200 ;
        RECT 2265.3200 137.8800 2266.9200 138.3600 ;
        RECT 2253.5600 132.4400 2256.5600 132.9200 ;
        RECT 2253.5600 137.8800 2256.5600 138.3600 ;
        RECT 2355.3200 116.1200 2356.9200 116.6000 ;
        RECT 2355.3200 121.5600 2356.9200 122.0400 ;
        RECT 2355.3200 127.0000 2356.9200 127.4800 ;
        RECT 2355.3200 105.2400 2356.9200 105.7200 ;
        RECT 2355.3200 110.6800 2356.9200 111.1600 ;
        RECT 2310.3200 116.1200 2311.9200 116.6000 ;
        RECT 2310.3200 121.5600 2311.9200 122.0400 ;
        RECT 2310.3200 127.0000 2311.9200 127.4800 ;
        RECT 2310.3200 105.2400 2311.9200 105.7200 ;
        RECT 2310.3200 110.6800 2311.9200 111.1600 ;
        RECT 2355.3200 88.9200 2356.9200 89.4000 ;
        RECT 2355.3200 94.3600 2356.9200 94.8400 ;
        RECT 2355.3200 99.8000 2356.9200 100.2800 ;
        RECT 2355.3200 83.4800 2356.9200 83.9600 ;
        RECT 2310.3200 88.9200 2311.9200 89.4000 ;
        RECT 2310.3200 94.3600 2311.9200 94.8400 ;
        RECT 2310.3200 99.8000 2311.9200 100.2800 ;
        RECT 2310.3200 83.4800 2311.9200 83.9600 ;
        RECT 2265.3200 116.1200 2266.9200 116.6000 ;
        RECT 2265.3200 121.5600 2266.9200 122.0400 ;
        RECT 2265.3200 127.0000 2266.9200 127.4800 ;
        RECT 2253.5600 116.1200 2256.5600 116.6000 ;
        RECT 2253.5600 121.5600 2256.5600 122.0400 ;
        RECT 2253.5600 127.0000 2256.5600 127.4800 ;
        RECT 2265.3200 105.2400 2266.9200 105.7200 ;
        RECT 2265.3200 110.6800 2266.9200 111.1600 ;
        RECT 2253.5600 105.2400 2256.5600 105.7200 ;
        RECT 2253.5600 110.6800 2256.5600 111.1600 ;
        RECT 2265.3200 88.9200 2266.9200 89.4000 ;
        RECT 2265.3200 94.3600 2266.9200 94.8400 ;
        RECT 2265.3200 99.8000 2266.9200 100.2800 ;
        RECT 2253.5600 88.9200 2256.5600 89.4000 ;
        RECT 2253.5600 94.3600 2256.5600 94.8400 ;
        RECT 2253.5600 99.8000 2256.5600 100.2800 ;
        RECT 2253.5600 83.4800 2256.5600 83.9600 ;
        RECT 2265.3200 83.4800 2266.9200 83.9600 ;
        RECT 2253.5600 288.3900 2460.6600 291.3900 ;
        RECT 2253.5600 75.2900 2460.6600 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 2254.5600 34.6700 2256.5600 61.6000 ;
        RECT 2457.6600 34.6700 2459.6600 61.6000 ;
      LAYER met3 ;
        RECT 2457.6600 51.3800 2459.6600 51.8600 ;
        RECT 2254.5600 51.3800 2256.5600 51.8600 ;
        RECT 2457.6600 45.9400 2459.6600 46.4200 ;
        RECT 2457.6600 40.5000 2459.6600 40.9800 ;
        RECT 2254.5600 45.9400 2256.5600 46.4200 ;
        RECT 2254.5600 40.5000 2256.5600 40.9800 ;
        RECT 2254.5600 59.6000 2459.6600 61.6000 ;
        RECT 2254.5600 34.6700 2459.6600 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 2601.3300 2446.9200 2817.4300 ;
        RECT 2400.3200 2601.3300 2401.9200 2817.4300 ;
        RECT 2355.3200 2601.3300 2356.9200 2817.4300 ;
        RECT 2310.3200 2601.3300 2311.9200 2817.4300 ;
        RECT 2265.3200 2601.3300 2266.9200 2817.4300 ;
        RECT 2457.6600 2601.3300 2460.6600 2817.4300 ;
        RECT 2253.5600 2601.3300 2256.5600 2817.4300 ;
      LAYER met3 ;
        RECT 2457.6600 2794.4800 2460.6600 2794.9600 ;
        RECT 2457.6600 2799.9200 2460.6600 2800.4000 ;
        RECT 2445.3200 2794.4800 2446.9200 2794.9600 ;
        RECT 2445.3200 2799.9200 2446.9200 2800.4000 ;
        RECT 2457.6600 2805.3600 2460.6600 2805.8400 ;
        RECT 2445.3200 2805.3600 2446.9200 2805.8400 ;
        RECT 2457.6600 2783.6000 2460.6600 2784.0800 ;
        RECT 2457.6600 2789.0400 2460.6600 2789.5200 ;
        RECT 2445.3200 2783.6000 2446.9200 2784.0800 ;
        RECT 2445.3200 2789.0400 2446.9200 2789.5200 ;
        RECT 2457.6600 2767.2800 2460.6600 2767.7600 ;
        RECT 2457.6600 2772.7200 2460.6600 2773.2000 ;
        RECT 2445.3200 2767.2800 2446.9200 2767.7600 ;
        RECT 2445.3200 2772.7200 2446.9200 2773.2000 ;
        RECT 2457.6600 2778.1600 2460.6600 2778.6400 ;
        RECT 2445.3200 2778.1600 2446.9200 2778.6400 ;
        RECT 2400.3200 2794.4800 2401.9200 2794.9600 ;
        RECT 2400.3200 2799.9200 2401.9200 2800.4000 ;
        RECT 2400.3200 2805.3600 2401.9200 2805.8400 ;
        RECT 2400.3200 2783.6000 2401.9200 2784.0800 ;
        RECT 2400.3200 2789.0400 2401.9200 2789.5200 ;
        RECT 2400.3200 2767.2800 2401.9200 2767.7600 ;
        RECT 2400.3200 2772.7200 2401.9200 2773.2000 ;
        RECT 2400.3200 2778.1600 2401.9200 2778.6400 ;
        RECT 2457.6600 2750.9600 2460.6600 2751.4400 ;
        RECT 2457.6600 2756.4000 2460.6600 2756.8800 ;
        RECT 2457.6600 2761.8400 2460.6600 2762.3200 ;
        RECT 2445.3200 2750.9600 2446.9200 2751.4400 ;
        RECT 2445.3200 2756.4000 2446.9200 2756.8800 ;
        RECT 2445.3200 2761.8400 2446.9200 2762.3200 ;
        RECT 2457.6600 2740.0800 2460.6600 2740.5600 ;
        RECT 2457.6600 2745.5200 2460.6600 2746.0000 ;
        RECT 2445.3200 2740.0800 2446.9200 2740.5600 ;
        RECT 2445.3200 2745.5200 2446.9200 2746.0000 ;
        RECT 2457.6600 2723.7600 2460.6600 2724.2400 ;
        RECT 2457.6600 2729.2000 2460.6600 2729.6800 ;
        RECT 2457.6600 2734.6400 2460.6600 2735.1200 ;
        RECT 2445.3200 2723.7600 2446.9200 2724.2400 ;
        RECT 2445.3200 2729.2000 2446.9200 2729.6800 ;
        RECT 2445.3200 2734.6400 2446.9200 2735.1200 ;
        RECT 2457.6600 2712.8800 2460.6600 2713.3600 ;
        RECT 2457.6600 2718.3200 2460.6600 2718.8000 ;
        RECT 2445.3200 2712.8800 2446.9200 2713.3600 ;
        RECT 2445.3200 2718.3200 2446.9200 2718.8000 ;
        RECT 2400.3200 2750.9600 2401.9200 2751.4400 ;
        RECT 2400.3200 2756.4000 2401.9200 2756.8800 ;
        RECT 2400.3200 2761.8400 2401.9200 2762.3200 ;
        RECT 2400.3200 2740.0800 2401.9200 2740.5600 ;
        RECT 2400.3200 2745.5200 2401.9200 2746.0000 ;
        RECT 2400.3200 2723.7600 2401.9200 2724.2400 ;
        RECT 2400.3200 2729.2000 2401.9200 2729.6800 ;
        RECT 2400.3200 2734.6400 2401.9200 2735.1200 ;
        RECT 2400.3200 2712.8800 2401.9200 2713.3600 ;
        RECT 2400.3200 2718.3200 2401.9200 2718.8000 ;
        RECT 2355.3200 2794.4800 2356.9200 2794.9600 ;
        RECT 2355.3200 2799.9200 2356.9200 2800.4000 ;
        RECT 2355.3200 2805.3600 2356.9200 2805.8400 ;
        RECT 2310.3200 2794.4800 2311.9200 2794.9600 ;
        RECT 2310.3200 2799.9200 2311.9200 2800.4000 ;
        RECT 2310.3200 2805.3600 2311.9200 2805.8400 ;
        RECT 2355.3200 2783.6000 2356.9200 2784.0800 ;
        RECT 2355.3200 2789.0400 2356.9200 2789.5200 ;
        RECT 2355.3200 2767.2800 2356.9200 2767.7600 ;
        RECT 2355.3200 2772.7200 2356.9200 2773.2000 ;
        RECT 2355.3200 2778.1600 2356.9200 2778.6400 ;
        RECT 2310.3200 2783.6000 2311.9200 2784.0800 ;
        RECT 2310.3200 2789.0400 2311.9200 2789.5200 ;
        RECT 2310.3200 2767.2800 2311.9200 2767.7600 ;
        RECT 2310.3200 2772.7200 2311.9200 2773.2000 ;
        RECT 2310.3200 2778.1600 2311.9200 2778.6400 ;
        RECT 2265.3200 2794.4800 2266.9200 2794.9600 ;
        RECT 2265.3200 2799.9200 2266.9200 2800.4000 ;
        RECT 2253.5600 2799.9200 2256.5600 2800.4000 ;
        RECT 2253.5600 2794.4800 2256.5600 2794.9600 ;
        RECT 2253.5600 2805.3600 2256.5600 2805.8400 ;
        RECT 2265.3200 2805.3600 2266.9200 2805.8400 ;
        RECT 2265.3200 2783.6000 2266.9200 2784.0800 ;
        RECT 2265.3200 2789.0400 2266.9200 2789.5200 ;
        RECT 2253.5600 2789.0400 2256.5600 2789.5200 ;
        RECT 2253.5600 2783.6000 2256.5600 2784.0800 ;
        RECT 2265.3200 2767.2800 2266.9200 2767.7600 ;
        RECT 2265.3200 2772.7200 2266.9200 2773.2000 ;
        RECT 2253.5600 2772.7200 2256.5600 2773.2000 ;
        RECT 2253.5600 2767.2800 2256.5600 2767.7600 ;
        RECT 2253.5600 2778.1600 2256.5600 2778.6400 ;
        RECT 2265.3200 2778.1600 2266.9200 2778.6400 ;
        RECT 2355.3200 2750.9600 2356.9200 2751.4400 ;
        RECT 2355.3200 2756.4000 2356.9200 2756.8800 ;
        RECT 2355.3200 2761.8400 2356.9200 2762.3200 ;
        RECT 2355.3200 2740.0800 2356.9200 2740.5600 ;
        RECT 2355.3200 2745.5200 2356.9200 2746.0000 ;
        RECT 2310.3200 2750.9600 2311.9200 2751.4400 ;
        RECT 2310.3200 2756.4000 2311.9200 2756.8800 ;
        RECT 2310.3200 2761.8400 2311.9200 2762.3200 ;
        RECT 2310.3200 2740.0800 2311.9200 2740.5600 ;
        RECT 2310.3200 2745.5200 2311.9200 2746.0000 ;
        RECT 2355.3200 2723.7600 2356.9200 2724.2400 ;
        RECT 2355.3200 2729.2000 2356.9200 2729.6800 ;
        RECT 2355.3200 2734.6400 2356.9200 2735.1200 ;
        RECT 2355.3200 2712.8800 2356.9200 2713.3600 ;
        RECT 2355.3200 2718.3200 2356.9200 2718.8000 ;
        RECT 2310.3200 2723.7600 2311.9200 2724.2400 ;
        RECT 2310.3200 2729.2000 2311.9200 2729.6800 ;
        RECT 2310.3200 2734.6400 2311.9200 2735.1200 ;
        RECT 2310.3200 2712.8800 2311.9200 2713.3600 ;
        RECT 2310.3200 2718.3200 2311.9200 2718.8000 ;
        RECT 2265.3200 2750.9600 2266.9200 2751.4400 ;
        RECT 2265.3200 2756.4000 2266.9200 2756.8800 ;
        RECT 2265.3200 2761.8400 2266.9200 2762.3200 ;
        RECT 2253.5600 2750.9600 2256.5600 2751.4400 ;
        RECT 2253.5600 2756.4000 2256.5600 2756.8800 ;
        RECT 2253.5600 2761.8400 2256.5600 2762.3200 ;
        RECT 2265.3200 2740.0800 2266.9200 2740.5600 ;
        RECT 2265.3200 2745.5200 2266.9200 2746.0000 ;
        RECT 2253.5600 2740.0800 2256.5600 2740.5600 ;
        RECT 2253.5600 2745.5200 2256.5600 2746.0000 ;
        RECT 2265.3200 2723.7600 2266.9200 2724.2400 ;
        RECT 2265.3200 2729.2000 2266.9200 2729.6800 ;
        RECT 2265.3200 2734.6400 2266.9200 2735.1200 ;
        RECT 2253.5600 2723.7600 2256.5600 2724.2400 ;
        RECT 2253.5600 2729.2000 2256.5600 2729.6800 ;
        RECT 2253.5600 2734.6400 2256.5600 2735.1200 ;
        RECT 2265.3200 2712.8800 2266.9200 2713.3600 ;
        RECT 2265.3200 2718.3200 2266.9200 2718.8000 ;
        RECT 2253.5600 2712.8800 2256.5600 2713.3600 ;
        RECT 2253.5600 2718.3200 2256.5600 2718.8000 ;
        RECT 2457.6600 2696.5600 2460.6600 2697.0400 ;
        RECT 2457.6600 2702.0000 2460.6600 2702.4800 ;
        RECT 2457.6600 2707.4400 2460.6600 2707.9200 ;
        RECT 2445.3200 2696.5600 2446.9200 2697.0400 ;
        RECT 2445.3200 2702.0000 2446.9200 2702.4800 ;
        RECT 2445.3200 2707.4400 2446.9200 2707.9200 ;
        RECT 2457.6600 2685.6800 2460.6600 2686.1600 ;
        RECT 2457.6600 2691.1200 2460.6600 2691.6000 ;
        RECT 2445.3200 2685.6800 2446.9200 2686.1600 ;
        RECT 2445.3200 2691.1200 2446.9200 2691.6000 ;
        RECT 2457.6600 2669.3600 2460.6600 2669.8400 ;
        RECT 2457.6600 2674.8000 2460.6600 2675.2800 ;
        RECT 2457.6600 2680.2400 2460.6600 2680.7200 ;
        RECT 2445.3200 2669.3600 2446.9200 2669.8400 ;
        RECT 2445.3200 2674.8000 2446.9200 2675.2800 ;
        RECT 2445.3200 2680.2400 2446.9200 2680.7200 ;
        RECT 2457.6600 2658.4800 2460.6600 2658.9600 ;
        RECT 2457.6600 2663.9200 2460.6600 2664.4000 ;
        RECT 2445.3200 2658.4800 2446.9200 2658.9600 ;
        RECT 2445.3200 2663.9200 2446.9200 2664.4000 ;
        RECT 2400.3200 2696.5600 2401.9200 2697.0400 ;
        RECT 2400.3200 2702.0000 2401.9200 2702.4800 ;
        RECT 2400.3200 2707.4400 2401.9200 2707.9200 ;
        RECT 2400.3200 2685.6800 2401.9200 2686.1600 ;
        RECT 2400.3200 2691.1200 2401.9200 2691.6000 ;
        RECT 2400.3200 2669.3600 2401.9200 2669.8400 ;
        RECT 2400.3200 2674.8000 2401.9200 2675.2800 ;
        RECT 2400.3200 2680.2400 2401.9200 2680.7200 ;
        RECT 2400.3200 2658.4800 2401.9200 2658.9600 ;
        RECT 2400.3200 2663.9200 2401.9200 2664.4000 ;
        RECT 2457.6600 2642.1600 2460.6600 2642.6400 ;
        RECT 2457.6600 2647.6000 2460.6600 2648.0800 ;
        RECT 2457.6600 2653.0400 2460.6600 2653.5200 ;
        RECT 2445.3200 2642.1600 2446.9200 2642.6400 ;
        RECT 2445.3200 2647.6000 2446.9200 2648.0800 ;
        RECT 2445.3200 2653.0400 2446.9200 2653.5200 ;
        RECT 2457.6600 2631.2800 2460.6600 2631.7600 ;
        RECT 2457.6600 2636.7200 2460.6600 2637.2000 ;
        RECT 2445.3200 2631.2800 2446.9200 2631.7600 ;
        RECT 2445.3200 2636.7200 2446.9200 2637.2000 ;
        RECT 2457.6600 2614.9600 2460.6600 2615.4400 ;
        RECT 2457.6600 2620.4000 2460.6600 2620.8800 ;
        RECT 2457.6600 2625.8400 2460.6600 2626.3200 ;
        RECT 2445.3200 2614.9600 2446.9200 2615.4400 ;
        RECT 2445.3200 2620.4000 2446.9200 2620.8800 ;
        RECT 2445.3200 2625.8400 2446.9200 2626.3200 ;
        RECT 2457.6600 2609.5200 2460.6600 2610.0000 ;
        RECT 2445.3200 2609.5200 2446.9200 2610.0000 ;
        RECT 2400.3200 2642.1600 2401.9200 2642.6400 ;
        RECT 2400.3200 2647.6000 2401.9200 2648.0800 ;
        RECT 2400.3200 2653.0400 2401.9200 2653.5200 ;
        RECT 2400.3200 2631.2800 2401.9200 2631.7600 ;
        RECT 2400.3200 2636.7200 2401.9200 2637.2000 ;
        RECT 2400.3200 2614.9600 2401.9200 2615.4400 ;
        RECT 2400.3200 2620.4000 2401.9200 2620.8800 ;
        RECT 2400.3200 2625.8400 2401.9200 2626.3200 ;
        RECT 2400.3200 2609.5200 2401.9200 2610.0000 ;
        RECT 2355.3200 2696.5600 2356.9200 2697.0400 ;
        RECT 2355.3200 2702.0000 2356.9200 2702.4800 ;
        RECT 2355.3200 2707.4400 2356.9200 2707.9200 ;
        RECT 2355.3200 2685.6800 2356.9200 2686.1600 ;
        RECT 2355.3200 2691.1200 2356.9200 2691.6000 ;
        RECT 2310.3200 2696.5600 2311.9200 2697.0400 ;
        RECT 2310.3200 2702.0000 2311.9200 2702.4800 ;
        RECT 2310.3200 2707.4400 2311.9200 2707.9200 ;
        RECT 2310.3200 2685.6800 2311.9200 2686.1600 ;
        RECT 2310.3200 2691.1200 2311.9200 2691.6000 ;
        RECT 2355.3200 2669.3600 2356.9200 2669.8400 ;
        RECT 2355.3200 2674.8000 2356.9200 2675.2800 ;
        RECT 2355.3200 2680.2400 2356.9200 2680.7200 ;
        RECT 2355.3200 2658.4800 2356.9200 2658.9600 ;
        RECT 2355.3200 2663.9200 2356.9200 2664.4000 ;
        RECT 2310.3200 2669.3600 2311.9200 2669.8400 ;
        RECT 2310.3200 2674.8000 2311.9200 2675.2800 ;
        RECT 2310.3200 2680.2400 2311.9200 2680.7200 ;
        RECT 2310.3200 2658.4800 2311.9200 2658.9600 ;
        RECT 2310.3200 2663.9200 2311.9200 2664.4000 ;
        RECT 2265.3200 2696.5600 2266.9200 2697.0400 ;
        RECT 2265.3200 2702.0000 2266.9200 2702.4800 ;
        RECT 2265.3200 2707.4400 2266.9200 2707.9200 ;
        RECT 2253.5600 2696.5600 2256.5600 2697.0400 ;
        RECT 2253.5600 2702.0000 2256.5600 2702.4800 ;
        RECT 2253.5600 2707.4400 2256.5600 2707.9200 ;
        RECT 2265.3200 2685.6800 2266.9200 2686.1600 ;
        RECT 2265.3200 2691.1200 2266.9200 2691.6000 ;
        RECT 2253.5600 2685.6800 2256.5600 2686.1600 ;
        RECT 2253.5600 2691.1200 2256.5600 2691.6000 ;
        RECT 2265.3200 2669.3600 2266.9200 2669.8400 ;
        RECT 2265.3200 2674.8000 2266.9200 2675.2800 ;
        RECT 2265.3200 2680.2400 2266.9200 2680.7200 ;
        RECT 2253.5600 2669.3600 2256.5600 2669.8400 ;
        RECT 2253.5600 2674.8000 2256.5600 2675.2800 ;
        RECT 2253.5600 2680.2400 2256.5600 2680.7200 ;
        RECT 2265.3200 2658.4800 2266.9200 2658.9600 ;
        RECT 2265.3200 2663.9200 2266.9200 2664.4000 ;
        RECT 2253.5600 2658.4800 2256.5600 2658.9600 ;
        RECT 2253.5600 2663.9200 2256.5600 2664.4000 ;
        RECT 2355.3200 2642.1600 2356.9200 2642.6400 ;
        RECT 2355.3200 2647.6000 2356.9200 2648.0800 ;
        RECT 2355.3200 2653.0400 2356.9200 2653.5200 ;
        RECT 2355.3200 2631.2800 2356.9200 2631.7600 ;
        RECT 2355.3200 2636.7200 2356.9200 2637.2000 ;
        RECT 2310.3200 2642.1600 2311.9200 2642.6400 ;
        RECT 2310.3200 2647.6000 2311.9200 2648.0800 ;
        RECT 2310.3200 2653.0400 2311.9200 2653.5200 ;
        RECT 2310.3200 2631.2800 2311.9200 2631.7600 ;
        RECT 2310.3200 2636.7200 2311.9200 2637.2000 ;
        RECT 2355.3200 2614.9600 2356.9200 2615.4400 ;
        RECT 2355.3200 2620.4000 2356.9200 2620.8800 ;
        RECT 2355.3200 2625.8400 2356.9200 2626.3200 ;
        RECT 2355.3200 2609.5200 2356.9200 2610.0000 ;
        RECT 2310.3200 2614.9600 2311.9200 2615.4400 ;
        RECT 2310.3200 2620.4000 2311.9200 2620.8800 ;
        RECT 2310.3200 2625.8400 2311.9200 2626.3200 ;
        RECT 2310.3200 2609.5200 2311.9200 2610.0000 ;
        RECT 2265.3200 2642.1600 2266.9200 2642.6400 ;
        RECT 2265.3200 2647.6000 2266.9200 2648.0800 ;
        RECT 2265.3200 2653.0400 2266.9200 2653.5200 ;
        RECT 2253.5600 2642.1600 2256.5600 2642.6400 ;
        RECT 2253.5600 2647.6000 2256.5600 2648.0800 ;
        RECT 2253.5600 2653.0400 2256.5600 2653.5200 ;
        RECT 2265.3200 2631.2800 2266.9200 2631.7600 ;
        RECT 2265.3200 2636.7200 2266.9200 2637.2000 ;
        RECT 2253.5600 2631.2800 2256.5600 2631.7600 ;
        RECT 2253.5600 2636.7200 2256.5600 2637.2000 ;
        RECT 2265.3200 2614.9600 2266.9200 2615.4400 ;
        RECT 2265.3200 2620.4000 2266.9200 2620.8800 ;
        RECT 2265.3200 2625.8400 2266.9200 2626.3200 ;
        RECT 2253.5600 2614.9600 2256.5600 2615.4400 ;
        RECT 2253.5600 2620.4000 2256.5600 2620.8800 ;
        RECT 2253.5600 2625.8400 2256.5600 2626.3200 ;
        RECT 2253.5600 2609.5200 2256.5600 2610.0000 ;
        RECT 2265.3200 2609.5200 2266.9200 2610.0000 ;
        RECT 2253.5600 2814.4300 2460.6600 2817.4300 ;
        RECT 2253.5600 2601.3300 2460.6600 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 2371.6900 2446.9200 2587.7900 ;
        RECT 2400.3200 2371.6900 2401.9200 2587.7900 ;
        RECT 2355.3200 2371.6900 2356.9200 2587.7900 ;
        RECT 2310.3200 2371.6900 2311.9200 2587.7900 ;
        RECT 2265.3200 2371.6900 2266.9200 2587.7900 ;
        RECT 2457.6600 2371.6900 2460.6600 2587.7900 ;
        RECT 2253.5600 2371.6900 2256.5600 2587.7900 ;
      LAYER met3 ;
        RECT 2457.6600 2564.8400 2460.6600 2565.3200 ;
        RECT 2457.6600 2570.2800 2460.6600 2570.7600 ;
        RECT 2445.3200 2564.8400 2446.9200 2565.3200 ;
        RECT 2445.3200 2570.2800 2446.9200 2570.7600 ;
        RECT 2457.6600 2575.7200 2460.6600 2576.2000 ;
        RECT 2445.3200 2575.7200 2446.9200 2576.2000 ;
        RECT 2457.6600 2553.9600 2460.6600 2554.4400 ;
        RECT 2457.6600 2559.4000 2460.6600 2559.8800 ;
        RECT 2445.3200 2553.9600 2446.9200 2554.4400 ;
        RECT 2445.3200 2559.4000 2446.9200 2559.8800 ;
        RECT 2457.6600 2537.6400 2460.6600 2538.1200 ;
        RECT 2457.6600 2543.0800 2460.6600 2543.5600 ;
        RECT 2445.3200 2537.6400 2446.9200 2538.1200 ;
        RECT 2445.3200 2543.0800 2446.9200 2543.5600 ;
        RECT 2457.6600 2548.5200 2460.6600 2549.0000 ;
        RECT 2445.3200 2548.5200 2446.9200 2549.0000 ;
        RECT 2400.3200 2564.8400 2401.9200 2565.3200 ;
        RECT 2400.3200 2570.2800 2401.9200 2570.7600 ;
        RECT 2400.3200 2575.7200 2401.9200 2576.2000 ;
        RECT 2400.3200 2553.9600 2401.9200 2554.4400 ;
        RECT 2400.3200 2559.4000 2401.9200 2559.8800 ;
        RECT 2400.3200 2537.6400 2401.9200 2538.1200 ;
        RECT 2400.3200 2543.0800 2401.9200 2543.5600 ;
        RECT 2400.3200 2548.5200 2401.9200 2549.0000 ;
        RECT 2457.6600 2521.3200 2460.6600 2521.8000 ;
        RECT 2457.6600 2526.7600 2460.6600 2527.2400 ;
        RECT 2457.6600 2532.2000 2460.6600 2532.6800 ;
        RECT 2445.3200 2521.3200 2446.9200 2521.8000 ;
        RECT 2445.3200 2526.7600 2446.9200 2527.2400 ;
        RECT 2445.3200 2532.2000 2446.9200 2532.6800 ;
        RECT 2457.6600 2510.4400 2460.6600 2510.9200 ;
        RECT 2457.6600 2515.8800 2460.6600 2516.3600 ;
        RECT 2445.3200 2510.4400 2446.9200 2510.9200 ;
        RECT 2445.3200 2515.8800 2446.9200 2516.3600 ;
        RECT 2457.6600 2494.1200 2460.6600 2494.6000 ;
        RECT 2457.6600 2499.5600 2460.6600 2500.0400 ;
        RECT 2457.6600 2505.0000 2460.6600 2505.4800 ;
        RECT 2445.3200 2494.1200 2446.9200 2494.6000 ;
        RECT 2445.3200 2499.5600 2446.9200 2500.0400 ;
        RECT 2445.3200 2505.0000 2446.9200 2505.4800 ;
        RECT 2457.6600 2483.2400 2460.6600 2483.7200 ;
        RECT 2457.6600 2488.6800 2460.6600 2489.1600 ;
        RECT 2445.3200 2483.2400 2446.9200 2483.7200 ;
        RECT 2445.3200 2488.6800 2446.9200 2489.1600 ;
        RECT 2400.3200 2521.3200 2401.9200 2521.8000 ;
        RECT 2400.3200 2526.7600 2401.9200 2527.2400 ;
        RECT 2400.3200 2532.2000 2401.9200 2532.6800 ;
        RECT 2400.3200 2510.4400 2401.9200 2510.9200 ;
        RECT 2400.3200 2515.8800 2401.9200 2516.3600 ;
        RECT 2400.3200 2494.1200 2401.9200 2494.6000 ;
        RECT 2400.3200 2499.5600 2401.9200 2500.0400 ;
        RECT 2400.3200 2505.0000 2401.9200 2505.4800 ;
        RECT 2400.3200 2483.2400 2401.9200 2483.7200 ;
        RECT 2400.3200 2488.6800 2401.9200 2489.1600 ;
        RECT 2355.3200 2564.8400 2356.9200 2565.3200 ;
        RECT 2355.3200 2570.2800 2356.9200 2570.7600 ;
        RECT 2355.3200 2575.7200 2356.9200 2576.2000 ;
        RECT 2310.3200 2564.8400 2311.9200 2565.3200 ;
        RECT 2310.3200 2570.2800 2311.9200 2570.7600 ;
        RECT 2310.3200 2575.7200 2311.9200 2576.2000 ;
        RECT 2355.3200 2553.9600 2356.9200 2554.4400 ;
        RECT 2355.3200 2559.4000 2356.9200 2559.8800 ;
        RECT 2355.3200 2537.6400 2356.9200 2538.1200 ;
        RECT 2355.3200 2543.0800 2356.9200 2543.5600 ;
        RECT 2355.3200 2548.5200 2356.9200 2549.0000 ;
        RECT 2310.3200 2553.9600 2311.9200 2554.4400 ;
        RECT 2310.3200 2559.4000 2311.9200 2559.8800 ;
        RECT 2310.3200 2537.6400 2311.9200 2538.1200 ;
        RECT 2310.3200 2543.0800 2311.9200 2543.5600 ;
        RECT 2310.3200 2548.5200 2311.9200 2549.0000 ;
        RECT 2265.3200 2564.8400 2266.9200 2565.3200 ;
        RECT 2265.3200 2570.2800 2266.9200 2570.7600 ;
        RECT 2253.5600 2570.2800 2256.5600 2570.7600 ;
        RECT 2253.5600 2564.8400 2256.5600 2565.3200 ;
        RECT 2253.5600 2575.7200 2256.5600 2576.2000 ;
        RECT 2265.3200 2575.7200 2266.9200 2576.2000 ;
        RECT 2265.3200 2553.9600 2266.9200 2554.4400 ;
        RECT 2265.3200 2559.4000 2266.9200 2559.8800 ;
        RECT 2253.5600 2559.4000 2256.5600 2559.8800 ;
        RECT 2253.5600 2553.9600 2256.5600 2554.4400 ;
        RECT 2265.3200 2537.6400 2266.9200 2538.1200 ;
        RECT 2265.3200 2543.0800 2266.9200 2543.5600 ;
        RECT 2253.5600 2543.0800 2256.5600 2543.5600 ;
        RECT 2253.5600 2537.6400 2256.5600 2538.1200 ;
        RECT 2253.5600 2548.5200 2256.5600 2549.0000 ;
        RECT 2265.3200 2548.5200 2266.9200 2549.0000 ;
        RECT 2355.3200 2521.3200 2356.9200 2521.8000 ;
        RECT 2355.3200 2526.7600 2356.9200 2527.2400 ;
        RECT 2355.3200 2532.2000 2356.9200 2532.6800 ;
        RECT 2355.3200 2510.4400 2356.9200 2510.9200 ;
        RECT 2355.3200 2515.8800 2356.9200 2516.3600 ;
        RECT 2310.3200 2521.3200 2311.9200 2521.8000 ;
        RECT 2310.3200 2526.7600 2311.9200 2527.2400 ;
        RECT 2310.3200 2532.2000 2311.9200 2532.6800 ;
        RECT 2310.3200 2510.4400 2311.9200 2510.9200 ;
        RECT 2310.3200 2515.8800 2311.9200 2516.3600 ;
        RECT 2355.3200 2494.1200 2356.9200 2494.6000 ;
        RECT 2355.3200 2499.5600 2356.9200 2500.0400 ;
        RECT 2355.3200 2505.0000 2356.9200 2505.4800 ;
        RECT 2355.3200 2483.2400 2356.9200 2483.7200 ;
        RECT 2355.3200 2488.6800 2356.9200 2489.1600 ;
        RECT 2310.3200 2494.1200 2311.9200 2494.6000 ;
        RECT 2310.3200 2499.5600 2311.9200 2500.0400 ;
        RECT 2310.3200 2505.0000 2311.9200 2505.4800 ;
        RECT 2310.3200 2483.2400 2311.9200 2483.7200 ;
        RECT 2310.3200 2488.6800 2311.9200 2489.1600 ;
        RECT 2265.3200 2521.3200 2266.9200 2521.8000 ;
        RECT 2265.3200 2526.7600 2266.9200 2527.2400 ;
        RECT 2265.3200 2532.2000 2266.9200 2532.6800 ;
        RECT 2253.5600 2521.3200 2256.5600 2521.8000 ;
        RECT 2253.5600 2526.7600 2256.5600 2527.2400 ;
        RECT 2253.5600 2532.2000 2256.5600 2532.6800 ;
        RECT 2265.3200 2510.4400 2266.9200 2510.9200 ;
        RECT 2265.3200 2515.8800 2266.9200 2516.3600 ;
        RECT 2253.5600 2510.4400 2256.5600 2510.9200 ;
        RECT 2253.5600 2515.8800 2256.5600 2516.3600 ;
        RECT 2265.3200 2494.1200 2266.9200 2494.6000 ;
        RECT 2265.3200 2499.5600 2266.9200 2500.0400 ;
        RECT 2265.3200 2505.0000 2266.9200 2505.4800 ;
        RECT 2253.5600 2494.1200 2256.5600 2494.6000 ;
        RECT 2253.5600 2499.5600 2256.5600 2500.0400 ;
        RECT 2253.5600 2505.0000 2256.5600 2505.4800 ;
        RECT 2265.3200 2483.2400 2266.9200 2483.7200 ;
        RECT 2265.3200 2488.6800 2266.9200 2489.1600 ;
        RECT 2253.5600 2483.2400 2256.5600 2483.7200 ;
        RECT 2253.5600 2488.6800 2256.5600 2489.1600 ;
        RECT 2457.6600 2466.9200 2460.6600 2467.4000 ;
        RECT 2457.6600 2472.3600 2460.6600 2472.8400 ;
        RECT 2457.6600 2477.8000 2460.6600 2478.2800 ;
        RECT 2445.3200 2466.9200 2446.9200 2467.4000 ;
        RECT 2445.3200 2472.3600 2446.9200 2472.8400 ;
        RECT 2445.3200 2477.8000 2446.9200 2478.2800 ;
        RECT 2457.6600 2456.0400 2460.6600 2456.5200 ;
        RECT 2457.6600 2461.4800 2460.6600 2461.9600 ;
        RECT 2445.3200 2456.0400 2446.9200 2456.5200 ;
        RECT 2445.3200 2461.4800 2446.9200 2461.9600 ;
        RECT 2457.6600 2439.7200 2460.6600 2440.2000 ;
        RECT 2457.6600 2445.1600 2460.6600 2445.6400 ;
        RECT 2457.6600 2450.6000 2460.6600 2451.0800 ;
        RECT 2445.3200 2439.7200 2446.9200 2440.2000 ;
        RECT 2445.3200 2445.1600 2446.9200 2445.6400 ;
        RECT 2445.3200 2450.6000 2446.9200 2451.0800 ;
        RECT 2457.6600 2428.8400 2460.6600 2429.3200 ;
        RECT 2457.6600 2434.2800 2460.6600 2434.7600 ;
        RECT 2445.3200 2428.8400 2446.9200 2429.3200 ;
        RECT 2445.3200 2434.2800 2446.9200 2434.7600 ;
        RECT 2400.3200 2466.9200 2401.9200 2467.4000 ;
        RECT 2400.3200 2472.3600 2401.9200 2472.8400 ;
        RECT 2400.3200 2477.8000 2401.9200 2478.2800 ;
        RECT 2400.3200 2456.0400 2401.9200 2456.5200 ;
        RECT 2400.3200 2461.4800 2401.9200 2461.9600 ;
        RECT 2400.3200 2439.7200 2401.9200 2440.2000 ;
        RECT 2400.3200 2445.1600 2401.9200 2445.6400 ;
        RECT 2400.3200 2450.6000 2401.9200 2451.0800 ;
        RECT 2400.3200 2428.8400 2401.9200 2429.3200 ;
        RECT 2400.3200 2434.2800 2401.9200 2434.7600 ;
        RECT 2457.6600 2412.5200 2460.6600 2413.0000 ;
        RECT 2457.6600 2417.9600 2460.6600 2418.4400 ;
        RECT 2457.6600 2423.4000 2460.6600 2423.8800 ;
        RECT 2445.3200 2412.5200 2446.9200 2413.0000 ;
        RECT 2445.3200 2417.9600 2446.9200 2418.4400 ;
        RECT 2445.3200 2423.4000 2446.9200 2423.8800 ;
        RECT 2457.6600 2401.6400 2460.6600 2402.1200 ;
        RECT 2457.6600 2407.0800 2460.6600 2407.5600 ;
        RECT 2445.3200 2401.6400 2446.9200 2402.1200 ;
        RECT 2445.3200 2407.0800 2446.9200 2407.5600 ;
        RECT 2457.6600 2385.3200 2460.6600 2385.8000 ;
        RECT 2457.6600 2390.7600 2460.6600 2391.2400 ;
        RECT 2457.6600 2396.2000 2460.6600 2396.6800 ;
        RECT 2445.3200 2385.3200 2446.9200 2385.8000 ;
        RECT 2445.3200 2390.7600 2446.9200 2391.2400 ;
        RECT 2445.3200 2396.2000 2446.9200 2396.6800 ;
        RECT 2457.6600 2379.8800 2460.6600 2380.3600 ;
        RECT 2445.3200 2379.8800 2446.9200 2380.3600 ;
        RECT 2400.3200 2412.5200 2401.9200 2413.0000 ;
        RECT 2400.3200 2417.9600 2401.9200 2418.4400 ;
        RECT 2400.3200 2423.4000 2401.9200 2423.8800 ;
        RECT 2400.3200 2401.6400 2401.9200 2402.1200 ;
        RECT 2400.3200 2407.0800 2401.9200 2407.5600 ;
        RECT 2400.3200 2385.3200 2401.9200 2385.8000 ;
        RECT 2400.3200 2390.7600 2401.9200 2391.2400 ;
        RECT 2400.3200 2396.2000 2401.9200 2396.6800 ;
        RECT 2400.3200 2379.8800 2401.9200 2380.3600 ;
        RECT 2355.3200 2466.9200 2356.9200 2467.4000 ;
        RECT 2355.3200 2472.3600 2356.9200 2472.8400 ;
        RECT 2355.3200 2477.8000 2356.9200 2478.2800 ;
        RECT 2355.3200 2456.0400 2356.9200 2456.5200 ;
        RECT 2355.3200 2461.4800 2356.9200 2461.9600 ;
        RECT 2310.3200 2466.9200 2311.9200 2467.4000 ;
        RECT 2310.3200 2472.3600 2311.9200 2472.8400 ;
        RECT 2310.3200 2477.8000 2311.9200 2478.2800 ;
        RECT 2310.3200 2456.0400 2311.9200 2456.5200 ;
        RECT 2310.3200 2461.4800 2311.9200 2461.9600 ;
        RECT 2355.3200 2439.7200 2356.9200 2440.2000 ;
        RECT 2355.3200 2445.1600 2356.9200 2445.6400 ;
        RECT 2355.3200 2450.6000 2356.9200 2451.0800 ;
        RECT 2355.3200 2428.8400 2356.9200 2429.3200 ;
        RECT 2355.3200 2434.2800 2356.9200 2434.7600 ;
        RECT 2310.3200 2439.7200 2311.9200 2440.2000 ;
        RECT 2310.3200 2445.1600 2311.9200 2445.6400 ;
        RECT 2310.3200 2450.6000 2311.9200 2451.0800 ;
        RECT 2310.3200 2428.8400 2311.9200 2429.3200 ;
        RECT 2310.3200 2434.2800 2311.9200 2434.7600 ;
        RECT 2265.3200 2466.9200 2266.9200 2467.4000 ;
        RECT 2265.3200 2472.3600 2266.9200 2472.8400 ;
        RECT 2265.3200 2477.8000 2266.9200 2478.2800 ;
        RECT 2253.5600 2466.9200 2256.5600 2467.4000 ;
        RECT 2253.5600 2472.3600 2256.5600 2472.8400 ;
        RECT 2253.5600 2477.8000 2256.5600 2478.2800 ;
        RECT 2265.3200 2456.0400 2266.9200 2456.5200 ;
        RECT 2265.3200 2461.4800 2266.9200 2461.9600 ;
        RECT 2253.5600 2456.0400 2256.5600 2456.5200 ;
        RECT 2253.5600 2461.4800 2256.5600 2461.9600 ;
        RECT 2265.3200 2439.7200 2266.9200 2440.2000 ;
        RECT 2265.3200 2445.1600 2266.9200 2445.6400 ;
        RECT 2265.3200 2450.6000 2266.9200 2451.0800 ;
        RECT 2253.5600 2439.7200 2256.5600 2440.2000 ;
        RECT 2253.5600 2445.1600 2256.5600 2445.6400 ;
        RECT 2253.5600 2450.6000 2256.5600 2451.0800 ;
        RECT 2265.3200 2428.8400 2266.9200 2429.3200 ;
        RECT 2265.3200 2434.2800 2266.9200 2434.7600 ;
        RECT 2253.5600 2428.8400 2256.5600 2429.3200 ;
        RECT 2253.5600 2434.2800 2256.5600 2434.7600 ;
        RECT 2355.3200 2412.5200 2356.9200 2413.0000 ;
        RECT 2355.3200 2417.9600 2356.9200 2418.4400 ;
        RECT 2355.3200 2423.4000 2356.9200 2423.8800 ;
        RECT 2355.3200 2401.6400 2356.9200 2402.1200 ;
        RECT 2355.3200 2407.0800 2356.9200 2407.5600 ;
        RECT 2310.3200 2412.5200 2311.9200 2413.0000 ;
        RECT 2310.3200 2417.9600 2311.9200 2418.4400 ;
        RECT 2310.3200 2423.4000 2311.9200 2423.8800 ;
        RECT 2310.3200 2401.6400 2311.9200 2402.1200 ;
        RECT 2310.3200 2407.0800 2311.9200 2407.5600 ;
        RECT 2355.3200 2385.3200 2356.9200 2385.8000 ;
        RECT 2355.3200 2390.7600 2356.9200 2391.2400 ;
        RECT 2355.3200 2396.2000 2356.9200 2396.6800 ;
        RECT 2355.3200 2379.8800 2356.9200 2380.3600 ;
        RECT 2310.3200 2385.3200 2311.9200 2385.8000 ;
        RECT 2310.3200 2390.7600 2311.9200 2391.2400 ;
        RECT 2310.3200 2396.2000 2311.9200 2396.6800 ;
        RECT 2310.3200 2379.8800 2311.9200 2380.3600 ;
        RECT 2265.3200 2412.5200 2266.9200 2413.0000 ;
        RECT 2265.3200 2417.9600 2266.9200 2418.4400 ;
        RECT 2265.3200 2423.4000 2266.9200 2423.8800 ;
        RECT 2253.5600 2412.5200 2256.5600 2413.0000 ;
        RECT 2253.5600 2417.9600 2256.5600 2418.4400 ;
        RECT 2253.5600 2423.4000 2256.5600 2423.8800 ;
        RECT 2265.3200 2401.6400 2266.9200 2402.1200 ;
        RECT 2265.3200 2407.0800 2266.9200 2407.5600 ;
        RECT 2253.5600 2401.6400 2256.5600 2402.1200 ;
        RECT 2253.5600 2407.0800 2256.5600 2407.5600 ;
        RECT 2265.3200 2385.3200 2266.9200 2385.8000 ;
        RECT 2265.3200 2390.7600 2266.9200 2391.2400 ;
        RECT 2265.3200 2396.2000 2266.9200 2396.6800 ;
        RECT 2253.5600 2385.3200 2256.5600 2385.8000 ;
        RECT 2253.5600 2390.7600 2256.5600 2391.2400 ;
        RECT 2253.5600 2396.2000 2256.5600 2396.6800 ;
        RECT 2253.5600 2379.8800 2256.5600 2380.3600 ;
        RECT 2265.3200 2379.8800 2266.9200 2380.3600 ;
        RECT 2253.5600 2584.7900 2460.6600 2587.7900 ;
        RECT 2253.5600 2371.6900 2460.6600 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 2142.0500 2446.9200 2358.1500 ;
        RECT 2400.3200 2142.0500 2401.9200 2358.1500 ;
        RECT 2355.3200 2142.0500 2356.9200 2358.1500 ;
        RECT 2310.3200 2142.0500 2311.9200 2358.1500 ;
        RECT 2265.3200 2142.0500 2266.9200 2358.1500 ;
        RECT 2457.6600 2142.0500 2460.6600 2358.1500 ;
        RECT 2253.5600 2142.0500 2256.5600 2358.1500 ;
      LAYER met3 ;
        RECT 2457.6600 2335.2000 2460.6600 2335.6800 ;
        RECT 2457.6600 2340.6400 2460.6600 2341.1200 ;
        RECT 2445.3200 2335.2000 2446.9200 2335.6800 ;
        RECT 2445.3200 2340.6400 2446.9200 2341.1200 ;
        RECT 2457.6600 2346.0800 2460.6600 2346.5600 ;
        RECT 2445.3200 2346.0800 2446.9200 2346.5600 ;
        RECT 2457.6600 2324.3200 2460.6600 2324.8000 ;
        RECT 2457.6600 2329.7600 2460.6600 2330.2400 ;
        RECT 2445.3200 2324.3200 2446.9200 2324.8000 ;
        RECT 2445.3200 2329.7600 2446.9200 2330.2400 ;
        RECT 2457.6600 2308.0000 2460.6600 2308.4800 ;
        RECT 2457.6600 2313.4400 2460.6600 2313.9200 ;
        RECT 2445.3200 2308.0000 2446.9200 2308.4800 ;
        RECT 2445.3200 2313.4400 2446.9200 2313.9200 ;
        RECT 2457.6600 2318.8800 2460.6600 2319.3600 ;
        RECT 2445.3200 2318.8800 2446.9200 2319.3600 ;
        RECT 2400.3200 2335.2000 2401.9200 2335.6800 ;
        RECT 2400.3200 2340.6400 2401.9200 2341.1200 ;
        RECT 2400.3200 2346.0800 2401.9200 2346.5600 ;
        RECT 2400.3200 2324.3200 2401.9200 2324.8000 ;
        RECT 2400.3200 2329.7600 2401.9200 2330.2400 ;
        RECT 2400.3200 2308.0000 2401.9200 2308.4800 ;
        RECT 2400.3200 2313.4400 2401.9200 2313.9200 ;
        RECT 2400.3200 2318.8800 2401.9200 2319.3600 ;
        RECT 2457.6600 2291.6800 2460.6600 2292.1600 ;
        RECT 2457.6600 2297.1200 2460.6600 2297.6000 ;
        RECT 2457.6600 2302.5600 2460.6600 2303.0400 ;
        RECT 2445.3200 2291.6800 2446.9200 2292.1600 ;
        RECT 2445.3200 2297.1200 2446.9200 2297.6000 ;
        RECT 2445.3200 2302.5600 2446.9200 2303.0400 ;
        RECT 2457.6600 2280.8000 2460.6600 2281.2800 ;
        RECT 2457.6600 2286.2400 2460.6600 2286.7200 ;
        RECT 2445.3200 2280.8000 2446.9200 2281.2800 ;
        RECT 2445.3200 2286.2400 2446.9200 2286.7200 ;
        RECT 2457.6600 2264.4800 2460.6600 2264.9600 ;
        RECT 2457.6600 2269.9200 2460.6600 2270.4000 ;
        RECT 2457.6600 2275.3600 2460.6600 2275.8400 ;
        RECT 2445.3200 2264.4800 2446.9200 2264.9600 ;
        RECT 2445.3200 2269.9200 2446.9200 2270.4000 ;
        RECT 2445.3200 2275.3600 2446.9200 2275.8400 ;
        RECT 2457.6600 2253.6000 2460.6600 2254.0800 ;
        RECT 2457.6600 2259.0400 2460.6600 2259.5200 ;
        RECT 2445.3200 2253.6000 2446.9200 2254.0800 ;
        RECT 2445.3200 2259.0400 2446.9200 2259.5200 ;
        RECT 2400.3200 2291.6800 2401.9200 2292.1600 ;
        RECT 2400.3200 2297.1200 2401.9200 2297.6000 ;
        RECT 2400.3200 2302.5600 2401.9200 2303.0400 ;
        RECT 2400.3200 2280.8000 2401.9200 2281.2800 ;
        RECT 2400.3200 2286.2400 2401.9200 2286.7200 ;
        RECT 2400.3200 2264.4800 2401.9200 2264.9600 ;
        RECT 2400.3200 2269.9200 2401.9200 2270.4000 ;
        RECT 2400.3200 2275.3600 2401.9200 2275.8400 ;
        RECT 2400.3200 2253.6000 2401.9200 2254.0800 ;
        RECT 2400.3200 2259.0400 2401.9200 2259.5200 ;
        RECT 2355.3200 2335.2000 2356.9200 2335.6800 ;
        RECT 2355.3200 2340.6400 2356.9200 2341.1200 ;
        RECT 2355.3200 2346.0800 2356.9200 2346.5600 ;
        RECT 2310.3200 2335.2000 2311.9200 2335.6800 ;
        RECT 2310.3200 2340.6400 2311.9200 2341.1200 ;
        RECT 2310.3200 2346.0800 2311.9200 2346.5600 ;
        RECT 2355.3200 2324.3200 2356.9200 2324.8000 ;
        RECT 2355.3200 2329.7600 2356.9200 2330.2400 ;
        RECT 2355.3200 2308.0000 2356.9200 2308.4800 ;
        RECT 2355.3200 2313.4400 2356.9200 2313.9200 ;
        RECT 2355.3200 2318.8800 2356.9200 2319.3600 ;
        RECT 2310.3200 2324.3200 2311.9200 2324.8000 ;
        RECT 2310.3200 2329.7600 2311.9200 2330.2400 ;
        RECT 2310.3200 2308.0000 2311.9200 2308.4800 ;
        RECT 2310.3200 2313.4400 2311.9200 2313.9200 ;
        RECT 2310.3200 2318.8800 2311.9200 2319.3600 ;
        RECT 2265.3200 2335.2000 2266.9200 2335.6800 ;
        RECT 2265.3200 2340.6400 2266.9200 2341.1200 ;
        RECT 2253.5600 2340.6400 2256.5600 2341.1200 ;
        RECT 2253.5600 2335.2000 2256.5600 2335.6800 ;
        RECT 2253.5600 2346.0800 2256.5600 2346.5600 ;
        RECT 2265.3200 2346.0800 2266.9200 2346.5600 ;
        RECT 2265.3200 2324.3200 2266.9200 2324.8000 ;
        RECT 2265.3200 2329.7600 2266.9200 2330.2400 ;
        RECT 2253.5600 2329.7600 2256.5600 2330.2400 ;
        RECT 2253.5600 2324.3200 2256.5600 2324.8000 ;
        RECT 2265.3200 2308.0000 2266.9200 2308.4800 ;
        RECT 2265.3200 2313.4400 2266.9200 2313.9200 ;
        RECT 2253.5600 2313.4400 2256.5600 2313.9200 ;
        RECT 2253.5600 2308.0000 2256.5600 2308.4800 ;
        RECT 2253.5600 2318.8800 2256.5600 2319.3600 ;
        RECT 2265.3200 2318.8800 2266.9200 2319.3600 ;
        RECT 2355.3200 2291.6800 2356.9200 2292.1600 ;
        RECT 2355.3200 2297.1200 2356.9200 2297.6000 ;
        RECT 2355.3200 2302.5600 2356.9200 2303.0400 ;
        RECT 2355.3200 2280.8000 2356.9200 2281.2800 ;
        RECT 2355.3200 2286.2400 2356.9200 2286.7200 ;
        RECT 2310.3200 2291.6800 2311.9200 2292.1600 ;
        RECT 2310.3200 2297.1200 2311.9200 2297.6000 ;
        RECT 2310.3200 2302.5600 2311.9200 2303.0400 ;
        RECT 2310.3200 2280.8000 2311.9200 2281.2800 ;
        RECT 2310.3200 2286.2400 2311.9200 2286.7200 ;
        RECT 2355.3200 2264.4800 2356.9200 2264.9600 ;
        RECT 2355.3200 2269.9200 2356.9200 2270.4000 ;
        RECT 2355.3200 2275.3600 2356.9200 2275.8400 ;
        RECT 2355.3200 2253.6000 2356.9200 2254.0800 ;
        RECT 2355.3200 2259.0400 2356.9200 2259.5200 ;
        RECT 2310.3200 2264.4800 2311.9200 2264.9600 ;
        RECT 2310.3200 2269.9200 2311.9200 2270.4000 ;
        RECT 2310.3200 2275.3600 2311.9200 2275.8400 ;
        RECT 2310.3200 2253.6000 2311.9200 2254.0800 ;
        RECT 2310.3200 2259.0400 2311.9200 2259.5200 ;
        RECT 2265.3200 2291.6800 2266.9200 2292.1600 ;
        RECT 2265.3200 2297.1200 2266.9200 2297.6000 ;
        RECT 2265.3200 2302.5600 2266.9200 2303.0400 ;
        RECT 2253.5600 2291.6800 2256.5600 2292.1600 ;
        RECT 2253.5600 2297.1200 2256.5600 2297.6000 ;
        RECT 2253.5600 2302.5600 2256.5600 2303.0400 ;
        RECT 2265.3200 2280.8000 2266.9200 2281.2800 ;
        RECT 2265.3200 2286.2400 2266.9200 2286.7200 ;
        RECT 2253.5600 2280.8000 2256.5600 2281.2800 ;
        RECT 2253.5600 2286.2400 2256.5600 2286.7200 ;
        RECT 2265.3200 2264.4800 2266.9200 2264.9600 ;
        RECT 2265.3200 2269.9200 2266.9200 2270.4000 ;
        RECT 2265.3200 2275.3600 2266.9200 2275.8400 ;
        RECT 2253.5600 2264.4800 2256.5600 2264.9600 ;
        RECT 2253.5600 2269.9200 2256.5600 2270.4000 ;
        RECT 2253.5600 2275.3600 2256.5600 2275.8400 ;
        RECT 2265.3200 2253.6000 2266.9200 2254.0800 ;
        RECT 2265.3200 2259.0400 2266.9200 2259.5200 ;
        RECT 2253.5600 2253.6000 2256.5600 2254.0800 ;
        RECT 2253.5600 2259.0400 2256.5600 2259.5200 ;
        RECT 2457.6600 2237.2800 2460.6600 2237.7600 ;
        RECT 2457.6600 2242.7200 2460.6600 2243.2000 ;
        RECT 2457.6600 2248.1600 2460.6600 2248.6400 ;
        RECT 2445.3200 2237.2800 2446.9200 2237.7600 ;
        RECT 2445.3200 2242.7200 2446.9200 2243.2000 ;
        RECT 2445.3200 2248.1600 2446.9200 2248.6400 ;
        RECT 2457.6600 2226.4000 2460.6600 2226.8800 ;
        RECT 2457.6600 2231.8400 2460.6600 2232.3200 ;
        RECT 2445.3200 2226.4000 2446.9200 2226.8800 ;
        RECT 2445.3200 2231.8400 2446.9200 2232.3200 ;
        RECT 2457.6600 2210.0800 2460.6600 2210.5600 ;
        RECT 2457.6600 2215.5200 2460.6600 2216.0000 ;
        RECT 2457.6600 2220.9600 2460.6600 2221.4400 ;
        RECT 2445.3200 2210.0800 2446.9200 2210.5600 ;
        RECT 2445.3200 2215.5200 2446.9200 2216.0000 ;
        RECT 2445.3200 2220.9600 2446.9200 2221.4400 ;
        RECT 2457.6600 2199.2000 2460.6600 2199.6800 ;
        RECT 2457.6600 2204.6400 2460.6600 2205.1200 ;
        RECT 2445.3200 2199.2000 2446.9200 2199.6800 ;
        RECT 2445.3200 2204.6400 2446.9200 2205.1200 ;
        RECT 2400.3200 2237.2800 2401.9200 2237.7600 ;
        RECT 2400.3200 2242.7200 2401.9200 2243.2000 ;
        RECT 2400.3200 2248.1600 2401.9200 2248.6400 ;
        RECT 2400.3200 2226.4000 2401.9200 2226.8800 ;
        RECT 2400.3200 2231.8400 2401.9200 2232.3200 ;
        RECT 2400.3200 2210.0800 2401.9200 2210.5600 ;
        RECT 2400.3200 2215.5200 2401.9200 2216.0000 ;
        RECT 2400.3200 2220.9600 2401.9200 2221.4400 ;
        RECT 2400.3200 2199.2000 2401.9200 2199.6800 ;
        RECT 2400.3200 2204.6400 2401.9200 2205.1200 ;
        RECT 2457.6600 2182.8800 2460.6600 2183.3600 ;
        RECT 2457.6600 2188.3200 2460.6600 2188.8000 ;
        RECT 2457.6600 2193.7600 2460.6600 2194.2400 ;
        RECT 2445.3200 2182.8800 2446.9200 2183.3600 ;
        RECT 2445.3200 2188.3200 2446.9200 2188.8000 ;
        RECT 2445.3200 2193.7600 2446.9200 2194.2400 ;
        RECT 2457.6600 2172.0000 2460.6600 2172.4800 ;
        RECT 2457.6600 2177.4400 2460.6600 2177.9200 ;
        RECT 2445.3200 2172.0000 2446.9200 2172.4800 ;
        RECT 2445.3200 2177.4400 2446.9200 2177.9200 ;
        RECT 2457.6600 2155.6800 2460.6600 2156.1600 ;
        RECT 2457.6600 2161.1200 2460.6600 2161.6000 ;
        RECT 2457.6600 2166.5600 2460.6600 2167.0400 ;
        RECT 2445.3200 2155.6800 2446.9200 2156.1600 ;
        RECT 2445.3200 2161.1200 2446.9200 2161.6000 ;
        RECT 2445.3200 2166.5600 2446.9200 2167.0400 ;
        RECT 2457.6600 2150.2400 2460.6600 2150.7200 ;
        RECT 2445.3200 2150.2400 2446.9200 2150.7200 ;
        RECT 2400.3200 2182.8800 2401.9200 2183.3600 ;
        RECT 2400.3200 2188.3200 2401.9200 2188.8000 ;
        RECT 2400.3200 2193.7600 2401.9200 2194.2400 ;
        RECT 2400.3200 2172.0000 2401.9200 2172.4800 ;
        RECT 2400.3200 2177.4400 2401.9200 2177.9200 ;
        RECT 2400.3200 2155.6800 2401.9200 2156.1600 ;
        RECT 2400.3200 2161.1200 2401.9200 2161.6000 ;
        RECT 2400.3200 2166.5600 2401.9200 2167.0400 ;
        RECT 2400.3200 2150.2400 2401.9200 2150.7200 ;
        RECT 2355.3200 2237.2800 2356.9200 2237.7600 ;
        RECT 2355.3200 2242.7200 2356.9200 2243.2000 ;
        RECT 2355.3200 2248.1600 2356.9200 2248.6400 ;
        RECT 2355.3200 2226.4000 2356.9200 2226.8800 ;
        RECT 2355.3200 2231.8400 2356.9200 2232.3200 ;
        RECT 2310.3200 2237.2800 2311.9200 2237.7600 ;
        RECT 2310.3200 2242.7200 2311.9200 2243.2000 ;
        RECT 2310.3200 2248.1600 2311.9200 2248.6400 ;
        RECT 2310.3200 2226.4000 2311.9200 2226.8800 ;
        RECT 2310.3200 2231.8400 2311.9200 2232.3200 ;
        RECT 2355.3200 2210.0800 2356.9200 2210.5600 ;
        RECT 2355.3200 2215.5200 2356.9200 2216.0000 ;
        RECT 2355.3200 2220.9600 2356.9200 2221.4400 ;
        RECT 2355.3200 2199.2000 2356.9200 2199.6800 ;
        RECT 2355.3200 2204.6400 2356.9200 2205.1200 ;
        RECT 2310.3200 2210.0800 2311.9200 2210.5600 ;
        RECT 2310.3200 2215.5200 2311.9200 2216.0000 ;
        RECT 2310.3200 2220.9600 2311.9200 2221.4400 ;
        RECT 2310.3200 2199.2000 2311.9200 2199.6800 ;
        RECT 2310.3200 2204.6400 2311.9200 2205.1200 ;
        RECT 2265.3200 2237.2800 2266.9200 2237.7600 ;
        RECT 2265.3200 2242.7200 2266.9200 2243.2000 ;
        RECT 2265.3200 2248.1600 2266.9200 2248.6400 ;
        RECT 2253.5600 2237.2800 2256.5600 2237.7600 ;
        RECT 2253.5600 2242.7200 2256.5600 2243.2000 ;
        RECT 2253.5600 2248.1600 2256.5600 2248.6400 ;
        RECT 2265.3200 2226.4000 2266.9200 2226.8800 ;
        RECT 2265.3200 2231.8400 2266.9200 2232.3200 ;
        RECT 2253.5600 2226.4000 2256.5600 2226.8800 ;
        RECT 2253.5600 2231.8400 2256.5600 2232.3200 ;
        RECT 2265.3200 2210.0800 2266.9200 2210.5600 ;
        RECT 2265.3200 2215.5200 2266.9200 2216.0000 ;
        RECT 2265.3200 2220.9600 2266.9200 2221.4400 ;
        RECT 2253.5600 2210.0800 2256.5600 2210.5600 ;
        RECT 2253.5600 2215.5200 2256.5600 2216.0000 ;
        RECT 2253.5600 2220.9600 2256.5600 2221.4400 ;
        RECT 2265.3200 2199.2000 2266.9200 2199.6800 ;
        RECT 2265.3200 2204.6400 2266.9200 2205.1200 ;
        RECT 2253.5600 2199.2000 2256.5600 2199.6800 ;
        RECT 2253.5600 2204.6400 2256.5600 2205.1200 ;
        RECT 2355.3200 2182.8800 2356.9200 2183.3600 ;
        RECT 2355.3200 2188.3200 2356.9200 2188.8000 ;
        RECT 2355.3200 2193.7600 2356.9200 2194.2400 ;
        RECT 2355.3200 2172.0000 2356.9200 2172.4800 ;
        RECT 2355.3200 2177.4400 2356.9200 2177.9200 ;
        RECT 2310.3200 2182.8800 2311.9200 2183.3600 ;
        RECT 2310.3200 2188.3200 2311.9200 2188.8000 ;
        RECT 2310.3200 2193.7600 2311.9200 2194.2400 ;
        RECT 2310.3200 2172.0000 2311.9200 2172.4800 ;
        RECT 2310.3200 2177.4400 2311.9200 2177.9200 ;
        RECT 2355.3200 2155.6800 2356.9200 2156.1600 ;
        RECT 2355.3200 2161.1200 2356.9200 2161.6000 ;
        RECT 2355.3200 2166.5600 2356.9200 2167.0400 ;
        RECT 2355.3200 2150.2400 2356.9200 2150.7200 ;
        RECT 2310.3200 2155.6800 2311.9200 2156.1600 ;
        RECT 2310.3200 2161.1200 2311.9200 2161.6000 ;
        RECT 2310.3200 2166.5600 2311.9200 2167.0400 ;
        RECT 2310.3200 2150.2400 2311.9200 2150.7200 ;
        RECT 2265.3200 2182.8800 2266.9200 2183.3600 ;
        RECT 2265.3200 2188.3200 2266.9200 2188.8000 ;
        RECT 2265.3200 2193.7600 2266.9200 2194.2400 ;
        RECT 2253.5600 2182.8800 2256.5600 2183.3600 ;
        RECT 2253.5600 2188.3200 2256.5600 2188.8000 ;
        RECT 2253.5600 2193.7600 2256.5600 2194.2400 ;
        RECT 2265.3200 2172.0000 2266.9200 2172.4800 ;
        RECT 2265.3200 2177.4400 2266.9200 2177.9200 ;
        RECT 2253.5600 2172.0000 2256.5600 2172.4800 ;
        RECT 2253.5600 2177.4400 2256.5600 2177.9200 ;
        RECT 2265.3200 2155.6800 2266.9200 2156.1600 ;
        RECT 2265.3200 2161.1200 2266.9200 2161.6000 ;
        RECT 2265.3200 2166.5600 2266.9200 2167.0400 ;
        RECT 2253.5600 2155.6800 2256.5600 2156.1600 ;
        RECT 2253.5600 2161.1200 2256.5600 2161.6000 ;
        RECT 2253.5600 2166.5600 2256.5600 2167.0400 ;
        RECT 2253.5600 2150.2400 2256.5600 2150.7200 ;
        RECT 2265.3200 2150.2400 2266.9200 2150.7200 ;
        RECT 2253.5600 2355.1500 2460.6600 2358.1500 ;
        RECT 2253.5600 2142.0500 2460.6600 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 1912.4100 2446.9200 2128.5100 ;
        RECT 2400.3200 1912.4100 2401.9200 2128.5100 ;
        RECT 2355.3200 1912.4100 2356.9200 2128.5100 ;
        RECT 2310.3200 1912.4100 2311.9200 2128.5100 ;
        RECT 2265.3200 1912.4100 2266.9200 2128.5100 ;
        RECT 2457.6600 1912.4100 2460.6600 2128.5100 ;
        RECT 2253.5600 1912.4100 2256.5600 2128.5100 ;
      LAYER met3 ;
        RECT 2457.6600 2105.5600 2460.6600 2106.0400 ;
        RECT 2457.6600 2111.0000 2460.6600 2111.4800 ;
        RECT 2445.3200 2105.5600 2446.9200 2106.0400 ;
        RECT 2445.3200 2111.0000 2446.9200 2111.4800 ;
        RECT 2457.6600 2116.4400 2460.6600 2116.9200 ;
        RECT 2445.3200 2116.4400 2446.9200 2116.9200 ;
        RECT 2457.6600 2094.6800 2460.6600 2095.1600 ;
        RECT 2457.6600 2100.1200 2460.6600 2100.6000 ;
        RECT 2445.3200 2094.6800 2446.9200 2095.1600 ;
        RECT 2445.3200 2100.1200 2446.9200 2100.6000 ;
        RECT 2457.6600 2078.3600 2460.6600 2078.8400 ;
        RECT 2457.6600 2083.8000 2460.6600 2084.2800 ;
        RECT 2445.3200 2078.3600 2446.9200 2078.8400 ;
        RECT 2445.3200 2083.8000 2446.9200 2084.2800 ;
        RECT 2457.6600 2089.2400 2460.6600 2089.7200 ;
        RECT 2445.3200 2089.2400 2446.9200 2089.7200 ;
        RECT 2400.3200 2105.5600 2401.9200 2106.0400 ;
        RECT 2400.3200 2111.0000 2401.9200 2111.4800 ;
        RECT 2400.3200 2116.4400 2401.9200 2116.9200 ;
        RECT 2400.3200 2094.6800 2401.9200 2095.1600 ;
        RECT 2400.3200 2100.1200 2401.9200 2100.6000 ;
        RECT 2400.3200 2078.3600 2401.9200 2078.8400 ;
        RECT 2400.3200 2083.8000 2401.9200 2084.2800 ;
        RECT 2400.3200 2089.2400 2401.9200 2089.7200 ;
        RECT 2457.6600 2062.0400 2460.6600 2062.5200 ;
        RECT 2457.6600 2067.4800 2460.6600 2067.9600 ;
        RECT 2457.6600 2072.9200 2460.6600 2073.4000 ;
        RECT 2445.3200 2062.0400 2446.9200 2062.5200 ;
        RECT 2445.3200 2067.4800 2446.9200 2067.9600 ;
        RECT 2445.3200 2072.9200 2446.9200 2073.4000 ;
        RECT 2457.6600 2051.1600 2460.6600 2051.6400 ;
        RECT 2457.6600 2056.6000 2460.6600 2057.0800 ;
        RECT 2445.3200 2051.1600 2446.9200 2051.6400 ;
        RECT 2445.3200 2056.6000 2446.9200 2057.0800 ;
        RECT 2457.6600 2034.8400 2460.6600 2035.3200 ;
        RECT 2457.6600 2040.2800 2460.6600 2040.7600 ;
        RECT 2457.6600 2045.7200 2460.6600 2046.2000 ;
        RECT 2445.3200 2034.8400 2446.9200 2035.3200 ;
        RECT 2445.3200 2040.2800 2446.9200 2040.7600 ;
        RECT 2445.3200 2045.7200 2446.9200 2046.2000 ;
        RECT 2457.6600 2023.9600 2460.6600 2024.4400 ;
        RECT 2457.6600 2029.4000 2460.6600 2029.8800 ;
        RECT 2445.3200 2023.9600 2446.9200 2024.4400 ;
        RECT 2445.3200 2029.4000 2446.9200 2029.8800 ;
        RECT 2400.3200 2062.0400 2401.9200 2062.5200 ;
        RECT 2400.3200 2067.4800 2401.9200 2067.9600 ;
        RECT 2400.3200 2072.9200 2401.9200 2073.4000 ;
        RECT 2400.3200 2051.1600 2401.9200 2051.6400 ;
        RECT 2400.3200 2056.6000 2401.9200 2057.0800 ;
        RECT 2400.3200 2034.8400 2401.9200 2035.3200 ;
        RECT 2400.3200 2040.2800 2401.9200 2040.7600 ;
        RECT 2400.3200 2045.7200 2401.9200 2046.2000 ;
        RECT 2400.3200 2023.9600 2401.9200 2024.4400 ;
        RECT 2400.3200 2029.4000 2401.9200 2029.8800 ;
        RECT 2355.3200 2105.5600 2356.9200 2106.0400 ;
        RECT 2355.3200 2111.0000 2356.9200 2111.4800 ;
        RECT 2355.3200 2116.4400 2356.9200 2116.9200 ;
        RECT 2310.3200 2105.5600 2311.9200 2106.0400 ;
        RECT 2310.3200 2111.0000 2311.9200 2111.4800 ;
        RECT 2310.3200 2116.4400 2311.9200 2116.9200 ;
        RECT 2355.3200 2094.6800 2356.9200 2095.1600 ;
        RECT 2355.3200 2100.1200 2356.9200 2100.6000 ;
        RECT 2355.3200 2078.3600 2356.9200 2078.8400 ;
        RECT 2355.3200 2083.8000 2356.9200 2084.2800 ;
        RECT 2355.3200 2089.2400 2356.9200 2089.7200 ;
        RECT 2310.3200 2094.6800 2311.9200 2095.1600 ;
        RECT 2310.3200 2100.1200 2311.9200 2100.6000 ;
        RECT 2310.3200 2078.3600 2311.9200 2078.8400 ;
        RECT 2310.3200 2083.8000 2311.9200 2084.2800 ;
        RECT 2310.3200 2089.2400 2311.9200 2089.7200 ;
        RECT 2265.3200 2105.5600 2266.9200 2106.0400 ;
        RECT 2265.3200 2111.0000 2266.9200 2111.4800 ;
        RECT 2253.5600 2111.0000 2256.5600 2111.4800 ;
        RECT 2253.5600 2105.5600 2256.5600 2106.0400 ;
        RECT 2253.5600 2116.4400 2256.5600 2116.9200 ;
        RECT 2265.3200 2116.4400 2266.9200 2116.9200 ;
        RECT 2265.3200 2094.6800 2266.9200 2095.1600 ;
        RECT 2265.3200 2100.1200 2266.9200 2100.6000 ;
        RECT 2253.5600 2100.1200 2256.5600 2100.6000 ;
        RECT 2253.5600 2094.6800 2256.5600 2095.1600 ;
        RECT 2265.3200 2078.3600 2266.9200 2078.8400 ;
        RECT 2265.3200 2083.8000 2266.9200 2084.2800 ;
        RECT 2253.5600 2083.8000 2256.5600 2084.2800 ;
        RECT 2253.5600 2078.3600 2256.5600 2078.8400 ;
        RECT 2253.5600 2089.2400 2256.5600 2089.7200 ;
        RECT 2265.3200 2089.2400 2266.9200 2089.7200 ;
        RECT 2355.3200 2062.0400 2356.9200 2062.5200 ;
        RECT 2355.3200 2067.4800 2356.9200 2067.9600 ;
        RECT 2355.3200 2072.9200 2356.9200 2073.4000 ;
        RECT 2355.3200 2051.1600 2356.9200 2051.6400 ;
        RECT 2355.3200 2056.6000 2356.9200 2057.0800 ;
        RECT 2310.3200 2062.0400 2311.9200 2062.5200 ;
        RECT 2310.3200 2067.4800 2311.9200 2067.9600 ;
        RECT 2310.3200 2072.9200 2311.9200 2073.4000 ;
        RECT 2310.3200 2051.1600 2311.9200 2051.6400 ;
        RECT 2310.3200 2056.6000 2311.9200 2057.0800 ;
        RECT 2355.3200 2034.8400 2356.9200 2035.3200 ;
        RECT 2355.3200 2040.2800 2356.9200 2040.7600 ;
        RECT 2355.3200 2045.7200 2356.9200 2046.2000 ;
        RECT 2355.3200 2023.9600 2356.9200 2024.4400 ;
        RECT 2355.3200 2029.4000 2356.9200 2029.8800 ;
        RECT 2310.3200 2034.8400 2311.9200 2035.3200 ;
        RECT 2310.3200 2040.2800 2311.9200 2040.7600 ;
        RECT 2310.3200 2045.7200 2311.9200 2046.2000 ;
        RECT 2310.3200 2023.9600 2311.9200 2024.4400 ;
        RECT 2310.3200 2029.4000 2311.9200 2029.8800 ;
        RECT 2265.3200 2062.0400 2266.9200 2062.5200 ;
        RECT 2265.3200 2067.4800 2266.9200 2067.9600 ;
        RECT 2265.3200 2072.9200 2266.9200 2073.4000 ;
        RECT 2253.5600 2062.0400 2256.5600 2062.5200 ;
        RECT 2253.5600 2067.4800 2256.5600 2067.9600 ;
        RECT 2253.5600 2072.9200 2256.5600 2073.4000 ;
        RECT 2265.3200 2051.1600 2266.9200 2051.6400 ;
        RECT 2265.3200 2056.6000 2266.9200 2057.0800 ;
        RECT 2253.5600 2051.1600 2256.5600 2051.6400 ;
        RECT 2253.5600 2056.6000 2256.5600 2057.0800 ;
        RECT 2265.3200 2034.8400 2266.9200 2035.3200 ;
        RECT 2265.3200 2040.2800 2266.9200 2040.7600 ;
        RECT 2265.3200 2045.7200 2266.9200 2046.2000 ;
        RECT 2253.5600 2034.8400 2256.5600 2035.3200 ;
        RECT 2253.5600 2040.2800 2256.5600 2040.7600 ;
        RECT 2253.5600 2045.7200 2256.5600 2046.2000 ;
        RECT 2265.3200 2023.9600 2266.9200 2024.4400 ;
        RECT 2265.3200 2029.4000 2266.9200 2029.8800 ;
        RECT 2253.5600 2023.9600 2256.5600 2024.4400 ;
        RECT 2253.5600 2029.4000 2256.5600 2029.8800 ;
        RECT 2457.6600 2007.6400 2460.6600 2008.1200 ;
        RECT 2457.6600 2013.0800 2460.6600 2013.5600 ;
        RECT 2457.6600 2018.5200 2460.6600 2019.0000 ;
        RECT 2445.3200 2007.6400 2446.9200 2008.1200 ;
        RECT 2445.3200 2013.0800 2446.9200 2013.5600 ;
        RECT 2445.3200 2018.5200 2446.9200 2019.0000 ;
        RECT 2457.6600 1996.7600 2460.6600 1997.2400 ;
        RECT 2457.6600 2002.2000 2460.6600 2002.6800 ;
        RECT 2445.3200 1996.7600 2446.9200 1997.2400 ;
        RECT 2445.3200 2002.2000 2446.9200 2002.6800 ;
        RECT 2457.6600 1980.4400 2460.6600 1980.9200 ;
        RECT 2457.6600 1985.8800 2460.6600 1986.3600 ;
        RECT 2457.6600 1991.3200 2460.6600 1991.8000 ;
        RECT 2445.3200 1980.4400 2446.9200 1980.9200 ;
        RECT 2445.3200 1985.8800 2446.9200 1986.3600 ;
        RECT 2445.3200 1991.3200 2446.9200 1991.8000 ;
        RECT 2457.6600 1969.5600 2460.6600 1970.0400 ;
        RECT 2457.6600 1975.0000 2460.6600 1975.4800 ;
        RECT 2445.3200 1969.5600 2446.9200 1970.0400 ;
        RECT 2445.3200 1975.0000 2446.9200 1975.4800 ;
        RECT 2400.3200 2007.6400 2401.9200 2008.1200 ;
        RECT 2400.3200 2013.0800 2401.9200 2013.5600 ;
        RECT 2400.3200 2018.5200 2401.9200 2019.0000 ;
        RECT 2400.3200 1996.7600 2401.9200 1997.2400 ;
        RECT 2400.3200 2002.2000 2401.9200 2002.6800 ;
        RECT 2400.3200 1980.4400 2401.9200 1980.9200 ;
        RECT 2400.3200 1985.8800 2401.9200 1986.3600 ;
        RECT 2400.3200 1991.3200 2401.9200 1991.8000 ;
        RECT 2400.3200 1969.5600 2401.9200 1970.0400 ;
        RECT 2400.3200 1975.0000 2401.9200 1975.4800 ;
        RECT 2457.6600 1953.2400 2460.6600 1953.7200 ;
        RECT 2457.6600 1958.6800 2460.6600 1959.1600 ;
        RECT 2457.6600 1964.1200 2460.6600 1964.6000 ;
        RECT 2445.3200 1953.2400 2446.9200 1953.7200 ;
        RECT 2445.3200 1958.6800 2446.9200 1959.1600 ;
        RECT 2445.3200 1964.1200 2446.9200 1964.6000 ;
        RECT 2457.6600 1942.3600 2460.6600 1942.8400 ;
        RECT 2457.6600 1947.8000 2460.6600 1948.2800 ;
        RECT 2445.3200 1942.3600 2446.9200 1942.8400 ;
        RECT 2445.3200 1947.8000 2446.9200 1948.2800 ;
        RECT 2457.6600 1926.0400 2460.6600 1926.5200 ;
        RECT 2457.6600 1931.4800 2460.6600 1931.9600 ;
        RECT 2457.6600 1936.9200 2460.6600 1937.4000 ;
        RECT 2445.3200 1926.0400 2446.9200 1926.5200 ;
        RECT 2445.3200 1931.4800 2446.9200 1931.9600 ;
        RECT 2445.3200 1936.9200 2446.9200 1937.4000 ;
        RECT 2457.6600 1920.6000 2460.6600 1921.0800 ;
        RECT 2445.3200 1920.6000 2446.9200 1921.0800 ;
        RECT 2400.3200 1953.2400 2401.9200 1953.7200 ;
        RECT 2400.3200 1958.6800 2401.9200 1959.1600 ;
        RECT 2400.3200 1964.1200 2401.9200 1964.6000 ;
        RECT 2400.3200 1942.3600 2401.9200 1942.8400 ;
        RECT 2400.3200 1947.8000 2401.9200 1948.2800 ;
        RECT 2400.3200 1926.0400 2401.9200 1926.5200 ;
        RECT 2400.3200 1931.4800 2401.9200 1931.9600 ;
        RECT 2400.3200 1936.9200 2401.9200 1937.4000 ;
        RECT 2400.3200 1920.6000 2401.9200 1921.0800 ;
        RECT 2355.3200 2007.6400 2356.9200 2008.1200 ;
        RECT 2355.3200 2013.0800 2356.9200 2013.5600 ;
        RECT 2355.3200 2018.5200 2356.9200 2019.0000 ;
        RECT 2355.3200 1996.7600 2356.9200 1997.2400 ;
        RECT 2355.3200 2002.2000 2356.9200 2002.6800 ;
        RECT 2310.3200 2007.6400 2311.9200 2008.1200 ;
        RECT 2310.3200 2013.0800 2311.9200 2013.5600 ;
        RECT 2310.3200 2018.5200 2311.9200 2019.0000 ;
        RECT 2310.3200 1996.7600 2311.9200 1997.2400 ;
        RECT 2310.3200 2002.2000 2311.9200 2002.6800 ;
        RECT 2355.3200 1980.4400 2356.9200 1980.9200 ;
        RECT 2355.3200 1985.8800 2356.9200 1986.3600 ;
        RECT 2355.3200 1991.3200 2356.9200 1991.8000 ;
        RECT 2355.3200 1969.5600 2356.9200 1970.0400 ;
        RECT 2355.3200 1975.0000 2356.9200 1975.4800 ;
        RECT 2310.3200 1980.4400 2311.9200 1980.9200 ;
        RECT 2310.3200 1985.8800 2311.9200 1986.3600 ;
        RECT 2310.3200 1991.3200 2311.9200 1991.8000 ;
        RECT 2310.3200 1969.5600 2311.9200 1970.0400 ;
        RECT 2310.3200 1975.0000 2311.9200 1975.4800 ;
        RECT 2265.3200 2007.6400 2266.9200 2008.1200 ;
        RECT 2265.3200 2013.0800 2266.9200 2013.5600 ;
        RECT 2265.3200 2018.5200 2266.9200 2019.0000 ;
        RECT 2253.5600 2007.6400 2256.5600 2008.1200 ;
        RECT 2253.5600 2013.0800 2256.5600 2013.5600 ;
        RECT 2253.5600 2018.5200 2256.5600 2019.0000 ;
        RECT 2265.3200 1996.7600 2266.9200 1997.2400 ;
        RECT 2265.3200 2002.2000 2266.9200 2002.6800 ;
        RECT 2253.5600 1996.7600 2256.5600 1997.2400 ;
        RECT 2253.5600 2002.2000 2256.5600 2002.6800 ;
        RECT 2265.3200 1980.4400 2266.9200 1980.9200 ;
        RECT 2265.3200 1985.8800 2266.9200 1986.3600 ;
        RECT 2265.3200 1991.3200 2266.9200 1991.8000 ;
        RECT 2253.5600 1980.4400 2256.5600 1980.9200 ;
        RECT 2253.5600 1985.8800 2256.5600 1986.3600 ;
        RECT 2253.5600 1991.3200 2256.5600 1991.8000 ;
        RECT 2265.3200 1969.5600 2266.9200 1970.0400 ;
        RECT 2265.3200 1975.0000 2266.9200 1975.4800 ;
        RECT 2253.5600 1969.5600 2256.5600 1970.0400 ;
        RECT 2253.5600 1975.0000 2256.5600 1975.4800 ;
        RECT 2355.3200 1953.2400 2356.9200 1953.7200 ;
        RECT 2355.3200 1958.6800 2356.9200 1959.1600 ;
        RECT 2355.3200 1964.1200 2356.9200 1964.6000 ;
        RECT 2355.3200 1942.3600 2356.9200 1942.8400 ;
        RECT 2355.3200 1947.8000 2356.9200 1948.2800 ;
        RECT 2310.3200 1953.2400 2311.9200 1953.7200 ;
        RECT 2310.3200 1958.6800 2311.9200 1959.1600 ;
        RECT 2310.3200 1964.1200 2311.9200 1964.6000 ;
        RECT 2310.3200 1942.3600 2311.9200 1942.8400 ;
        RECT 2310.3200 1947.8000 2311.9200 1948.2800 ;
        RECT 2355.3200 1926.0400 2356.9200 1926.5200 ;
        RECT 2355.3200 1931.4800 2356.9200 1931.9600 ;
        RECT 2355.3200 1936.9200 2356.9200 1937.4000 ;
        RECT 2355.3200 1920.6000 2356.9200 1921.0800 ;
        RECT 2310.3200 1926.0400 2311.9200 1926.5200 ;
        RECT 2310.3200 1931.4800 2311.9200 1931.9600 ;
        RECT 2310.3200 1936.9200 2311.9200 1937.4000 ;
        RECT 2310.3200 1920.6000 2311.9200 1921.0800 ;
        RECT 2265.3200 1953.2400 2266.9200 1953.7200 ;
        RECT 2265.3200 1958.6800 2266.9200 1959.1600 ;
        RECT 2265.3200 1964.1200 2266.9200 1964.6000 ;
        RECT 2253.5600 1953.2400 2256.5600 1953.7200 ;
        RECT 2253.5600 1958.6800 2256.5600 1959.1600 ;
        RECT 2253.5600 1964.1200 2256.5600 1964.6000 ;
        RECT 2265.3200 1942.3600 2266.9200 1942.8400 ;
        RECT 2265.3200 1947.8000 2266.9200 1948.2800 ;
        RECT 2253.5600 1942.3600 2256.5600 1942.8400 ;
        RECT 2253.5600 1947.8000 2256.5600 1948.2800 ;
        RECT 2265.3200 1926.0400 2266.9200 1926.5200 ;
        RECT 2265.3200 1931.4800 2266.9200 1931.9600 ;
        RECT 2265.3200 1936.9200 2266.9200 1937.4000 ;
        RECT 2253.5600 1926.0400 2256.5600 1926.5200 ;
        RECT 2253.5600 1931.4800 2256.5600 1931.9600 ;
        RECT 2253.5600 1936.9200 2256.5600 1937.4000 ;
        RECT 2253.5600 1920.6000 2256.5600 1921.0800 ;
        RECT 2265.3200 1920.6000 2266.9200 1921.0800 ;
        RECT 2253.5600 2125.5100 2460.6600 2128.5100 ;
        RECT 2253.5600 1912.4100 2460.6600 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 1682.7700 2446.9200 1898.8700 ;
        RECT 2400.3200 1682.7700 2401.9200 1898.8700 ;
        RECT 2355.3200 1682.7700 2356.9200 1898.8700 ;
        RECT 2310.3200 1682.7700 2311.9200 1898.8700 ;
        RECT 2265.3200 1682.7700 2266.9200 1898.8700 ;
        RECT 2457.6600 1682.7700 2460.6600 1898.8700 ;
        RECT 2253.5600 1682.7700 2256.5600 1898.8700 ;
      LAYER met3 ;
        RECT 2457.6600 1875.9200 2460.6600 1876.4000 ;
        RECT 2457.6600 1881.3600 2460.6600 1881.8400 ;
        RECT 2445.3200 1875.9200 2446.9200 1876.4000 ;
        RECT 2445.3200 1881.3600 2446.9200 1881.8400 ;
        RECT 2457.6600 1886.8000 2460.6600 1887.2800 ;
        RECT 2445.3200 1886.8000 2446.9200 1887.2800 ;
        RECT 2457.6600 1865.0400 2460.6600 1865.5200 ;
        RECT 2457.6600 1870.4800 2460.6600 1870.9600 ;
        RECT 2445.3200 1865.0400 2446.9200 1865.5200 ;
        RECT 2445.3200 1870.4800 2446.9200 1870.9600 ;
        RECT 2457.6600 1848.7200 2460.6600 1849.2000 ;
        RECT 2457.6600 1854.1600 2460.6600 1854.6400 ;
        RECT 2445.3200 1848.7200 2446.9200 1849.2000 ;
        RECT 2445.3200 1854.1600 2446.9200 1854.6400 ;
        RECT 2457.6600 1859.6000 2460.6600 1860.0800 ;
        RECT 2445.3200 1859.6000 2446.9200 1860.0800 ;
        RECT 2400.3200 1875.9200 2401.9200 1876.4000 ;
        RECT 2400.3200 1881.3600 2401.9200 1881.8400 ;
        RECT 2400.3200 1886.8000 2401.9200 1887.2800 ;
        RECT 2400.3200 1865.0400 2401.9200 1865.5200 ;
        RECT 2400.3200 1870.4800 2401.9200 1870.9600 ;
        RECT 2400.3200 1848.7200 2401.9200 1849.2000 ;
        RECT 2400.3200 1854.1600 2401.9200 1854.6400 ;
        RECT 2400.3200 1859.6000 2401.9200 1860.0800 ;
        RECT 2457.6600 1832.4000 2460.6600 1832.8800 ;
        RECT 2457.6600 1837.8400 2460.6600 1838.3200 ;
        RECT 2457.6600 1843.2800 2460.6600 1843.7600 ;
        RECT 2445.3200 1832.4000 2446.9200 1832.8800 ;
        RECT 2445.3200 1837.8400 2446.9200 1838.3200 ;
        RECT 2445.3200 1843.2800 2446.9200 1843.7600 ;
        RECT 2457.6600 1821.5200 2460.6600 1822.0000 ;
        RECT 2457.6600 1826.9600 2460.6600 1827.4400 ;
        RECT 2445.3200 1821.5200 2446.9200 1822.0000 ;
        RECT 2445.3200 1826.9600 2446.9200 1827.4400 ;
        RECT 2457.6600 1805.2000 2460.6600 1805.6800 ;
        RECT 2457.6600 1810.6400 2460.6600 1811.1200 ;
        RECT 2457.6600 1816.0800 2460.6600 1816.5600 ;
        RECT 2445.3200 1805.2000 2446.9200 1805.6800 ;
        RECT 2445.3200 1810.6400 2446.9200 1811.1200 ;
        RECT 2445.3200 1816.0800 2446.9200 1816.5600 ;
        RECT 2457.6600 1794.3200 2460.6600 1794.8000 ;
        RECT 2457.6600 1799.7600 2460.6600 1800.2400 ;
        RECT 2445.3200 1794.3200 2446.9200 1794.8000 ;
        RECT 2445.3200 1799.7600 2446.9200 1800.2400 ;
        RECT 2400.3200 1832.4000 2401.9200 1832.8800 ;
        RECT 2400.3200 1837.8400 2401.9200 1838.3200 ;
        RECT 2400.3200 1843.2800 2401.9200 1843.7600 ;
        RECT 2400.3200 1821.5200 2401.9200 1822.0000 ;
        RECT 2400.3200 1826.9600 2401.9200 1827.4400 ;
        RECT 2400.3200 1805.2000 2401.9200 1805.6800 ;
        RECT 2400.3200 1810.6400 2401.9200 1811.1200 ;
        RECT 2400.3200 1816.0800 2401.9200 1816.5600 ;
        RECT 2400.3200 1794.3200 2401.9200 1794.8000 ;
        RECT 2400.3200 1799.7600 2401.9200 1800.2400 ;
        RECT 2355.3200 1875.9200 2356.9200 1876.4000 ;
        RECT 2355.3200 1881.3600 2356.9200 1881.8400 ;
        RECT 2355.3200 1886.8000 2356.9200 1887.2800 ;
        RECT 2310.3200 1875.9200 2311.9200 1876.4000 ;
        RECT 2310.3200 1881.3600 2311.9200 1881.8400 ;
        RECT 2310.3200 1886.8000 2311.9200 1887.2800 ;
        RECT 2355.3200 1865.0400 2356.9200 1865.5200 ;
        RECT 2355.3200 1870.4800 2356.9200 1870.9600 ;
        RECT 2355.3200 1848.7200 2356.9200 1849.2000 ;
        RECT 2355.3200 1854.1600 2356.9200 1854.6400 ;
        RECT 2355.3200 1859.6000 2356.9200 1860.0800 ;
        RECT 2310.3200 1865.0400 2311.9200 1865.5200 ;
        RECT 2310.3200 1870.4800 2311.9200 1870.9600 ;
        RECT 2310.3200 1848.7200 2311.9200 1849.2000 ;
        RECT 2310.3200 1854.1600 2311.9200 1854.6400 ;
        RECT 2310.3200 1859.6000 2311.9200 1860.0800 ;
        RECT 2265.3200 1875.9200 2266.9200 1876.4000 ;
        RECT 2265.3200 1881.3600 2266.9200 1881.8400 ;
        RECT 2253.5600 1881.3600 2256.5600 1881.8400 ;
        RECT 2253.5600 1875.9200 2256.5600 1876.4000 ;
        RECT 2253.5600 1886.8000 2256.5600 1887.2800 ;
        RECT 2265.3200 1886.8000 2266.9200 1887.2800 ;
        RECT 2265.3200 1865.0400 2266.9200 1865.5200 ;
        RECT 2265.3200 1870.4800 2266.9200 1870.9600 ;
        RECT 2253.5600 1870.4800 2256.5600 1870.9600 ;
        RECT 2253.5600 1865.0400 2256.5600 1865.5200 ;
        RECT 2265.3200 1848.7200 2266.9200 1849.2000 ;
        RECT 2265.3200 1854.1600 2266.9200 1854.6400 ;
        RECT 2253.5600 1854.1600 2256.5600 1854.6400 ;
        RECT 2253.5600 1848.7200 2256.5600 1849.2000 ;
        RECT 2253.5600 1859.6000 2256.5600 1860.0800 ;
        RECT 2265.3200 1859.6000 2266.9200 1860.0800 ;
        RECT 2355.3200 1832.4000 2356.9200 1832.8800 ;
        RECT 2355.3200 1837.8400 2356.9200 1838.3200 ;
        RECT 2355.3200 1843.2800 2356.9200 1843.7600 ;
        RECT 2355.3200 1821.5200 2356.9200 1822.0000 ;
        RECT 2355.3200 1826.9600 2356.9200 1827.4400 ;
        RECT 2310.3200 1832.4000 2311.9200 1832.8800 ;
        RECT 2310.3200 1837.8400 2311.9200 1838.3200 ;
        RECT 2310.3200 1843.2800 2311.9200 1843.7600 ;
        RECT 2310.3200 1821.5200 2311.9200 1822.0000 ;
        RECT 2310.3200 1826.9600 2311.9200 1827.4400 ;
        RECT 2355.3200 1805.2000 2356.9200 1805.6800 ;
        RECT 2355.3200 1810.6400 2356.9200 1811.1200 ;
        RECT 2355.3200 1816.0800 2356.9200 1816.5600 ;
        RECT 2355.3200 1794.3200 2356.9200 1794.8000 ;
        RECT 2355.3200 1799.7600 2356.9200 1800.2400 ;
        RECT 2310.3200 1805.2000 2311.9200 1805.6800 ;
        RECT 2310.3200 1810.6400 2311.9200 1811.1200 ;
        RECT 2310.3200 1816.0800 2311.9200 1816.5600 ;
        RECT 2310.3200 1794.3200 2311.9200 1794.8000 ;
        RECT 2310.3200 1799.7600 2311.9200 1800.2400 ;
        RECT 2265.3200 1832.4000 2266.9200 1832.8800 ;
        RECT 2265.3200 1837.8400 2266.9200 1838.3200 ;
        RECT 2265.3200 1843.2800 2266.9200 1843.7600 ;
        RECT 2253.5600 1832.4000 2256.5600 1832.8800 ;
        RECT 2253.5600 1837.8400 2256.5600 1838.3200 ;
        RECT 2253.5600 1843.2800 2256.5600 1843.7600 ;
        RECT 2265.3200 1821.5200 2266.9200 1822.0000 ;
        RECT 2265.3200 1826.9600 2266.9200 1827.4400 ;
        RECT 2253.5600 1821.5200 2256.5600 1822.0000 ;
        RECT 2253.5600 1826.9600 2256.5600 1827.4400 ;
        RECT 2265.3200 1805.2000 2266.9200 1805.6800 ;
        RECT 2265.3200 1810.6400 2266.9200 1811.1200 ;
        RECT 2265.3200 1816.0800 2266.9200 1816.5600 ;
        RECT 2253.5600 1805.2000 2256.5600 1805.6800 ;
        RECT 2253.5600 1810.6400 2256.5600 1811.1200 ;
        RECT 2253.5600 1816.0800 2256.5600 1816.5600 ;
        RECT 2265.3200 1794.3200 2266.9200 1794.8000 ;
        RECT 2265.3200 1799.7600 2266.9200 1800.2400 ;
        RECT 2253.5600 1794.3200 2256.5600 1794.8000 ;
        RECT 2253.5600 1799.7600 2256.5600 1800.2400 ;
        RECT 2457.6600 1778.0000 2460.6600 1778.4800 ;
        RECT 2457.6600 1783.4400 2460.6600 1783.9200 ;
        RECT 2457.6600 1788.8800 2460.6600 1789.3600 ;
        RECT 2445.3200 1778.0000 2446.9200 1778.4800 ;
        RECT 2445.3200 1783.4400 2446.9200 1783.9200 ;
        RECT 2445.3200 1788.8800 2446.9200 1789.3600 ;
        RECT 2457.6600 1767.1200 2460.6600 1767.6000 ;
        RECT 2457.6600 1772.5600 2460.6600 1773.0400 ;
        RECT 2445.3200 1767.1200 2446.9200 1767.6000 ;
        RECT 2445.3200 1772.5600 2446.9200 1773.0400 ;
        RECT 2457.6600 1750.8000 2460.6600 1751.2800 ;
        RECT 2457.6600 1756.2400 2460.6600 1756.7200 ;
        RECT 2457.6600 1761.6800 2460.6600 1762.1600 ;
        RECT 2445.3200 1750.8000 2446.9200 1751.2800 ;
        RECT 2445.3200 1756.2400 2446.9200 1756.7200 ;
        RECT 2445.3200 1761.6800 2446.9200 1762.1600 ;
        RECT 2457.6600 1739.9200 2460.6600 1740.4000 ;
        RECT 2457.6600 1745.3600 2460.6600 1745.8400 ;
        RECT 2445.3200 1739.9200 2446.9200 1740.4000 ;
        RECT 2445.3200 1745.3600 2446.9200 1745.8400 ;
        RECT 2400.3200 1778.0000 2401.9200 1778.4800 ;
        RECT 2400.3200 1783.4400 2401.9200 1783.9200 ;
        RECT 2400.3200 1788.8800 2401.9200 1789.3600 ;
        RECT 2400.3200 1767.1200 2401.9200 1767.6000 ;
        RECT 2400.3200 1772.5600 2401.9200 1773.0400 ;
        RECT 2400.3200 1750.8000 2401.9200 1751.2800 ;
        RECT 2400.3200 1756.2400 2401.9200 1756.7200 ;
        RECT 2400.3200 1761.6800 2401.9200 1762.1600 ;
        RECT 2400.3200 1739.9200 2401.9200 1740.4000 ;
        RECT 2400.3200 1745.3600 2401.9200 1745.8400 ;
        RECT 2457.6600 1723.6000 2460.6600 1724.0800 ;
        RECT 2457.6600 1729.0400 2460.6600 1729.5200 ;
        RECT 2457.6600 1734.4800 2460.6600 1734.9600 ;
        RECT 2445.3200 1723.6000 2446.9200 1724.0800 ;
        RECT 2445.3200 1729.0400 2446.9200 1729.5200 ;
        RECT 2445.3200 1734.4800 2446.9200 1734.9600 ;
        RECT 2457.6600 1712.7200 2460.6600 1713.2000 ;
        RECT 2457.6600 1718.1600 2460.6600 1718.6400 ;
        RECT 2445.3200 1712.7200 2446.9200 1713.2000 ;
        RECT 2445.3200 1718.1600 2446.9200 1718.6400 ;
        RECT 2457.6600 1696.4000 2460.6600 1696.8800 ;
        RECT 2457.6600 1701.8400 2460.6600 1702.3200 ;
        RECT 2457.6600 1707.2800 2460.6600 1707.7600 ;
        RECT 2445.3200 1696.4000 2446.9200 1696.8800 ;
        RECT 2445.3200 1701.8400 2446.9200 1702.3200 ;
        RECT 2445.3200 1707.2800 2446.9200 1707.7600 ;
        RECT 2457.6600 1690.9600 2460.6600 1691.4400 ;
        RECT 2445.3200 1690.9600 2446.9200 1691.4400 ;
        RECT 2400.3200 1723.6000 2401.9200 1724.0800 ;
        RECT 2400.3200 1729.0400 2401.9200 1729.5200 ;
        RECT 2400.3200 1734.4800 2401.9200 1734.9600 ;
        RECT 2400.3200 1712.7200 2401.9200 1713.2000 ;
        RECT 2400.3200 1718.1600 2401.9200 1718.6400 ;
        RECT 2400.3200 1696.4000 2401.9200 1696.8800 ;
        RECT 2400.3200 1701.8400 2401.9200 1702.3200 ;
        RECT 2400.3200 1707.2800 2401.9200 1707.7600 ;
        RECT 2400.3200 1690.9600 2401.9200 1691.4400 ;
        RECT 2355.3200 1778.0000 2356.9200 1778.4800 ;
        RECT 2355.3200 1783.4400 2356.9200 1783.9200 ;
        RECT 2355.3200 1788.8800 2356.9200 1789.3600 ;
        RECT 2355.3200 1767.1200 2356.9200 1767.6000 ;
        RECT 2355.3200 1772.5600 2356.9200 1773.0400 ;
        RECT 2310.3200 1778.0000 2311.9200 1778.4800 ;
        RECT 2310.3200 1783.4400 2311.9200 1783.9200 ;
        RECT 2310.3200 1788.8800 2311.9200 1789.3600 ;
        RECT 2310.3200 1767.1200 2311.9200 1767.6000 ;
        RECT 2310.3200 1772.5600 2311.9200 1773.0400 ;
        RECT 2355.3200 1750.8000 2356.9200 1751.2800 ;
        RECT 2355.3200 1756.2400 2356.9200 1756.7200 ;
        RECT 2355.3200 1761.6800 2356.9200 1762.1600 ;
        RECT 2355.3200 1739.9200 2356.9200 1740.4000 ;
        RECT 2355.3200 1745.3600 2356.9200 1745.8400 ;
        RECT 2310.3200 1750.8000 2311.9200 1751.2800 ;
        RECT 2310.3200 1756.2400 2311.9200 1756.7200 ;
        RECT 2310.3200 1761.6800 2311.9200 1762.1600 ;
        RECT 2310.3200 1739.9200 2311.9200 1740.4000 ;
        RECT 2310.3200 1745.3600 2311.9200 1745.8400 ;
        RECT 2265.3200 1778.0000 2266.9200 1778.4800 ;
        RECT 2265.3200 1783.4400 2266.9200 1783.9200 ;
        RECT 2265.3200 1788.8800 2266.9200 1789.3600 ;
        RECT 2253.5600 1778.0000 2256.5600 1778.4800 ;
        RECT 2253.5600 1783.4400 2256.5600 1783.9200 ;
        RECT 2253.5600 1788.8800 2256.5600 1789.3600 ;
        RECT 2265.3200 1767.1200 2266.9200 1767.6000 ;
        RECT 2265.3200 1772.5600 2266.9200 1773.0400 ;
        RECT 2253.5600 1767.1200 2256.5600 1767.6000 ;
        RECT 2253.5600 1772.5600 2256.5600 1773.0400 ;
        RECT 2265.3200 1750.8000 2266.9200 1751.2800 ;
        RECT 2265.3200 1756.2400 2266.9200 1756.7200 ;
        RECT 2265.3200 1761.6800 2266.9200 1762.1600 ;
        RECT 2253.5600 1750.8000 2256.5600 1751.2800 ;
        RECT 2253.5600 1756.2400 2256.5600 1756.7200 ;
        RECT 2253.5600 1761.6800 2256.5600 1762.1600 ;
        RECT 2265.3200 1739.9200 2266.9200 1740.4000 ;
        RECT 2265.3200 1745.3600 2266.9200 1745.8400 ;
        RECT 2253.5600 1739.9200 2256.5600 1740.4000 ;
        RECT 2253.5600 1745.3600 2256.5600 1745.8400 ;
        RECT 2355.3200 1723.6000 2356.9200 1724.0800 ;
        RECT 2355.3200 1729.0400 2356.9200 1729.5200 ;
        RECT 2355.3200 1734.4800 2356.9200 1734.9600 ;
        RECT 2355.3200 1712.7200 2356.9200 1713.2000 ;
        RECT 2355.3200 1718.1600 2356.9200 1718.6400 ;
        RECT 2310.3200 1723.6000 2311.9200 1724.0800 ;
        RECT 2310.3200 1729.0400 2311.9200 1729.5200 ;
        RECT 2310.3200 1734.4800 2311.9200 1734.9600 ;
        RECT 2310.3200 1712.7200 2311.9200 1713.2000 ;
        RECT 2310.3200 1718.1600 2311.9200 1718.6400 ;
        RECT 2355.3200 1696.4000 2356.9200 1696.8800 ;
        RECT 2355.3200 1701.8400 2356.9200 1702.3200 ;
        RECT 2355.3200 1707.2800 2356.9200 1707.7600 ;
        RECT 2355.3200 1690.9600 2356.9200 1691.4400 ;
        RECT 2310.3200 1696.4000 2311.9200 1696.8800 ;
        RECT 2310.3200 1701.8400 2311.9200 1702.3200 ;
        RECT 2310.3200 1707.2800 2311.9200 1707.7600 ;
        RECT 2310.3200 1690.9600 2311.9200 1691.4400 ;
        RECT 2265.3200 1723.6000 2266.9200 1724.0800 ;
        RECT 2265.3200 1729.0400 2266.9200 1729.5200 ;
        RECT 2265.3200 1734.4800 2266.9200 1734.9600 ;
        RECT 2253.5600 1723.6000 2256.5600 1724.0800 ;
        RECT 2253.5600 1729.0400 2256.5600 1729.5200 ;
        RECT 2253.5600 1734.4800 2256.5600 1734.9600 ;
        RECT 2265.3200 1712.7200 2266.9200 1713.2000 ;
        RECT 2265.3200 1718.1600 2266.9200 1718.6400 ;
        RECT 2253.5600 1712.7200 2256.5600 1713.2000 ;
        RECT 2253.5600 1718.1600 2256.5600 1718.6400 ;
        RECT 2265.3200 1696.4000 2266.9200 1696.8800 ;
        RECT 2265.3200 1701.8400 2266.9200 1702.3200 ;
        RECT 2265.3200 1707.2800 2266.9200 1707.7600 ;
        RECT 2253.5600 1696.4000 2256.5600 1696.8800 ;
        RECT 2253.5600 1701.8400 2256.5600 1702.3200 ;
        RECT 2253.5600 1707.2800 2256.5600 1707.7600 ;
        RECT 2253.5600 1690.9600 2256.5600 1691.4400 ;
        RECT 2265.3200 1690.9600 2266.9200 1691.4400 ;
        RECT 2253.5600 1895.8700 2460.6600 1898.8700 ;
        RECT 2253.5600 1682.7700 2460.6600 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 1453.1300 2446.9200 1669.2300 ;
        RECT 2400.3200 1453.1300 2401.9200 1669.2300 ;
        RECT 2355.3200 1453.1300 2356.9200 1669.2300 ;
        RECT 2310.3200 1453.1300 2311.9200 1669.2300 ;
        RECT 2265.3200 1453.1300 2266.9200 1669.2300 ;
        RECT 2457.6600 1453.1300 2460.6600 1669.2300 ;
        RECT 2253.5600 1453.1300 2256.5600 1669.2300 ;
      LAYER met3 ;
        RECT 2457.6600 1646.2800 2460.6600 1646.7600 ;
        RECT 2457.6600 1651.7200 2460.6600 1652.2000 ;
        RECT 2445.3200 1646.2800 2446.9200 1646.7600 ;
        RECT 2445.3200 1651.7200 2446.9200 1652.2000 ;
        RECT 2457.6600 1657.1600 2460.6600 1657.6400 ;
        RECT 2445.3200 1657.1600 2446.9200 1657.6400 ;
        RECT 2457.6600 1635.4000 2460.6600 1635.8800 ;
        RECT 2457.6600 1640.8400 2460.6600 1641.3200 ;
        RECT 2445.3200 1635.4000 2446.9200 1635.8800 ;
        RECT 2445.3200 1640.8400 2446.9200 1641.3200 ;
        RECT 2457.6600 1619.0800 2460.6600 1619.5600 ;
        RECT 2457.6600 1624.5200 2460.6600 1625.0000 ;
        RECT 2445.3200 1619.0800 2446.9200 1619.5600 ;
        RECT 2445.3200 1624.5200 2446.9200 1625.0000 ;
        RECT 2457.6600 1629.9600 2460.6600 1630.4400 ;
        RECT 2445.3200 1629.9600 2446.9200 1630.4400 ;
        RECT 2400.3200 1646.2800 2401.9200 1646.7600 ;
        RECT 2400.3200 1651.7200 2401.9200 1652.2000 ;
        RECT 2400.3200 1657.1600 2401.9200 1657.6400 ;
        RECT 2400.3200 1635.4000 2401.9200 1635.8800 ;
        RECT 2400.3200 1640.8400 2401.9200 1641.3200 ;
        RECT 2400.3200 1619.0800 2401.9200 1619.5600 ;
        RECT 2400.3200 1624.5200 2401.9200 1625.0000 ;
        RECT 2400.3200 1629.9600 2401.9200 1630.4400 ;
        RECT 2457.6600 1602.7600 2460.6600 1603.2400 ;
        RECT 2457.6600 1608.2000 2460.6600 1608.6800 ;
        RECT 2457.6600 1613.6400 2460.6600 1614.1200 ;
        RECT 2445.3200 1602.7600 2446.9200 1603.2400 ;
        RECT 2445.3200 1608.2000 2446.9200 1608.6800 ;
        RECT 2445.3200 1613.6400 2446.9200 1614.1200 ;
        RECT 2457.6600 1591.8800 2460.6600 1592.3600 ;
        RECT 2457.6600 1597.3200 2460.6600 1597.8000 ;
        RECT 2445.3200 1591.8800 2446.9200 1592.3600 ;
        RECT 2445.3200 1597.3200 2446.9200 1597.8000 ;
        RECT 2457.6600 1575.5600 2460.6600 1576.0400 ;
        RECT 2457.6600 1581.0000 2460.6600 1581.4800 ;
        RECT 2457.6600 1586.4400 2460.6600 1586.9200 ;
        RECT 2445.3200 1575.5600 2446.9200 1576.0400 ;
        RECT 2445.3200 1581.0000 2446.9200 1581.4800 ;
        RECT 2445.3200 1586.4400 2446.9200 1586.9200 ;
        RECT 2457.6600 1564.6800 2460.6600 1565.1600 ;
        RECT 2457.6600 1570.1200 2460.6600 1570.6000 ;
        RECT 2445.3200 1564.6800 2446.9200 1565.1600 ;
        RECT 2445.3200 1570.1200 2446.9200 1570.6000 ;
        RECT 2400.3200 1602.7600 2401.9200 1603.2400 ;
        RECT 2400.3200 1608.2000 2401.9200 1608.6800 ;
        RECT 2400.3200 1613.6400 2401.9200 1614.1200 ;
        RECT 2400.3200 1591.8800 2401.9200 1592.3600 ;
        RECT 2400.3200 1597.3200 2401.9200 1597.8000 ;
        RECT 2400.3200 1575.5600 2401.9200 1576.0400 ;
        RECT 2400.3200 1581.0000 2401.9200 1581.4800 ;
        RECT 2400.3200 1586.4400 2401.9200 1586.9200 ;
        RECT 2400.3200 1564.6800 2401.9200 1565.1600 ;
        RECT 2400.3200 1570.1200 2401.9200 1570.6000 ;
        RECT 2355.3200 1646.2800 2356.9200 1646.7600 ;
        RECT 2355.3200 1651.7200 2356.9200 1652.2000 ;
        RECT 2355.3200 1657.1600 2356.9200 1657.6400 ;
        RECT 2310.3200 1646.2800 2311.9200 1646.7600 ;
        RECT 2310.3200 1651.7200 2311.9200 1652.2000 ;
        RECT 2310.3200 1657.1600 2311.9200 1657.6400 ;
        RECT 2355.3200 1635.4000 2356.9200 1635.8800 ;
        RECT 2355.3200 1640.8400 2356.9200 1641.3200 ;
        RECT 2355.3200 1619.0800 2356.9200 1619.5600 ;
        RECT 2355.3200 1624.5200 2356.9200 1625.0000 ;
        RECT 2355.3200 1629.9600 2356.9200 1630.4400 ;
        RECT 2310.3200 1635.4000 2311.9200 1635.8800 ;
        RECT 2310.3200 1640.8400 2311.9200 1641.3200 ;
        RECT 2310.3200 1619.0800 2311.9200 1619.5600 ;
        RECT 2310.3200 1624.5200 2311.9200 1625.0000 ;
        RECT 2310.3200 1629.9600 2311.9200 1630.4400 ;
        RECT 2265.3200 1646.2800 2266.9200 1646.7600 ;
        RECT 2265.3200 1651.7200 2266.9200 1652.2000 ;
        RECT 2253.5600 1651.7200 2256.5600 1652.2000 ;
        RECT 2253.5600 1646.2800 2256.5600 1646.7600 ;
        RECT 2253.5600 1657.1600 2256.5600 1657.6400 ;
        RECT 2265.3200 1657.1600 2266.9200 1657.6400 ;
        RECT 2265.3200 1635.4000 2266.9200 1635.8800 ;
        RECT 2265.3200 1640.8400 2266.9200 1641.3200 ;
        RECT 2253.5600 1640.8400 2256.5600 1641.3200 ;
        RECT 2253.5600 1635.4000 2256.5600 1635.8800 ;
        RECT 2265.3200 1619.0800 2266.9200 1619.5600 ;
        RECT 2265.3200 1624.5200 2266.9200 1625.0000 ;
        RECT 2253.5600 1624.5200 2256.5600 1625.0000 ;
        RECT 2253.5600 1619.0800 2256.5600 1619.5600 ;
        RECT 2253.5600 1629.9600 2256.5600 1630.4400 ;
        RECT 2265.3200 1629.9600 2266.9200 1630.4400 ;
        RECT 2355.3200 1602.7600 2356.9200 1603.2400 ;
        RECT 2355.3200 1608.2000 2356.9200 1608.6800 ;
        RECT 2355.3200 1613.6400 2356.9200 1614.1200 ;
        RECT 2355.3200 1591.8800 2356.9200 1592.3600 ;
        RECT 2355.3200 1597.3200 2356.9200 1597.8000 ;
        RECT 2310.3200 1602.7600 2311.9200 1603.2400 ;
        RECT 2310.3200 1608.2000 2311.9200 1608.6800 ;
        RECT 2310.3200 1613.6400 2311.9200 1614.1200 ;
        RECT 2310.3200 1591.8800 2311.9200 1592.3600 ;
        RECT 2310.3200 1597.3200 2311.9200 1597.8000 ;
        RECT 2355.3200 1575.5600 2356.9200 1576.0400 ;
        RECT 2355.3200 1581.0000 2356.9200 1581.4800 ;
        RECT 2355.3200 1586.4400 2356.9200 1586.9200 ;
        RECT 2355.3200 1564.6800 2356.9200 1565.1600 ;
        RECT 2355.3200 1570.1200 2356.9200 1570.6000 ;
        RECT 2310.3200 1575.5600 2311.9200 1576.0400 ;
        RECT 2310.3200 1581.0000 2311.9200 1581.4800 ;
        RECT 2310.3200 1586.4400 2311.9200 1586.9200 ;
        RECT 2310.3200 1564.6800 2311.9200 1565.1600 ;
        RECT 2310.3200 1570.1200 2311.9200 1570.6000 ;
        RECT 2265.3200 1602.7600 2266.9200 1603.2400 ;
        RECT 2265.3200 1608.2000 2266.9200 1608.6800 ;
        RECT 2265.3200 1613.6400 2266.9200 1614.1200 ;
        RECT 2253.5600 1602.7600 2256.5600 1603.2400 ;
        RECT 2253.5600 1608.2000 2256.5600 1608.6800 ;
        RECT 2253.5600 1613.6400 2256.5600 1614.1200 ;
        RECT 2265.3200 1591.8800 2266.9200 1592.3600 ;
        RECT 2265.3200 1597.3200 2266.9200 1597.8000 ;
        RECT 2253.5600 1591.8800 2256.5600 1592.3600 ;
        RECT 2253.5600 1597.3200 2256.5600 1597.8000 ;
        RECT 2265.3200 1575.5600 2266.9200 1576.0400 ;
        RECT 2265.3200 1581.0000 2266.9200 1581.4800 ;
        RECT 2265.3200 1586.4400 2266.9200 1586.9200 ;
        RECT 2253.5600 1575.5600 2256.5600 1576.0400 ;
        RECT 2253.5600 1581.0000 2256.5600 1581.4800 ;
        RECT 2253.5600 1586.4400 2256.5600 1586.9200 ;
        RECT 2265.3200 1564.6800 2266.9200 1565.1600 ;
        RECT 2265.3200 1570.1200 2266.9200 1570.6000 ;
        RECT 2253.5600 1564.6800 2256.5600 1565.1600 ;
        RECT 2253.5600 1570.1200 2256.5600 1570.6000 ;
        RECT 2457.6600 1548.3600 2460.6600 1548.8400 ;
        RECT 2457.6600 1553.8000 2460.6600 1554.2800 ;
        RECT 2457.6600 1559.2400 2460.6600 1559.7200 ;
        RECT 2445.3200 1548.3600 2446.9200 1548.8400 ;
        RECT 2445.3200 1553.8000 2446.9200 1554.2800 ;
        RECT 2445.3200 1559.2400 2446.9200 1559.7200 ;
        RECT 2457.6600 1537.4800 2460.6600 1537.9600 ;
        RECT 2457.6600 1542.9200 2460.6600 1543.4000 ;
        RECT 2445.3200 1537.4800 2446.9200 1537.9600 ;
        RECT 2445.3200 1542.9200 2446.9200 1543.4000 ;
        RECT 2457.6600 1521.1600 2460.6600 1521.6400 ;
        RECT 2457.6600 1526.6000 2460.6600 1527.0800 ;
        RECT 2457.6600 1532.0400 2460.6600 1532.5200 ;
        RECT 2445.3200 1521.1600 2446.9200 1521.6400 ;
        RECT 2445.3200 1526.6000 2446.9200 1527.0800 ;
        RECT 2445.3200 1532.0400 2446.9200 1532.5200 ;
        RECT 2457.6600 1510.2800 2460.6600 1510.7600 ;
        RECT 2457.6600 1515.7200 2460.6600 1516.2000 ;
        RECT 2445.3200 1510.2800 2446.9200 1510.7600 ;
        RECT 2445.3200 1515.7200 2446.9200 1516.2000 ;
        RECT 2400.3200 1548.3600 2401.9200 1548.8400 ;
        RECT 2400.3200 1553.8000 2401.9200 1554.2800 ;
        RECT 2400.3200 1559.2400 2401.9200 1559.7200 ;
        RECT 2400.3200 1537.4800 2401.9200 1537.9600 ;
        RECT 2400.3200 1542.9200 2401.9200 1543.4000 ;
        RECT 2400.3200 1521.1600 2401.9200 1521.6400 ;
        RECT 2400.3200 1526.6000 2401.9200 1527.0800 ;
        RECT 2400.3200 1532.0400 2401.9200 1532.5200 ;
        RECT 2400.3200 1510.2800 2401.9200 1510.7600 ;
        RECT 2400.3200 1515.7200 2401.9200 1516.2000 ;
        RECT 2457.6600 1493.9600 2460.6600 1494.4400 ;
        RECT 2457.6600 1499.4000 2460.6600 1499.8800 ;
        RECT 2457.6600 1504.8400 2460.6600 1505.3200 ;
        RECT 2445.3200 1493.9600 2446.9200 1494.4400 ;
        RECT 2445.3200 1499.4000 2446.9200 1499.8800 ;
        RECT 2445.3200 1504.8400 2446.9200 1505.3200 ;
        RECT 2457.6600 1483.0800 2460.6600 1483.5600 ;
        RECT 2457.6600 1488.5200 2460.6600 1489.0000 ;
        RECT 2445.3200 1483.0800 2446.9200 1483.5600 ;
        RECT 2445.3200 1488.5200 2446.9200 1489.0000 ;
        RECT 2457.6600 1466.7600 2460.6600 1467.2400 ;
        RECT 2457.6600 1472.2000 2460.6600 1472.6800 ;
        RECT 2457.6600 1477.6400 2460.6600 1478.1200 ;
        RECT 2445.3200 1466.7600 2446.9200 1467.2400 ;
        RECT 2445.3200 1472.2000 2446.9200 1472.6800 ;
        RECT 2445.3200 1477.6400 2446.9200 1478.1200 ;
        RECT 2457.6600 1461.3200 2460.6600 1461.8000 ;
        RECT 2445.3200 1461.3200 2446.9200 1461.8000 ;
        RECT 2400.3200 1493.9600 2401.9200 1494.4400 ;
        RECT 2400.3200 1499.4000 2401.9200 1499.8800 ;
        RECT 2400.3200 1504.8400 2401.9200 1505.3200 ;
        RECT 2400.3200 1483.0800 2401.9200 1483.5600 ;
        RECT 2400.3200 1488.5200 2401.9200 1489.0000 ;
        RECT 2400.3200 1466.7600 2401.9200 1467.2400 ;
        RECT 2400.3200 1472.2000 2401.9200 1472.6800 ;
        RECT 2400.3200 1477.6400 2401.9200 1478.1200 ;
        RECT 2400.3200 1461.3200 2401.9200 1461.8000 ;
        RECT 2355.3200 1548.3600 2356.9200 1548.8400 ;
        RECT 2355.3200 1553.8000 2356.9200 1554.2800 ;
        RECT 2355.3200 1559.2400 2356.9200 1559.7200 ;
        RECT 2355.3200 1537.4800 2356.9200 1537.9600 ;
        RECT 2355.3200 1542.9200 2356.9200 1543.4000 ;
        RECT 2310.3200 1548.3600 2311.9200 1548.8400 ;
        RECT 2310.3200 1553.8000 2311.9200 1554.2800 ;
        RECT 2310.3200 1559.2400 2311.9200 1559.7200 ;
        RECT 2310.3200 1537.4800 2311.9200 1537.9600 ;
        RECT 2310.3200 1542.9200 2311.9200 1543.4000 ;
        RECT 2355.3200 1521.1600 2356.9200 1521.6400 ;
        RECT 2355.3200 1526.6000 2356.9200 1527.0800 ;
        RECT 2355.3200 1532.0400 2356.9200 1532.5200 ;
        RECT 2355.3200 1510.2800 2356.9200 1510.7600 ;
        RECT 2355.3200 1515.7200 2356.9200 1516.2000 ;
        RECT 2310.3200 1521.1600 2311.9200 1521.6400 ;
        RECT 2310.3200 1526.6000 2311.9200 1527.0800 ;
        RECT 2310.3200 1532.0400 2311.9200 1532.5200 ;
        RECT 2310.3200 1510.2800 2311.9200 1510.7600 ;
        RECT 2310.3200 1515.7200 2311.9200 1516.2000 ;
        RECT 2265.3200 1548.3600 2266.9200 1548.8400 ;
        RECT 2265.3200 1553.8000 2266.9200 1554.2800 ;
        RECT 2265.3200 1559.2400 2266.9200 1559.7200 ;
        RECT 2253.5600 1548.3600 2256.5600 1548.8400 ;
        RECT 2253.5600 1553.8000 2256.5600 1554.2800 ;
        RECT 2253.5600 1559.2400 2256.5600 1559.7200 ;
        RECT 2265.3200 1537.4800 2266.9200 1537.9600 ;
        RECT 2265.3200 1542.9200 2266.9200 1543.4000 ;
        RECT 2253.5600 1537.4800 2256.5600 1537.9600 ;
        RECT 2253.5600 1542.9200 2256.5600 1543.4000 ;
        RECT 2265.3200 1521.1600 2266.9200 1521.6400 ;
        RECT 2265.3200 1526.6000 2266.9200 1527.0800 ;
        RECT 2265.3200 1532.0400 2266.9200 1532.5200 ;
        RECT 2253.5600 1521.1600 2256.5600 1521.6400 ;
        RECT 2253.5600 1526.6000 2256.5600 1527.0800 ;
        RECT 2253.5600 1532.0400 2256.5600 1532.5200 ;
        RECT 2265.3200 1510.2800 2266.9200 1510.7600 ;
        RECT 2265.3200 1515.7200 2266.9200 1516.2000 ;
        RECT 2253.5600 1510.2800 2256.5600 1510.7600 ;
        RECT 2253.5600 1515.7200 2256.5600 1516.2000 ;
        RECT 2355.3200 1493.9600 2356.9200 1494.4400 ;
        RECT 2355.3200 1499.4000 2356.9200 1499.8800 ;
        RECT 2355.3200 1504.8400 2356.9200 1505.3200 ;
        RECT 2355.3200 1483.0800 2356.9200 1483.5600 ;
        RECT 2355.3200 1488.5200 2356.9200 1489.0000 ;
        RECT 2310.3200 1493.9600 2311.9200 1494.4400 ;
        RECT 2310.3200 1499.4000 2311.9200 1499.8800 ;
        RECT 2310.3200 1504.8400 2311.9200 1505.3200 ;
        RECT 2310.3200 1483.0800 2311.9200 1483.5600 ;
        RECT 2310.3200 1488.5200 2311.9200 1489.0000 ;
        RECT 2355.3200 1466.7600 2356.9200 1467.2400 ;
        RECT 2355.3200 1472.2000 2356.9200 1472.6800 ;
        RECT 2355.3200 1477.6400 2356.9200 1478.1200 ;
        RECT 2355.3200 1461.3200 2356.9200 1461.8000 ;
        RECT 2310.3200 1466.7600 2311.9200 1467.2400 ;
        RECT 2310.3200 1472.2000 2311.9200 1472.6800 ;
        RECT 2310.3200 1477.6400 2311.9200 1478.1200 ;
        RECT 2310.3200 1461.3200 2311.9200 1461.8000 ;
        RECT 2265.3200 1493.9600 2266.9200 1494.4400 ;
        RECT 2265.3200 1499.4000 2266.9200 1499.8800 ;
        RECT 2265.3200 1504.8400 2266.9200 1505.3200 ;
        RECT 2253.5600 1493.9600 2256.5600 1494.4400 ;
        RECT 2253.5600 1499.4000 2256.5600 1499.8800 ;
        RECT 2253.5600 1504.8400 2256.5600 1505.3200 ;
        RECT 2265.3200 1483.0800 2266.9200 1483.5600 ;
        RECT 2265.3200 1488.5200 2266.9200 1489.0000 ;
        RECT 2253.5600 1483.0800 2256.5600 1483.5600 ;
        RECT 2253.5600 1488.5200 2256.5600 1489.0000 ;
        RECT 2265.3200 1466.7600 2266.9200 1467.2400 ;
        RECT 2265.3200 1472.2000 2266.9200 1472.6800 ;
        RECT 2265.3200 1477.6400 2266.9200 1478.1200 ;
        RECT 2253.5600 1466.7600 2256.5600 1467.2400 ;
        RECT 2253.5600 1472.2000 2256.5600 1472.6800 ;
        RECT 2253.5600 1477.6400 2256.5600 1478.1200 ;
        RECT 2253.5600 1461.3200 2256.5600 1461.8000 ;
        RECT 2265.3200 1461.3200 2266.9200 1461.8000 ;
        RECT 2253.5600 1666.2300 2460.6600 1669.2300 ;
        RECT 2253.5600 1453.1300 2460.6600 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 1223.4900 2446.9200 1439.5900 ;
        RECT 2400.3200 1223.4900 2401.9200 1439.5900 ;
        RECT 2355.3200 1223.4900 2356.9200 1439.5900 ;
        RECT 2310.3200 1223.4900 2311.9200 1439.5900 ;
        RECT 2265.3200 1223.4900 2266.9200 1439.5900 ;
        RECT 2457.6600 1223.4900 2460.6600 1439.5900 ;
        RECT 2253.5600 1223.4900 2256.5600 1439.5900 ;
      LAYER met3 ;
        RECT 2457.6600 1416.6400 2460.6600 1417.1200 ;
        RECT 2457.6600 1422.0800 2460.6600 1422.5600 ;
        RECT 2445.3200 1416.6400 2446.9200 1417.1200 ;
        RECT 2445.3200 1422.0800 2446.9200 1422.5600 ;
        RECT 2457.6600 1427.5200 2460.6600 1428.0000 ;
        RECT 2445.3200 1427.5200 2446.9200 1428.0000 ;
        RECT 2457.6600 1405.7600 2460.6600 1406.2400 ;
        RECT 2457.6600 1411.2000 2460.6600 1411.6800 ;
        RECT 2445.3200 1405.7600 2446.9200 1406.2400 ;
        RECT 2445.3200 1411.2000 2446.9200 1411.6800 ;
        RECT 2457.6600 1389.4400 2460.6600 1389.9200 ;
        RECT 2457.6600 1394.8800 2460.6600 1395.3600 ;
        RECT 2445.3200 1389.4400 2446.9200 1389.9200 ;
        RECT 2445.3200 1394.8800 2446.9200 1395.3600 ;
        RECT 2457.6600 1400.3200 2460.6600 1400.8000 ;
        RECT 2445.3200 1400.3200 2446.9200 1400.8000 ;
        RECT 2400.3200 1416.6400 2401.9200 1417.1200 ;
        RECT 2400.3200 1422.0800 2401.9200 1422.5600 ;
        RECT 2400.3200 1427.5200 2401.9200 1428.0000 ;
        RECT 2400.3200 1405.7600 2401.9200 1406.2400 ;
        RECT 2400.3200 1411.2000 2401.9200 1411.6800 ;
        RECT 2400.3200 1389.4400 2401.9200 1389.9200 ;
        RECT 2400.3200 1394.8800 2401.9200 1395.3600 ;
        RECT 2400.3200 1400.3200 2401.9200 1400.8000 ;
        RECT 2457.6600 1373.1200 2460.6600 1373.6000 ;
        RECT 2457.6600 1378.5600 2460.6600 1379.0400 ;
        RECT 2457.6600 1384.0000 2460.6600 1384.4800 ;
        RECT 2445.3200 1373.1200 2446.9200 1373.6000 ;
        RECT 2445.3200 1378.5600 2446.9200 1379.0400 ;
        RECT 2445.3200 1384.0000 2446.9200 1384.4800 ;
        RECT 2457.6600 1362.2400 2460.6600 1362.7200 ;
        RECT 2457.6600 1367.6800 2460.6600 1368.1600 ;
        RECT 2445.3200 1362.2400 2446.9200 1362.7200 ;
        RECT 2445.3200 1367.6800 2446.9200 1368.1600 ;
        RECT 2457.6600 1345.9200 2460.6600 1346.4000 ;
        RECT 2457.6600 1351.3600 2460.6600 1351.8400 ;
        RECT 2457.6600 1356.8000 2460.6600 1357.2800 ;
        RECT 2445.3200 1345.9200 2446.9200 1346.4000 ;
        RECT 2445.3200 1351.3600 2446.9200 1351.8400 ;
        RECT 2445.3200 1356.8000 2446.9200 1357.2800 ;
        RECT 2457.6600 1335.0400 2460.6600 1335.5200 ;
        RECT 2457.6600 1340.4800 2460.6600 1340.9600 ;
        RECT 2445.3200 1335.0400 2446.9200 1335.5200 ;
        RECT 2445.3200 1340.4800 2446.9200 1340.9600 ;
        RECT 2400.3200 1373.1200 2401.9200 1373.6000 ;
        RECT 2400.3200 1378.5600 2401.9200 1379.0400 ;
        RECT 2400.3200 1384.0000 2401.9200 1384.4800 ;
        RECT 2400.3200 1362.2400 2401.9200 1362.7200 ;
        RECT 2400.3200 1367.6800 2401.9200 1368.1600 ;
        RECT 2400.3200 1345.9200 2401.9200 1346.4000 ;
        RECT 2400.3200 1351.3600 2401.9200 1351.8400 ;
        RECT 2400.3200 1356.8000 2401.9200 1357.2800 ;
        RECT 2400.3200 1335.0400 2401.9200 1335.5200 ;
        RECT 2400.3200 1340.4800 2401.9200 1340.9600 ;
        RECT 2355.3200 1416.6400 2356.9200 1417.1200 ;
        RECT 2355.3200 1422.0800 2356.9200 1422.5600 ;
        RECT 2355.3200 1427.5200 2356.9200 1428.0000 ;
        RECT 2310.3200 1416.6400 2311.9200 1417.1200 ;
        RECT 2310.3200 1422.0800 2311.9200 1422.5600 ;
        RECT 2310.3200 1427.5200 2311.9200 1428.0000 ;
        RECT 2355.3200 1405.7600 2356.9200 1406.2400 ;
        RECT 2355.3200 1411.2000 2356.9200 1411.6800 ;
        RECT 2355.3200 1389.4400 2356.9200 1389.9200 ;
        RECT 2355.3200 1394.8800 2356.9200 1395.3600 ;
        RECT 2355.3200 1400.3200 2356.9200 1400.8000 ;
        RECT 2310.3200 1405.7600 2311.9200 1406.2400 ;
        RECT 2310.3200 1411.2000 2311.9200 1411.6800 ;
        RECT 2310.3200 1389.4400 2311.9200 1389.9200 ;
        RECT 2310.3200 1394.8800 2311.9200 1395.3600 ;
        RECT 2310.3200 1400.3200 2311.9200 1400.8000 ;
        RECT 2265.3200 1416.6400 2266.9200 1417.1200 ;
        RECT 2265.3200 1422.0800 2266.9200 1422.5600 ;
        RECT 2253.5600 1422.0800 2256.5600 1422.5600 ;
        RECT 2253.5600 1416.6400 2256.5600 1417.1200 ;
        RECT 2253.5600 1427.5200 2256.5600 1428.0000 ;
        RECT 2265.3200 1427.5200 2266.9200 1428.0000 ;
        RECT 2265.3200 1405.7600 2266.9200 1406.2400 ;
        RECT 2265.3200 1411.2000 2266.9200 1411.6800 ;
        RECT 2253.5600 1411.2000 2256.5600 1411.6800 ;
        RECT 2253.5600 1405.7600 2256.5600 1406.2400 ;
        RECT 2265.3200 1389.4400 2266.9200 1389.9200 ;
        RECT 2265.3200 1394.8800 2266.9200 1395.3600 ;
        RECT 2253.5600 1394.8800 2256.5600 1395.3600 ;
        RECT 2253.5600 1389.4400 2256.5600 1389.9200 ;
        RECT 2253.5600 1400.3200 2256.5600 1400.8000 ;
        RECT 2265.3200 1400.3200 2266.9200 1400.8000 ;
        RECT 2355.3200 1373.1200 2356.9200 1373.6000 ;
        RECT 2355.3200 1378.5600 2356.9200 1379.0400 ;
        RECT 2355.3200 1384.0000 2356.9200 1384.4800 ;
        RECT 2355.3200 1362.2400 2356.9200 1362.7200 ;
        RECT 2355.3200 1367.6800 2356.9200 1368.1600 ;
        RECT 2310.3200 1373.1200 2311.9200 1373.6000 ;
        RECT 2310.3200 1378.5600 2311.9200 1379.0400 ;
        RECT 2310.3200 1384.0000 2311.9200 1384.4800 ;
        RECT 2310.3200 1362.2400 2311.9200 1362.7200 ;
        RECT 2310.3200 1367.6800 2311.9200 1368.1600 ;
        RECT 2355.3200 1345.9200 2356.9200 1346.4000 ;
        RECT 2355.3200 1351.3600 2356.9200 1351.8400 ;
        RECT 2355.3200 1356.8000 2356.9200 1357.2800 ;
        RECT 2355.3200 1335.0400 2356.9200 1335.5200 ;
        RECT 2355.3200 1340.4800 2356.9200 1340.9600 ;
        RECT 2310.3200 1345.9200 2311.9200 1346.4000 ;
        RECT 2310.3200 1351.3600 2311.9200 1351.8400 ;
        RECT 2310.3200 1356.8000 2311.9200 1357.2800 ;
        RECT 2310.3200 1335.0400 2311.9200 1335.5200 ;
        RECT 2310.3200 1340.4800 2311.9200 1340.9600 ;
        RECT 2265.3200 1373.1200 2266.9200 1373.6000 ;
        RECT 2265.3200 1378.5600 2266.9200 1379.0400 ;
        RECT 2265.3200 1384.0000 2266.9200 1384.4800 ;
        RECT 2253.5600 1373.1200 2256.5600 1373.6000 ;
        RECT 2253.5600 1378.5600 2256.5600 1379.0400 ;
        RECT 2253.5600 1384.0000 2256.5600 1384.4800 ;
        RECT 2265.3200 1362.2400 2266.9200 1362.7200 ;
        RECT 2265.3200 1367.6800 2266.9200 1368.1600 ;
        RECT 2253.5600 1362.2400 2256.5600 1362.7200 ;
        RECT 2253.5600 1367.6800 2256.5600 1368.1600 ;
        RECT 2265.3200 1345.9200 2266.9200 1346.4000 ;
        RECT 2265.3200 1351.3600 2266.9200 1351.8400 ;
        RECT 2265.3200 1356.8000 2266.9200 1357.2800 ;
        RECT 2253.5600 1345.9200 2256.5600 1346.4000 ;
        RECT 2253.5600 1351.3600 2256.5600 1351.8400 ;
        RECT 2253.5600 1356.8000 2256.5600 1357.2800 ;
        RECT 2265.3200 1335.0400 2266.9200 1335.5200 ;
        RECT 2265.3200 1340.4800 2266.9200 1340.9600 ;
        RECT 2253.5600 1335.0400 2256.5600 1335.5200 ;
        RECT 2253.5600 1340.4800 2256.5600 1340.9600 ;
        RECT 2457.6600 1318.7200 2460.6600 1319.2000 ;
        RECT 2457.6600 1324.1600 2460.6600 1324.6400 ;
        RECT 2457.6600 1329.6000 2460.6600 1330.0800 ;
        RECT 2445.3200 1318.7200 2446.9200 1319.2000 ;
        RECT 2445.3200 1324.1600 2446.9200 1324.6400 ;
        RECT 2445.3200 1329.6000 2446.9200 1330.0800 ;
        RECT 2457.6600 1307.8400 2460.6600 1308.3200 ;
        RECT 2457.6600 1313.2800 2460.6600 1313.7600 ;
        RECT 2445.3200 1307.8400 2446.9200 1308.3200 ;
        RECT 2445.3200 1313.2800 2446.9200 1313.7600 ;
        RECT 2457.6600 1291.5200 2460.6600 1292.0000 ;
        RECT 2457.6600 1296.9600 2460.6600 1297.4400 ;
        RECT 2457.6600 1302.4000 2460.6600 1302.8800 ;
        RECT 2445.3200 1291.5200 2446.9200 1292.0000 ;
        RECT 2445.3200 1296.9600 2446.9200 1297.4400 ;
        RECT 2445.3200 1302.4000 2446.9200 1302.8800 ;
        RECT 2457.6600 1280.6400 2460.6600 1281.1200 ;
        RECT 2457.6600 1286.0800 2460.6600 1286.5600 ;
        RECT 2445.3200 1280.6400 2446.9200 1281.1200 ;
        RECT 2445.3200 1286.0800 2446.9200 1286.5600 ;
        RECT 2400.3200 1318.7200 2401.9200 1319.2000 ;
        RECT 2400.3200 1324.1600 2401.9200 1324.6400 ;
        RECT 2400.3200 1329.6000 2401.9200 1330.0800 ;
        RECT 2400.3200 1307.8400 2401.9200 1308.3200 ;
        RECT 2400.3200 1313.2800 2401.9200 1313.7600 ;
        RECT 2400.3200 1291.5200 2401.9200 1292.0000 ;
        RECT 2400.3200 1296.9600 2401.9200 1297.4400 ;
        RECT 2400.3200 1302.4000 2401.9200 1302.8800 ;
        RECT 2400.3200 1280.6400 2401.9200 1281.1200 ;
        RECT 2400.3200 1286.0800 2401.9200 1286.5600 ;
        RECT 2457.6600 1264.3200 2460.6600 1264.8000 ;
        RECT 2457.6600 1269.7600 2460.6600 1270.2400 ;
        RECT 2457.6600 1275.2000 2460.6600 1275.6800 ;
        RECT 2445.3200 1264.3200 2446.9200 1264.8000 ;
        RECT 2445.3200 1269.7600 2446.9200 1270.2400 ;
        RECT 2445.3200 1275.2000 2446.9200 1275.6800 ;
        RECT 2457.6600 1253.4400 2460.6600 1253.9200 ;
        RECT 2457.6600 1258.8800 2460.6600 1259.3600 ;
        RECT 2445.3200 1253.4400 2446.9200 1253.9200 ;
        RECT 2445.3200 1258.8800 2446.9200 1259.3600 ;
        RECT 2457.6600 1237.1200 2460.6600 1237.6000 ;
        RECT 2457.6600 1242.5600 2460.6600 1243.0400 ;
        RECT 2457.6600 1248.0000 2460.6600 1248.4800 ;
        RECT 2445.3200 1237.1200 2446.9200 1237.6000 ;
        RECT 2445.3200 1242.5600 2446.9200 1243.0400 ;
        RECT 2445.3200 1248.0000 2446.9200 1248.4800 ;
        RECT 2457.6600 1231.6800 2460.6600 1232.1600 ;
        RECT 2445.3200 1231.6800 2446.9200 1232.1600 ;
        RECT 2400.3200 1264.3200 2401.9200 1264.8000 ;
        RECT 2400.3200 1269.7600 2401.9200 1270.2400 ;
        RECT 2400.3200 1275.2000 2401.9200 1275.6800 ;
        RECT 2400.3200 1253.4400 2401.9200 1253.9200 ;
        RECT 2400.3200 1258.8800 2401.9200 1259.3600 ;
        RECT 2400.3200 1237.1200 2401.9200 1237.6000 ;
        RECT 2400.3200 1242.5600 2401.9200 1243.0400 ;
        RECT 2400.3200 1248.0000 2401.9200 1248.4800 ;
        RECT 2400.3200 1231.6800 2401.9200 1232.1600 ;
        RECT 2355.3200 1318.7200 2356.9200 1319.2000 ;
        RECT 2355.3200 1324.1600 2356.9200 1324.6400 ;
        RECT 2355.3200 1329.6000 2356.9200 1330.0800 ;
        RECT 2355.3200 1307.8400 2356.9200 1308.3200 ;
        RECT 2355.3200 1313.2800 2356.9200 1313.7600 ;
        RECT 2310.3200 1318.7200 2311.9200 1319.2000 ;
        RECT 2310.3200 1324.1600 2311.9200 1324.6400 ;
        RECT 2310.3200 1329.6000 2311.9200 1330.0800 ;
        RECT 2310.3200 1307.8400 2311.9200 1308.3200 ;
        RECT 2310.3200 1313.2800 2311.9200 1313.7600 ;
        RECT 2355.3200 1291.5200 2356.9200 1292.0000 ;
        RECT 2355.3200 1296.9600 2356.9200 1297.4400 ;
        RECT 2355.3200 1302.4000 2356.9200 1302.8800 ;
        RECT 2355.3200 1280.6400 2356.9200 1281.1200 ;
        RECT 2355.3200 1286.0800 2356.9200 1286.5600 ;
        RECT 2310.3200 1291.5200 2311.9200 1292.0000 ;
        RECT 2310.3200 1296.9600 2311.9200 1297.4400 ;
        RECT 2310.3200 1302.4000 2311.9200 1302.8800 ;
        RECT 2310.3200 1280.6400 2311.9200 1281.1200 ;
        RECT 2310.3200 1286.0800 2311.9200 1286.5600 ;
        RECT 2265.3200 1318.7200 2266.9200 1319.2000 ;
        RECT 2265.3200 1324.1600 2266.9200 1324.6400 ;
        RECT 2265.3200 1329.6000 2266.9200 1330.0800 ;
        RECT 2253.5600 1318.7200 2256.5600 1319.2000 ;
        RECT 2253.5600 1324.1600 2256.5600 1324.6400 ;
        RECT 2253.5600 1329.6000 2256.5600 1330.0800 ;
        RECT 2265.3200 1307.8400 2266.9200 1308.3200 ;
        RECT 2265.3200 1313.2800 2266.9200 1313.7600 ;
        RECT 2253.5600 1307.8400 2256.5600 1308.3200 ;
        RECT 2253.5600 1313.2800 2256.5600 1313.7600 ;
        RECT 2265.3200 1291.5200 2266.9200 1292.0000 ;
        RECT 2265.3200 1296.9600 2266.9200 1297.4400 ;
        RECT 2265.3200 1302.4000 2266.9200 1302.8800 ;
        RECT 2253.5600 1291.5200 2256.5600 1292.0000 ;
        RECT 2253.5600 1296.9600 2256.5600 1297.4400 ;
        RECT 2253.5600 1302.4000 2256.5600 1302.8800 ;
        RECT 2265.3200 1280.6400 2266.9200 1281.1200 ;
        RECT 2265.3200 1286.0800 2266.9200 1286.5600 ;
        RECT 2253.5600 1280.6400 2256.5600 1281.1200 ;
        RECT 2253.5600 1286.0800 2256.5600 1286.5600 ;
        RECT 2355.3200 1264.3200 2356.9200 1264.8000 ;
        RECT 2355.3200 1269.7600 2356.9200 1270.2400 ;
        RECT 2355.3200 1275.2000 2356.9200 1275.6800 ;
        RECT 2355.3200 1253.4400 2356.9200 1253.9200 ;
        RECT 2355.3200 1258.8800 2356.9200 1259.3600 ;
        RECT 2310.3200 1264.3200 2311.9200 1264.8000 ;
        RECT 2310.3200 1269.7600 2311.9200 1270.2400 ;
        RECT 2310.3200 1275.2000 2311.9200 1275.6800 ;
        RECT 2310.3200 1253.4400 2311.9200 1253.9200 ;
        RECT 2310.3200 1258.8800 2311.9200 1259.3600 ;
        RECT 2355.3200 1237.1200 2356.9200 1237.6000 ;
        RECT 2355.3200 1242.5600 2356.9200 1243.0400 ;
        RECT 2355.3200 1248.0000 2356.9200 1248.4800 ;
        RECT 2355.3200 1231.6800 2356.9200 1232.1600 ;
        RECT 2310.3200 1237.1200 2311.9200 1237.6000 ;
        RECT 2310.3200 1242.5600 2311.9200 1243.0400 ;
        RECT 2310.3200 1248.0000 2311.9200 1248.4800 ;
        RECT 2310.3200 1231.6800 2311.9200 1232.1600 ;
        RECT 2265.3200 1264.3200 2266.9200 1264.8000 ;
        RECT 2265.3200 1269.7600 2266.9200 1270.2400 ;
        RECT 2265.3200 1275.2000 2266.9200 1275.6800 ;
        RECT 2253.5600 1264.3200 2256.5600 1264.8000 ;
        RECT 2253.5600 1269.7600 2256.5600 1270.2400 ;
        RECT 2253.5600 1275.2000 2256.5600 1275.6800 ;
        RECT 2265.3200 1253.4400 2266.9200 1253.9200 ;
        RECT 2265.3200 1258.8800 2266.9200 1259.3600 ;
        RECT 2253.5600 1253.4400 2256.5600 1253.9200 ;
        RECT 2253.5600 1258.8800 2256.5600 1259.3600 ;
        RECT 2265.3200 1237.1200 2266.9200 1237.6000 ;
        RECT 2265.3200 1242.5600 2266.9200 1243.0400 ;
        RECT 2265.3200 1248.0000 2266.9200 1248.4800 ;
        RECT 2253.5600 1237.1200 2256.5600 1237.6000 ;
        RECT 2253.5600 1242.5600 2256.5600 1243.0400 ;
        RECT 2253.5600 1248.0000 2256.5600 1248.4800 ;
        RECT 2253.5600 1231.6800 2256.5600 1232.1600 ;
        RECT 2265.3200 1231.6800 2266.9200 1232.1600 ;
        RECT 2253.5600 1436.5900 2460.6600 1439.5900 ;
        RECT 2253.5600 1223.4900 2460.6600 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 993.8500 2446.9200 1209.9500 ;
        RECT 2400.3200 993.8500 2401.9200 1209.9500 ;
        RECT 2355.3200 993.8500 2356.9200 1209.9500 ;
        RECT 2310.3200 993.8500 2311.9200 1209.9500 ;
        RECT 2265.3200 993.8500 2266.9200 1209.9500 ;
        RECT 2457.6600 993.8500 2460.6600 1209.9500 ;
        RECT 2253.5600 993.8500 2256.5600 1209.9500 ;
      LAYER met3 ;
        RECT 2457.6600 1187.0000 2460.6600 1187.4800 ;
        RECT 2457.6600 1192.4400 2460.6600 1192.9200 ;
        RECT 2445.3200 1187.0000 2446.9200 1187.4800 ;
        RECT 2445.3200 1192.4400 2446.9200 1192.9200 ;
        RECT 2457.6600 1197.8800 2460.6600 1198.3600 ;
        RECT 2445.3200 1197.8800 2446.9200 1198.3600 ;
        RECT 2457.6600 1176.1200 2460.6600 1176.6000 ;
        RECT 2457.6600 1181.5600 2460.6600 1182.0400 ;
        RECT 2445.3200 1176.1200 2446.9200 1176.6000 ;
        RECT 2445.3200 1181.5600 2446.9200 1182.0400 ;
        RECT 2457.6600 1159.8000 2460.6600 1160.2800 ;
        RECT 2457.6600 1165.2400 2460.6600 1165.7200 ;
        RECT 2445.3200 1159.8000 2446.9200 1160.2800 ;
        RECT 2445.3200 1165.2400 2446.9200 1165.7200 ;
        RECT 2457.6600 1170.6800 2460.6600 1171.1600 ;
        RECT 2445.3200 1170.6800 2446.9200 1171.1600 ;
        RECT 2400.3200 1187.0000 2401.9200 1187.4800 ;
        RECT 2400.3200 1192.4400 2401.9200 1192.9200 ;
        RECT 2400.3200 1197.8800 2401.9200 1198.3600 ;
        RECT 2400.3200 1176.1200 2401.9200 1176.6000 ;
        RECT 2400.3200 1181.5600 2401.9200 1182.0400 ;
        RECT 2400.3200 1159.8000 2401.9200 1160.2800 ;
        RECT 2400.3200 1165.2400 2401.9200 1165.7200 ;
        RECT 2400.3200 1170.6800 2401.9200 1171.1600 ;
        RECT 2457.6600 1143.4800 2460.6600 1143.9600 ;
        RECT 2457.6600 1148.9200 2460.6600 1149.4000 ;
        RECT 2457.6600 1154.3600 2460.6600 1154.8400 ;
        RECT 2445.3200 1143.4800 2446.9200 1143.9600 ;
        RECT 2445.3200 1148.9200 2446.9200 1149.4000 ;
        RECT 2445.3200 1154.3600 2446.9200 1154.8400 ;
        RECT 2457.6600 1132.6000 2460.6600 1133.0800 ;
        RECT 2457.6600 1138.0400 2460.6600 1138.5200 ;
        RECT 2445.3200 1132.6000 2446.9200 1133.0800 ;
        RECT 2445.3200 1138.0400 2446.9200 1138.5200 ;
        RECT 2457.6600 1116.2800 2460.6600 1116.7600 ;
        RECT 2457.6600 1121.7200 2460.6600 1122.2000 ;
        RECT 2457.6600 1127.1600 2460.6600 1127.6400 ;
        RECT 2445.3200 1116.2800 2446.9200 1116.7600 ;
        RECT 2445.3200 1121.7200 2446.9200 1122.2000 ;
        RECT 2445.3200 1127.1600 2446.9200 1127.6400 ;
        RECT 2457.6600 1105.4000 2460.6600 1105.8800 ;
        RECT 2457.6600 1110.8400 2460.6600 1111.3200 ;
        RECT 2445.3200 1105.4000 2446.9200 1105.8800 ;
        RECT 2445.3200 1110.8400 2446.9200 1111.3200 ;
        RECT 2400.3200 1143.4800 2401.9200 1143.9600 ;
        RECT 2400.3200 1148.9200 2401.9200 1149.4000 ;
        RECT 2400.3200 1154.3600 2401.9200 1154.8400 ;
        RECT 2400.3200 1132.6000 2401.9200 1133.0800 ;
        RECT 2400.3200 1138.0400 2401.9200 1138.5200 ;
        RECT 2400.3200 1116.2800 2401.9200 1116.7600 ;
        RECT 2400.3200 1121.7200 2401.9200 1122.2000 ;
        RECT 2400.3200 1127.1600 2401.9200 1127.6400 ;
        RECT 2400.3200 1105.4000 2401.9200 1105.8800 ;
        RECT 2400.3200 1110.8400 2401.9200 1111.3200 ;
        RECT 2355.3200 1187.0000 2356.9200 1187.4800 ;
        RECT 2355.3200 1192.4400 2356.9200 1192.9200 ;
        RECT 2355.3200 1197.8800 2356.9200 1198.3600 ;
        RECT 2310.3200 1187.0000 2311.9200 1187.4800 ;
        RECT 2310.3200 1192.4400 2311.9200 1192.9200 ;
        RECT 2310.3200 1197.8800 2311.9200 1198.3600 ;
        RECT 2355.3200 1176.1200 2356.9200 1176.6000 ;
        RECT 2355.3200 1181.5600 2356.9200 1182.0400 ;
        RECT 2355.3200 1159.8000 2356.9200 1160.2800 ;
        RECT 2355.3200 1165.2400 2356.9200 1165.7200 ;
        RECT 2355.3200 1170.6800 2356.9200 1171.1600 ;
        RECT 2310.3200 1176.1200 2311.9200 1176.6000 ;
        RECT 2310.3200 1181.5600 2311.9200 1182.0400 ;
        RECT 2310.3200 1159.8000 2311.9200 1160.2800 ;
        RECT 2310.3200 1165.2400 2311.9200 1165.7200 ;
        RECT 2310.3200 1170.6800 2311.9200 1171.1600 ;
        RECT 2265.3200 1187.0000 2266.9200 1187.4800 ;
        RECT 2265.3200 1192.4400 2266.9200 1192.9200 ;
        RECT 2253.5600 1192.4400 2256.5600 1192.9200 ;
        RECT 2253.5600 1187.0000 2256.5600 1187.4800 ;
        RECT 2253.5600 1197.8800 2256.5600 1198.3600 ;
        RECT 2265.3200 1197.8800 2266.9200 1198.3600 ;
        RECT 2265.3200 1176.1200 2266.9200 1176.6000 ;
        RECT 2265.3200 1181.5600 2266.9200 1182.0400 ;
        RECT 2253.5600 1181.5600 2256.5600 1182.0400 ;
        RECT 2253.5600 1176.1200 2256.5600 1176.6000 ;
        RECT 2265.3200 1159.8000 2266.9200 1160.2800 ;
        RECT 2265.3200 1165.2400 2266.9200 1165.7200 ;
        RECT 2253.5600 1165.2400 2256.5600 1165.7200 ;
        RECT 2253.5600 1159.8000 2256.5600 1160.2800 ;
        RECT 2253.5600 1170.6800 2256.5600 1171.1600 ;
        RECT 2265.3200 1170.6800 2266.9200 1171.1600 ;
        RECT 2355.3200 1143.4800 2356.9200 1143.9600 ;
        RECT 2355.3200 1148.9200 2356.9200 1149.4000 ;
        RECT 2355.3200 1154.3600 2356.9200 1154.8400 ;
        RECT 2355.3200 1132.6000 2356.9200 1133.0800 ;
        RECT 2355.3200 1138.0400 2356.9200 1138.5200 ;
        RECT 2310.3200 1143.4800 2311.9200 1143.9600 ;
        RECT 2310.3200 1148.9200 2311.9200 1149.4000 ;
        RECT 2310.3200 1154.3600 2311.9200 1154.8400 ;
        RECT 2310.3200 1132.6000 2311.9200 1133.0800 ;
        RECT 2310.3200 1138.0400 2311.9200 1138.5200 ;
        RECT 2355.3200 1116.2800 2356.9200 1116.7600 ;
        RECT 2355.3200 1121.7200 2356.9200 1122.2000 ;
        RECT 2355.3200 1127.1600 2356.9200 1127.6400 ;
        RECT 2355.3200 1105.4000 2356.9200 1105.8800 ;
        RECT 2355.3200 1110.8400 2356.9200 1111.3200 ;
        RECT 2310.3200 1116.2800 2311.9200 1116.7600 ;
        RECT 2310.3200 1121.7200 2311.9200 1122.2000 ;
        RECT 2310.3200 1127.1600 2311.9200 1127.6400 ;
        RECT 2310.3200 1105.4000 2311.9200 1105.8800 ;
        RECT 2310.3200 1110.8400 2311.9200 1111.3200 ;
        RECT 2265.3200 1143.4800 2266.9200 1143.9600 ;
        RECT 2265.3200 1148.9200 2266.9200 1149.4000 ;
        RECT 2265.3200 1154.3600 2266.9200 1154.8400 ;
        RECT 2253.5600 1143.4800 2256.5600 1143.9600 ;
        RECT 2253.5600 1148.9200 2256.5600 1149.4000 ;
        RECT 2253.5600 1154.3600 2256.5600 1154.8400 ;
        RECT 2265.3200 1132.6000 2266.9200 1133.0800 ;
        RECT 2265.3200 1138.0400 2266.9200 1138.5200 ;
        RECT 2253.5600 1132.6000 2256.5600 1133.0800 ;
        RECT 2253.5600 1138.0400 2256.5600 1138.5200 ;
        RECT 2265.3200 1116.2800 2266.9200 1116.7600 ;
        RECT 2265.3200 1121.7200 2266.9200 1122.2000 ;
        RECT 2265.3200 1127.1600 2266.9200 1127.6400 ;
        RECT 2253.5600 1116.2800 2256.5600 1116.7600 ;
        RECT 2253.5600 1121.7200 2256.5600 1122.2000 ;
        RECT 2253.5600 1127.1600 2256.5600 1127.6400 ;
        RECT 2265.3200 1105.4000 2266.9200 1105.8800 ;
        RECT 2265.3200 1110.8400 2266.9200 1111.3200 ;
        RECT 2253.5600 1105.4000 2256.5600 1105.8800 ;
        RECT 2253.5600 1110.8400 2256.5600 1111.3200 ;
        RECT 2457.6600 1089.0800 2460.6600 1089.5600 ;
        RECT 2457.6600 1094.5200 2460.6600 1095.0000 ;
        RECT 2457.6600 1099.9600 2460.6600 1100.4400 ;
        RECT 2445.3200 1089.0800 2446.9200 1089.5600 ;
        RECT 2445.3200 1094.5200 2446.9200 1095.0000 ;
        RECT 2445.3200 1099.9600 2446.9200 1100.4400 ;
        RECT 2457.6600 1078.2000 2460.6600 1078.6800 ;
        RECT 2457.6600 1083.6400 2460.6600 1084.1200 ;
        RECT 2445.3200 1078.2000 2446.9200 1078.6800 ;
        RECT 2445.3200 1083.6400 2446.9200 1084.1200 ;
        RECT 2457.6600 1061.8800 2460.6600 1062.3600 ;
        RECT 2457.6600 1067.3200 2460.6600 1067.8000 ;
        RECT 2457.6600 1072.7600 2460.6600 1073.2400 ;
        RECT 2445.3200 1061.8800 2446.9200 1062.3600 ;
        RECT 2445.3200 1067.3200 2446.9200 1067.8000 ;
        RECT 2445.3200 1072.7600 2446.9200 1073.2400 ;
        RECT 2457.6600 1051.0000 2460.6600 1051.4800 ;
        RECT 2457.6600 1056.4400 2460.6600 1056.9200 ;
        RECT 2445.3200 1051.0000 2446.9200 1051.4800 ;
        RECT 2445.3200 1056.4400 2446.9200 1056.9200 ;
        RECT 2400.3200 1089.0800 2401.9200 1089.5600 ;
        RECT 2400.3200 1094.5200 2401.9200 1095.0000 ;
        RECT 2400.3200 1099.9600 2401.9200 1100.4400 ;
        RECT 2400.3200 1078.2000 2401.9200 1078.6800 ;
        RECT 2400.3200 1083.6400 2401.9200 1084.1200 ;
        RECT 2400.3200 1061.8800 2401.9200 1062.3600 ;
        RECT 2400.3200 1067.3200 2401.9200 1067.8000 ;
        RECT 2400.3200 1072.7600 2401.9200 1073.2400 ;
        RECT 2400.3200 1051.0000 2401.9200 1051.4800 ;
        RECT 2400.3200 1056.4400 2401.9200 1056.9200 ;
        RECT 2457.6600 1034.6800 2460.6600 1035.1600 ;
        RECT 2457.6600 1040.1200 2460.6600 1040.6000 ;
        RECT 2457.6600 1045.5600 2460.6600 1046.0400 ;
        RECT 2445.3200 1034.6800 2446.9200 1035.1600 ;
        RECT 2445.3200 1040.1200 2446.9200 1040.6000 ;
        RECT 2445.3200 1045.5600 2446.9200 1046.0400 ;
        RECT 2457.6600 1023.8000 2460.6600 1024.2800 ;
        RECT 2457.6600 1029.2400 2460.6600 1029.7200 ;
        RECT 2445.3200 1023.8000 2446.9200 1024.2800 ;
        RECT 2445.3200 1029.2400 2446.9200 1029.7200 ;
        RECT 2457.6600 1007.4800 2460.6600 1007.9600 ;
        RECT 2457.6600 1012.9200 2460.6600 1013.4000 ;
        RECT 2457.6600 1018.3600 2460.6600 1018.8400 ;
        RECT 2445.3200 1007.4800 2446.9200 1007.9600 ;
        RECT 2445.3200 1012.9200 2446.9200 1013.4000 ;
        RECT 2445.3200 1018.3600 2446.9200 1018.8400 ;
        RECT 2457.6600 1002.0400 2460.6600 1002.5200 ;
        RECT 2445.3200 1002.0400 2446.9200 1002.5200 ;
        RECT 2400.3200 1034.6800 2401.9200 1035.1600 ;
        RECT 2400.3200 1040.1200 2401.9200 1040.6000 ;
        RECT 2400.3200 1045.5600 2401.9200 1046.0400 ;
        RECT 2400.3200 1023.8000 2401.9200 1024.2800 ;
        RECT 2400.3200 1029.2400 2401.9200 1029.7200 ;
        RECT 2400.3200 1007.4800 2401.9200 1007.9600 ;
        RECT 2400.3200 1012.9200 2401.9200 1013.4000 ;
        RECT 2400.3200 1018.3600 2401.9200 1018.8400 ;
        RECT 2400.3200 1002.0400 2401.9200 1002.5200 ;
        RECT 2355.3200 1089.0800 2356.9200 1089.5600 ;
        RECT 2355.3200 1094.5200 2356.9200 1095.0000 ;
        RECT 2355.3200 1099.9600 2356.9200 1100.4400 ;
        RECT 2355.3200 1078.2000 2356.9200 1078.6800 ;
        RECT 2355.3200 1083.6400 2356.9200 1084.1200 ;
        RECT 2310.3200 1089.0800 2311.9200 1089.5600 ;
        RECT 2310.3200 1094.5200 2311.9200 1095.0000 ;
        RECT 2310.3200 1099.9600 2311.9200 1100.4400 ;
        RECT 2310.3200 1078.2000 2311.9200 1078.6800 ;
        RECT 2310.3200 1083.6400 2311.9200 1084.1200 ;
        RECT 2355.3200 1061.8800 2356.9200 1062.3600 ;
        RECT 2355.3200 1067.3200 2356.9200 1067.8000 ;
        RECT 2355.3200 1072.7600 2356.9200 1073.2400 ;
        RECT 2355.3200 1051.0000 2356.9200 1051.4800 ;
        RECT 2355.3200 1056.4400 2356.9200 1056.9200 ;
        RECT 2310.3200 1061.8800 2311.9200 1062.3600 ;
        RECT 2310.3200 1067.3200 2311.9200 1067.8000 ;
        RECT 2310.3200 1072.7600 2311.9200 1073.2400 ;
        RECT 2310.3200 1051.0000 2311.9200 1051.4800 ;
        RECT 2310.3200 1056.4400 2311.9200 1056.9200 ;
        RECT 2265.3200 1089.0800 2266.9200 1089.5600 ;
        RECT 2265.3200 1094.5200 2266.9200 1095.0000 ;
        RECT 2265.3200 1099.9600 2266.9200 1100.4400 ;
        RECT 2253.5600 1089.0800 2256.5600 1089.5600 ;
        RECT 2253.5600 1094.5200 2256.5600 1095.0000 ;
        RECT 2253.5600 1099.9600 2256.5600 1100.4400 ;
        RECT 2265.3200 1078.2000 2266.9200 1078.6800 ;
        RECT 2265.3200 1083.6400 2266.9200 1084.1200 ;
        RECT 2253.5600 1078.2000 2256.5600 1078.6800 ;
        RECT 2253.5600 1083.6400 2256.5600 1084.1200 ;
        RECT 2265.3200 1061.8800 2266.9200 1062.3600 ;
        RECT 2265.3200 1067.3200 2266.9200 1067.8000 ;
        RECT 2265.3200 1072.7600 2266.9200 1073.2400 ;
        RECT 2253.5600 1061.8800 2256.5600 1062.3600 ;
        RECT 2253.5600 1067.3200 2256.5600 1067.8000 ;
        RECT 2253.5600 1072.7600 2256.5600 1073.2400 ;
        RECT 2265.3200 1051.0000 2266.9200 1051.4800 ;
        RECT 2265.3200 1056.4400 2266.9200 1056.9200 ;
        RECT 2253.5600 1051.0000 2256.5600 1051.4800 ;
        RECT 2253.5600 1056.4400 2256.5600 1056.9200 ;
        RECT 2355.3200 1034.6800 2356.9200 1035.1600 ;
        RECT 2355.3200 1040.1200 2356.9200 1040.6000 ;
        RECT 2355.3200 1045.5600 2356.9200 1046.0400 ;
        RECT 2355.3200 1023.8000 2356.9200 1024.2800 ;
        RECT 2355.3200 1029.2400 2356.9200 1029.7200 ;
        RECT 2310.3200 1034.6800 2311.9200 1035.1600 ;
        RECT 2310.3200 1040.1200 2311.9200 1040.6000 ;
        RECT 2310.3200 1045.5600 2311.9200 1046.0400 ;
        RECT 2310.3200 1023.8000 2311.9200 1024.2800 ;
        RECT 2310.3200 1029.2400 2311.9200 1029.7200 ;
        RECT 2355.3200 1007.4800 2356.9200 1007.9600 ;
        RECT 2355.3200 1012.9200 2356.9200 1013.4000 ;
        RECT 2355.3200 1018.3600 2356.9200 1018.8400 ;
        RECT 2355.3200 1002.0400 2356.9200 1002.5200 ;
        RECT 2310.3200 1007.4800 2311.9200 1007.9600 ;
        RECT 2310.3200 1012.9200 2311.9200 1013.4000 ;
        RECT 2310.3200 1018.3600 2311.9200 1018.8400 ;
        RECT 2310.3200 1002.0400 2311.9200 1002.5200 ;
        RECT 2265.3200 1034.6800 2266.9200 1035.1600 ;
        RECT 2265.3200 1040.1200 2266.9200 1040.6000 ;
        RECT 2265.3200 1045.5600 2266.9200 1046.0400 ;
        RECT 2253.5600 1034.6800 2256.5600 1035.1600 ;
        RECT 2253.5600 1040.1200 2256.5600 1040.6000 ;
        RECT 2253.5600 1045.5600 2256.5600 1046.0400 ;
        RECT 2265.3200 1023.8000 2266.9200 1024.2800 ;
        RECT 2265.3200 1029.2400 2266.9200 1029.7200 ;
        RECT 2253.5600 1023.8000 2256.5600 1024.2800 ;
        RECT 2253.5600 1029.2400 2256.5600 1029.7200 ;
        RECT 2265.3200 1007.4800 2266.9200 1007.9600 ;
        RECT 2265.3200 1012.9200 2266.9200 1013.4000 ;
        RECT 2265.3200 1018.3600 2266.9200 1018.8400 ;
        RECT 2253.5600 1007.4800 2256.5600 1007.9600 ;
        RECT 2253.5600 1012.9200 2256.5600 1013.4000 ;
        RECT 2253.5600 1018.3600 2256.5600 1018.8400 ;
        RECT 2253.5600 1002.0400 2256.5600 1002.5200 ;
        RECT 2265.3200 1002.0400 2266.9200 1002.5200 ;
        RECT 2253.5600 1206.9500 2460.6600 1209.9500 ;
        RECT 2253.5600 993.8500 2460.6600 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2445.3200 764.2100 2446.9200 980.3100 ;
        RECT 2400.3200 764.2100 2401.9200 980.3100 ;
        RECT 2355.3200 764.2100 2356.9200 980.3100 ;
        RECT 2310.3200 764.2100 2311.9200 980.3100 ;
        RECT 2265.3200 764.2100 2266.9200 980.3100 ;
        RECT 2457.6600 764.2100 2460.6600 980.3100 ;
        RECT 2253.5600 764.2100 2256.5600 980.3100 ;
      LAYER met3 ;
        RECT 2457.6600 957.3600 2460.6600 957.8400 ;
        RECT 2457.6600 962.8000 2460.6600 963.2800 ;
        RECT 2445.3200 957.3600 2446.9200 957.8400 ;
        RECT 2445.3200 962.8000 2446.9200 963.2800 ;
        RECT 2457.6600 968.2400 2460.6600 968.7200 ;
        RECT 2445.3200 968.2400 2446.9200 968.7200 ;
        RECT 2457.6600 946.4800 2460.6600 946.9600 ;
        RECT 2457.6600 951.9200 2460.6600 952.4000 ;
        RECT 2445.3200 946.4800 2446.9200 946.9600 ;
        RECT 2445.3200 951.9200 2446.9200 952.4000 ;
        RECT 2457.6600 930.1600 2460.6600 930.6400 ;
        RECT 2457.6600 935.6000 2460.6600 936.0800 ;
        RECT 2445.3200 930.1600 2446.9200 930.6400 ;
        RECT 2445.3200 935.6000 2446.9200 936.0800 ;
        RECT 2457.6600 941.0400 2460.6600 941.5200 ;
        RECT 2445.3200 941.0400 2446.9200 941.5200 ;
        RECT 2400.3200 957.3600 2401.9200 957.8400 ;
        RECT 2400.3200 962.8000 2401.9200 963.2800 ;
        RECT 2400.3200 968.2400 2401.9200 968.7200 ;
        RECT 2400.3200 946.4800 2401.9200 946.9600 ;
        RECT 2400.3200 951.9200 2401.9200 952.4000 ;
        RECT 2400.3200 930.1600 2401.9200 930.6400 ;
        RECT 2400.3200 935.6000 2401.9200 936.0800 ;
        RECT 2400.3200 941.0400 2401.9200 941.5200 ;
        RECT 2457.6600 913.8400 2460.6600 914.3200 ;
        RECT 2457.6600 919.2800 2460.6600 919.7600 ;
        RECT 2457.6600 924.7200 2460.6600 925.2000 ;
        RECT 2445.3200 913.8400 2446.9200 914.3200 ;
        RECT 2445.3200 919.2800 2446.9200 919.7600 ;
        RECT 2445.3200 924.7200 2446.9200 925.2000 ;
        RECT 2457.6600 902.9600 2460.6600 903.4400 ;
        RECT 2457.6600 908.4000 2460.6600 908.8800 ;
        RECT 2445.3200 902.9600 2446.9200 903.4400 ;
        RECT 2445.3200 908.4000 2446.9200 908.8800 ;
        RECT 2457.6600 886.6400 2460.6600 887.1200 ;
        RECT 2457.6600 892.0800 2460.6600 892.5600 ;
        RECT 2457.6600 897.5200 2460.6600 898.0000 ;
        RECT 2445.3200 886.6400 2446.9200 887.1200 ;
        RECT 2445.3200 892.0800 2446.9200 892.5600 ;
        RECT 2445.3200 897.5200 2446.9200 898.0000 ;
        RECT 2457.6600 875.7600 2460.6600 876.2400 ;
        RECT 2457.6600 881.2000 2460.6600 881.6800 ;
        RECT 2445.3200 875.7600 2446.9200 876.2400 ;
        RECT 2445.3200 881.2000 2446.9200 881.6800 ;
        RECT 2400.3200 913.8400 2401.9200 914.3200 ;
        RECT 2400.3200 919.2800 2401.9200 919.7600 ;
        RECT 2400.3200 924.7200 2401.9200 925.2000 ;
        RECT 2400.3200 902.9600 2401.9200 903.4400 ;
        RECT 2400.3200 908.4000 2401.9200 908.8800 ;
        RECT 2400.3200 886.6400 2401.9200 887.1200 ;
        RECT 2400.3200 892.0800 2401.9200 892.5600 ;
        RECT 2400.3200 897.5200 2401.9200 898.0000 ;
        RECT 2400.3200 875.7600 2401.9200 876.2400 ;
        RECT 2400.3200 881.2000 2401.9200 881.6800 ;
        RECT 2355.3200 957.3600 2356.9200 957.8400 ;
        RECT 2355.3200 962.8000 2356.9200 963.2800 ;
        RECT 2355.3200 968.2400 2356.9200 968.7200 ;
        RECT 2310.3200 957.3600 2311.9200 957.8400 ;
        RECT 2310.3200 962.8000 2311.9200 963.2800 ;
        RECT 2310.3200 968.2400 2311.9200 968.7200 ;
        RECT 2355.3200 946.4800 2356.9200 946.9600 ;
        RECT 2355.3200 951.9200 2356.9200 952.4000 ;
        RECT 2355.3200 930.1600 2356.9200 930.6400 ;
        RECT 2355.3200 935.6000 2356.9200 936.0800 ;
        RECT 2355.3200 941.0400 2356.9200 941.5200 ;
        RECT 2310.3200 946.4800 2311.9200 946.9600 ;
        RECT 2310.3200 951.9200 2311.9200 952.4000 ;
        RECT 2310.3200 930.1600 2311.9200 930.6400 ;
        RECT 2310.3200 935.6000 2311.9200 936.0800 ;
        RECT 2310.3200 941.0400 2311.9200 941.5200 ;
        RECT 2265.3200 957.3600 2266.9200 957.8400 ;
        RECT 2265.3200 962.8000 2266.9200 963.2800 ;
        RECT 2253.5600 962.8000 2256.5600 963.2800 ;
        RECT 2253.5600 957.3600 2256.5600 957.8400 ;
        RECT 2253.5600 968.2400 2256.5600 968.7200 ;
        RECT 2265.3200 968.2400 2266.9200 968.7200 ;
        RECT 2265.3200 946.4800 2266.9200 946.9600 ;
        RECT 2265.3200 951.9200 2266.9200 952.4000 ;
        RECT 2253.5600 951.9200 2256.5600 952.4000 ;
        RECT 2253.5600 946.4800 2256.5600 946.9600 ;
        RECT 2265.3200 930.1600 2266.9200 930.6400 ;
        RECT 2265.3200 935.6000 2266.9200 936.0800 ;
        RECT 2253.5600 935.6000 2256.5600 936.0800 ;
        RECT 2253.5600 930.1600 2256.5600 930.6400 ;
        RECT 2253.5600 941.0400 2256.5600 941.5200 ;
        RECT 2265.3200 941.0400 2266.9200 941.5200 ;
        RECT 2355.3200 913.8400 2356.9200 914.3200 ;
        RECT 2355.3200 919.2800 2356.9200 919.7600 ;
        RECT 2355.3200 924.7200 2356.9200 925.2000 ;
        RECT 2355.3200 902.9600 2356.9200 903.4400 ;
        RECT 2355.3200 908.4000 2356.9200 908.8800 ;
        RECT 2310.3200 913.8400 2311.9200 914.3200 ;
        RECT 2310.3200 919.2800 2311.9200 919.7600 ;
        RECT 2310.3200 924.7200 2311.9200 925.2000 ;
        RECT 2310.3200 902.9600 2311.9200 903.4400 ;
        RECT 2310.3200 908.4000 2311.9200 908.8800 ;
        RECT 2355.3200 886.6400 2356.9200 887.1200 ;
        RECT 2355.3200 892.0800 2356.9200 892.5600 ;
        RECT 2355.3200 897.5200 2356.9200 898.0000 ;
        RECT 2355.3200 875.7600 2356.9200 876.2400 ;
        RECT 2355.3200 881.2000 2356.9200 881.6800 ;
        RECT 2310.3200 886.6400 2311.9200 887.1200 ;
        RECT 2310.3200 892.0800 2311.9200 892.5600 ;
        RECT 2310.3200 897.5200 2311.9200 898.0000 ;
        RECT 2310.3200 875.7600 2311.9200 876.2400 ;
        RECT 2310.3200 881.2000 2311.9200 881.6800 ;
        RECT 2265.3200 913.8400 2266.9200 914.3200 ;
        RECT 2265.3200 919.2800 2266.9200 919.7600 ;
        RECT 2265.3200 924.7200 2266.9200 925.2000 ;
        RECT 2253.5600 913.8400 2256.5600 914.3200 ;
        RECT 2253.5600 919.2800 2256.5600 919.7600 ;
        RECT 2253.5600 924.7200 2256.5600 925.2000 ;
        RECT 2265.3200 902.9600 2266.9200 903.4400 ;
        RECT 2265.3200 908.4000 2266.9200 908.8800 ;
        RECT 2253.5600 902.9600 2256.5600 903.4400 ;
        RECT 2253.5600 908.4000 2256.5600 908.8800 ;
        RECT 2265.3200 886.6400 2266.9200 887.1200 ;
        RECT 2265.3200 892.0800 2266.9200 892.5600 ;
        RECT 2265.3200 897.5200 2266.9200 898.0000 ;
        RECT 2253.5600 886.6400 2256.5600 887.1200 ;
        RECT 2253.5600 892.0800 2256.5600 892.5600 ;
        RECT 2253.5600 897.5200 2256.5600 898.0000 ;
        RECT 2265.3200 875.7600 2266.9200 876.2400 ;
        RECT 2265.3200 881.2000 2266.9200 881.6800 ;
        RECT 2253.5600 875.7600 2256.5600 876.2400 ;
        RECT 2253.5600 881.2000 2256.5600 881.6800 ;
        RECT 2457.6600 859.4400 2460.6600 859.9200 ;
        RECT 2457.6600 864.8800 2460.6600 865.3600 ;
        RECT 2457.6600 870.3200 2460.6600 870.8000 ;
        RECT 2445.3200 859.4400 2446.9200 859.9200 ;
        RECT 2445.3200 864.8800 2446.9200 865.3600 ;
        RECT 2445.3200 870.3200 2446.9200 870.8000 ;
        RECT 2457.6600 848.5600 2460.6600 849.0400 ;
        RECT 2457.6600 854.0000 2460.6600 854.4800 ;
        RECT 2445.3200 848.5600 2446.9200 849.0400 ;
        RECT 2445.3200 854.0000 2446.9200 854.4800 ;
        RECT 2457.6600 832.2400 2460.6600 832.7200 ;
        RECT 2457.6600 837.6800 2460.6600 838.1600 ;
        RECT 2457.6600 843.1200 2460.6600 843.6000 ;
        RECT 2445.3200 832.2400 2446.9200 832.7200 ;
        RECT 2445.3200 837.6800 2446.9200 838.1600 ;
        RECT 2445.3200 843.1200 2446.9200 843.6000 ;
        RECT 2457.6600 821.3600 2460.6600 821.8400 ;
        RECT 2457.6600 826.8000 2460.6600 827.2800 ;
        RECT 2445.3200 821.3600 2446.9200 821.8400 ;
        RECT 2445.3200 826.8000 2446.9200 827.2800 ;
        RECT 2400.3200 859.4400 2401.9200 859.9200 ;
        RECT 2400.3200 864.8800 2401.9200 865.3600 ;
        RECT 2400.3200 870.3200 2401.9200 870.8000 ;
        RECT 2400.3200 848.5600 2401.9200 849.0400 ;
        RECT 2400.3200 854.0000 2401.9200 854.4800 ;
        RECT 2400.3200 832.2400 2401.9200 832.7200 ;
        RECT 2400.3200 837.6800 2401.9200 838.1600 ;
        RECT 2400.3200 843.1200 2401.9200 843.6000 ;
        RECT 2400.3200 821.3600 2401.9200 821.8400 ;
        RECT 2400.3200 826.8000 2401.9200 827.2800 ;
        RECT 2457.6600 805.0400 2460.6600 805.5200 ;
        RECT 2457.6600 810.4800 2460.6600 810.9600 ;
        RECT 2457.6600 815.9200 2460.6600 816.4000 ;
        RECT 2445.3200 805.0400 2446.9200 805.5200 ;
        RECT 2445.3200 810.4800 2446.9200 810.9600 ;
        RECT 2445.3200 815.9200 2446.9200 816.4000 ;
        RECT 2457.6600 794.1600 2460.6600 794.6400 ;
        RECT 2457.6600 799.6000 2460.6600 800.0800 ;
        RECT 2445.3200 794.1600 2446.9200 794.6400 ;
        RECT 2445.3200 799.6000 2446.9200 800.0800 ;
        RECT 2457.6600 777.8400 2460.6600 778.3200 ;
        RECT 2457.6600 783.2800 2460.6600 783.7600 ;
        RECT 2457.6600 788.7200 2460.6600 789.2000 ;
        RECT 2445.3200 777.8400 2446.9200 778.3200 ;
        RECT 2445.3200 783.2800 2446.9200 783.7600 ;
        RECT 2445.3200 788.7200 2446.9200 789.2000 ;
        RECT 2457.6600 772.4000 2460.6600 772.8800 ;
        RECT 2445.3200 772.4000 2446.9200 772.8800 ;
        RECT 2400.3200 805.0400 2401.9200 805.5200 ;
        RECT 2400.3200 810.4800 2401.9200 810.9600 ;
        RECT 2400.3200 815.9200 2401.9200 816.4000 ;
        RECT 2400.3200 794.1600 2401.9200 794.6400 ;
        RECT 2400.3200 799.6000 2401.9200 800.0800 ;
        RECT 2400.3200 777.8400 2401.9200 778.3200 ;
        RECT 2400.3200 783.2800 2401.9200 783.7600 ;
        RECT 2400.3200 788.7200 2401.9200 789.2000 ;
        RECT 2400.3200 772.4000 2401.9200 772.8800 ;
        RECT 2355.3200 859.4400 2356.9200 859.9200 ;
        RECT 2355.3200 864.8800 2356.9200 865.3600 ;
        RECT 2355.3200 870.3200 2356.9200 870.8000 ;
        RECT 2355.3200 848.5600 2356.9200 849.0400 ;
        RECT 2355.3200 854.0000 2356.9200 854.4800 ;
        RECT 2310.3200 859.4400 2311.9200 859.9200 ;
        RECT 2310.3200 864.8800 2311.9200 865.3600 ;
        RECT 2310.3200 870.3200 2311.9200 870.8000 ;
        RECT 2310.3200 848.5600 2311.9200 849.0400 ;
        RECT 2310.3200 854.0000 2311.9200 854.4800 ;
        RECT 2355.3200 832.2400 2356.9200 832.7200 ;
        RECT 2355.3200 837.6800 2356.9200 838.1600 ;
        RECT 2355.3200 843.1200 2356.9200 843.6000 ;
        RECT 2355.3200 821.3600 2356.9200 821.8400 ;
        RECT 2355.3200 826.8000 2356.9200 827.2800 ;
        RECT 2310.3200 832.2400 2311.9200 832.7200 ;
        RECT 2310.3200 837.6800 2311.9200 838.1600 ;
        RECT 2310.3200 843.1200 2311.9200 843.6000 ;
        RECT 2310.3200 821.3600 2311.9200 821.8400 ;
        RECT 2310.3200 826.8000 2311.9200 827.2800 ;
        RECT 2265.3200 859.4400 2266.9200 859.9200 ;
        RECT 2265.3200 864.8800 2266.9200 865.3600 ;
        RECT 2265.3200 870.3200 2266.9200 870.8000 ;
        RECT 2253.5600 859.4400 2256.5600 859.9200 ;
        RECT 2253.5600 864.8800 2256.5600 865.3600 ;
        RECT 2253.5600 870.3200 2256.5600 870.8000 ;
        RECT 2265.3200 848.5600 2266.9200 849.0400 ;
        RECT 2265.3200 854.0000 2266.9200 854.4800 ;
        RECT 2253.5600 848.5600 2256.5600 849.0400 ;
        RECT 2253.5600 854.0000 2256.5600 854.4800 ;
        RECT 2265.3200 832.2400 2266.9200 832.7200 ;
        RECT 2265.3200 837.6800 2266.9200 838.1600 ;
        RECT 2265.3200 843.1200 2266.9200 843.6000 ;
        RECT 2253.5600 832.2400 2256.5600 832.7200 ;
        RECT 2253.5600 837.6800 2256.5600 838.1600 ;
        RECT 2253.5600 843.1200 2256.5600 843.6000 ;
        RECT 2265.3200 821.3600 2266.9200 821.8400 ;
        RECT 2265.3200 826.8000 2266.9200 827.2800 ;
        RECT 2253.5600 821.3600 2256.5600 821.8400 ;
        RECT 2253.5600 826.8000 2256.5600 827.2800 ;
        RECT 2355.3200 805.0400 2356.9200 805.5200 ;
        RECT 2355.3200 810.4800 2356.9200 810.9600 ;
        RECT 2355.3200 815.9200 2356.9200 816.4000 ;
        RECT 2355.3200 794.1600 2356.9200 794.6400 ;
        RECT 2355.3200 799.6000 2356.9200 800.0800 ;
        RECT 2310.3200 805.0400 2311.9200 805.5200 ;
        RECT 2310.3200 810.4800 2311.9200 810.9600 ;
        RECT 2310.3200 815.9200 2311.9200 816.4000 ;
        RECT 2310.3200 794.1600 2311.9200 794.6400 ;
        RECT 2310.3200 799.6000 2311.9200 800.0800 ;
        RECT 2355.3200 777.8400 2356.9200 778.3200 ;
        RECT 2355.3200 783.2800 2356.9200 783.7600 ;
        RECT 2355.3200 788.7200 2356.9200 789.2000 ;
        RECT 2355.3200 772.4000 2356.9200 772.8800 ;
        RECT 2310.3200 777.8400 2311.9200 778.3200 ;
        RECT 2310.3200 783.2800 2311.9200 783.7600 ;
        RECT 2310.3200 788.7200 2311.9200 789.2000 ;
        RECT 2310.3200 772.4000 2311.9200 772.8800 ;
        RECT 2265.3200 805.0400 2266.9200 805.5200 ;
        RECT 2265.3200 810.4800 2266.9200 810.9600 ;
        RECT 2265.3200 815.9200 2266.9200 816.4000 ;
        RECT 2253.5600 805.0400 2256.5600 805.5200 ;
        RECT 2253.5600 810.4800 2256.5600 810.9600 ;
        RECT 2253.5600 815.9200 2256.5600 816.4000 ;
        RECT 2265.3200 794.1600 2266.9200 794.6400 ;
        RECT 2265.3200 799.6000 2266.9200 800.0800 ;
        RECT 2253.5600 794.1600 2256.5600 794.6400 ;
        RECT 2253.5600 799.6000 2256.5600 800.0800 ;
        RECT 2265.3200 777.8400 2266.9200 778.3200 ;
        RECT 2265.3200 783.2800 2266.9200 783.7600 ;
        RECT 2265.3200 788.7200 2266.9200 789.2000 ;
        RECT 2253.5600 777.8400 2256.5600 778.3200 ;
        RECT 2253.5600 783.2800 2256.5600 783.7600 ;
        RECT 2253.5600 788.7200 2256.5600 789.2000 ;
        RECT 2253.5600 772.4000 2256.5600 772.8800 ;
        RECT 2265.3200 772.4000 2266.9200 772.8800 ;
        RECT 2253.5600 977.3100 2460.6600 980.3100 ;
        RECT 2253.5600 764.2100 2460.6600 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 2474.7800 2830.6100 2476.7800 2857.5400 ;
        RECT 2677.8800 2830.6100 2679.8800 2857.5400 ;
      LAYER met3 ;
        RECT 2677.8800 2847.3200 2679.8800 2847.8000 ;
        RECT 2474.7800 2847.3200 2476.7800 2847.8000 ;
        RECT 2677.8800 2841.8800 2679.8800 2842.3600 ;
        RECT 2677.8800 2836.4400 2679.8800 2836.9200 ;
        RECT 2474.7800 2841.8800 2476.7800 2842.3600 ;
        RECT 2474.7800 2836.4400 2476.7800 2836.9200 ;
        RECT 2474.7800 2855.5400 2679.8800 2857.5400 ;
        RECT 2474.7800 2830.6100 2679.8800 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 534.5700 2667.1400 750.6700 ;
        RECT 2620.5400 534.5700 2622.1400 750.6700 ;
        RECT 2575.5400 534.5700 2577.1400 750.6700 ;
        RECT 2530.5400 534.5700 2532.1400 750.6700 ;
        RECT 2485.5400 534.5700 2487.1400 750.6700 ;
        RECT 2677.8800 534.5700 2680.8800 750.6700 ;
        RECT 2473.7800 534.5700 2476.7800 750.6700 ;
      LAYER met3 ;
        RECT 2677.8800 727.7200 2680.8800 728.2000 ;
        RECT 2677.8800 733.1600 2680.8800 733.6400 ;
        RECT 2665.5400 727.7200 2667.1400 728.2000 ;
        RECT 2665.5400 733.1600 2667.1400 733.6400 ;
        RECT 2677.8800 738.6000 2680.8800 739.0800 ;
        RECT 2665.5400 738.6000 2667.1400 739.0800 ;
        RECT 2677.8800 716.8400 2680.8800 717.3200 ;
        RECT 2677.8800 722.2800 2680.8800 722.7600 ;
        RECT 2665.5400 716.8400 2667.1400 717.3200 ;
        RECT 2665.5400 722.2800 2667.1400 722.7600 ;
        RECT 2677.8800 700.5200 2680.8800 701.0000 ;
        RECT 2677.8800 705.9600 2680.8800 706.4400 ;
        RECT 2665.5400 700.5200 2667.1400 701.0000 ;
        RECT 2665.5400 705.9600 2667.1400 706.4400 ;
        RECT 2677.8800 711.4000 2680.8800 711.8800 ;
        RECT 2665.5400 711.4000 2667.1400 711.8800 ;
        RECT 2620.5400 727.7200 2622.1400 728.2000 ;
        RECT 2620.5400 733.1600 2622.1400 733.6400 ;
        RECT 2620.5400 738.6000 2622.1400 739.0800 ;
        RECT 2620.5400 716.8400 2622.1400 717.3200 ;
        RECT 2620.5400 722.2800 2622.1400 722.7600 ;
        RECT 2620.5400 700.5200 2622.1400 701.0000 ;
        RECT 2620.5400 705.9600 2622.1400 706.4400 ;
        RECT 2620.5400 711.4000 2622.1400 711.8800 ;
        RECT 2677.8800 684.2000 2680.8800 684.6800 ;
        RECT 2677.8800 689.6400 2680.8800 690.1200 ;
        RECT 2677.8800 695.0800 2680.8800 695.5600 ;
        RECT 2665.5400 684.2000 2667.1400 684.6800 ;
        RECT 2665.5400 689.6400 2667.1400 690.1200 ;
        RECT 2665.5400 695.0800 2667.1400 695.5600 ;
        RECT 2677.8800 673.3200 2680.8800 673.8000 ;
        RECT 2677.8800 678.7600 2680.8800 679.2400 ;
        RECT 2665.5400 673.3200 2667.1400 673.8000 ;
        RECT 2665.5400 678.7600 2667.1400 679.2400 ;
        RECT 2677.8800 657.0000 2680.8800 657.4800 ;
        RECT 2677.8800 662.4400 2680.8800 662.9200 ;
        RECT 2677.8800 667.8800 2680.8800 668.3600 ;
        RECT 2665.5400 657.0000 2667.1400 657.4800 ;
        RECT 2665.5400 662.4400 2667.1400 662.9200 ;
        RECT 2665.5400 667.8800 2667.1400 668.3600 ;
        RECT 2677.8800 646.1200 2680.8800 646.6000 ;
        RECT 2677.8800 651.5600 2680.8800 652.0400 ;
        RECT 2665.5400 646.1200 2667.1400 646.6000 ;
        RECT 2665.5400 651.5600 2667.1400 652.0400 ;
        RECT 2620.5400 684.2000 2622.1400 684.6800 ;
        RECT 2620.5400 689.6400 2622.1400 690.1200 ;
        RECT 2620.5400 695.0800 2622.1400 695.5600 ;
        RECT 2620.5400 673.3200 2622.1400 673.8000 ;
        RECT 2620.5400 678.7600 2622.1400 679.2400 ;
        RECT 2620.5400 657.0000 2622.1400 657.4800 ;
        RECT 2620.5400 662.4400 2622.1400 662.9200 ;
        RECT 2620.5400 667.8800 2622.1400 668.3600 ;
        RECT 2620.5400 646.1200 2622.1400 646.6000 ;
        RECT 2620.5400 651.5600 2622.1400 652.0400 ;
        RECT 2575.5400 727.7200 2577.1400 728.2000 ;
        RECT 2575.5400 733.1600 2577.1400 733.6400 ;
        RECT 2575.5400 738.6000 2577.1400 739.0800 ;
        RECT 2530.5400 727.7200 2532.1400 728.2000 ;
        RECT 2530.5400 733.1600 2532.1400 733.6400 ;
        RECT 2530.5400 738.6000 2532.1400 739.0800 ;
        RECT 2575.5400 716.8400 2577.1400 717.3200 ;
        RECT 2575.5400 722.2800 2577.1400 722.7600 ;
        RECT 2575.5400 700.5200 2577.1400 701.0000 ;
        RECT 2575.5400 705.9600 2577.1400 706.4400 ;
        RECT 2575.5400 711.4000 2577.1400 711.8800 ;
        RECT 2530.5400 716.8400 2532.1400 717.3200 ;
        RECT 2530.5400 722.2800 2532.1400 722.7600 ;
        RECT 2530.5400 700.5200 2532.1400 701.0000 ;
        RECT 2530.5400 705.9600 2532.1400 706.4400 ;
        RECT 2530.5400 711.4000 2532.1400 711.8800 ;
        RECT 2485.5400 727.7200 2487.1400 728.2000 ;
        RECT 2485.5400 733.1600 2487.1400 733.6400 ;
        RECT 2473.7800 733.1600 2476.7800 733.6400 ;
        RECT 2473.7800 727.7200 2476.7800 728.2000 ;
        RECT 2473.7800 738.6000 2476.7800 739.0800 ;
        RECT 2485.5400 738.6000 2487.1400 739.0800 ;
        RECT 2485.5400 716.8400 2487.1400 717.3200 ;
        RECT 2485.5400 722.2800 2487.1400 722.7600 ;
        RECT 2473.7800 722.2800 2476.7800 722.7600 ;
        RECT 2473.7800 716.8400 2476.7800 717.3200 ;
        RECT 2485.5400 700.5200 2487.1400 701.0000 ;
        RECT 2485.5400 705.9600 2487.1400 706.4400 ;
        RECT 2473.7800 705.9600 2476.7800 706.4400 ;
        RECT 2473.7800 700.5200 2476.7800 701.0000 ;
        RECT 2473.7800 711.4000 2476.7800 711.8800 ;
        RECT 2485.5400 711.4000 2487.1400 711.8800 ;
        RECT 2575.5400 684.2000 2577.1400 684.6800 ;
        RECT 2575.5400 689.6400 2577.1400 690.1200 ;
        RECT 2575.5400 695.0800 2577.1400 695.5600 ;
        RECT 2575.5400 673.3200 2577.1400 673.8000 ;
        RECT 2575.5400 678.7600 2577.1400 679.2400 ;
        RECT 2530.5400 684.2000 2532.1400 684.6800 ;
        RECT 2530.5400 689.6400 2532.1400 690.1200 ;
        RECT 2530.5400 695.0800 2532.1400 695.5600 ;
        RECT 2530.5400 673.3200 2532.1400 673.8000 ;
        RECT 2530.5400 678.7600 2532.1400 679.2400 ;
        RECT 2575.5400 657.0000 2577.1400 657.4800 ;
        RECT 2575.5400 662.4400 2577.1400 662.9200 ;
        RECT 2575.5400 667.8800 2577.1400 668.3600 ;
        RECT 2575.5400 646.1200 2577.1400 646.6000 ;
        RECT 2575.5400 651.5600 2577.1400 652.0400 ;
        RECT 2530.5400 657.0000 2532.1400 657.4800 ;
        RECT 2530.5400 662.4400 2532.1400 662.9200 ;
        RECT 2530.5400 667.8800 2532.1400 668.3600 ;
        RECT 2530.5400 646.1200 2532.1400 646.6000 ;
        RECT 2530.5400 651.5600 2532.1400 652.0400 ;
        RECT 2485.5400 684.2000 2487.1400 684.6800 ;
        RECT 2485.5400 689.6400 2487.1400 690.1200 ;
        RECT 2485.5400 695.0800 2487.1400 695.5600 ;
        RECT 2473.7800 684.2000 2476.7800 684.6800 ;
        RECT 2473.7800 689.6400 2476.7800 690.1200 ;
        RECT 2473.7800 695.0800 2476.7800 695.5600 ;
        RECT 2485.5400 673.3200 2487.1400 673.8000 ;
        RECT 2485.5400 678.7600 2487.1400 679.2400 ;
        RECT 2473.7800 673.3200 2476.7800 673.8000 ;
        RECT 2473.7800 678.7600 2476.7800 679.2400 ;
        RECT 2485.5400 657.0000 2487.1400 657.4800 ;
        RECT 2485.5400 662.4400 2487.1400 662.9200 ;
        RECT 2485.5400 667.8800 2487.1400 668.3600 ;
        RECT 2473.7800 657.0000 2476.7800 657.4800 ;
        RECT 2473.7800 662.4400 2476.7800 662.9200 ;
        RECT 2473.7800 667.8800 2476.7800 668.3600 ;
        RECT 2485.5400 646.1200 2487.1400 646.6000 ;
        RECT 2485.5400 651.5600 2487.1400 652.0400 ;
        RECT 2473.7800 646.1200 2476.7800 646.6000 ;
        RECT 2473.7800 651.5600 2476.7800 652.0400 ;
        RECT 2677.8800 629.8000 2680.8800 630.2800 ;
        RECT 2677.8800 635.2400 2680.8800 635.7200 ;
        RECT 2677.8800 640.6800 2680.8800 641.1600 ;
        RECT 2665.5400 629.8000 2667.1400 630.2800 ;
        RECT 2665.5400 635.2400 2667.1400 635.7200 ;
        RECT 2665.5400 640.6800 2667.1400 641.1600 ;
        RECT 2677.8800 618.9200 2680.8800 619.4000 ;
        RECT 2677.8800 624.3600 2680.8800 624.8400 ;
        RECT 2665.5400 618.9200 2667.1400 619.4000 ;
        RECT 2665.5400 624.3600 2667.1400 624.8400 ;
        RECT 2677.8800 602.6000 2680.8800 603.0800 ;
        RECT 2677.8800 608.0400 2680.8800 608.5200 ;
        RECT 2677.8800 613.4800 2680.8800 613.9600 ;
        RECT 2665.5400 602.6000 2667.1400 603.0800 ;
        RECT 2665.5400 608.0400 2667.1400 608.5200 ;
        RECT 2665.5400 613.4800 2667.1400 613.9600 ;
        RECT 2677.8800 591.7200 2680.8800 592.2000 ;
        RECT 2677.8800 597.1600 2680.8800 597.6400 ;
        RECT 2665.5400 591.7200 2667.1400 592.2000 ;
        RECT 2665.5400 597.1600 2667.1400 597.6400 ;
        RECT 2620.5400 629.8000 2622.1400 630.2800 ;
        RECT 2620.5400 635.2400 2622.1400 635.7200 ;
        RECT 2620.5400 640.6800 2622.1400 641.1600 ;
        RECT 2620.5400 618.9200 2622.1400 619.4000 ;
        RECT 2620.5400 624.3600 2622.1400 624.8400 ;
        RECT 2620.5400 602.6000 2622.1400 603.0800 ;
        RECT 2620.5400 608.0400 2622.1400 608.5200 ;
        RECT 2620.5400 613.4800 2622.1400 613.9600 ;
        RECT 2620.5400 591.7200 2622.1400 592.2000 ;
        RECT 2620.5400 597.1600 2622.1400 597.6400 ;
        RECT 2677.8800 575.4000 2680.8800 575.8800 ;
        RECT 2677.8800 580.8400 2680.8800 581.3200 ;
        RECT 2677.8800 586.2800 2680.8800 586.7600 ;
        RECT 2665.5400 575.4000 2667.1400 575.8800 ;
        RECT 2665.5400 580.8400 2667.1400 581.3200 ;
        RECT 2665.5400 586.2800 2667.1400 586.7600 ;
        RECT 2677.8800 564.5200 2680.8800 565.0000 ;
        RECT 2677.8800 569.9600 2680.8800 570.4400 ;
        RECT 2665.5400 564.5200 2667.1400 565.0000 ;
        RECT 2665.5400 569.9600 2667.1400 570.4400 ;
        RECT 2677.8800 548.2000 2680.8800 548.6800 ;
        RECT 2677.8800 553.6400 2680.8800 554.1200 ;
        RECT 2677.8800 559.0800 2680.8800 559.5600 ;
        RECT 2665.5400 548.2000 2667.1400 548.6800 ;
        RECT 2665.5400 553.6400 2667.1400 554.1200 ;
        RECT 2665.5400 559.0800 2667.1400 559.5600 ;
        RECT 2677.8800 542.7600 2680.8800 543.2400 ;
        RECT 2665.5400 542.7600 2667.1400 543.2400 ;
        RECT 2620.5400 575.4000 2622.1400 575.8800 ;
        RECT 2620.5400 580.8400 2622.1400 581.3200 ;
        RECT 2620.5400 586.2800 2622.1400 586.7600 ;
        RECT 2620.5400 564.5200 2622.1400 565.0000 ;
        RECT 2620.5400 569.9600 2622.1400 570.4400 ;
        RECT 2620.5400 548.2000 2622.1400 548.6800 ;
        RECT 2620.5400 553.6400 2622.1400 554.1200 ;
        RECT 2620.5400 559.0800 2622.1400 559.5600 ;
        RECT 2620.5400 542.7600 2622.1400 543.2400 ;
        RECT 2575.5400 629.8000 2577.1400 630.2800 ;
        RECT 2575.5400 635.2400 2577.1400 635.7200 ;
        RECT 2575.5400 640.6800 2577.1400 641.1600 ;
        RECT 2575.5400 618.9200 2577.1400 619.4000 ;
        RECT 2575.5400 624.3600 2577.1400 624.8400 ;
        RECT 2530.5400 629.8000 2532.1400 630.2800 ;
        RECT 2530.5400 635.2400 2532.1400 635.7200 ;
        RECT 2530.5400 640.6800 2532.1400 641.1600 ;
        RECT 2530.5400 618.9200 2532.1400 619.4000 ;
        RECT 2530.5400 624.3600 2532.1400 624.8400 ;
        RECT 2575.5400 602.6000 2577.1400 603.0800 ;
        RECT 2575.5400 608.0400 2577.1400 608.5200 ;
        RECT 2575.5400 613.4800 2577.1400 613.9600 ;
        RECT 2575.5400 591.7200 2577.1400 592.2000 ;
        RECT 2575.5400 597.1600 2577.1400 597.6400 ;
        RECT 2530.5400 602.6000 2532.1400 603.0800 ;
        RECT 2530.5400 608.0400 2532.1400 608.5200 ;
        RECT 2530.5400 613.4800 2532.1400 613.9600 ;
        RECT 2530.5400 591.7200 2532.1400 592.2000 ;
        RECT 2530.5400 597.1600 2532.1400 597.6400 ;
        RECT 2485.5400 629.8000 2487.1400 630.2800 ;
        RECT 2485.5400 635.2400 2487.1400 635.7200 ;
        RECT 2485.5400 640.6800 2487.1400 641.1600 ;
        RECT 2473.7800 629.8000 2476.7800 630.2800 ;
        RECT 2473.7800 635.2400 2476.7800 635.7200 ;
        RECT 2473.7800 640.6800 2476.7800 641.1600 ;
        RECT 2485.5400 618.9200 2487.1400 619.4000 ;
        RECT 2485.5400 624.3600 2487.1400 624.8400 ;
        RECT 2473.7800 618.9200 2476.7800 619.4000 ;
        RECT 2473.7800 624.3600 2476.7800 624.8400 ;
        RECT 2485.5400 602.6000 2487.1400 603.0800 ;
        RECT 2485.5400 608.0400 2487.1400 608.5200 ;
        RECT 2485.5400 613.4800 2487.1400 613.9600 ;
        RECT 2473.7800 602.6000 2476.7800 603.0800 ;
        RECT 2473.7800 608.0400 2476.7800 608.5200 ;
        RECT 2473.7800 613.4800 2476.7800 613.9600 ;
        RECT 2485.5400 591.7200 2487.1400 592.2000 ;
        RECT 2485.5400 597.1600 2487.1400 597.6400 ;
        RECT 2473.7800 591.7200 2476.7800 592.2000 ;
        RECT 2473.7800 597.1600 2476.7800 597.6400 ;
        RECT 2575.5400 575.4000 2577.1400 575.8800 ;
        RECT 2575.5400 580.8400 2577.1400 581.3200 ;
        RECT 2575.5400 586.2800 2577.1400 586.7600 ;
        RECT 2575.5400 564.5200 2577.1400 565.0000 ;
        RECT 2575.5400 569.9600 2577.1400 570.4400 ;
        RECT 2530.5400 575.4000 2532.1400 575.8800 ;
        RECT 2530.5400 580.8400 2532.1400 581.3200 ;
        RECT 2530.5400 586.2800 2532.1400 586.7600 ;
        RECT 2530.5400 564.5200 2532.1400 565.0000 ;
        RECT 2530.5400 569.9600 2532.1400 570.4400 ;
        RECT 2575.5400 548.2000 2577.1400 548.6800 ;
        RECT 2575.5400 553.6400 2577.1400 554.1200 ;
        RECT 2575.5400 559.0800 2577.1400 559.5600 ;
        RECT 2575.5400 542.7600 2577.1400 543.2400 ;
        RECT 2530.5400 548.2000 2532.1400 548.6800 ;
        RECT 2530.5400 553.6400 2532.1400 554.1200 ;
        RECT 2530.5400 559.0800 2532.1400 559.5600 ;
        RECT 2530.5400 542.7600 2532.1400 543.2400 ;
        RECT 2485.5400 575.4000 2487.1400 575.8800 ;
        RECT 2485.5400 580.8400 2487.1400 581.3200 ;
        RECT 2485.5400 586.2800 2487.1400 586.7600 ;
        RECT 2473.7800 575.4000 2476.7800 575.8800 ;
        RECT 2473.7800 580.8400 2476.7800 581.3200 ;
        RECT 2473.7800 586.2800 2476.7800 586.7600 ;
        RECT 2485.5400 564.5200 2487.1400 565.0000 ;
        RECT 2485.5400 569.9600 2487.1400 570.4400 ;
        RECT 2473.7800 564.5200 2476.7800 565.0000 ;
        RECT 2473.7800 569.9600 2476.7800 570.4400 ;
        RECT 2485.5400 548.2000 2487.1400 548.6800 ;
        RECT 2485.5400 553.6400 2487.1400 554.1200 ;
        RECT 2485.5400 559.0800 2487.1400 559.5600 ;
        RECT 2473.7800 548.2000 2476.7800 548.6800 ;
        RECT 2473.7800 553.6400 2476.7800 554.1200 ;
        RECT 2473.7800 559.0800 2476.7800 559.5600 ;
        RECT 2473.7800 542.7600 2476.7800 543.2400 ;
        RECT 2485.5400 542.7600 2487.1400 543.2400 ;
        RECT 2473.7800 747.6700 2680.8800 750.6700 ;
        RECT 2473.7800 534.5700 2680.8800 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 304.9300 2667.1400 521.0300 ;
        RECT 2620.5400 304.9300 2622.1400 521.0300 ;
        RECT 2575.5400 304.9300 2577.1400 521.0300 ;
        RECT 2530.5400 304.9300 2532.1400 521.0300 ;
        RECT 2485.5400 304.9300 2487.1400 521.0300 ;
        RECT 2677.8800 304.9300 2680.8800 521.0300 ;
        RECT 2473.7800 304.9300 2476.7800 521.0300 ;
      LAYER met3 ;
        RECT 2677.8800 498.0800 2680.8800 498.5600 ;
        RECT 2677.8800 503.5200 2680.8800 504.0000 ;
        RECT 2665.5400 498.0800 2667.1400 498.5600 ;
        RECT 2665.5400 503.5200 2667.1400 504.0000 ;
        RECT 2677.8800 508.9600 2680.8800 509.4400 ;
        RECT 2665.5400 508.9600 2667.1400 509.4400 ;
        RECT 2677.8800 487.2000 2680.8800 487.6800 ;
        RECT 2677.8800 492.6400 2680.8800 493.1200 ;
        RECT 2665.5400 487.2000 2667.1400 487.6800 ;
        RECT 2665.5400 492.6400 2667.1400 493.1200 ;
        RECT 2677.8800 470.8800 2680.8800 471.3600 ;
        RECT 2677.8800 476.3200 2680.8800 476.8000 ;
        RECT 2665.5400 470.8800 2667.1400 471.3600 ;
        RECT 2665.5400 476.3200 2667.1400 476.8000 ;
        RECT 2677.8800 481.7600 2680.8800 482.2400 ;
        RECT 2665.5400 481.7600 2667.1400 482.2400 ;
        RECT 2620.5400 498.0800 2622.1400 498.5600 ;
        RECT 2620.5400 503.5200 2622.1400 504.0000 ;
        RECT 2620.5400 508.9600 2622.1400 509.4400 ;
        RECT 2620.5400 487.2000 2622.1400 487.6800 ;
        RECT 2620.5400 492.6400 2622.1400 493.1200 ;
        RECT 2620.5400 470.8800 2622.1400 471.3600 ;
        RECT 2620.5400 476.3200 2622.1400 476.8000 ;
        RECT 2620.5400 481.7600 2622.1400 482.2400 ;
        RECT 2677.8800 454.5600 2680.8800 455.0400 ;
        RECT 2677.8800 460.0000 2680.8800 460.4800 ;
        RECT 2677.8800 465.4400 2680.8800 465.9200 ;
        RECT 2665.5400 454.5600 2667.1400 455.0400 ;
        RECT 2665.5400 460.0000 2667.1400 460.4800 ;
        RECT 2665.5400 465.4400 2667.1400 465.9200 ;
        RECT 2677.8800 443.6800 2680.8800 444.1600 ;
        RECT 2677.8800 449.1200 2680.8800 449.6000 ;
        RECT 2665.5400 443.6800 2667.1400 444.1600 ;
        RECT 2665.5400 449.1200 2667.1400 449.6000 ;
        RECT 2677.8800 427.3600 2680.8800 427.8400 ;
        RECT 2677.8800 432.8000 2680.8800 433.2800 ;
        RECT 2677.8800 438.2400 2680.8800 438.7200 ;
        RECT 2665.5400 427.3600 2667.1400 427.8400 ;
        RECT 2665.5400 432.8000 2667.1400 433.2800 ;
        RECT 2665.5400 438.2400 2667.1400 438.7200 ;
        RECT 2677.8800 416.4800 2680.8800 416.9600 ;
        RECT 2677.8800 421.9200 2680.8800 422.4000 ;
        RECT 2665.5400 416.4800 2667.1400 416.9600 ;
        RECT 2665.5400 421.9200 2667.1400 422.4000 ;
        RECT 2620.5400 454.5600 2622.1400 455.0400 ;
        RECT 2620.5400 460.0000 2622.1400 460.4800 ;
        RECT 2620.5400 465.4400 2622.1400 465.9200 ;
        RECT 2620.5400 443.6800 2622.1400 444.1600 ;
        RECT 2620.5400 449.1200 2622.1400 449.6000 ;
        RECT 2620.5400 427.3600 2622.1400 427.8400 ;
        RECT 2620.5400 432.8000 2622.1400 433.2800 ;
        RECT 2620.5400 438.2400 2622.1400 438.7200 ;
        RECT 2620.5400 416.4800 2622.1400 416.9600 ;
        RECT 2620.5400 421.9200 2622.1400 422.4000 ;
        RECT 2575.5400 498.0800 2577.1400 498.5600 ;
        RECT 2575.5400 503.5200 2577.1400 504.0000 ;
        RECT 2575.5400 508.9600 2577.1400 509.4400 ;
        RECT 2530.5400 498.0800 2532.1400 498.5600 ;
        RECT 2530.5400 503.5200 2532.1400 504.0000 ;
        RECT 2530.5400 508.9600 2532.1400 509.4400 ;
        RECT 2575.5400 487.2000 2577.1400 487.6800 ;
        RECT 2575.5400 492.6400 2577.1400 493.1200 ;
        RECT 2575.5400 470.8800 2577.1400 471.3600 ;
        RECT 2575.5400 476.3200 2577.1400 476.8000 ;
        RECT 2575.5400 481.7600 2577.1400 482.2400 ;
        RECT 2530.5400 487.2000 2532.1400 487.6800 ;
        RECT 2530.5400 492.6400 2532.1400 493.1200 ;
        RECT 2530.5400 470.8800 2532.1400 471.3600 ;
        RECT 2530.5400 476.3200 2532.1400 476.8000 ;
        RECT 2530.5400 481.7600 2532.1400 482.2400 ;
        RECT 2485.5400 498.0800 2487.1400 498.5600 ;
        RECT 2485.5400 503.5200 2487.1400 504.0000 ;
        RECT 2473.7800 503.5200 2476.7800 504.0000 ;
        RECT 2473.7800 498.0800 2476.7800 498.5600 ;
        RECT 2473.7800 508.9600 2476.7800 509.4400 ;
        RECT 2485.5400 508.9600 2487.1400 509.4400 ;
        RECT 2485.5400 487.2000 2487.1400 487.6800 ;
        RECT 2485.5400 492.6400 2487.1400 493.1200 ;
        RECT 2473.7800 492.6400 2476.7800 493.1200 ;
        RECT 2473.7800 487.2000 2476.7800 487.6800 ;
        RECT 2485.5400 470.8800 2487.1400 471.3600 ;
        RECT 2485.5400 476.3200 2487.1400 476.8000 ;
        RECT 2473.7800 476.3200 2476.7800 476.8000 ;
        RECT 2473.7800 470.8800 2476.7800 471.3600 ;
        RECT 2473.7800 481.7600 2476.7800 482.2400 ;
        RECT 2485.5400 481.7600 2487.1400 482.2400 ;
        RECT 2575.5400 454.5600 2577.1400 455.0400 ;
        RECT 2575.5400 460.0000 2577.1400 460.4800 ;
        RECT 2575.5400 465.4400 2577.1400 465.9200 ;
        RECT 2575.5400 443.6800 2577.1400 444.1600 ;
        RECT 2575.5400 449.1200 2577.1400 449.6000 ;
        RECT 2530.5400 454.5600 2532.1400 455.0400 ;
        RECT 2530.5400 460.0000 2532.1400 460.4800 ;
        RECT 2530.5400 465.4400 2532.1400 465.9200 ;
        RECT 2530.5400 443.6800 2532.1400 444.1600 ;
        RECT 2530.5400 449.1200 2532.1400 449.6000 ;
        RECT 2575.5400 427.3600 2577.1400 427.8400 ;
        RECT 2575.5400 432.8000 2577.1400 433.2800 ;
        RECT 2575.5400 438.2400 2577.1400 438.7200 ;
        RECT 2575.5400 416.4800 2577.1400 416.9600 ;
        RECT 2575.5400 421.9200 2577.1400 422.4000 ;
        RECT 2530.5400 427.3600 2532.1400 427.8400 ;
        RECT 2530.5400 432.8000 2532.1400 433.2800 ;
        RECT 2530.5400 438.2400 2532.1400 438.7200 ;
        RECT 2530.5400 416.4800 2532.1400 416.9600 ;
        RECT 2530.5400 421.9200 2532.1400 422.4000 ;
        RECT 2485.5400 454.5600 2487.1400 455.0400 ;
        RECT 2485.5400 460.0000 2487.1400 460.4800 ;
        RECT 2485.5400 465.4400 2487.1400 465.9200 ;
        RECT 2473.7800 454.5600 2476.7800 455.0400 ;
        RECT 2473.7800 460.0000 2476.7800 460.4800 ;
        RECT 2473.7800 465.4400 2476.7800 465.9200 ;
        RECT 2485.5400 443.6800 2487.1400 444.1600 ;
        RECT 2485.5400 449.1200 2487.1400 449.6000 ;
        RECT 2473.7800 443.6800 2476.7800 444.1600 ;
        RECT 2473.7800 449.1200 2476.7800 449.6000 ;
        RECT 2485.5400 427.3600 2487.1400 427.8400 ;
        RECT 2485.5400 432.8000 2487.1400 433.2800 ;
        RECT 2485.5400 438.2400 2487.1400 438.7200 ;
        RECT 2473.7800 427.3600 2476.7800 427.8400 ;
        RECT 2473.7800 432.8000 2476.7800 433.2800 ;
        RECT 2473.7800 438.2400 2476.7800 438.7200 ;
        RECT 2485.5400 416.4800 2487.1400 416.9600 ;
        RECT 2485.5400 421.9200 2487.1400 422.4000 ;
        RECT 2473.7800 416.4800 2476.7800 416.9600 ;
        RECT 2473.7800 421.9200 2476.7800 422.4000 ;
        RECT 2677.8800 400.1600 2680.8800 400.6400 ;
        RECT 2677.8800 405.6000 2680.8800 406.0800 ;
        RECT 2677.8800 411.0400 2680.8800 411.5200 ;
        RECT 2665.5400 400.1600 2667.1400 400.6400 ;
        RECT 2665.5400 405.6000 2667.1400 406.0800 ;
        RECT 2665.5400 411.0400 2667.1400 411.5200 ;
        RECT 2677.8800 389.2800 2680.8800 389.7600 ;
        RECT 2677.8800 394.7200 2680.8800 395.2000 ;
        RECT 2665.5400 389.2800 2667.1400 389.7600 ;
        RECT 2665.5400 394.7200 2667.1400 395.2000 ;
        RECT 2677.8800 372.9600 2680.8800 373.4400 ;
        RECT 2677.8800 378.4000 2680.8800 378.8800 ;
        RECT 2677.8800 383.8400 2680.8800 384.3200 ;
        RECT 2665.5400 372.9600 2667.1400 373.4400 ;
        RECT 2665.5400 378.4000 2667.1400 378.8800 ;
        RECT 2665.5400 383.8400 2667.1400 384.3200 ;
        RECT 2677.8800 362.0800 2680.8800 362.5600 ;
        RECT 2677.8800 367.5200 2680.8800 368.0000 ;
        RECT 2665.5400 362.0800 2667.1400 362.5600 ;
        RECT 2665.5400 367.5200 2667.1400 368.0000 ;
        RECT 2620.5400 400.1600 2622.1400 400.6400 ;
        RECT 2620.5400 405.6000 2622.1400 406.0800 ;
        RECT 2620.5400 411.0400 2622.1400 411.5200 ;
        RECT 2620.5400 389.2800 2622.1400 389.7600 ;
        RECT 2620.5400 394.7200 2622.1400 395.2000 ;
        RECT 2620.5400 372.9600 2622.1400 373.4400 ;
        RECT 2620.5400 378.4000 2622.1400 378.8800 ;
        RECT 2620.5400 383.8400 2622.1400 384.3200 ;
        RECT 2620.5400 362.0800 2622.1400 362.5600 ;
        RECT 2620.5400 367.5200 2622.1400 368.0000 ;
        RECT 2677.8800 345.7600 2680.8800 346.2400 ;
        RECT 2677.8800 351.2000 2680.8800 351.6800 ;
        RECT 2677.8800 356.6400 2680.8800 357.1200 ;
        RECT 2665.5400 345.7600 2667.1400 346.2400 ;
        RECT 2665.5400 351.2000 2667.1400 351.6800 ;
        RECT 2665.5400 356.6400 2667.1400 357.1200 ;
        RECT 2677.8800 334.8800 2680.8800 335.3600 ;
        RECT 2677.8800 340.3200 2680.8800 340.8000 ;
        RECT 2665.5400 334.8800 2667.1400 335.3600 ;
        RECT 2665.5400 340.3200 2667.1400 340.8000 ;
        RECT 2677.8800 318.5600 2680.8800 319.0400 ;
        RECT 2677.8800 324.0000 2680.8800 324.4800 ;
        RECT 2677.8800 329.4400 2680.8800 329.9200 ;
        RECT 2665.5400 318.5600 2667.1400 319.0400 ;
        RECT 2665.5400 324.0000 2667.1400 324.4800 ;
        RECT 2665.5400 329.4400 2667.1400 329.9200 ;
        RECT 2677.8800 313.1200 2680.8800 313.6000 ;
        RECT 2665.5400 313.1200 2667.1400 313.6000 ;
        RECT 2620.5400 345.7600 2622.1400 346.2400 ;
        RECT 2620.5400 351.2000 2622.1400 351.6800 ;
        RECT 2620.5400 356.6400 2622.1400 357.1200 ;
        RECT 2620.5400 334.8800 2622.1400 335.3600 ;
        RECT 2620.5400 340.3200 2622.1400 340.8000 ;
        RECT 2620.5400 318.5600 2622.1400 319.0400 ;
        RECT 2620.5400 324.0000 2622.1400 324.4800 ;
        RECT 2620.5400 329.4400 2622.1400 329.9200 ;
        RECT 2620.5400 313.1200 2622.1400 313.6000 ;
        RECT 2575.5400 400.1600 2577.1400 400.6400 ;
        RECT 2575.5400 405.6000 2577.1400 406.0800 ;
        RECT 2575.5400 411.0400 2577.1400 411.5200 ;
        RECT 2575.5400 389.2800 2577.1400 389.7600 ;
        RECT 2575.5400 394.7200 2577.1400 395.2000 ;
        RECT 2530.5400 400.1600 2532.1400 400.6400 ;
        RECT 2530.5400 405.6000 2532.1400 406.0800 ;
        RECT 2530.5400 411.0400 2532.1400 411.5200 ;
        RECT 2530.5400 389.2800 2532.1400 389.7600 ;
        RECT 2530.5400 394.7200 2532.1400 395.2000 ;
        RECT 2575.5400 372.9600 2577.1400 373.4400 ;
        RECT 2575.5400 378.4000 2577.1400 378.8800 ;
        RECT 2575.5400 383.8400 2577.1400 384.3200 ;
        RECT 2575.5400 362.0800 2577.1400 362.5600 ;
        RECT 2575.5400 367.5200 2577.1400 368.0000 ;
        RECT 2530.5400 372.9600 2532.1400 373.4400 ;
        RECT 2530.5400 378.4000 2532.1400 378.8800 ;
        RECT 2530.5400 383.8400 2532.1400 384.3200 ;
        RECT 2530.5400 362.0800 2532.1400 362.5600 ;
        RECT 2530.5400 367.5200 2532.1400 368.0000 ;
        RECT 2485.5400 400.1600 2487.1400 400.6400 ;
        RECT 2485.5400 405.6000 2487.1400 406.0800 ;
        RECT 2485.5400 411.0400 2487.1400 411.5200 ;
        RECT 2473.7800 400.1600 2476.7800 400.6400 ;
        RECT 2473.7800 405.6000 2476.7800 406.0800 ;
        RECT 2473.7800 411.0400 2476.7800 411.5200 ;
        RECT 2485.5400 389.2800 2487.1400 389.7600 ;
        RECT 2485.5400 394.7200 2487.1400 395.2000 ;
        RECT 2473.7800 389.2800 2476.7800 389.7600 ;
        RECT 2473.7800 394.7200 2476.7800 395.2000 ;
        RECT 2485.5400 372.9600 2487.1400 373.4400 ;
        RECT 2485.5400 378.4000 2487.1400 378.8800 ;
        RECT 2485.5400 383.8400 2487.1400 384.3200 ;
        RECT 2473.7800 372.9600 2476.7800 373.4400 ;
        RECT 2473.7800 378.4000 2476.7800 378.8800 ;
        RECT 2473.7800 383.8400 2476.7800 384.3200 ;
        RECT 2485.5400 362.0800 2487.1400 362.5600 ;
        RECT 2485.5400 367.5200 2487.1400 368.0000 ;
        RECT 2473.7800 362.0800 2476.7800 362.5600 ;
        RECT 2473.7800 367.5200 2476.7800 368.0000 ;
        RECT 2575.5400 345.7600 2577.1400 346.2400 ;
        RECT 2575.5400 351.2000 2577.1400 351.6800 ;
        RECT 2575.5400 356.6400 2577.1400 357.1200 ;
        RECT 2575.5400 334.8800 2577.1400 335.3600 ;
        RECT 2575.5400 340.3200 2577.1400 340.8000 ;
        RECT 2530.5400 345.7600 2532.1400 346.2400 ;
        RECT 2530.5400 351.2000 2532.1400 351.6800 ;
        RECT 2530.5400 356.6400 2532.1400 357.1200 ;
        RECT 2530.5400 334.8800 2532.1400 335.3600 ;
        RECT 2530.5400 340.3200 2532.1400 340.8000 ;
        RECT 2575.5400 318.5600 2577.1400 319.0400 ;
        RECT 2575.5400 324.0000 2577.1400 324.4800 ;
        RECT 2575.5400 329.4400 2577.1400 329.9200 ;
        RECT 2575.5400 313.1200 2577.1400 313.6000 ;
        RECT 2530.5400 318.5600 2532.1400 319.0400 ;
        RECT 2530.5400 324.0000 2532.1400 324.4800 ;
        RECT 2530.5400 329.4400 2532.1400 329.9200 ;
        RECT 2530.5400 313.1200 2532.1400 313.6000 ;
        RECT 2485.5400 345.7600 2487.1400 346.2400 ;
        RECT 2485.5400 351.2000 2487.1400 351.6800 ;
        RECT 2485.5400 356.6400 2487.1400 357.1200 ;
        RECT 2473.7800 345.7600 2476.7800 346.2400 ;
        RECT 2473.7800 351.2000 2476.7800 351.6800 ;
        RECT 2473.7800 356.6400 2476.7800 357.1200 ;
        RECT 2485.5400 334.8800 2487.1400 335.3600 ;
        RECT 2485.5400 340.3200 2487.1400 340.8000 ;
        RECT 2473.7800 334.8800 2476.7800 335.3600 ;
        RECT 2473.7800 340.3200 2476.7800 340.8000 ;
        RECT 2485.5400 318.5600 2487.1400 319.0400 ;
        RECT 2485.5400 324.0000 2487.1400 324.4800 ;
        RECT 2485.5400 329.4400 2487.1400 329.9200 ;
        RECT 2473.7800 318.5600 2476.7800 319.0400 ;
        RECT 2473.7800 324.0000 2476.7800 324.4800 ;
        RECT 2473.7800 329.4400 2476.7800 329.9200 ;
        RECT 2473.7800 313.1200 2476.7800 313.6000 ;
        RECT 2485.5400 313.1200 2487.1400 313.6000 ;
        RECT 2473.7800 518.0300 2680.8800 521.0300 ;
        RECT 2473.7800 304.9300 2680.8800 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 75.2900 2667.1400 291.3900 ;
        RECT 2620.5400 75.2900 2622.1400 291.3900 ;
        RECT 2575.5400 75.2900 2577.1400 291.3900 ;
        RECT 2530.5400 75.2900 2532.1400 291.3900 ;
        RECT 2485.5400 75.2900 2487.1400 291.3900 ;
        RECT 2677.8800 75.2900 2680.8800 291.3900 ;
        RECT 2473.7800 75.2900 2476.7800 291.3900 ;
      LAYER met3 ;
        RECT 2677.8800 268.4400 2680.8800 268.9200 ;
        RECT 2677.8800 273.8800 2680.8800 274.3600 ;
        RECT 2665.5400 268.4400 2667.1400 268.9200 ;
        RECT 2665.5400 273.8800 2667.1400 274.3600 ;
        RECT 2677.8800 279.3200 2680.8800 279.8000 ;
        RECT 2665.5400 279.3200 2667.1400 279.8000 ;
        RECT 2677.8800 257.5600 2680.8800 258.0400 ;
        RECT 2677.8800 263.0000 2680.8800 263.4800 ;
        RECT 2665.5400 257.5600 2667.1400 258.0400 ;
        RECT 2665.5400 263.0000 2667.1400 263.4800 ;
        RECT 2677.8800 241.2400 2680.8800 241.7200 ;
        RECT 2677.8800 246.6800 2680.8800 247.1600 ;
        RECT 2665.5400 241.2400 2667.1400 241.7200 ;
        RECT 2665.5400 246.6800 2667.1400 247.1600 ;
        RECT 2677.8800 252.1200 2680.8800 252.6000 ;
        RECT 2665.5400 252.1200 2667.1400 252.6000 ;
        RECT 2620.5400 268.4400 2622.1400 268.9200 ;
        RECT 2620.5400 273.8800 2622.1400 274.3600 ;
        RECT 2620.5400 279.3200 2622.1400 279.8000 ;
        RECT 2620.5400 257.5600 2622.1400 258.0400 ;
        RECT 2620.5400 263.0000 2622.1400 263.4800 ;
        RECT 2620.5400 241.2400 2622.1400 241.7200 ;
        RECT 2620.5400 246.6800 2622.1400 247.1600 ;
        RECT 2620.5400 252.1200 2622.1400 252.6000 ;
        RECT 2677.8800 224.9200 2680.8800 225.4000 ;
        RECT 2677.8800 230.3600 2680.8800 230.8400 ;
        RECT 2677.8800 235.8000 2680.8800 236.2800 ;
        RECT 2665.5400 224.9200 2667.1400 225.4000 ;
        RECT 2665.5400 230.3600 2667.1400 230.8400 ;
        RECT 2665.5400 235.8000 2667.1400 236.2800 ;
        RECT 2677.8800 214.0400 2680.8800 214.5200 ;
        RECT 2677.8800 219.4800 2680.8800 219.9600 ;
        RECT 2665.5400 214.0400 2667.1400 214.5200 ;
        RECT 2665.5400 219.4800 2667.1400 219.9600 ;
        RECT 2677.8800 197.7200 2680.8800 198.2000 ;
        RECT 2677.8800 203.1600 2680.8800 203.6400 ;
        RECT 2677.8800 208.6000 2680.8800 209.0800 ;
        RECT 2665.5400 197.7200 2667.1400 198.2000 ;
        RECT 2665.5400 203.1600 2667.1400 203.6400 ;
        RECT 2665.5400 208.6000 2667.1400 209.0800 ;
        RECT 2677.8800 186.8400 2680.8800 187.3200 ;
        RECT 2677.8800 192.2800 2680.8800 192.7600 ;
        RECT 2665.5400 186.8400 2667.1400 187.3200 ;
        RECT 2665.5400 192.2800 2667.1400 192.7600 ;
        RECT 2620.5400 224.9200 2622.1400 225.4000 ;
        RECT 2620.5400 230.3600 2622.1400 230.8400 ;
        RECT 2620.5400 235.8000 2622.1400 236.2800 ;
        RECT 2620.5400 214.0400 2622.1400 214.5200 ;
        RECT 2620.5400 219.4800 2622.1400 219.9600 ;
        RECT 2620.5400 197.7200 2622.1400 198.2000 ;
        RECT 2620.5400 203.1600 2622.1400 203.6400 ;
        RECT 2620.5400 208.6000 2622.1400 209.0800 ;
        RECT 2620.5400 186.8400 2622.1400 187.3200 ;
        RECT 2620.5400 192.2800 2622.1400 192.7600 ;
        RECT 2575.5400 268.4400 2577.1400 268.9200 ;
        RECT 2575.5400 273.8800 2577.1400 274.3600 ;
        RECT 2575.5400 279.3200 2577.1400 279.8000 ;
        RECT 2530.5400 268.4400 2532.1400 268.9200 ;
        RECT 2530.5400 273.8800 2532.1400 274.3600 ;
        RECT 2530.5400 279.3200 2532.1400 279.8000 ;
        RECT 2575.5400 257.5600 2577.1400 258.0400 ;
        RECT 2575.5400 263.0000 2577.1400 263.4800 ;
        RECT 2575.5400 241.2400 2577.1400 241.7200 ;
        RECT 2575.5400 246.6800 2577.1400 247.1600 ;
        RECT 2575.5400 252.1200 2577.1400 252.6000 ;
        RECT 2530.5400 257.5600 2532.1400 258.0400 ;
        RECT 2530.5400 263.0000 2532.1400 263.4800 ;
        RECT 2530.5400 241.2400 2532.1400 241.7200 ;
        RECT 2530.5400 246.6800 2532.1400 247.1600 ;
        RECT 2530.5400 252.1200 2532.1400 252.6000 ;
        RECT 2485.5400 268.4400 2487.1400 268.9200 ;
        RECT 2485.5400 273.8800 2487.1400 274.3600 ;
        RECT 2473.7800 273.8800 2476.7800 274.3600 ;
        RECT 2473.7800 268.4400 2476.7800 268.9200 ;
        RECT 2473.7800 279.3200 2476.7800 279.8000 ;
        RECT 2485.5400 279.3200 2487.1400 279.8000 ;
        RECT 2485.5400 257.5600 2487.1400 258.0400 ;
        RECT 2485.5400 263.0000 2487.1400 263.4800 ;
        RECT 2473.7800 263.0000 2476.7800 263.4800 ;
        RECT 2473.7800 257.5600 2476.7800 258.0400 ;
        RECT 2485.5400 241.2400 2487.1400 241.7200 ;
        RECT 2485.5400 246.6800 2487.1400 247.1600 ;
        RECT 2473.7800 246.6800 2476.7800 247.1600 ;
        RECT 2473.7800 241.2400 2476.7800 241.7200 ;
        RECT 2473.7800 252.1200 2476.7800 252.6000 ;
        RECT 2485.5400 252.1200 2487.1400 252.6000 ;
        RECT 2575.5400 224.9200 2577.1400 225.4000 ;
        RECT 2575.5400 230.3600 2577.1400 230.8400 ;
        RECT 2575.5400 235.8000 2577.1400 236.2800 ;
        RECT 2575.5400 214.0400 2577.1400 214.5200 ;
        RECT 2575.5400 219.4800 2577.1400 219.9600 ;
        RECT 2530.5400 224.9200 2532.1400 225.4000 ;
        RECT 2530.5400 230.3600 2532.1400 230.8400 ;
        RECT 2530.5400 235.8000 2532.1400 236.2800 ;
        RECT 2530.5400 214.0400 2532.1400 214.5200 ;
        RECT 2530.5400 219.4800 2532.1400 219.9600 ;
        RECT 2575.5400 197.7200 2577.1400 198.2000 ;
        RECT 2575.5400 203.1600 2577.1400 203.6400 ;
        RECT 2575.5400 208.6000 2577.1400 209.0800 ;
        RECT 2575.5400 186.8400 2577.1400 187.3200 ;
        RECT 2575.5400 192.2800 2577.1400 192.7600 ;
        RECT 2530.5400 197.7200 2532.1400 198.2000 ;
        RECT 2530.5400 203.1600 2532.1400 203.6400 ;
        RECT 2530.5400 208.6000 2532.1400 209.0800 ;
        RECT 2530.5400 186.8400 2532.1400 187.3200 ;
        RECT 2530.5400 192.2800 2532.1400 192.7600 ;
        RECT 2485.5400 224.9200 2487.1400 225.4000 ;
        RECT 2485.5400 230.3600 2487.1400 230.8400 ;
        RECT 2485.5400 235.8000 2487.1400 236.2800 ;
        RECT 2473.7800 224.9200 2476.7800 225.4000 ;
        RECT 2473.7800 230.3600 2476.7800 230.8400 ;
        RECT 2473.7800 235.8000 2476.7800 236.2800 ;
        RECT 2485.5400 214.0400 2487.1400 214.5200 ;
        RECT 2485.5400 219.4800 2487.1400 219.9600 ;
        RECT 2473.7800 214.0400 2476.7800 214.5200 ;
        RECT 2473.7800 219.4800 2476.7800 219.9600 ;
        RECT 2485.5400 197.7200 2487.1400 198.2000 ;
        RECT 2485.5400 203.1600 2487.1400 203.6400 ;
        RECT 2485.5400 208.6000 2487.1400 209.0800 ;
        RECT 2473.7800 197.7200 2476.7800 198.2000 ;
        RECT 2473.7800 203.1600 2476.7800 203.6400 ;
        RECT 2473.7800 208.6000 2476.7800 209.0800 ;
        RECT 2485.5400 186.8400 2487.1400 187.3200 ;
        RECT 2485.5400 192.2800 2487.1400 192.7600 ;
        RECT 2473.7800 186.8400 2476.7800 187.3200 ;
        RECT 2473.7800 192.2800 2476.7800 192.7600 ;
        RECT 2677.8800 170.5200 2680.8800 171.0000 ;
        RECT 2677.8800 175.9600 2680.8800 176.4400 ;
        RECT 2677.8800 181.4000 2680.8800 181.8800 ;
        RECT 2665.5400 170.5200 2667.1400 171.0000 ;
        RECT 2665.5400 175.9600 2667.1400 176.4400 ;
        RECT 2665.5400 181.4000 2667.1400 181.8800 ;
        RECT 2677.8800 159.6400 2680.8800 160.1200 ;
        RECT 2677.8800 165.0800 2680.8800 165.5600 ;
        RECT 2665.5400 159.6400 2667.1400 160.1200 ;
        RECT 2665.5400 165.0800 2667.1400 165.5600 ;
        RECT 2677.8800 143.3200 2680.8800 143.8000 ;
        RECT 2677.8800 148.7600 2680.8800 149.2400 ;
        RECT 2677.8800 154.2000 2680.8800 154.6800 ;
        RECT 2665.5400 143.3200 2667.1400 143.8000 ;
        RECT 2665.5400 148.7600 2667.1400 149.2400 ;
        RECT 2665.5400 154.2000 2667.1400 154.6800 ;
        RECT 2677.8800 132.4400 2680.8800 132.9200 ;
        RECT 2677.8800 137.8800 2680.8800 138.3600 ;
        RECT 2665.5400 132.4400 2667.1400 132.9200 ;
        RECT 2665.5400 137.8800 2667.1400 138.3600 ;
        RECT 2620.5400 170.5200 2622.1400 171.0000 ;
        RECT 2620.5400 175.9600 2622.1400 176.4400 ;
        RECT 2620.5400 181.4000 2622.1400 181.8800 ;
        RECT 2620.5400 159.6400 2622.1400 160.1200 ;
        RECT 2620.5400 165.0800 2622.1400 165.5600 ;
        RECT 2620.5400 143.3200 2622.1400 143.8000 ;
        RECT 2620.5400 148.7600 2622.1400 149.2400 ;
        RECT 2620.5400 154.2000 2622.1400 154.6800 ;
        RECT 2620.5400 132.4400 2622.1400 132.9200 ;
        RECT 2620.5400 137.8800 2622.1400 138.3600 ;
        RECT 2677.8800 116.1200 2680.8800 116.6000 ;
        RECT 2677.8800 121.5600 2680.8800 122.0400 ;
        RECT 2677.8800 127.0000 2680.8800 127.4800 ;
        RECT 2665.5400 116.1200 2667.1400 116.6000 ;
        RECT 2665.5400 121.5600 2667.1400 122.0400 ;
        RECT 2665.5400 127.0000 2667.1400 127.4800 ;
        RECT 2677.8800 105.2400 2680.8800 105.7200 ;
        RECT 2677.8800 110.6800 2680.8800 111.1600 ;
        RECT 2665.5400 105.2400 2667.1400 105.7200 ;
        RECT 2665.5400 110.6800 2667.1400 111.1600 ;
        RECT 2677.8800 88.9200 2680.8800 89.4000 ;
        RECT 2677.8800 94.3600 2680.8800 94.8400 ;
        RECT 2677.8800 99.8000 2680.8800 100.2800 ;
        RECT 2665.5400 88.9200 2667.1400 89.4000 ;
        RECT 2665.5400 94.3600 2667.1400 94.8400 ;
        RECT 2665.5400 99.8000 2667.1400 100.2800 ;
        RECT 2677.8800 83.4800 2680.8800 83.9600 ;
        RECT 2665.5400 83.4800 2667.1400 83.9600 ;
        RECT 2620.5400 116.1200 2622.1400 116.6000 ;
        RECT 2620.5400 121.5600 2622.1400 122.0400 ;
        RECT 2620.5400 127.0000 2622.1400 127.4800 ;
        RECT 2620.5400 105.2400 2622.1400 105.7200 ;
        RECT 2620.5400 110.6800 2622.1400 111.1600 ;
        RECT 2620.5400 88.9200 2622.1400 89.4000 ;
        RECT 2620.5400 94.3600 2622.1400 94.8400 ;
        RECT 2620.5400 99.8000 2622.1400 100.2800 ;
        RECT 2620.5400 83.4800 2622.1400 83.9600 ;
        RECT 2575.5400 170.5200 2577.1400 171.0000 ;
        RECT 2575.5400 175.9600 2577.1400 176.4400 ;
        RECT 2575.5400 181.4000 2577.1400 181.8800 ;
        RECT 2575.5400 159.6400 2577.1400 160.1200 ;
        RECT 2575.5400 165.0800 2577.1400 165.5600 ;
        RECT 2530.5400 170.5200 2532.1400 171.0000 ;
        RECT 2530.5400 175.9600 2532.1400 176.4400 ;
        RECT 2530.5400 181.4000 2532.1400 181.8800 ;
        RECT 2530.5400 159.6400 2532.1400 160.1200 ;
        RECT 2530.5400 165.0800 2532.1400 165.5600 ;
        RECT 2575.5400 143.3200 2577.1400 143.8000 ;
        RECT 2575.5400 148.7600 2577.1400 149.2400 ;
        RECT 2575.5400 154.2000 2577.1400 154.6800 ;
        RECT 2575.5400 132.4400 2577.1400 132.9200 ;
        RECT 2575.5400 137.8800 2577.1400 138.3600 ;
        RECT 2530.5400 143.3200 2532.1400 143.8000 ;
        RECT 2530.5400 148.7600 2532.1400 149.2400 ;
        RECT 2530.5400 154.2000 2532.1400 154.6800 ;
        RECT 2530.5400 132.4400 2532.1400 132.9200 ;
        RECT 2530.5400 137.8800 2532.1400 138.3600 ;
        RECT 2485.5400 170.5200 2487.1400 171.0000 ;
        RECT 2485.5400 175.9600 2487.1400 176.4400 ;
        RECT 2485.5400 181.4000 2487.1400 181.8800 ;
        RECT 2473.7800 170.5200 2476.7800 171.0000 ;
        RECT 2473.7800 175.9600 2476.7800 176.4400 ;
        RECT 2473.7800 181.4000 2476.7800 181.8800 ;
        RECT 2485.5400 159.6400 2487.1400 160.1200 ;
        RECT 2485.5400 165.0800 2487.1400 165.5600 ;
        RECT 2473.7800 159.6400 2476.7800 160.1200 ;
        RECT 2473.7800 165.0800 2476.7800 165.5600 ;
        RECT 2485.5400 143.3200 2487.1400 143.8000 ;
        RECT 2485.5400 148.7600 2487.1400 149.2400 ;
        RECT 2485.5400 154.2000 2487.1400 154.6800 ;
        RECT 2473.7800 143.3200 2476.7800 143.8000 ;
        RECT 2473.7800 148.7600 2476.7800 149.2400 ;
        RECT 2473.7800 154.2000 2476.7800 154.6800 ;
        RECT 2485.5400 132.4400 2487.1400 132.9200 ;
        RECT 2485.5400 137.8800 2487.1400 138.3600 ;
        RECT 2473.7800 132.4400 2476.7800 132.9200 ;
        RECT 2473.7800 137.8800 2476.7800 138.3600 ;
        RECT 2575.5400 116.1200 2577.1400 116.6000 ;
        RECT 2575.5400 121.5600 2577.1400 122.0400 ;
        RECT 2575.5400 127.0000 2577.1400 127.4800 ;
        RECT 2575.5400 105.2400 2577.1400 105.7200 ;
        RECT 2575.5400 110.6800 2577.1400 111.1600 ;
        RECT 2530.5400 116.1200 2532.1400 116.6000 ;
        RECT 2530.5400 121.5600 2532.1400 122.0400 ;
        RECT 2530.5400 127.0000 2532.1400 127.4800 ;
        RECT 2530.5400 105.2400 2532.1400 105.7200 ;
        RECT 2530.5400 110.6800 2532.1400 111.1600 ;
        RECT 2575.5400 88.9200 2577.1400 89.4000 ;
        RECT 2575.5400 94.3600 2577.1400 94.8400 ;
        RECT 2575.5400 99.8000 2577.1400 100.2800 ;
        RECT 2575.5400 83.4800 2577.1400 83.9600 ;
        RECT 2530.5400 88.9200 2532.1400 89.4000 ;
        RECT 2530.5400 94.3600 2532.1400 94.8400 ;
        RECT 2530.5400 99.8000 2532.1400 100.2800 ;
        RECT 2530.5400 83.4800 2532.1400 83.9600 ;
        RECT 2485.5400 116.1200 2487.1400 116.6000 ;
        RECT 2485.5400 121.5600 2487.1400 122.0400 ;
        RECT 2485.5400 127.0000 2487.1400 127.4800 ;
        RECT 2473.7800 116.1200 2476.7800 116.6000 ;
        RECT 2473.7800 121.5600 2476.7800 122.0400 ;
        RECT 2473.7800 127.0000 2476.7800 127.4800 ;
        RECT 2485.5400 105.2400 2487.1400 105.7200 ;
        RECT 2485.5400 110.6800 2487.1400 111.1600 ;
        RECT 2473.7800 105.2400 2476.7800 105.7200 ;
        RECT 2473.7800 110.6800 2476.7800 111.1600 ;
        RECT 2485.5400 88.9200 2487.1400 89.4000 ;
        RECT 2485.5400 94.3600 2487.1400 94.8400 ;
        RECT 2485.5400 99.8000 2487.1400 100.2800 ;
        RECT 2473.7800 88.9200 2476.7800 89.4000 ;
        RECT 2473.7800 94.3600 2476.7800 94.8400 ;
        RECT 2473.7800 99.8000 2476.7800 100.2800 ;
        RECT 2473.7800 83.4800 2476.7800 83.9600 ;
        RECT 2485.5400 83.4800 2487.1400 83.9600 ;
        RECT 2473.7800 288.3900 2680.8800 291.3900 ;
        RECT 2473.7800 75.2900 2680.8800 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 2474.7800 34.6700 2476.7800 61.6000 ;
        RECT 2677.8800 34.6700 2679.8800 61.6000 ;
      LAYER met3 ;
        RECT 2677.8800 51.3800 2679.8800 51.8600 ;
        RECT 2474.7800 51.3800 2476.7800 51.8600 ;
        RECT 2677.8800 45.9400 2679.8800 46.4200 ;
        RECT 2677.8800 40.5000 2679.8800 40.9800 ;
        RECT 2474.7800 45.9400 2476.7800 46.4200 ;
        RECT 2474.7800 40.5000 2476.7800 40.9800 ;
        RECT 2474.7800 59.6000 2679.8800 61.6000 ;
        RECT 2474.7800 34.6700 2679.8800 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 2601.3300 2667.1400 2817.4300 ;
        RECT 2620.5400 2601.3300 2622.1400 2817.4300 ;
        RECT 2575.5400 2601.3300 2577.1400 2817.4300 ;
        RECT 2530.5400 2601.3300 2532.1400 2817.4300 ;
        RECT 2485.5400 2601.3300 2487.1400 2817.4300 ;
        RECT 2677.8800 2601.3300 2680.8800 2817.4300 ;
        RECT 2473.7800 2601.3300 2476.7800 2817.4300 ;
      LAYER met3 ;
        RECT 2677.8800 2794.4800 2680.8800 2794.9600 ;
        RECT 2677.8800 2799.9200 2680.8800 2800.4000 ;
        RECT 2665.5400 2794.4800 2667.1400 2794.9600 ;
        RECT 2665.5400 2799.9200 2667.1400 2800.4000 ;
        RECT 2677.8800 2805.3600 2680.8800 2805.8400 ;
        RECT 2665.5400 2805.3600 2667.1400 2805.8400 ;
        RECT 2677.8800 2783.6000 2680.8800 2784.0800 ;
        RECT 2677.8800 2789.0400 2680.8800 2789.5200 ;
        RECT 2665.5400 2783.6000 2667.1400 2784.0800 ;
        RECT 2665.5400 2789.0400 2667.1400 2789.5200 ;
        RECT 2677.8800 2767.2800 2680.8800 2767.7600 ;
        RECT 2677.8800 2772.7200 2680.8800 2773.2000 ;
        RECT 2665.5400 2767.2800 2667.1400 2767.7600 ;
        RECT 2665.5400 2772.7200 2667.1400 2773.2000 ;
        RECT 2677.8800 2778.1600 2680.8800 2778.6400 ;
        RECT 2665.5400 2778.1600 2667.1400 2778.6400 ;
        RECT 2620.5400 2794.4800 2622.1400 2794.9600 ;
        RECT 2620.5400 2799.9200 2622.1400 2800.4000 ;
        RECT 2620.5400 2805.3600 2622.1400 2805.8400 ;
        RECT 2620.5400 2783.6000 2622.1400 2784.0800 ;
        RECT 2620.5400 2789.0400 2622.1400 2789.5200 ;
        RECT 2620.5400 2767.2800 2622.1400 2767.7600 ;
        RECT 2620.5400 2772.7200 2622.1400 2773.2000 ;
        RECT 2620.5400 2778.1600 2622.1400 2778.6400 ;
        RECT 2677.8800 2750.9600 2680.8800 2751.4400 ;
        RECT 2677.8800 2756.4000 2680.8800 2756.8800 ;
        RECT 2677.8800 2761.8400 2680.8800 2762.3200 ;
        RECT 2665.5400 2750.9600 2667.1400 2751.4400 ;
        RECT 2665.5400 2756.4000 2667.1400 2756.8800 ;
        RECT 2665.5400 2761.8400 2667.1400 2762.3200 ;
        RECT 2677.8800 2740.0800 2680.8800 2740.5600 ;
        RECT 2677.8800 2745.5200 2680.8800 2746.0000 ;
        RECT 2665.5400 2740.0800 2667.1400 2740.5600 ;
        RECT 2665.5400 2745.5200 2667.1400 2746.0000 ;
        RECT 2677.8800 2723.7600 2680.8800 2724.2400 ;
        RECT 2677.8800 2729.2000 2680.8800 2729.6800 ;
        RECT 2677.8800 2734.6400 2680.8800 2735.1200 ;
        RECT 2665.5400 2723.7600 2667.1400 2724.2400 ;
        RECT 2665.5400 2729.2000 2667.1400 2729.6800 ;
        RECT 2665.5400 2734.6400 2667.1400 2735.1200 ;
        RECT 2677.8800 2712.8800 2680.8800 2713.3600 ;
        RECT 2677.8800 2718.3200 2680.8800 2718.8000 ;
        RECT 2665.5400 2712.8800 2667.1400 2713.3600 ;
        RECT 2665.5400 2718.3200 2667.1400 2718.8000 ;
        RECT 2620.5400 2750.9600 2622.1400 2751.4400 ;
        RECT 2620.5400 2756.4000 2622.1400 2756.8800 ;
        RECT 2620.5400 2761.8400 2622.1400 2762.3200 ;
        RECT 2620.5400 2740.0800 2622.1400 2740.5600 ;
        RECT 2620.5400 2745.5200 2622.1400 2746.0000 ;
        RECT 2620.5400 2723.7600 2622.1400 2724.2400 ;
        RECT 2620.5400 2729.2000 2622.1400 2729.6800 ;
        RECT 2620.5400 2734.6400 2622.1400 2735.1200 ;
        RECT 2620.5400 2712.8800 2622.1400 2713.3600 ;
        RECT 2620.5400 2718.3200 2622.1400 2718.8000 ;
        RECT 2575.5400 2794.4800 2577.1400 2794.9600 ;
        RECT 2575.5400 2799.9200 2577.1400 2800.4000 ;
        RECT 2575.5400 2805.3600 2577.1400 2805.8400 ;
        RECT 2530.5400 2794.4800 2532.1400 2794.9600 ;
        RECT 2530.5400 2799.9200 2532.1400 2800.4000 ;
        RECT 2530.5400 2805.3600 2532.1400 2805.8400 ;
        RECT 2575.5400 2783.6000 2577.1400 2784.0800 ;
        RECT 2575.5400 2789.0400 2577.1400 2789.5200 ;
        RECT 2575.5400 2767.2800 2577.1400 2767.7600 ;
        RECT 2575.5400 2772.7200 2577.1400 2773.2000 ;
        RECT 2575.5400 2778.1600 2577.1400 2778.6400 ;
        RECT 2530.5400 2783.6000 2532.1400 2784.0800 ;
        RECT 2530.5400 2789.0400 2532.1400 2789.5200 ;
        RECT 2530.5400 2767.2800 2532.1400 2767.7600 ;
        RECT 2530.5400 2772.7200 2532.1400 2773.2000 ;
        RECT 2530.5400 2778.1600 2532.1400 2778.6400 ;
        RECT 2485.5400 2794.4800 2487.1400 2794.9600 ;
        RECT 2485.5400 2799.9200 2487.1400 2800.4000 ;
        RECT 2473.7800 2799.9200 2476.7800 2800.4000 ;
        RECT 2473.7800 2794.4800 2476.7800 2794.9600 ;
        RECT 2473.7800 2805.3600 2476.7800 2805.8400 ;
        RECT 2485.5400 2805.3600 2487.1400 2805.8400 ;
        RECT 2485.5400 2783.6000 2487.1400 2784.0800 ;
        RECT 2485.5400 2789.0400 2487.1400 2789.5200 ;
        RECT 2473.7800 2789.0400 2476.7800 2789.5200 ;
        RECT 2473.7800 2783.6000 2476.7800 2784.0800 ;
        RECT 2485.5400 2767.2800 2487.1400 2767.7600 ;
        RECT 2485.5400 2772.7200 2487.1400 2773.2000 ;
        RECT 2473.7800 2772.7200 2476.7800 2773.2000 ;
        RECT 2473.7800 2767.2800 2476.7800 2767.7600 ;
        RECT 2473.7800 2778.1600 2476.7800 2778.6400 ;
        RECT 2485.5400 2778.1600 2487.1400 2778.6400 ;
        RECT 2575.5400 2750.9600 2577.1400 2751.4400 ;
        RECT 2575.5400 2756.4000 2577.1400 2756.8800 ;
        RECT 2575.5400 2761.8400 2577.1400 2762.3200 ;
        RECT 2575.5400 2740.0800 2577.1400 2740.5600 ;
        RECT 2575.5400 2745.5200 2577.1400 2746.0000 ;
        RECT 2530.5400 2750.9600 2532.1400 2751.4400 ;
        RECT 2530.5400 2756.4000 2532.1400 2756.8800 ;
        RECT 2530.5400 2761.8400 2532.1400 2762.3200 ;
        RECT 2530.5400 2740.0800 2532.1400 2740.5600 ;
        RECT 2530.5400 2745.5200 2532.1400 2746.0000 ;
        RECT 2575.5400 2723.7600 2577.1400 2724.2400 ;
        RECT 2575.5400 2729.2000 2577.1400 2729.6800 ;
        RECT 2575.5400 2734.6400 2577.1400 2735.1200 ;
        RECT 2575.5400 2712.8800 2577.1400 2713.3600 ;
        RECT 2575.5400 2718.3200 2577.1400 2718.8000 ;
        RECT 2530.5400 2723.7600 2532.1400 2724.2400 ;
        RECT 2530.5400 2729.2000 2532.1400 2729.6800 ;
        RECT 2530.5400 2734.6400 2532.1400 2735.1200 ;
        RECT 2530.5400 2712.8800 2532.1400 2713.3600 ;
        RECT 2530.5400 2718.3200 2532.1400 2718.8000 ;
        RECT 2485.5400 2750.9600 2487.1400 2751.4400 ;
        RECT 2485.5400 2756.4000 2487.1400 2756.8800 ;
        RECT 2485.5400 2761.8400 2487.1400 2762.3200 ;
        RECT 2473.7800 2750.9600 2476.7800 2751.4400 ;
        RECT 2473.7800 2756.4000 2476.7800 2756.8800 ;
        RECT 2473.7800 2761.8400 2476.7800 2762.3200 ;
        RECT 2485.5400 2740.0800 2487.1400 2740.5600 ;
        RECT 2485.5400 2745.5200 2487.1400 2746.0000 ;
        RECT 2473.7800 2740.0800 2476.7800 2740.5600 ;
        RECT 2473.7800 2745.5200 2476.7800 2746.0000 ;
        RECT 2485.5400 2723.7600 2487.1400 2724.2400 ;
        RECT 2485.5400 2729.2000 2487.1400 2729.6800 ;
        RECT 2485.5400 2734.6400 2487.1400 2735.1200 ;
        RECT 2473.7800 2723.7600 2476.7800 2724.2400 ;
        RECT 2473.7800 2729.2000 2476.7800 2729.6800 ;
        RECT 2473.7800 2734.6400 2476.7800 2735.1200 ;
        RECT 2485.5400 2712.8800 2487.1400 2713.3600 ;
        RECT 2485.5400 2718.3200 2487.1400 2718.8000 ;
        RECT 2473.7800 2712.8800 2476.7800 2713.3600 ;
        RECT 2473.7800 2718.3200 2476.7800 2718.8000 ;
        RECT 2677.8800 2696.5600 2680.8800 2697.0400 ;
        RECT 2677.8800 2702.0000 2680.8800 2702.4800 ;
        RECT 2677.8800 2707.4400 2680.8800 2707.9200 ;
        RECT 2665.5400 2696.5600 2667.1400 2697.0400 ;
        RECT 2665.5400 2702.0000 2667.1400 2702.4800 ;
        RECT 2665.5400 2707.4400 2667.1400 2707.9200 ;
        RECT 2677.8800 2685.6800 2680.8800 2686.1600 ;
        RECT 2677.8800 2691.1200 2680.8800 2691.6000 ;
        RECT 2665.5400 2685.6800 2667.1400 2686.1600 ;
        RECT 2665.5400 2691.1200 2667.1400 2691.6000 ;
        RECT 2677.8800 2669.3600 2680.8800 2669.8400 ;
        RECT 2677.8800 2674.8000 2680.8800 2675.2800 ;
        RECT 2677.8800 2680.2400 2680.8800 2680.7200 ;
        RECT 2665.5400 2669.3600 2667.1400 2669.8400 ;
        RECT 2665.5400 2674.8000 2667.1400 2675.2800 ;
        RECT 2665.5400 2680.2400 2667.1400 2680.7200 ;
        RECT 2677.8800 2658.4800 2680.8800 2658.9600 ;
        RECT 2677.8800 2663.9200 2680.8800 2664.4000 ;
        RECT 2665.5400 2658.4800 2667.1400 2658.9600 ;
        RECT 2665.5400 2663.9200 2667.1400 2664.4000 ;
        RECT 2620.5400 2696.5600 2622.1400 2697.0400 ;
        RECT 2620.5400 2702.0000 2622.1400 2702.4800 ;
        RECT 2620.5400 2707.4400 2622.1400 2707.9200 ;
        RECT 2620.5400 2685.6800 2622.1400 2686.1600 ;
        RECT 2620.5400 2691.1200 2622.1400 2691.6000 ;
        RECT 2620.5400 2669.3600 2622.1400 2669.8400 ;
        RECT 2620.5400 2674.8000 2622.1400 2675.2800 ;
        RECT 2620.5400 2680.2400 2622.1400 2680.7200 ;
        RECT 2620.5400 2658.4800 2622.1400 2658.9600 ;
        RECT 2620.5400 2663.9200 2622.1400 2664.4000 ;
        RECT 2677.8800 2642.1600 2680.8800 2642.6400 ;
        RECT 2677.8800 2647.6000 2680.8800 2648.0800 ;
        RECT 2677.8800 2653.0400 2680.8800 2653.5200 ;
        RECT 2665.5400 2642.1600 2667.1400 2642.6400 ;
        RECT 2665.5400 2647.6000 2667.1400 2648.0800 ;
        RECT 2665.5400 2653.0400 2667.1400 2653.5200 ;
        RECT 2677.8800 2631.2800 2680.8800 2631.7600 ;
        RECT 2677.8800 2636.7200 2680.8800 2637.2000 ;
        RECT 2665.5400 2631.2800 2667.1400 2631.7600 ;
        RECT 2665.5400 2636.7200 2667.1400 2637.2000 ;
        RECT 2677.8800 2614.9600 2680.8800 2615.4400 ;
        RECT 2677.8800 2620.4000 2680.8800 2620.8800 ;
        RECT 2677.8800 2625.8400 2680.8800 2626.3200 ;
        RECT 2665.5400 2614.9600 2667.1400 2615.4400 ;
        RECT 2665.5400 2620.4000 2667.1400 2620.8800 ;
        RECT 2665.5400 2625.8400 2667.1400 2626.3200 ;
        RECT 2677.8800 2609.5200 2680.8800 2610.0000 ;
        RECT 2665.5400 2609.5200 2667.1400 2610.0000 ;
        RECT 2620.5400 2642.1600 2622.1400 2642.6400 ;
        RECT 2620.5400 2647.6000 2622.1400 2648.0800 ;
        RECT 2620.5400 2653.0400 2622.1400 2653.5200 ;
        RECT 2620.5400 2631.2800 2622.1400 2631.7600 ;
        RECT 2620.5400 2636.7200 2622.1400 2637.2000 ;
        RECT 2620.5400 2614.9600 2622.1400 2615.4400 ;
        RECT 2620.5400 2620.4000 2622.1400 2620.8800 ;
        RECT 2620.5400 2625.8400 2622.1400 2626.3200 ;
        RECT 2620.5400 2609.5200 2622.1400 2610.0000 ;
        RECT 2575.5400 2696.5600 2577.1400 2697.0400 ;
        RECT 2575.5400 2702.0000 2577.1400 2702.4800 ;
        RECT 2575.5400 2707.4400 2577.1400 2707.9200 ;
        RECT 2575.5400 2685.6800 2577.1400 2686.1600 ;
        RECT 2575.5400 2691.1200 2577.1400 2691.6000 ;
        RECT 2530.5400 2696.5600 2532.1400 2697.0400 ;
        RECT 2530.5400 2702.0000 2532.1400 2702.4800 ;
        RECT 2530.5400 2707.4400 2532.1400 2707.9200 ;
        RECT 2530.5400 2685.6800 2532.1400 2686.1600 ;
        RECT 2530.5400 2691.1200 2532.1400 2691.6000 ;
        RECT 2575.5400 2669.3600 2577.1400 2669.8400 ;
        RECT 2575.5400 2674.8000 2577.1400 2675.2800 ;
        RECT 2575.5400 2680.2400 2577.1400 2680.7200 ;
        RECT 2575.5400 2658.4800 2577.1400 2658.9600 ;
        RECT 2575.5400 2663.9200 2577.1400 2664.4000 ;
        RECT 2530.5400 2669.3600 2532.1400 2669.8400 ;
        RECT 2530.5400 2674.8000 2532.1400 2675.2800 ;
        RECT 2530.5400 2680.2400 2532.1400 2680.7200 ;
        RECT 2530.5400 2658.4800 2532.1400 2658.9600 ;
        RECT 2530.5400 2663.9200 2532.1400 2664.4000 ;
        RECT 2485.5400 2696.5600 2487.1400 2697.0400 ;
        RECT 2485.5400 2702.0000 2487.1400 2702.4800 ;
        RECT 2485.5400 2707.4400 2487.1400 2707.9200 ;
        RECT 2473.7800 2696.5600 2476.7800 2697.0400 ;
        RECT 2473.7800 2702.0000 2476.7800 2702.4800 ;
        RECT 2473.7800 2707.4400 2476.7800 2707.9200 ;
        RECT 2485.5400 2685.6800 2487.1400 2686.1600 ;
        RECT 2485.5400 2691.1200 2487.1400 2691.6000 ;
        RECT 2473.7800 2685.6800 2476.7800 2686.1600 ;
        RECT 2473.7800 2691.1200 2476.7800 2691.6000 ;
        RECT 2485.5400 2669.3600 2487.1400 2669.8400 ;
        RECT 2485.5400 2674.8000 2487.1400 2675.2800 ;
        RECT 2485.5400 2680.2400 2487.1400 2680.7200 ;
        RECT 2473.7800 2669.3600 2476.7800 2669.8400 ;
        RECT 2473.7800 2674.8000 2476.7800 2675.2800 ;
        RECT 2473.7800 2680.2400 2476.7800 2680.7200 ;
        RECT 2485.5400 2658.4800 2487.1400 2658.9600 ;
        RECT 2485.5400 2663.9200 2487.1400 2664.4000 ;
        RECT 2473.7800 2658.4800 2476.7800 2658.9600 ;
        RECT 2473.7800 2663.9200 2476.7800 2664.4000 ;
        RECT 2575.5400 2642.1600 2577.1400 2642.6400 ;
        RECT 2575.5400 2647.6000 2577.1400 2648.0800 ;
        RECT 2575.5400 2653.0400 2577.1400 2653.5200 ;
        RECT 2575.5400 2631.2800 2577.1400 2631.7600 ;
        RECT 2575.5400 2636.7200 2577.1400 2637.2000 ;
        RECT 2530.5400 2642.1600 2532.1400 2642.6400 ;
        RECT 2530.5400 2647.6000 2532.1400 2648.0800 ;
        RECT 2530.5400 2653.0400 2532.1400 2653.5200 ;
        RECT 2530.5400 2631.2800 2532.1400 2631.7600 ;
        RECT 2530.5400 2636.7200 2532.1400 2637.2000 ;
        RECT 2575.5400 2614.9600 2577.1400 2615.4400 ;
        RECT 2575.5400 2620.4000 2577.1400 2620.8800 ;
        RECT 2575.5400 2625.8400 2577.1400 2626.3200 ;
        RECT 2575.5400 2609.5200 2577.1400 2610.0000 ;
        RECT 2530.5400 2614.9600 2532.1400 2615.4400 ;
        RECT 2530.5400 2620.4000 2532.1400 2620.8800 ;
        RECT 2530.5400 2625.8400 2532.1400 2626.3200 ;
        RECT 2530.5400 2609.5200 2532.1400 2610.0000 ;
        RECT 2485.5400 2642.1600 2487.1400 2642.6400 ;
        RECT 2485.5400 2647.6000 2487.1400 2648.0800 ;
        RECT 2485.5400 2653.0400 2487.1400 2653.5200 ;
        RECT 2473.7800 2642.1600 2476.7800 2642.6400 ;
        RECT 2473.7800 2647.6000 2476.7800 2648.0800 ;
        RECT 2473.7800 2653.0400 2476.7800 2653.5200 ;
        RECT 2485.5400 2631.2800 2487.1400 2631.7600 ;
        RECT 2485.5400 2636.7200 2487.1400 2637.2000 ;
        RECT 2473.7800 2631.2800 2476.7800 2631.7600 ;
        RECT 2473.7800 2636.7200 2476.7800 2637.2000 ;
        RECT 2485.5400 2614.9600 2487.1400 2615.4400 ;
        RECT 2485.5400 2620.4000 2487.1400 2620.8800 ;
        RECT 2485.5400 2625.8400 2487.1400 2626.3200 ;
        RECT 2473.7800 2614.9600 2476.7800 2615.4400 ;
        RECT 2473.7800 2620.4000 2476.7800 2620.8800 ;
        RECT 2473.7800 2625.8400 2476.7800 2626.3200 ;
        RECT 2473.7800 2609.5200 2476.7800 2610.0000 ;
        RECT 2485.5400 2609.5200 2487.1400 2610.0000 ;
        RECT 2473.7800 2814.4300 2680.8800 2817.4300 ;
        RECT 2473.7800 2601.3300 2680.8800 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 2371.6900 2667.1400 2587.7900 ;
        RECT 2620.5400 2371.6900 2622.1400 2587.7900 ;
        RECT 2575.5400 2371.6900 2577.1400 2587.7900 ;
        RECT 2530.5400 2371.6900 2532.1400 2587.7900 ;
        RECT 2485.5400 2371.6900 2487.1400 2587.7900 ;
        RECT 2677.8800 2371.6900 2680.8800 2587.7900 ;
        RECT 2473.7800 2371.6900 2476.7800 2587.7900 ;
      LAYER met3 ;
        RECT 2677.8800 2564.8400 2680.8800 2565.3200 ;
        RECT 2677.8800 2570.2800 2680.8800 2570.7600 ;
        RECT 2665.5400 2564.8400 2667.1400 2565.3200 ;
        RECT 2665.5400 2570.2800 2667.1400 2570.7600 ;
        RECT 2677.8800 2575.7200 2680.8800 2576.2000 ;
        RECT 2665.5400 2575.7200 2667.1400 2576.2000 ;
        RECT 2677.8800 2553.9600 2680.8800 2554.4400 ;
        RECT 2677.8800 2559.4000 2680.8800 2559.8800 ;
        RECT 2665.5400 2553.9600 2667.1400 2554.4400 ;
        RECT 2665.5400 2559.4000 2667.1400 2559.8800 ;
        RECT 2677.8800 2537.6400 2680.8800 2538.1200 ;
        RECT 2677.8800 2543.0800 2680.8800 2543.5600 ;
        RECT 2665.5400 2537.6400 2667.1400 2538.1200 ;
        RECT 2665.5400 2543.0800 2667.1400 2543.5600 ;
        RECT 2677.8800 2548.5200 2680.8800 2549.0000 ;
        RECT 2665.5400 2548.5200 2667.1400 2549.0000 ;
        RECT 2620.5400 2564.8400 2622.1400 2565.3200 ;
        RECT 2620.5400 2570.2800 2622.1400 2570.7600 ;
        RECT 2620.5400 2575.7200 2622.1400 2576.2000 ;
        RECT 2620.5400 2553.9600 2622.1400 2554.4400 ;
        RECT 2620.5400 2559.4000 2622.1400 2559.8800 ;
        RECT 2620.5400 2537.6400 2622.1400 2538.1200 ;
        RECT 2620.5400 2543.0800 2622.1400 2543.5600 ;
        RECT 2620.5400 2548.5200 2622.1400 2549.0000 ;
        RECT 2677.8800 2521.3200 2680.8800 2521.8000 ;
        RECT 2677.8800 2526.7600 2680.8800 2527.2400 ;
        RECT 2677.8800 2532.2000 2680.8800 2532.6800 ;
        RECT 2665.5400 2521.3200 2667.1400 2521.8000 ;
        RECT 2665.5400 2526.7600 2667.1400 2527.2400 ;
        RECT 2665.5400 2532.2000 2667.1400 2532.6800 ;
        RECT 2677.8800 2510.4400 2680.8800 2510.9200 ;
        RECT 2677.8800 2515.8800 2680.8800 2516.3600 ;
        RECT 2665.5400 2510.4400 2667.1400 2510.9200 ;
        RECT 2665.5400 2515.8800 2667.1400 2516.3600 ;
        RECT 2677.8800 2494.1200 2680.8800 2494.6000 ;
        RECT 2677.8800 2499.5600 2680.8800 2500.0400 ;
        RECT 2677.8800 2505.0000 2680.8800 2505.4800 ;
        RECT 2665.5400 2494.1200 2667.1400 2494.6000 ;
        RECT 2665.5400 2499.5600 2667.1400 2500.0400 ;
        RECT 2665.5400 2505.0000 2667.1400 2505.4800 ;
        RECT 2677.8800 2483.2400 2680.8800 2483.7200 ;
        RECT 2677.8800 2488.6800 2680.8800 2489.1600 ;
        RECT 2665.5400 2483.2400 2667.1400 2483.7200 ;
        RECT 2665.5400 2488.6800 2667.1400 2489.1600 ;
        RECT 2620.5400 2521.3200 2622.1400 2521.8000 ;
        RECT 2620.5400 2526.7600 2622.1400 2527.2400 ;
        RECT 2620.5400 2532.2000 2622.1400 2532.6800 ;
        RECT 2620.5400 2510.4400 2622.1400 2510.9200 ;
        RECT 2620.5400 2515.8800 2622.1400 2516.3600 ;
        RECT 2620.5400 2494.1200 2622.1400 2494.6000 ;
        RECT 2620.5400 2499.5600 2622.1400 2500.0400 ;
        RECT 2620.5400 2505.0000 2622.1400 2505.4800 ;
        RECT 2620.5400 2483.2400 2622.1400 2483.7200 ;
        RECT 2620.5400 2488.6800 2622.1400 2489.1600 ;
        RECT 2575.5400 2564.8400 2577.1400 2565.3200 ;
        RECT 2575.5400 2570.2800 2577.1400 2570.7600 ;
        RECT 2575.5400 2575.7200 2577.1400 2576.2000 ;
        RECT 2530.5400 2564.8400 2532.1400 2565.3200 ;
        RECT 2530.5400 2570.2800 2532.1400 2570.7600 ;
        RECT 2530.5400 2575.7200 2532.1400 2576.2000 ;
        RECT 2575.5400 2553.9600 2577.1400 2554.4400 ;
        RECT 2575.5400 2559.4000 2577.1400 2559.8800 ;
        RECT 2575.5400 2537.6400 2577.1400 2538.1200 ;
        RECT 2575.5400 2543.0800 2577.1400 2543.5600 ;
        RECT 2575.5400 2548.5200 2577.1400 2549.0000 ;
        RECT 2530.5400 2553.9600 2532.1400 2554.4400 ;
        RECT 2530.5400 2559.4000 2532.1400 2559.8800 ;
        RECT 2530.5400 2537.6400 2532.1400 2538.1200 ;
        RECT 2530.5400 2543.0800 2532.1400 2543.5600 ;
        RECT 2530.5400 2548.5200 2532.1400 2549.0000 ;
        RECT 2485.5400 2564.8400 2487.1400 2565.3200 ;
        RECT 2485.5400 2570.2800 2487.1400 2570.7600 ;
        RECT 2473.7800 2570.2800 2476.7800 2570.7600 ;
        RECT 2473.7800 2564.8400 2476.7800 2565.3200 ;
        RECT 2473.7800 2575.7200 2476.7800 2576.2000 ;
        RECT 2485.5400 2575.7200 2487.1400 2576.2000 ;
        RECT 2485.5400 2553.9600 2487.1400 2554.4400 ;
        RECT 2485.5400 2559.4000 2487.1400 2559.8800 ;
        RECT 2473.7800 2559.4000 2476.7800 2559.8800 ;
        RECT 2473.7800 2553.9600 2476.7800 2554.4400 ;
        RECT 2485.5400 2537.6400 2487.1400 2538.1200 ;
        RECT 2485.5400 2543.0800 2487.1400 2543.5600 ;
        RECT 2473.7800 2543.0800 2476.7800 2543.5600 ;
        RECT 2473.7800 2537.6400 2476.7800 2538.1200 ;
        RECT 2473.7800 2548.5200 2476.7800 2549.0000 ;
        RECT 2485.5400 2548.5200 2487.1400 2549.0000 ;
        RECT 2575.5400 2521.3200 2577.1400 2521.8000 ;
        RECT 2575.5400 2526.7600 2577.1400 2527.2400 ;
        RECT 2575.5400 2532.2000 2577.1400 2532.6800 ;
        RECT 2575.5400 2510.4400 2577.1400 2510.9200 ;
        RECT 2575.5400 2515.8800 2577.1400 2516.3600 ;
        RECT 2530.5400 2521.3200 2532.1400 2521.8000 ;
        RECT 2530.5400 2526.7600 2532.1400 2527.2400 ;
        RECT 2530.5400 2532.2000 2532.1400 2532.6800 ;
        RECT 2530.5400 2510.4400 2532.1400 2510.9200 ;
        RECT 2530.5400 2515.8800 2532.1400 2516.3600 ;
        RECT 2575.5400 2494.1200 2577.1400 2494.6000 ;
        RECT 2575.5400 2499.5600 2577.1400 2500.0400 ;
        RECT 2575.5400 2505.0000 2577.1400 2505.4800 ;
        RECT 2575.5400 2483.2400 2577.1400 2483.7200 ;
        RECT 2575.5400 2488.6800 2577.1400 2489.1600 ;
        RECT 2530.5400 2494.1200 2532.1400 2494.6000 ;
        RECT 2530.5400 2499.5600 2532.1400 2500.0400 ;
        RECT 2530.5400 2505.0000 2532.1400 2505.4800 ;
        RECT 2530.5400 2483.2400 2532.1400 2483.7200 ;
        RECT 2530.5400 2488.6800 2532.1400 2489.1600 ;
        RECT 2485.5400 2521.3200 2487.1400 2521.8000 ;
        RECT 2485.5400 2526.7600 2487.1400 2527.2400 ;
        RECT 2485.5400 2532.2000 2487.1400 2532.6800 ;
        RECT 2473.7800 2521.3200 2476.7800 2521.8000 ;
        RECT 2473.7800 2526.7600 2476.7800 2527.2400 ;
        RECT 2473.7800 2532.2000 2476.7800 2532.6800 ;
        RECT 2485.5400 2510.4400 2487.1400 2510.9200 ;
        RECT 2485.5400 2515.8800 2487.1400 2516.3600 ;
        RECT 2473.7800 2510.4400 2476.7800 2510.9200 ;
        RECT 2473.7800 2515.8800 2476.7800 2516.3600 ;
        RECT 2485.5400 2494.1200 2487.1400 2494.6000 ;
        RECT 2485.5400 2499.5600 2487.1400 2500.0400 ;
        RECT 2485.5400 2505.0000 2487.1400 2505.4800 ;
        RECT 2473.7800 2494.1200 2476.7800 2494.6000 ;
        RECT 2473.7800 2499.5600 2476.7800 2500.0400 ;
        RECT 2473.7800 2505.0000 2476.7800 2505.4800 ;
        RECT 2485.5400 2483.2400 2487.1400 2483.7200 ;
        RECT 2485.5400 2488.6800 2487.1400 2489.1600 ;
        RECT 2473.7800 2483.2400 2476.7800 2483.7200 ;
        RECT 2473.7800 2488.6800 2476.7800 2489.1600 ;
        RECT 2677.8800 2466.9200 2680.8800 2467.4000 ;
        RECT 2677.8800 2472.3600 2680.8800 2472.8400 ;
        RECT 2677.8800 2477.8000 2680.8800 2478.2800 ;
        RECT 2665.5400 2466.9200 2667.1400 2467.4000 ;
        RECT 2665.5400 2472.3600 2667.1400 2472.8400 ;
        RECT 2665.5400 2477.8000 2667.1400 2478.2800 ;
        RECT 2677.8800 2456.0400 2680.8800 2456.5200 ;
        RECT 2677.8800 2461.4800 2680.8800 2461.9600 ;
        RECT 2665.5400 2456.0400 2667.1400 2456.5200 ;
        RECT 2665.5400 2461.4800 2667.1400 2461.9600 ;
        RECT 2677.8800 2439.7200 2680.8800 2440.2000 ;
        RECT 2677.8800 2445.1600 2680.8800 2445.6400 ;
        RECT 2677.8800 2450.6000 2680.8800 2451.0800 ;
        RECT 2665.5400 2439.7200 2667.1400 2440.2000 ;
        RECT 2665.5400 2445.1600 2667.1400 2445.6400 ;
        RECT 2665.5400 2450.6000 2667.1400 2451.0800 ;
        RECT 2677.8800 2428.8400 2680.8800 2429.3200 ;
        RECT 2677.8800 2434.2800 2680.8800 2434.7600 ;
        RECT 2665.5400 2428.8400 2667.1400 2429.3200 ;
        RECT 2665.5400 2434.2800 2667.1400 2434.7600 ;
        RECT 2620.5400 2466.9200 2622.1400 2467.4000 ;
        RECT 2620.5400 2472.3600 2622.1400 2472.8400 ;
        RECT 2620.5400 2477.8000 2622.1400 2478.2800 ;
        RECT 2620.5400 2456.0400 2622.1400 2456.5200 ;
        RECT 2620.5400 2461.4800 2622.1400 2461.9600 ;
        RECT 2620.5400 2439.7200 2622.1400 2440.2000 ;
        RECT 2620.5400 2445.1600 2622.1400 2445.6400 ;
        RECT 2620.5400 2450.6000 2622.1400 2451.0800 ;
        RECT 2620.5400 2428.8400 2622.1400 2429.3200 ;
        RECT 2620.5400 2434.2800 2622.1400 2434.7600 ;
        RECT 2677.8800 2412.5200 2680.8800 2413.0000 ;
        RECT 2677.8800 2417.9600 2680.8800 2418.4400 ;
        RECT 2677.8800 2423.4000 2680.8800 2423.8800 ;
        RECT 2665.5400 2412.5200 2667.1400 2413.0000 ;
        RECT 2665.5400 2417.9600 2667.1400 2418.4400 ;
        RECT 2665.5400 2423.4000 2667.1400 2423.8800 ;
        RECT 2677.8800 2401.6400 2680.8800 2402.1200 ;
        RECT 2677.8800 2407.0800 2680.8800 2407.5600 ;
        RECT 2665.5400 2401.6400 2667.1400 2402.1200 ;
        RECT 2665.5400 2407.0800 2667.1400 2407.5600 ;
        RECT 2677.8800 2385.3200 2680.8800 2385.8000 ;
        RECT 2677.8800 2390.7600 2680.8800 2391.2400 ;
        RECT 2677.8800 2396.2000 2680.8800 2396.6800 ;
        RECT 2665.5400 2385.3200 2667.1400 2385.8000 ;
        RECT 2665.5400 2390.7600 2667.1400 2391.2400 ;
        RECT 2665.5400 2396.2000 2667.1400 2396.6800 ;
        RECT 2677.8800 2379.8800 2680.8800 2380.3600 ;
        RECT 2665.5400 2379.8800 2667.1400 2380.3600 ;
        RECT 2620.5400 2412.5200 2622.1400 2413.0000 ;
        RECT 2620.5400 2417.9600 2622.1400 2418.4400 ;
        RECT 2620.5400 2423.4000 2622.1400 2423.8800 ;
        RECT 2620.5400 2401.6400 2622.1400 2402.1200 ;
        RECT 2620.5400 2407.0800 2622.1400 2407.5600 ;
        RECT 2620.5400 2385.3200 2622.1400 2385.8000 ;
        RECT 2620.5400 2390.7600 2622.1400 2391.2400 ;
        RECT 2620.5400 2396.2000 2622.1400 2396.6800 ;
        RECT 2620.5400 2379.8800 2622.1400 2380.3600 ;
        RECT 2575.5400 2466.9200 2577.1400 2467.4000 ;
        RECT 2575.5400 2472.3600 2577.1400 2472.8400 ;
        RECT 2575.5400 2477.8000 2577.1400 2478.2800 ;
        RECT 2575.5400 2456.0400 2577.1400 2456.5200 ;
        RECT 2575.5400 2461.4800 2577.1400 2461.9600 ;
        RECT 2530.5400 2466.9200 2532.1400 2467.4000 ;
        RECT 2530.5400 2472.3600 2532.1400 2472.8400 ;
        RECT 2530.5400 2477.8000 2532.1400 2478.2800 ;
        RECT 2530.5400 2456.0400 2532.1400 2456.5200 ;
        RECT 2530.5400 2461.4800 2532.1400 2461.9600 ;
        RECT 2575.5400 2439.7200 2577.1400 2440.2000 ;
        RECT 2575.5400 2445.1600 2577.1400 2445.6400 ;
        RECT 2575.5400 2450.6000 2577.1400 2451.0800 ;
        RECT 2575.5400 2428.8400 2577.1400 2429.3200 ;
        RECT 2575.5400 2434.2800 2577.1400 2434.7600 ;
        RECT 2530.5400 2439.7200 2532.1400 2440.2000 ;
        RECT 2530.5400 2445.1600 2532.1400 2445.6400 ;
        RECT 2530.5400 2450.6000 2532.1400 2451.0800 ;
        RECT 2530.5400 2428.8400 2532.1400 2429.3200 ;
        RECT 2530.5400 2434.2800 2532.1400 2434.7600 ;
        RECT 2485.5400 2466.9200 2487.1400 2467.4000 ;
        RECT 2485.5400 2472.3600 2487.1400 2472.8400 ;
        RECT 2485.5400 2477.8000 2487.1400 2478.2800 ;
        RECT 2473.7800 2466.9200 2476.7800 2467.4000 ;
        RECT 2473.7800 2472.3600 2476.7800 2472.8400 ;
        RECT 2473.7800 2477.8000 2476.7800 2478.2800 ;
        RECT 2485.5400 2456.0400 2487.1400 2456.5200 ;
        RECT 2485.5400 2461.4800 2487.1400 2461.9600 ;
        RECT 2473.7800 2456.0400 2476.7800 2456.5200 ;
        RECT 2473.7800 2461.4800 2476.7800 2461.9600 ;
        RECT 2485.5400 2439.7200 2487.1400 2440.2000 ;
        RECT 2485.5400 2445.1600 2487.1400 2445.6400 ;
        RECT 2485.5400 2450.6000 2487.1400 2451.0800 ;
        RECT 2473.7800 2439.7200 2476.7800 2440.2000 ;
        RECT 2473.7800 2445.1600 2476.7800 2445.6400 ;
        RECT 2473.7800 2450.6000 2476.7800 2451.0800 ;
        RECT 2485.5400 2428.8400 2487.1400 2429.3200 ;
        RECT 2485.5400 2434.2800 2487.1400 2434.7600 ;
        RECT 2473.7800 2428.8400 2476.7800 2429.3200 ;
        RECT 2473.7800 2434.2800 2476.7800 2434.7600 ;
        RECT 2575.5400 2412.5200 2577.1400 2413.0000 ;
        RECT 2575.5400 2417.9600 2577.1400 2418.4400 ;
        RECT 2575.5400 2423.4000 2577.1400 2423.8800 ;
        RECT 2575.5400 2401.6400 2577.1400 2402.1200 ;
        RECT 2575.5400 2407.0800 2577.1400 2407.5600 ;
        RECT 2530.5400 2412.5200 2532.1400 2413.0000 ;
        RECT 2530.5400 2417.9600 2532.1400 2418.4400 ;
        RECT 2530.5400 2423.4000 2532.1400 2423.8800 ;
        RECT 2530.5400 2401.6400 2532.1400 2402.1200 ;
        RECT 2530.5400 2407.0800 2532.1400 2407.5600 ;
        RECT 2575.5400 2385.3200 2577.1400 2385.8000 ;
        RECT 2575.5400 2390.7600 2577.1400 2391.2400 ;
        RECT 2575.5400 2396.2000 2577.1400 2396.6800 ;
        RECT 2575.5400 2379.8800 2577.1400 2380.3600 ;
        RECT 2530.5400 2385.3200 2532.1400 2385.8000 ;
        RECT 2530.5400 2390.7600 2532.1400 2391.2400 ;
        RECT 2530.5400 2396.2000 2532.1400 2396.6800 ;
        RECT 2530.5400 2379.8800 2532.1400 2380.3600 ;
        RECT 2485.5400 2412.5200 2487.1400 2413.0000 ;
        RECT 2485.5400 2417.9600 2487.1400 2418.4400 ;
        RECT 2485.5400 2423.4000 2487.1400 2423.8800 ;
        RECT 2473.7800 2412.5200 2476.7800 2413.0000 ;
        RECT 2473.7800 2417.9600 2476.7800 2418.4400 ;
        RECT 2473.7800 2423.4000 2476.7800 2423.8800 ;
        RECT 2485.5400 2401.6400 2487.1400 2402.1200 ;
        RECT 2485.5400 2407.0800 2487.1400 2407.5600 ;
        RECT 2473.7800 2401.6400 2476.7800 2402.1200 ;
        RECT 2473.7800 2407.0800 2476.7800 2407.5600 ;
        RECT 2485.5400 2385.3200 2487.1400 2385.8000 ;
        RECT 2485.5400 2390.7600 2487.1400 2391.2400 ;
        RECT 2485.5400 2396.2000 2487.1400 2396.6800 ;
        RECT 2473.7800 2385.3200 2476.7800 2385.8000 ;
        RECT 2473.7800 2390.7600 2476.7800 2391.2400 ;
        RECT 2473.7800 2396.2000 2476.7800 2396.6800 ;
        RECT 2473.7800 2379.8800 2476.7800 2380.3600 ;
        RECT 2485.5400 2379.8800 2487.1400 2380.3600 ;
        RECT 2473.7800 2584.7900 2680.8800 2587.7900 ;
        RECT 2473.7800 2371.6900 2680.8800 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 2142.0500 2667.1400 2358.1500 ;
        RECT 2620.5400 2142.0500 2622.1400 2358.1500 ;
        RECT 2575.5400 2142.0500 2577.1400 2358.1500 ;
        RECT 2530.5400 2142.0500 2532.1400 2358.1500 ;
        RECT 2485.5400 2142.0500 2487.1400 2358.1500 ;
        RECT 2677.8800 2142.0500 2680.8800 2358.1500 ;
        RECT 2473.7800 2142.0500 2476.7800 2358.1500 ;
      LAYER met3 ;
        RECT 2677.8800 2335.2000 2680.8800 2335.6800 ;
        RECT 2677.8800 2340.6400 2680.8800 2341.1200 ;
        RECT 2665.5400 2335.2000 2667.1400 2335.6800 ;
        RECT 2665.5400 2340.6400 2667.1400 2341.1200 ;
        RECT 2677.8800 2346.0800 2680.8800 2346.5600 ;
        RECT 2665.5400 2346.0800 2667.1400 2346.5600 ;
        RECT 2677.8800 2324.3200 2680.8800 2324.8000 ;
        RECT 2677.8800 2329.7600 2680.8800 2330.2400 ;
        RECT 2665.5400 2324.3200 2667.1400 2324.8000 ;
        RECT 2665.5400 2329.7600 2667.1400 2330.2400 ;
        RECT 2677.8800 2308.0000 2680.8800 2308.4800 ;
        RECT 2677.8800 2313.4400 2680.8800 2313.9200 ;
        RECT 2665.5400 2308.0000 2667.1400 2308.4800 ;
        RECT 2665.5400 2313.4400 2667.1400 2313.9200 ;
        RECT 2677.8800 2318.8800 2680.8800 2319.3600 ;
        RECT 2665.5400 2318.8800 2667.1400 2319.3600 ;
        RECT 2620.5400 2335.2000 2622.1400 2335.6800 ;
        RECT 2620.5400 2340.6400 2622.1400 2341.1200 ;
        RECT 2620.5400 2346.0800 2622.1400 2346.5600 ;
        RECT 2620.5400 2324.3200 2622.1400 2324.8000 ;
        RECT 2620.5400 2329.7600 2622.1400 2330.2400 ;
        RECT 2620.5400 2308.0000 2622.1400 2308.4800 ;
        RECT 2620.5400 2313.4400 2622.1400 2313.9200 ;
        RECT 2620.5400 2318.8800 2622.1400 2319.3600 ;
        RECT 2677.8800 2291.6800 2680.8800 2292.1600 ;
        RECT 2677.8800 2297.1200 2680.8800 2297.6000 ;
        RECT 2677.8800 2302.5600 2680.8800 2303.0400 ;
        RECT 2665.5400 2291.6800 2667.1400 2292.1600 ;
        RECT 2665.5400 2297.1200 2667.1400 2297.6000 ;
        RECT 2665.5400 2302.5600 2667.1400 2303.0400 ;
        RECT 2677.8800 2280.8000 2680.8800 2281.2800 ;
        RECT 2677.8800 2286.2400 2680.8800 2286.7200 ;
        RECT 2665.5400 2280.8000 2667.1400 2281.2800 ;
        RECT 2665.5400 2286.2400 2667.1400 2286.7200 ;
        RECT 2677.8800 2264.4800 2680.8800 2264.9600 ;
        RECT 2677.8800 2269.9200 2680.8800 2270.4000 ;
        RECT 2677.8800 2275.3600 2680.8800 2275.8400 ;
        RECT 2665.5400 2264.4800 2667.1400 2264.9600 ;
        RECT 2665.5400 2269.9200 2667.1400 2270.4000 ;
        RECT 2665.5400 2275.3600 2667.1400 2275.8400 ;
        RECT 2677.8800 2253.6000 2680.8800 2254.0800 ;
        RECT 2677.8800 2259.0400 2680.8800 2259.5200 ;
        RECT 2665.5400 2253.6000 2667.1400 2254.0800 ;
        RECT 2665.5400 2259.0400 2667.1400 2259.5200 ;
        RECT 2620.5400 2291.6800 2622.1400 2292.1600 ;
        RECT 2620.5400 2297.1200 2622.1400 2297.6000 ;
        RECT 2620.5400 2302.5600 2622.1400 2303.0400 ;
        RECT 2620.5400 2280.8000 2622.1400 2281.2800 ;
        RECT 2620.5400 2286.2400 2622.1400 2286.7200 ;
        RECT 2620.5400 2264.4800 2622.1400 2264.9600 ;
        RECT 2620.5400 2269.9200 2622.1400 2270.4000 ;
        RECT 2620.5400 2275.3600 2622.1400 2275.8400 ;
        RECT 2620.5400 2253.6000 2622.1400 2254.0800 ;
        RECT 2620.5400 2259.0400 2622.1400 2259.5200 ;
        RECT 2575.5400 2335.2000 2577.1400 2335.6800 ;
        RECT 2575.5400 2340.6400 2577.1400 2341.1200 ;
        RECT 2575.5400 2346.0800 2577.1400 2346.5600 ;
        RECT 2530.5400 2335.2000 2532.1400 2335.6800 ;
        RECT 2530.5400 2340.6400 2532.1400 2341.1200 ;
        RECT 2530.5400 2346.0800 2532.1400 2346.5600 ;
        RECT 2575.5400 2324.3200 2577.1400 2324.8000 ;
        RECT 2575.5400 2329.7600 2577.1400 2330.2400 ;
        RECT 2575.5400 2308.0000 2577.1400 2308.4800 ;
        RECT 2575.5400 2313.4400 2577.1400 2313.9200 ;
        RECT 2575.5400 2318.8800 2577.1400 2319.3600 ;
        RECT 2530.5400 2324.3200 2532.1400 2324.8000 ;
        RECT 2530.5400 2329.7600 2532.1400 2330.2400 ;
        RECT 2530.5400 2308.0000 2532.1400 2308.4800 ;
        RECT 2530.5400 2313.4400 2532.1400 2313.9200 ;
        RECT 2530.5400 2318.8800 2532.1400 2319.3600 ;
        RECT 2485.5400 2335.2000 2487.1400 2335.6800 ;
        RECT 2485.5400 2340.6400 2487.1400 2341.1200 ;
        RECT 2473.7800 2340.6400 2476.7800 2341.1200 ;
        RECT 2473.7800 2335.2000 2476.7800 2335.6800 ;
        RECT 2473.7800 2346.0800 2476.7800 2346.5600 ;
        RECT 2485.5400 2346.0800 2487.1400 2346.5600 ;
        RECT 2485.5400 2324.3200 2487.1400 2324.8000 ;
        RECT 2485.5400 2329.7600 2487.1400 2330.2400 ;
        RECT 2473.7800 2329.7600 2476.7800 2330.2400 ;
        RECT 2473.7800 2324.3200 2476.7800 2324.8000 ;
        RECT 2485.5400 2308.0000 2487.1400 2308.4800 ;
        RECT 2485.5400 2313.4400 2487.1400 2313.9200 ;
        RECT 2473.7800 2313.4400 2476.7800 2313.9200 ;
        RECT 2473.7800 2308.0000 2476.7800 2308.4800 ;
        RECT 2473.7800 2318.8800 2476.7800 2319.3600 ;
        RECT 2485.5400 2318.8800 2487.1400 2319.3600 ;
        RECT 2575.5400 2291.6800 2577.1400 2292.1600 ;
        RECT 2575.5400 2297.1200 2577.1400 2297.6000 ;
        RECT 2575.5400 2302.5600 2577.1400 2303.0400 ;
        RECT 2575.5400 2280.8000 2577.1400 2281.2800 ;
        RECT 2575.5400 2286.2400 2577.1400 2286.7200 ;
        RECT 2530.5400 2291.6800 2532.1400 2292.1600 ;
        RECT 2530.5400 2297.1200 2532.1400 2297.6000 ;
        RECT 2530.5400 2302.5600 2532.1400 2303.0400 ;
        RECT 2530.5400 2280.8000 2532.1400 2281.2800 ;
        RECT 2530.5400 2286.2400 2532.1400 2286.7200 ;
        RECT 2575.5400 2264.4800 2577.1400 2264.9600 ;
        RECT 2575.5400 2269.9200 2577.1400 2270.4000 ;
        RECT 2575.5400 2275.3600 2577.1400 2275.8400 ;
        RECT 2575.5400 2253.6000 2577.1400 2254.0800 ;
        RECT 2575.5400 2259.0400 2577.1400 2259.5200 ;
        RECT 2530.5400 2264.4800 2532.1400 2264.9600 ;
        RECT 2530.5400 2269.9200 2532.1400 2270.4000 ;
        RECT 2530.5400 2275.3600 2532.1400 2275.8400 ;
        RECT 2530.5400 2253.6000 2532.1400 2254.0800 ;
        RECT 2530.5400 2259.0400 2532.1400 2259.5200 ;
        RECT 2485.5400 2291.6800 2487.1400 2292.1600 ;
        RECT 2485.5400 2297.1200 2487.1400 2297.6000 ;
        RECT 2485.5400 2302.5600 2487.1400 2303.0400 ;
        RECT 2473.7800 2291.6800 2476.7800 2292.1600 ;
        RECT 2473.7800 2297.1200 2476.7800 2297.6000 ;
        RECT 2473.7800 2302.5600 2476.7800 2303.0400 ;
        RECT 2485.5400 2280.8000 2487.1400 2281.2800 ;
        RECT 2485.5400 2286.2400 2487.1400 2286.7200 ;
        RECT 2473.7800 2280.8000 2476.7800 2281.2800 ;
        RECT 2473.7800 2286.2400 2476.7800 2286.7200 ;
        RECT 2485.5400 2264.4800 2487.1400 2264.9600 ;
        RECT 2485.5400 2269.9200 2487.1400 2270.4000 ;
        RECT 2485.5400 2275.3600 2487.1400 2275.8400 ;
        RECT 2473.7800 2264.4800 2476.7800 2264.9600 ;
        RECT 2473.7800 2269.9200 2476.7800 2270.4000 ;
        RECT 2473.7800 2275.3600 2476.7800 2275.8400 ;
        RECT 2485.5400 2253.6000 2487.1400 2254.0800 ;
        RECT 2485.5400 2259.0400 2487.1400 2259.5200 ;
        RECT 2473.7800 2253.6000 2476.7800 2254.0800 ;
        RECT 2473.7800 2259.0400 2476.7800 2259.5200 ;
        RECT 2677.8800 2237.2800 2680.8800 2237.7600 ;
        RECT 2677.8800 2242.7200 2680.8800 2243.2000 ;
        RECT 2677.8800 2248.1600 2680.8800 2248.6400 ;
        RECT 2665.5400 2237.2800 2667.1400 2237.7600 ;
        RECT 2665.5400 2242.7200 2667.1400 2243.2000 ;
        RECT 2665.5400 2248.1600 2667.1400 2248.6400 ;
        RECT 2677.8800 2226.4000 2680.8800 2226.8800 ;
        RECT 2677.8800 2231.8400 2680.8800 2232.3200 ;
        RECT 2665.5400 2226.4000 2667.1400 2226.8800 ;
        RECT 2665.5400 2231.8400 2667.1400 2232.3200 ;
        RECT 2677.8800 2210.0800 2680.8800 2210.5600 ;
        RECT 2677.8800 2215.5200 2680.8800 2216.0000 ;
        RECT 2677.8800 2220.9600 2680.8800 2221.4400 ;
        RECT 2665.5400 2210.0800 2667.1400 2210.5600 ;
        RECT 2665.5400 2215.5200 2667.1400 2216.0000 ;
        RECT 2665.5400 2220.9600 2667.1400 2221.4400 ;
        RECT 2677.8800 2199.2000 2680.8800 2199.6800 ;
        RECT 2677.8800 2204.6400 2680.8800 2205.1200 ;
        RECT 2665.5400 2199.2000 2667.1400 2199.6800 ;
        RECT 2665.5400 2204.6400 2667.1400 2205.1200 ;
        RECT 2620.5400 2237.2800 2622.1400 2237.7600 ;
        RECT 2620.5400 2242.7200 2622.1400 2243.2000 ;
        RECT 2620.5400 2248.1600 2622.1400 2248.6400 ;
        RECT 2620.5400 2226.4000 2622.1400 2226.8800 ;
        RECT 2620.5400 2231.8400 2622.1400 2232.3200 ;
        RECT 2620.5400 2210.0800 2622.1400 2210.5600 ;
        RECT 2620.5400 2215.5200 2622.1400 2216.0000 ;
        RECT 2620.5400 2220.9600 2622.1400 2221.4400 ;
        RECT 2620.5400 2199.2000 2622.1400 2199.6800 ;
        RECT 2620.5400 2204.6400 2622.1400 2205.1200 ;
        RECT 2677.8800 2182.8800 2680.8800 2183.3600 ;
        RECT 2677.8800 2188.3200 2680.8800 2188.8000 ;
        RECT 2677.8800 2193.7600 2680.8800 2194.2400 ;
        RECT 2665.5400 2182.8800 2667.1400 2183.3600 ;
        RECT 2665.5400 2188.3200 2667.1400 2188.8000 ;
        RECT 2665.5400 2193.7600 2667.1400 2194.2400 ;
        RECT 2677.8800 2172.0000 2680.8800 2172.4800 ;
        RECT 2677.8800 2177.4400 2680.8800 2177.9200 ;
        RECT 2665.5400 2172.0000 2667.1400 2172.4800 ;
        RECT 2665.5400 2177.4400 2667.1400 2177.9200 ;
        RECT 2677.8800 2155.6800 2680.8800 2156.1600 ;
        RECT 2677.8800 2161.1200 2680.8800 2161.6000 ;
        RECT 2677.8800 2166.5600 2680.8800 2167.0400 ;
        RECT 2665.5400 2155.6800 2667.1400 2156.1600 ;
        RECT 2665.5400 2161.1200 2667.1400 2161.6000 ;
        RECT 2665.5400 2166.5600 2667.1400 2167.0400 ;
        RECT 2677.8800 2150.2400 2680.8800 2150.7200 ;
        RECT 2665.5400 2150.2400 2667.1400 2150.7200 ;
        RECT 2620.5400 2182.8800 2622.1400 2183.3600 ;
        RECT 2620.5400 2188.3200 2622.1400 2188.8000 ;
        RECT 2620.5400 2193.7600 2622.1400 2194.2400 ;
        RECT 2620.5400 2172.0000 2622.1400 2172.4800 ;
        RECT 2620.5400 2177.4400 2622.1400 2177.9200 ;
        RECT 2620.5400 2155.6800 2622.1400 2156.1600 ;
        RECT 2620.5400 2161.1200 2622.1400 2161.6000 ;
        RECT 2620.5400 2166.5600 2622.1400 2167.0400 ;
        RECT 2620.5400 2150.2400 2622.1400 2150.7200 ;
        RECT 2575.5400 2237.2800 2577.1400 2237.7600 ;
        RECT 2575.5400 2242.7200 2577.1400 2243.2000 ;
        RECT 2575.5400 2248.1600 2577.1400 2248.6400 ;
        RECT 2575.5400 2226.4000 2577.1400 2226.8800 ;
        RECT 2575.5400 2231.8400 2577.1400 2232.3200 ;
        RECT 2530.5400 2237.2800 2532.1400 2237.7600 ;
        RECT 2530.5400 2242.7200 2532.1400 2243.2000 ;
        RECT 2530.5400 2248.1600 2532.1400 2248.6400 ;
        RECT 2530.5400 2226.4000 2532.1400 2226.8800 ;
        RECT 2530.5400 2231.8400 2532.1400 2232.3200 ;
        RECT 2575.5400 2210.0800 2577.1400 2210.5600 ;
        RECT 2575.5400 2215.5200 2577.1400 2216.0000 ;
        RECT 2575.5400 2220.9600 2577.1400 2221.4400 ;
        RECT 2575.5400 2199.2000 2577.1400 2199.6800 ;
        RECT 2575.5400 2204.6400 2577.1400 2205.1200 ;
        RECT 2530.5400 2210.0800 2532.1400 2210.5600 ;
        RECT 2530.5400 2215.5200 2532.1400 2216.0000 ;
        RECT 2530.5400 2220.9600 2532.1400 2221.4400 ;
        RECT 2530.5400 2199.2000 2532.1400 2199.6800 ;
        RECT 2530.5400 2204.6400 2532.1400 2205.1200 ;
        RECT 2485.5400 2237.2800 2487.1400 2237.7600 ;
        RECT 2485.5400 2242.7200 2487.1400 2243.2000 ;
        RECT 2485.5400 2248.1600 2487.1400 2248.6400 ;
        RECT 2473.7800 2237.2800 2476.7800 2237.7600 ;
        RECT 2473.7800 2242.7200 2476.7800 2243.2000 ;
        RECT 2473.7800 2248.1600 2476.7800 2248.6400 ;
        RECT 2485.5400 2226.4000 2487.1400 2226.8800 ;
        RECT 2485.5400 2231.8400 2487.1400 2232.3200 ;
        RECT 2473.7800 2226.4000 2476.7800 2226.8800 ;
        RECT 2473.7800 2231.8400 2476.7800 2232.3200 ;
        RECT 2485.5400 2210.0800 2487.1400 2210.5600 ;
        RECT 2485.5400 2215.5200 2487.1400 2216.0000 ;
        RECT 2485.5400 2220.9600 2487.1400 2221.4400 ;
        RECT 2473.7800 2210.0800 2476.7800 2210.5600 ;
        RECT 2473.7800 2215.5200 2476.7800 2216.0000 ;
        RECT 2473.7800 2220.9600 2476.7800 2221.4400 ;
        RECT 2485.5400 2199.2000 2487.1400 2199.6800 ;
        RECT 2485.5400 2204.6400 2487.1400 2205.1200 ;
        RECT 2473.7800 2199.2000 2476.7800 2199.6800 ;
        RECT 2473.7800 2204.6400 2476.7800 2205.1200 ;
        RECT 2575.5400 2182.8800 2577.1400 2183.3600 ;
        RECT 2575.5400 2188.3200 2577.1400 2188.8000 ;
        RECT 2575.5400 2193.7600 2577.1400 2194.2400 ;
        RECT 2575.5400 2172.0000 2577.1400 2172.4800 ;
        RECT 2575.5400 2177.4400 2577.1400 2177.9200 ;
        RECT 2530.5400 2182.8800 2532.1400 2183.3600 ;
        RECT 2530.5400 2188.3200 2532.1400 2188.8000 ;
        RECT 2530.5400 2193.7600 2532.1400 2194.2400 ;
        RECT 2530.5400 2172.0000 2532.1400 2172.4800 ;
        RECT 2530.5400 2177.4400 2532.1400 2177.9200 ;
        RECT 2575.5400 2155.6800 2577.1400 2156.1600 ;
        RECT 2575.5400 2161.1200 2577.1400 2161.6000 ;
        RECT 2575.5400 2166.5600 2577.1400 2167.0400 ;
        RECT 2575.5400 2150.2400 2577.1400 2150.7200 ;
        RECT 2530.5400 2155.6800 2532.1400 2156.1600 ;
        RECT 2530.5400 2161.1200 2532.1400 2161.6000 ;
        RECT 2530.5400 2166.5600 2532.1400 2167.0400 ;
        RECT 2530.5400 2150.2400 2532.1400 2150.7200 ;
        RECT 2485.5400 2182.8800 2487.1400 2183.3600 ;
        RECT 2485.5400 2188.3200 2487.1400 2188.8000 ;
        RECT 2485.5400 2193.7600 2487.1400 2194.2400 ;
        RECT 2473.7800 2182.8800 2476.7800 2183.3600 ;
        RECT 2473.7800 2188.3200 2476.7800 2188.8000 ;
        RECT 2473.7800 2193.7600 2476.7800 2194.2400 ;
        RECT 2485.5400 2172.0000 2487.1400 2172.4800 ;
        RECT 2485.5400 2177.4400 2487.1400 2177.9200 ;
        RECT 2473.7800 2172.0000 2476.7800 2172.4800 ;
        RECT 2473.7800 2177.4400 2476.7800 2177.9200 ;
        RECT 2485.5400 2155.6800 2487.1400 2156.1600 ;
        RECT 2485.5400 2161.1200 2487.1400 2161.6000 ;
        RECT 2485.5400 2166.5600 2487.1400 2167.0400 ;
        RECT 2473.7800 2155.6800 2476.7800 2156.1600 ;
        RECT 2473.7800 2161.1200 2476.7800 2161.6000 ;
        RECT 2473.7800 2166.5600 2476.7800 2167.0400 ;
        RECT 2473.7800 2150.2400 2476.7800 2150.7200 ;
        RECT 2485.5400 2150.2400 2487.1400 2150.7200 ;
        RECT 2473.7800 2355.1500 2680.8800 2358.1500 ;
        RECT 2473.7800 2142.0500 2680.8800 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 1912.4100 2667.1400 2128.5100 ;
        RECT 2620.5400 1912.4100 2622.1400 2128.5100 ;
        RECT 2575.5400 1912.4100 2577.1400 2128.5100 ;
        RECT 2530.5400 1912.4100 2532.1400 2128.5100 ;
        RECT 2485.5400 1912.4100 2487.1400 2128.5100 ;
        RECT 2677.8800 1912.4100 2680.8800 2128.5100 ;
        RECT 2473.7800 1912.4100 2476.7800 2128.5100 ;
      LAYER met3 ;
        RECT 2677.8800 2105.5600 2680.8800 2106.0400 ;
        RECT 2677.8800 2111.0000 2680.8800 2111.4800 ;
        RECT 2665.5400 2105.5600 2667.1400 2106.0400 ;
        RECT 2665.5400 2111.0000 2667.1400 2111.4800 ;
        RECT 2677.8800 2116.4400 2680.8800 2116.9200 ;
        RECT 2665.5400 2116.4400 2667.1400 2116.9200 ;
        RECT 2677.8800 2094.6800 2680.8800 2095.1600 ;
        RECT 2677.8800 2100.1200 2680.8800 2100.6000 ;
        RECT 2665.5400 2094.6800 2667.1400 2095.1600 ;
        RECT 2665.5400 2100.1200 2667.1400 2100.6000 ;
        RECT 2677.8800 2078.3600 2680.8800 2078.8400 ;
        RECT 2677.8800 2083.8000 2680.8800 2084.2800 ;
        RECT 2665.5400 2078.3600 2667.1400 2078.8400 ;
        RECT 2665.5400 2083.8000 2667.1400 2084.2800 ;
        RECT 2677.8800 2089.2400 2680.8800 2089.7200 ;
        RECT 2665.5400 2089.2400 2667.1400 2089.7200 ;
        RECT 2620.5400 2105.5600 2622.1400 2106.0400 ;
        RECT 2620.5400 2111.0000 2622.1400 2111.4800 ;
        RECT 2620.5400 2116.4400 2622.1400 2116.9200 ;
        RECT 2620.5400 2094.6800 2622.1400 2095.1600 ;
        RECT 2620.5400 2100.1200 2622.1400 2100.6000 ;
        RECT 2620.5400 2078.3600 2622.1400 2078.8400 ;
        RECT 2620.5400 2083.8000 2622.1400 2084.2800 ;
        RECT 2620.5400 2089.2400 2622.1400 2089.7200 ;
        RECT 2677.8800 2062.0400 2680.8800 2062.5200 ;
        RECT 2677.8800 2067.4800 2680.8800 2067.9600 ;
        RECT 2677.8800 2072.9200 2680.8800 2073.4000 ;
        RECT 2665.5400 2062.0400 2667.1400 2062.5200 ;
        RECT 2665.5400 2067.4800 2667.1400 2067.9600 ;
        RECT 2665.5400 2072.9200 2667.1400 2073.4000 ;
        RECT 2677.8800 2051.1600 2680.8800 2051.6400 ;
        RECT 2677.8800 2056.6000 2680.8800 2057.0800 ;
        RECT 2665.5400 2051.1600 2667.1400 2051.6400 ;
        RECT 2665.5400 2056.6000 2667.1400 2057.0800 ;
        RECT 2677.8800 2034.8400 2680.8800 2035.3200 ;
        RECT 2677.8800 2040.2800 2680.8800 2040.7600 ;
        RECT 2677.8800 2045.7200 2680.8800 2046.2000 ;
        RECT 2665.5400 2034.8400 2667.1400 2035.3200 ;
        RECT 2665.5400 2040.2800 2667.1400 2040.7600 ;
        RECT 2665.5400 2045.7200 2667.1400 2046.2000 ;
        RECT 2677.8800 2023.9600 2680.8800 2024.4400 ;
        RECT 2677.8800 2029.4000 2680.8800 2029.8800 ;
        RECT 2665.5400 2023.9600 2667.1400 2024.4400 ;
        RECT 2665.5400 2029.4000 2667.1400 2029.8800 ;
        RECT 2620.5400 2062.0400 2622.1400 2062.5200 ;
        RECT 2620.5400 2067.4800 2622.1400 2067.9600 ;
        RECT 2620.5400 2072.9200 2622.1400 2073.4000 ;
        RECT 2620.5400 2051.1600 2622.1400 2051.6400 ;
        RECT 2620.5400 2056.6000 2622.1400 2057.0800 ;
        RECT 2620.5400 2034.8400 2622.1400 2035.3200 ;
        RECT 2620.5400 2040.2800 2622.1400 2040.7600 ;
        RECT 2620.5400 2045.7200 2622.1400 2046.2000 ;
        RECT 2620.5400 2023.9600 2622.1400 2024.4400 ;
        RECT 2620.5400 2029.4000 2622.1400 2029.8800 ;
        RECT 2575.5400 2105.5600 2577.1400 2106.0400 ;
        RECT 2575.5400 2111.0000 2577.1400 2111.4800 ;
        RECT 2575.5400 2116.4400 2577.1400 2116.9200 ;
        RECT 2530.5400 2105.5600 2532.1400 2106.0400 ;
        RECT 2530.5400 2111.0000 2532.1400 2111.4800 ;
        RECT 2530.5400 2116.4400 2532.1400 2116.9200 ;
        RECT 2575.5400 2094.6800 2577.1400 2095.1600 ;
        RECT 2575.5400 2100.1200 2577.1400 2100.6000 ;
        RECT 2575.5400 2078.3600 2577.1400 2078.8400 ;
        RECT 2575.5400 2083.8000 2577.1400 2084.2800 ;
        RECT 2575.5400 2089.2400 2577.1400 2089.7200 ;
        RECT 2530.5400 2094.6800 2532.1400 2095.1600 ;
        RECT 2530.5400 2100.1200 2532.1400 2100.6000 ;
        RECT 2530.5400 2078.3600 2532.1400 2078.8400 ;
        RECT 2530.5400 2083.8000 2532.1400 2084.2800 ;
        RECT 2530.5400 2089.2400 2532.1400 2089.7200 ;
        RECT 2485.5400 2105.5600 2487.1400 2106.0400 ;
        RECT 2485.5400 2111.0000 2487.1400 2111.4800 ;
        RECT 2473.7800 2111.0000 2476.7800 2111.4800 ;
        RECT 2473.7800 2105.5600 2476.7800 2106.0400 ;
        RECT 2473.7800 2116.4400 2476.7800 2116.9200 ;
        RECT 2485.5400 2116.4400 2487.1400 2116.9200 ;
        RECT 2485.5400 2094.6800 2487.1400 2095.1600 ;
        RECT 2485.5400 2100.1200 2487.1400 2100.6000 ;
        RECT 2473.7800 2100.1200 2476.7800 2100.6000 ;
        RECT 2473.7800 2094.6800 2476.7800 2095.1600 ;
        RECT 2485.5400 2078.3600 2487.1400 2078.8400 ;
        RECT 2485.5400 2083.8000 2487.1400 2084.2800 ;
        RECT 2473.7800 2083.8000 2476.7800 2084.2800 ;
        RECT 2473.7800 2078.3600 2476.7800 2078.8400 ;
        RECT 2473.7800 2089.2400 2476.7800 2089.7200 ;
        RECT 2485.5400 2089.2400 2487.1400 2089.7200 ;
        RECT 2575.5400 2062.0400 2577.1400 2062.5200 ;
        RECT 2575.5400 2067.4800 2577.1400 2067.9600 ;
        RECT 2575.5400 2072.9200 2577.1400 2073.4000 ;
        RECT 2575.5400 2051.1600 2577.1400 2051.6400 ;
        RECT 2575.5400 2056.6000 2577.1400 2057.0800 ;
        RECT 2530.5400 2062.0400 2532.1400 2062.5200 ;
        RECT 2530.5400 2067.4800 2532.1400 2067.9600 ;
        RECT 2530.5400 2072.9200 2532.1400 2073.4000 ;
        RECT 2530.5400 2051.1600 2532.1400 2051.6400 ;
        RECT 2530.5400 2056.6000 2532.1400 2057.0800 ;
        RECT 2575.5400 2034.8400 2577.1400 2035.3200 ;
        RECT 2575.5400 2040.2800 2577.1400 2040.7600 ;
        RECT 2575.5400 2045.7200 2577.1400 2046.2000 ;
        RECT 2575.5400 2023.9600 2577.1400 2024.4400 ;
        RECT 2575.5400 2029.4000 2577.1400 2029.8800 ;
        RECT 2530.5400 2034.8400 2532.1400 2035.3200 ;
        RECT 2530.5400 2040.2800 2532.1400 2040.7600 ;
        RECT 2530.5400 2045.7200 2532.1400 2046.2000 ;
        RECT 2530.5400 2023.9600 2532.1400 2024.4400 ;
        RECT 2530.5400 2029.4000 2532.1400 2029.8800 ;
        RECT 2485.5400 2062.0400 2487.1400 2062.5200 ;
        RECT 2485.5400 2067.4800 2487.1400 2067.9600 ;
        RECT 2485.5400 2072.9200 2487.1400 2073.4000 ;
        RECT 2473.7800 2062.0400 2476.7800 2062.5200 ;
        RECT 2473.7800 2067.4800 2476.7800 2067.9600 ;
        RECT 2473.7800 2072.9200 2476.7800 2073.4000 ;
        RECT 2485.5400 2051.1600 2487.1400 2051.6400 ;
        RECT 2485.5400 2056.6000 2487.1400 2057.0800 ;
        RECT 2473.7800 2051.1600 2476.7800 2051.6400 ;
        RECT 2473.7800 2056.6000 2476.7800 2057.0800 ;
        RECT 2485.5400 2034.8400 2487.1400 2035.3200 ;
        RECT 2485.5400 2040.2800 2487.1400 2040.7600 ;
        RECT 2485.5400 2045.7200 2487.1400 2046.2000 ;
        RECT 2473.7800 2034.8400 2476.7800 2035.3200 ;
        RECT 2473.7800 2040.2800 2476.7800 2040.7600 ;
        RECT 2473.7800 2045.7200 2476.7800 2046.2000 ;
        RECT 2485.5400 2023.9600 2487.1400 2024.4400 ;
        RECT 2485.5400 2029.4000 2487.1400 2029.8800 ;
        RECT 2473.7800 2023.9600 2476.7800 2024.4400 ;
        RECT 2473.7800 2029.4000 2476.7800 2029.8800 ;
        RECT 2677.8800 2007.6400 2680.8800 2008.1200 ;
        RECT 2677.8800 2013.0800 2680.8800 2013.5600 ;
        RECT 2677.8800 2018.5200 2680.8800 2019.0000 ;
        RECT 2665.5400 2007.6400 2667.1400 2008.1200 ;
        RECT 2665.5400 2013.0800 2667.1400 2013.5600 ;
        RECT 2665.5400 2018.5200 2667.1400 2019.0000 ;
        RECT 2677.8800 1996.7600 2680.8800 1997.2400 ;
        RECT 2677.8800 2002.2000 2680.8800 2002.6800 ;
        RECT 2665.5400 1996.7600 2667.1400 1997.2400 ;
        RECT 2665.5400 2002.2000 2667.1400 2002.6800 ;
        RECT 2677.8800 1980.4400 2680.8800 1980.9200 ;
        RECT 2677.8800 1985.8800 2680.8800 1986.3600 ;
        RECT 2677.8800 1991.3200 2680.8800 1991.8000 ;
        RECT 2665.5400 1980.4400 2667.1400 1980.9200 ;
        RECT 2665.5400 1985.8800 2667.1400 1986.3600 ;
        RECT 2665.5400 1991.3200 2667.1400 1991.8000 ;
        RECT 2677.8800 1969.5600 2680.8800 1970.0400 ;
        RECT 2677.8800 1975.0000 2680.8800 1975.4800 ;
        RECT 2665.5400 1969.5600 2667.1400 1970.0400 ;
        RECT 2665.5400 1975.0000 2667.1400 1975.4800 ;
        RECT 2620.5400 2007.6400 2622.1400 2008.1200 ;
        RECT 2620.5400 2013.0800 2622.1400 2013.5600 ;
        RECT 2620.5400 2018.5200 2622.1400 2019.0000 ;
        RECT 2620.5400 1996.7600 2622.1400 1997.2400 ;
        RECT 2620.5400 2002.2000 2622.1400 2002.6800 ;
        RECT 2620.5400 1980.4400 2622.1400 1980.9200 ;
        RECT 2620.5400 1985.8800 2622.1400 1986.3600 ;
        RECT 2620.5400 1991.3200 2622.1400 1991.8000 ;
        RECT 2620.5400 1969.5600 2622.1400 1970.0400 ;
        RECT 2620.5400 1975.0000 2622.1400 1975.4800 ;
        RECT 2677.8800 1953.2400 2680.8800 1953.7200 ;
        RECT 2677.8800 1958.6800 2680.8800 1959.1600 ;
        RECT 2677.8800 1964.1200 2680.8800 1964.6000 ;
        RECT 2665.5400 1953.2400 2667.1400 1953.7200 ;
        RECT 2665.5400 1958.6800 2667.1400 1959.1600 ;
        RECT 2665.5400 1964.1200 2667.1400 1964.6000 ;
        RECT 2677.8800 1942.3600 2680.8800 1942.8400 ;
        RECT 2677.8800 1947.8000 2680.8800 1948.2800 ;
        RECT 2665.5400 1942.3600 2667.1400 1942.8400 ;
        RECT 2665.5400 1947.8000 2667.1400 1948.2800 ;
        RECT 2677.8800 1926.0400 2680.8800 1926.5200 ;
        RECT 2677.8800 1931.4800 2680.8800 1931.9600 ;
        RECT 2677.8800 1936.9200 2680.8800 1937.4000 ;
        RECT 2665.5400 1926.0400 2667.1400 1926.5200 ;
        RECT 2665.5400 1931.4800 2667.1400 1931.9600 ;
        RECT 2665.5400 1936.9200 2667.1400 1937.4000 ;
        RECT 2677.8800 1920.6000 2680.8800 1921.0800 ;
        RECT 2665.5400 1920.6000 2667.1400 1921.0800 ;
        RECT 2620.5400 1953.2400 2622.1400 1953.7200 ;
        RECT 2620.5400 1958.6800 2622.1400 1959.1600 ;
        RECT 2620.5400 1964.1200 2622.1400 1964.6000 ;
        RECT 2620.5400 1942.3600 2622.1400 1942.8400 ;
        RECT 2620.5400 1947.8000 2622.1400 1948.2800 ;
        RECT 2620.5400 1926.0400 2622.1400 1926.5200 ;
        RECT 2620.5400 1931.4800 2622.1400 1931.9600 ;
        RECT 2620.5400 1936.9200 2622.1400 1937.4000 ;
        RECT 2620.5400 1920.6000 2622.1400 1921.0800 ;
        RECT 2575.5400 2007.6400 2577.1400 2008.1200 ;
        RECT 2575.5400 2013.0800 2577.1400 2013.5600 ;
        RECT 2575.5400 2018.5200 2577.1400 2019.0000 ;
        RECT 2575.5400 1996.7600 2577.1400 1997.2400 ;
        RECT 2575.5400 2002.2000 2577.1400 2002.6800 ;
        RECT 2530.5400 2007.6400 2532.1400 2008.1200 ;
        RECT 2530.5400 2013.0800 2532.1400 2013.5600 ;
        RECT 2530.5400 2018.5200 2532.1400 2019.0000 ;
        RECT 2530.5400 1996.7600 2532.1400 1997.2400 ;
        RECT 2530.5400 2002.2000 2532.1400 2002.6800 ;
        RECT 2575.5400 1980.4400 2577.1400 1980.9200 ;
        RECT 2575.5400 1985.8800 2577.1400 1986.3600 ;
        RECT 2575.5400 1991.3200 2577.1400 1991.8000 ;
        RECT 2575.5400 1969.5600 2577.1400 1970.0400 ;
        RECT 2575.5400 1975.0000 2577.1400 1975.4800 ;
        RECT 2530.5400 1980.4400 2532.1400 1980.9200 ;
        RECT 2530.5400 1985.8800 2532.1400 1986.3600 ;
        RECT 2530.5400 1991.3200 2532.1400 1991.8000 ;
        RECT 2530.5400 1969.5600 2532.1400 1970.0400 ;
        RECT 2530.5400 1975.0000 2532.1400 1975.4800 ;
        RECT 2485.5400 2007.6400 2487.1400 2008.1200 ;
        RECT 2485.5400 2013.0800 2487.1400 2013.5600 ;
        RECT 2485.5400 2018.5200 2487.1400 2019.0000 ;
        RECT 2473.7800 2007.6400 2476.7800 2008.1200 ;
        RECT 2473.7800 2013.0800 2476.7800 2013.5600 ;
        RECT 2473.7800 2018.5200 2476.7800 2019.0000 ;
        RECT 2485.5400 1996.7600 2487.1400 1997.2400 ;
        RECT 2485.5400 2002.2000 2487.1400 2002.6800 ;
        RECT 2473.7800 1996.7600 2476.7800 1997.2400 ;
        RECT 2473.7800 2002.2000 2476.7800 2002.6800 ;
        RECT 2485.5400 1980.4400 2487.1400 1980.9200 ;
        RECT 2485.5400 1985.8800 2487.1400 1986.3600 ;
        RECT 2485.5400 1991.3200 2487.1400 1991.8000 ;
        RECT 2473.7800 1980.4400 2476.7800 1980.9200 ;
        RECT 2473.7800 1985.8800 2476.7800 1986.3600 ;
        RECT 2473.7800 1991.3200 2476.7800 1991.8000 ;
        RECT 2485.5400 1969.5600 2487.1400 1970.0400 ;
        RECT 2485.5400 1975.0000 2487.1400 1975.4800 ;
        RECT 2473.7800 1969.5600 2476.7800 1970.0400 ;
        RECT 2473.7800 1975.0000 2476.7800 1975.4800 ;
        RECT 2575.5400 1953.2400 2577.1400 1953.7200 ;
        RECT 2575.5400 1958.6800 2577.1400 1959.1600 ;
        RECT 2575.5400 1964.1200 2577.1400 1964.6000 ;
        RECT 2575.5400 1942.3600 2577.1400 1942.8400 ;
        RECT 2575.5400 1947.8000 2577.1400 1948.2800 ;
        RECT 2530.5400 1953.2400 2532.1400 1953.7200 ;
        RECT 2530.5400 1958.6800 2532.1400 1959.1600 ;
        RECT 2530.5400 1964.1200 2532.1400 1964.6000 ;
        RECT 2530.5400 1942.3600 2532.1400 1942.8400 ;
        RECT 2530.5400 1947.8000 2532.1400 1948.2800 ;
        RECT 2575.5400 1926.0400 2577.1400 1926.5200 ;
        RECT 2575.5400 1931.4800 2577.1400 1931.9600 ;
        RECT 2575.5400 1936.9200 2577.1400 1937.4000 ;
        RECT 2575.5400 1920.6000 2577.1400 1921.0800 ;
        RECT 2530.5400 1926.0400 2532.1400 1926.5200 ;
        RECT 2530.5400 1931.4800 2532.1400 1931.9600 ;
        RECT 2530.5400 1936.9200 2532.1400 1937.4000 ;
        RECT 2530.5400 1920.6000 2532.1400 1921.0800 ;
        RECT 2485.5400 1953.2400 2487.1400 1953.7200 ;
        RECT 2485.5400 1958.6800 2487.1400 1959.1600 ;
        RECT 2485.5400 1964.1200 2487.1400 1964.6000 ;
        RECT 2473.7800 1953.2400 2476.7800 1953.7200 ;
        RECT 2473.7800 1958.6800 2476.7800 1959.1600 ;
        RECT 2473.7800 1964.1200 2476.7800 1964.6000 ;
        RECT 2485.5400 1942.3600 2487.1400 1942.8400 ;
        RECT 2485.5400 1947.8000 2487.1400 1948.2800 ;
        RECT 2473.7800 1942.3600 2476.7800 1942.8400 ;
        RECT 2473.7800 1947.8000 2476.7800 1948.2800 ;
        RECT 2485.5400 1926.0400 2487.1400 1926.5200 ;
        RECT 2485.5400 1931.4800 2487.1400 1931.9600 ;
        RECT 2485.5400 1936.9200 2487.1400 1937.4000 ;
        RECT 2473.7800 1926.0400 2476.7800 1926.5200 ;
        RECT 2473.7800 1931.4800 2476.7800 1931.9600 ;
        RECT 2473.7800 1936.9200 2476.7800 1937.4000 ;
        RECT 2473.7800 1920.6000 2476.7800 1921.0800 ;
        RECT 2485.5400 1920.6000 2487.1400 1921.0800 ;
        RECT 2473.7800 2125.5100 2680.8800 2128.5100 ;
        RECT 2473.7800 1912.4100 2680.8800 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 1682.7700 2667.1400 1898.8700 ;
        RECT 2620.5400 1682.7700 2622.1400 1898.8700 ;
        RECT 2575.5400 1682.7700 2577.1400 1898.8700 ;
        RECT 2530.5400 1682.7700 2532.1400 1898.8700 ;
        RECT 2485.5400 1682.7700 2487.1400 1898.8700 ;
        RECT 2677.8800 1682.7700 2680.8800 1898.8700 ;
        RECT 2473.7800 1682.7700 2476.7800 1898.8700 ;
      LAYER met3 ;
        RECT 2677.8800 1875.9200 2680.8800 1876.4000 ;
        RECT 2677.8800 1881.3600 2680.8800 1881.8400 ;
        RECT 2665.5400 1875.9200 2667.1400 1876.4000 ;
        RECT 2665.5400 1881.3600 2667.1400 1881.8400 ;
        RECT 2677.8800 1886.8000 2680.8800 1887.2800 ;
        RECT 2665.5400 1886.8000 2667.1400 1887.2800 ;
        RECT 2677.8800 1865.0400 2680.8800 1865.5200 ;
        RECT 2677.8800 1870.4800 2680.8800 1870.9600 ;
        RECT 2665.5400 1865.0400 2667.1400 1865.5200 ;
        RECT 2665.5400 1870.4800 2667.1400 1870.9600 ;
        RECT 2677.8800 1848.7200 2680.8800 1849.2000 ;
        RECT 2677.8800 1854.1600 2680.8800 1854.6400 ;
        RECT 2665.5400 1848.7200 2667.1400 1849.2000 ;
        RECT 2665.5400 1854.1600 2667.1400 1854.6400 ;
        RECT 2677.8800 1859.6000 2680.8800 1860.0800 ;
        RECT 2665.5400 1859.6000 2667.1400 1860.0800 ;
        RECT 2620.5400 1875.9200 2622.1400 1876.4000 ;
        RECT 2620.5400 1881.3600 2622.1400 1881.8400 ;
        RECT 2620.5400 1886.8000 2622.1400 1887.2800 ;
        RECT 2620.5400 1865.0400 2622.1400 1865.5200 ;
        RECT 2620.5400 1870.4800 2622.1400 1870.9600 ;
        RECT 2620.5400 1848.7200 2622.1400 1849.2000 ;
        RECT 2620.5400 1854.1600 2622.1400 1854.6400 ;
        RECT 2620.5400 1859.6000 2622.1400 1860.0800 ;
        RECT 2677.8800 1832.4000 2680.8800 1832.8800 ;
        RECT 2677.8800 1837.8400 2680.8800 1838.3200 ;
        RECT 2677.8800 1843.2800 2680.8800 1843.7600 ;
        RECT 2665.5400 1832.4000 2667.1400 1832.8800 ;
        RECT 2665.5400 1837.8400 2667.1400 1838.3200 ;
        RECT 2665.5400 1843.2800 2667.1400 1843.7600 ;
        RECT 2677.8800 1821.5200 2680.8800 1822.0000 ;
        RECT 2677.8800 1826.9600 2680.8800 1827.4400 ;
        RECT 2665.5400 1821.5200 2667.1400 1822.0000 ;
        RECT 2665.5400 1826.9600 2667.1400 1827.4400 ;
        RECT 2677.8800 1805.2000 2680.8800 1805.6800 ;
        RECT 2677.8800 1810.6400 2680.8800 1811.1200 ;
        RECT 2677.8800 1816.0800 2680.8800 1816.5600 ;
        RECT 2665.5400 1805.2000 2667.1400 1805.6800 ;
        RECT 2665.5400 1810.6400 2667.1400 1811.1200 ;
        RECT 2665.5400 1816.0800 2667.1400 1816.5600 ;
        RECT 2677.8800 1794.3200 2680.8800 1794.8000 ;
        RECT 2677.8800 1799.7600 2680.8800 1800.2400 ;
        RECT 2665.5400 1794.3200 2667.1400 1794.8000 ;
        RECT 2665.5400 1799.7600 2667.1400 1800.2400 ;
        RECT 2620.5400 1832.4000 2622.1400 1832.8800 ;
        RECT 2620.5400 1837.8400 2622.1400 1838.3200 ;
        RECT 2620.5400 1843.2800 2622.1400 1843.7600 ;
        RECT 2620.5400 1821.5200 2622.1400 1822.0000 ;
        RECT 2620.5400 1826.9600 2622.1400 1827.4400 ;
        RECT 2620.5400 1805.2000 2622.1400 1805.6800 ;
        RECT 2620.5400 1810.6400 2622.1400 1811.1200 ;
        RECT 2620.5400 1816.0800 2622.1400 1816.5600 ;
        RECT 2620.5400 1794.3200 2622.1400 1794.8000 ;
        RECT 2620.5400 1799.7600 2622.1400 1800.2400 ;
        RECT 2575.5400 1875.9200 2577.1400 1876.4000 ;
        RECT 2575.5400 1881.3600 2577.1400 1881.8400 ;
        RECT 2575.5400 1886.8000 2577.1400 1887.2800 ;
        RECT 2530.5400 1875.9200 2532.1400 1876.4000 ;
        RECT 2530.5400 1881.3600 2532.1400 1881.8400 ;
        RECT 2530.5400 1886.8000 2532.1400 1887.2800 ;
        RECT 2575.5400 1865.0400 2577.1400 1865.5200 ;
        RECT 2575.5400 1870.4800 2577.1400 1870.9600 ;
        RECT 2575.5400 1848.7200 2577.1400 1849.2000 ;
        RECT 2575.5400 1854.1600 2577.1400 1854.6400 ;
        RECT 2575.5400 1859.6000 2577.1400 1860.0800 ;
        RECT 2530.5400 1865.0400 2532.1400 1865.5200 ;
        RECT 2530.5400 1870.4800 2532.1400 1870.9600 ;
        RECT 2530.5400 1848.7200 2532.1400 1849.2000 ;
        RECT 2530.5400 1854.1600 2532.1400 1854.6400 ;
        RECT 2530.5400 1859.6000 2532.1400 1860.0800 ;
        RECT 2485.5400 1875.9200 2487.1400 1876.4000 ;
        RECT 2485.5400 1881.3600 2487.1400 1881.8400 ;
        RECT 2473.7800 1881.3600 2476.7800 1881.8400 ;
        RECT 2473.7800 1875.9200 2476.7800 1876.4000 ;
        RECT 2473.7800 1886.8000 2476.7800 1887.2800 ;
        RECT 2485.5400 1886.8000 2487.1400 1887.2800 ;
        RECT 2485.5400 1865.0400 2487.1400 1865.5200 ;
        RECT 2485.5400 1870.4800 2487.1400 1870.9600 ;
        RECT 2473.7800 1870.4800 2476.7800 1870.9600 ;
        RECT 2473.7800 1865.0400 2476.7800 1865.5200 ;
        RECT 2485.5400 1848.7200 2487.1400 1849.2000 ;
        RECT 2485.5400 1854.1600 2487.1400 1854.6400 ;
        RECT 2473.7800 1854.1600 2476.7800 1854.6400 ;
        RECT 2473.7800 1848.7200 2476.7800 1849.2000 ;
        RECT 2473.7800 1859.6000 2476.7800 1860.0800 ;
        RECT 2485.5400 1859.6000 2487.1400 1860.0800 ;
        RECT 2575.5400 1832.4000 2577.1400 1832.8800 ;
        RECT 2575.5400 1837.8400 2577.1400 1838.3200 ;
        RECT 2575.5400 1843.2800 2577.1400 1843.7600 ;
        RECT 2575.5400 1821.5200 2577.1400 1822.0000 ;
        RECT 2575.5400 1826.9600 2577.1400 1827.4400 ;
        RECT 2530.5400 1832.4000 2532.1400 1832.8800 ;
        RECT 2530.5400 1837.8400 2532.1400 1838.3200 ;
        RECT 2530.5400 1843.2800 2532.1400 1843.7600 ;
        RECT 2530.5400 1821.5200 2532.1400 1822.0000 ;
        RECT 2530.5400 1826.9600 2532.1400 1827.4400 ;
        RECT 2575.5400 1805.2000 2577.1400 1805.6800 ;
        RECT 2575.5400 1810.6400 2577.1400 1811.1200 ;
        RECT 2575.5400 1816.0800 2577.1400 1816.5600 ;
        RECT 2575.5400 1794.3200 2577.1400 1794.8000 ;
        RECT 2575.5400 1799.7600 2577.1400 1800.2400 ;
        RECT 2530.5400 1805.2000 2532.1400 1805.6800 ;
        RECT 2530.5400 1810.6400 2532.1400 1811.1200 ;
        RECT 2530.5400 1816.0800 2532.1400 1816.5600 ;
        RECT 2530.5400 1794.3200 2532.1400 1794.8000 ;
        RECT 2530.5400 1799.7600 2532.1400 1800.2400 ;
        RECT 2485.5400 1832.4000 2487.1400 1832.8800 ;
        RECT 2485.5400 1837.8400 2487.1400 1838.3200 ;
        RECT 2485.5400 1843.2800 2487.1400 1843.7600 ;
        RECT 2473.7800 1832.4000 2476.7800 1832.8800 ;
        RECT 2473.7800 1837.8400 2476.7800 1838.3200 ;
        RECT 2473.7800 1843.2800 2476.7800 1843.7600 ;
        RECT 2485.5400 1821.5200 2487.1400 1822.0000 ;
        RECT 2485.5400 1826.9600 2487.1400 1827.4400 ;
        RECT 2473.7800 1821.5200 2476.7800 1822.0000 ;
        RECT 2473.7800 1826.9600 2476.7800 1827.4400 ;
        RECT 2485.5400 1805.2000 2487.1400 1805.6800 ;
        RECT 2485.5400 1810.6400 2487.1400 1811.1200 ;
        RECT 2485.5400 1816.0800 2487.1400 1816.5600 ;
        RECT 2473.7800 1805.2000 2476.7800 1805.6800 ;
        RECT 2473.7800 1810.6400 2476.7800 1811.1200 ;
        RECT 2473.7800 1816.0800 2476.7800 1816.5600 ;
        RECT 2485.5400 1794.3200 2487.1400 1794.8000 ;
        RECT 2485.5400 1799.7600 2487.1400 1800.2400 ;
        RECT 2473.7800 1794.3200 2476.7800 1794.8000 ;
        RECT 2473.7800 1799.7600 2476.7800 1800.2400 ;
        RECT 2677.8800 1778.0000 2680.8800 1778.4800 ;
        RECT 2677.8800 1783.4400 2680.8800 1783.9200 ;
        RECT 2677.8800 1788.8800 2680.8800 1789.3600 ;
        RECT 2665.5400 1778.0000 2667.1400 1778.4800 ;
        RECT 2665.5400 1783.4400 2667.1400 1783.9200 ;
        RECT 2665.5400 1788.8800 2667.1400 1789.3600 ;
        RECT 2677.8800 1767.1200 2680.8800 1767.6000 ;
        RECT 2677.8800 1772.5600 2680.8800 1773.0400 ;
        RECT 2665.5400 1767.1200 2667.1400 1767.6000 ;
        RECT 2665.5400 1772.5600 2667.1400 1773.0400 ;
        RECT 2677.8800 1750.8000 2680.8800 1751.2800 ;
        RECT 2677.8800 1756.2400 2680.8800 1756.7200 ;
        RECT 2677.8800 1761.6800 2680.8800 1762.1600 ;
        RECT 2665.5400 1750.8000 2667.1400 1751.2800 ;
        RECT 2665.5400 1756.2400 2667.1400 1756.7200 ;
        RECT 2665.5400 1761.6800 2667.1400 1762.1600 ;
        RECT 2677.8800 1739.9200 2680.8800 1740.4000 ;
        RECT 2677.8800 1745.3600 2680.8800 1745.8400 ;
        RECT 2665.5400 1739.9200 2667.1400 1740.4000 ;
        RECT 2665.5400 1745.3600 2667.1400 1745.8400 ;
        RECT 2620.5400 1778.0000 2622.1400 1778.4800 ;
        RECT 2620.5400 1783.4400 2622.1400 1783.9200 ;
        RECT 2620.5400 1788.8800 2622.1400 1789.3600 ;
        RECT 2620.5400 1767.1200 2622.1400 1767.6000 ;
        RECT 2620.5400 1772.5600 2622.1400 1773.0400 ;
        RECT 2620.5400 1750.8000 2622.1400 1751.2800 ;
        RECT 2620.5400 1756.2400 2622.1400 1756.7200 ;
        RECT 2620.5400 1761.6800 2622.1400 1762.1600 ;
        RECT 2620.5400 1739.9200 2622.1400 1740.4000 ;
        RECT 2620.5400 1745.3600 2622.1400 1745.8400 ;
        RECT 2677.8800 1723.6000 2680.8800 1724.0800 ;
        RECT 2677.8800 1729.0400 2680.8800 1729.5200 ;
        RECT 2677.8800 1734.4800 2680.8800 1734.9600 ;
        RECT 2665.5400 1723.6000 2667.1400 1724.0800 ;
        RECT 2665.5400 1729.0400 2667.1400 1729.5200 ;
        RECT 2665.5400 1734.4800 2667.1400 1734.9600 ;
        RECT 2677.8800 1712.7200 2680.8800 1713.2000 ;
        RECT 2677.8800 1718.1600 2680.8800 1718.6400 ;
        RECT 2665.5400 1712.7200 2667.1400 1713.2000 ;
        RECT 2665.5400 1718.1600 2667.1400 1718.6400 ;
        RECT 2677.8800 1696.4000 2680.8800 1696.8800 ;
        RECT 2677.8800 1701.8400 2680.8800 1702.3200 ;
        RECT 2677.8800 1707.2800 2680.8800 1707.7600 ;
        RECT 2665.5400 1696.4000 2667.1400 1696.8800 ;
        RECT 2665.5400 1701.8400 2667.1400 1702.3200 ;
        RECT 2665.5400 1707.2800 2667.1400 1707.7600 ;
        RECT 2677.8800 1690.9600 2680.8800 1691.4400 ;
        RECT 2665.5400 1690.9600 2667.1400 1691.4400 ;
        RECT 2620.5400 1723.6000 2622.1400 1724.0800 ;
        RECT 2620.5400 1729.0400 2622.1400 1729.5200 ;
        RECT 2620.5400 1734.4800 2622.1400 1734.9600 ;
        RECT 2620.5400 1712.7200 2622.1400 1713.2000 ;
        RECT 2620.5400 1718.1600 2622.1400 1718.6400 ;
        RECT 2620.5400 1696.4000 2622.1400 1696.8800 ;
        RECT 2620.5400 1701.8400 2622.1400 1702.3200 ;
        RECT 2620.5400 1707.2800 2622.1400 1707.7600 ;
        RECT 2620.5400 1690.9600 2622.1400 1691.4400 ;
        RECT 2575.5400 1778.0000 2577.1400 1778.4800 ;
        RECT 2575.5400 1783.4400 2577.1400 1783.9200 ;
        RECT 2575.5400 1788.8800 2577.1400 1789.3600 ;
        RECT 2575.5400 1767.1200 2577.1400 1767.6000 ;
        RECT 2575.5400 1772.5600 2577.1400 1773.0400 ;
        RECT 2530.5400 1778.0000 2532.1400 1778.4800 ;
        RECT 2530.5400 1783.4400 2532.1400 1783.9200 ;
        RECT 2530.5400 1788.8800 2532.1400 1789.3600 ;
        RECT 2530.5400 1767.1200 2532.1400 1767.6000 ;
        RECT 2530.5400 1772.5600 2532.1400 1773.0400 ;
        RECT 2575.5400 1750.8000 2577.1400 1751.2800 ;
        RECT 2575.5400 1756.2400 2577.1400 1756.7200 ;
        RECT 2575.5400 1761.6800 2577.1400 1762.1600 ;
        RECT 2575.5400 1739.9200 2577.1400 1740.4000 ;
        RECT 2575.5400 1745.3600 2577.1400 1745.8400 ;
        RECT 2530.5400 1750.8000 2532.1400 1751.2800 ;
        RECT 2530.5400 1756.2400 2532.1400 1756.7200 ;
        RECT 2530.5400 1761.6800 2532.1400 1762.1600 ;
        RECT 2530.5400 1739.9200 2532.1400 1740.4000 ;
        RECT 2530.5400 1745.3600 2532.1400 1745.8400 ;
        RECT 2485.5400 1778.0000 2487.1400 1778.4800 ;
        RECT 2485.5400 1783.4400 2487.1400 1783.9200 ;
        RECT 2485.5400 1788.8800 2487.1400 1789.3600 ;
        RECT 2473.7800 1778.0000 2476.7800 1778.4800 ;
        RECT 2473.7800 1783.4400 2476.7800 1783.9200 ;
        RECT 2473.7800 1788.8800 2476.7800 1789.3600 ;
        RECT 2485.5400 1767.1200 2487.1400 1767.6000 ;
        RECT 2485.5400 1772.5600 2487.1400 1773.0400 ;
        RECT 2473.7800 1767.1200 2476.7800 1767.6000 ;
        RECT 2473.7800 1772.5600 2476.7800 1773.0400 ;
        RECT 2485.5400 1750.8000 2487.1400 1751.2800 ;
        RECT 2485.5400 1756.2400 2487.1400 1756.7200 ;
        RECT 2485.5400 1761.6800 2487.1400 1762.1600 ;
        RECT 2473.7800 1750.8000 2476.7800 1751.2800 ;
        RECT 2473.7800 1756.2400 2476.7800 1756.7200 ;
        RECT 2473.7800 1761.6800 2476.7800 1762.1600 ;
        RECT 2485.5400 1739.9200 2487.1400 1740.4000 ;
        RECT 2485.5400 1745.3600 2487.1400 1745.8400 ;
        RECT 2473.7800 1739.9200 2476.7800 1740.4000 ;
        RECT 2473.7800 1745.3600 2476.7800 1745.8400 ;
        RECT 2575.5400 1723.6000 2577.1400 1724.0800 ;
        RECT 2575.5400 1729.0400 2577.1400 1729.5200 ;
        RECT 2575.5400 1734.4800 2577.1400 1734.9600 ;
        RECT 2575.5400 1712.7200 2577.1400 1713.2000 ;
        RECT 2575.5400 1718.1600 2577.1400 1718.6400 ;
        RECT 2530.5400 1723.6000 2532.1400 1724.0800 ;
        RECT 2530.5400 1729.0400 2532.1400 1729.5200 ;
        RECT 2530.5400 1734.4800 2532.1400 1734.9600 ;
        RECT 2530.5400 1712.7200 2532.1400 1713.2000 ;
        RECT 2530.5400 1718.1600 2532.1400 1718.6400 ;
        RECT 2575.5400 1696.4000 2577.1400 1696.8800 ;
        RECT 2575.5400 1701.8400 2577.1400 1702.3200 ;
        RECT 2575.5400 1707.2800 2577.1400 1707.7600 ;
        RECT 2575.5400 1690.9600 2577.1400 1691.4400 ;
        RECT 2530.5400 1696.4000 2532.1400 1696.8800 ;
        RECT 2530.5400 1701.8400 2532.1400 1702.3200 ;
        RECT 2530.5400 1707.2800 2532.1400 1707.7600 ;
        RECT 2530.5400 1690.9600 2532.1400 1691.4400 ;
        RECT 2485.5400 1723.6000 2487.1400 1724.0800 ;
        RECT 2485.5400 1729.0400 2487.1400 1729.5200 ;
        RECT 2485.5400 1734.4800 2487.1400 1734.9600 ;
        RECT 2473.7800 1723.6000 2476.7800 1724.0800 ;
        RECT 2473.7800 1729.0400 2476.7800 1729.5200 ;
        RECT 2473.7800 1734.4800 2476.7800 1734.9600 ;
        RECT 2485.5400 1712.7200 2487.1400 1713.2000 ;
        RECT 2485.5400 1718.1600 2487.1400 1718.6400 ;
        RECT 2473.7800 1712.7200 2476.7800 1713.2000 ;
        RECT 2473.7800 1718.1600 2476.7800 1718.6400 ;
        RECT 2485.5400 1696.4000 2487.1400 1696.8800 ;
        RECT 2485.5400 1701.8400 2487.1400 1702.3200 ;
        RECT 2485.5400 1707.2800 2487.1400 1707.7600 ;
        RECT 2473.7800 1696.4000 2476.7800 1696.8800 ;
        RECT 2473.7800 1701.8400 2476.7800 1702.3200 ;
        RECT 2473.7800 1707.2800 2476.7800 1707.7600 ;
        RECT 2473.7800 1690.9600 2476.7800 1691.4400 ;
        RECT 2485.5400 1690.9600 2487.1400 1691.4400 ;
        RECT 2473.7800 1895.8700 2680.8800 1898.8700 ;
        RECT 2473.7800 1682.7700 2680.8800 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 1453.1300 2667.1400 1669.2300 ;
        RECT 2620.5400 1453.1300 2622.1400 1669.2300 ;
        RECT 2575.5400 1453.1300 2577.1400 1669.2300 ;
        RECT 2530.5400 1453.1300 2532.1400 1669.2300 ;
        RECT 2485.5400 1453.1300 2487.1400 1669.2300 ;
        RECT 2677.8800 1453.1300 2680.8800 1669.2300 ;
        RECT 2473.7800 1453.1300 2476.7800 1669.2300 ;
      LAYER met3 ;
        RECT 2677.8800 1646.2800 2680.8800 1646.7600 ;
        RECT 2677.8800 1651.7200 2680.8800 1652.2000 ;
        RECT 2665.5400 1646.2800 2667.1400 1646.7600 ;
        RECT 2665.5400 1651.7200 2667.1400 1652.2000 ;
        RECT 2677.8800 1657.1600 2680.8800 1657.6400 ;
        RECT 2665.5400 1657.1600 2667.1400 1657.6400 ;
        RECT 2677.8800 1635.4000 2680.8800 1635.8800 ;
        RECT 2677.8800 1640.8400 2680.8800 1641.3200 ;
        RECT 2665.5400 1635.4000 2667.1400 1635.8800 ;
        RECT 2665.5400 1640.8400 2667.1400 1641.3200 ;
        RECT 2677.8800 1619.0800 2680.8800 1619.5600 ;
        RECT 2677.8800 1624.5200 2680.8800 1625.0000 ;
        RECT 2665.5400 1619.0800 2667.1400 1619.5600 ;
        RECT 2665.5400 1624.5200 2667.1400 1625.0000 ;
        RECT 2677.8800 1629.9600 2680.8800 1630.4400 ;
        RECT 2665.5400 1629.9600 2667.1400 1630.4400 ;
        RECT 2620.5400 1646.2800 2622.1400 1646.7600 ;
        RECT 2620.5400 1651.7200 2622.1400 1652.2000 ;
        RECT 2620.5400 1657.1600 2622.1400 1657.6400 ;
        RECT 2620.5400 1635.4000 2622.1400 1635.8800 ;
        RECT 2620.5400 1640.8400 2622.1400 1641.3200 ;
        RECT 2620.5400 1619.0800 2622.1400 1619.5600 ;
        RECT 2620.5400 1624.5200 2622.1400 1625.0000 ;
        RECT 2620.5400 1629.9600 2622.1400 1630.4400 ;
        RECT 2677.8800 1602.7600 2680.8800 1603.2400 ;
        RECT 2677.8800 1608.2000 2680.8800 1608.6800 ;
        RECT 2677.8800 1613.6400 2680.8800 1614.1200 ;
        RECT 2665.5400 1602.7600 2667.1400 1603.2400 ;
        RECT 2665.5400 1608.2000 2667.1400 1608.6800 ;
        RECT 2665.5400 1613.6400 2667.1400 1614.1200 ;
        RECT 2677.8800 1591.8800 2680.8800 1592.3600 ;
        RECT 2677.8800 1597.3200 2680.8800 1597.8000 ;
        RECT 2665.5400 1591.8800 2667.1400 1592.3600 ;
        RECT 2665.5400 1597.3200 2667.1400 1597.8000 ;
        RECT 2677.8800 1575.5600 2680.8800 1576.0400 ;
        RECT 2677.8800 1581.0000 2680.8800 1581.4800 ;
        RECT 2677.8800 1586.4400 2680.8800 1586.9200 ;
        RECT 2665.5400 1575.5600 2667.1400 1576.0400 ;
        RECT 2665.5400 1581.0000 2667.1400 1581.4800 ;
        RECT 2665.5400 1586.4400 2667.1400 1586.9200 ;
        RECT 2677.8800 1564.6800 2680.8800 1565.1600 ;
        RECT 2677.8800 1570.1200 2680.8800 1570.6000 ;
        RECT 2665.5400 1564.6800 2667.1400 1565.1600 ;
        RECT 2665.5400 1570.1200 2667.1400 1570.6000 ;
        RECT 2620.5400 1602.7600 2622.1400 1603.2400 ;
        RECT 2620.5400 1608.2000 2622.1400 1608.6800 ;
        RECT 2620.5400 1613.6400 2622.1400 1614.1200 ;
        RECT 2620.5400 1591.8800 2622.1400 1592.3600 ;
        RECT 2620.5400 1597.3200 2622.1400 1597.8000 ;
        RECT 2620.5400 1575.5600 2622.1400 1576.0400 ;
        RECT 2620.5400 1581.0000 2622.1400 1581.4800 ;
        RECT 2620.5400 1586.4400 2622.1400 1586.9200 ;
        RECT 2620.5400 1564.6800 2622.1400 1565.1600 ;
        RECT 2620.5400 1570.1200 2622.1400 1570.6000 ;
        RECT 2575.5400 1646.2800 2577.1400 1646.7600 ;
        RECT 2575.5400 1651.7200 2577.1400 1652.2000 ;
        RECT 2575.5400 1657.1600 2577.1400 1657.6400 ;
        RECT 2530.5400 1646.2800 2532.1400 1646.7600 ;
        RECT 2530.5400 1651.7200 2532.1400 1652.2000 ;
        RECT 2530.5400 1657.1600 2532.1400 1657.6400 ;
        RECT 2575.5400 1635.4000 2577.1400 1635.8800 ;
        RECT 2575.5400 1640.8400 2577.1400 1641.3200 ;
        RECT 2575.5400 1619.0800 2577.1400 1619.5600 ;
        RECT 2575.5400 1624.5200 2577.1400 1625.0000 ;
        RECT 2575.5400 1629.9600 2577.1400 1630.4400 ;
        RECT 2530.5400 1635.4000 2532.1400 1635.8800 ;
        RECT 2530.5400 1640.8400 2532.1400 1641.3200 ;
        RECT 2530.5400 1619.0800 2532.1400 1619.5600 ;
        RECT 2530.5400 1624.5200 2532.1400 1625.0000 ;
        RECT 2530.5400 1629.9600 2532.1400 1630.4400 ;
        RECT 2485.5400 1646.2800 2487.1400 1646.7600 ;
        RECT 2485.5400 1651.7200 2487.1400 1652.2000 ;
        RECT 2473.7800 1651.7200 2476.7800 1652.2000 ;
        RECT 2473.7800 1646.2800 2476.7800 1646.7600 ;
        RECT 2473.7800 1657.1600 2476.7800 1657.6400 ;
        RECT 2485.5400 1657.1600 2487.1400 1657.6400 ;
        RECT 2485.5400 1635.4000 2487.1400 1635.8800 ;
        RECT 2485.5400 1640.8400 2487.1400 1641.3200 ;
        RECT 2473.7800 1640.8400 2476.7800 1641.3200 ;
        RECT 2473.7800 1635.4000 2476.7800 1635.8800 ;
        RECT 2485.5400 1619.0800 2487.1400 1619.5600 ;
        RECT 2485.5400 1624.5200 2487.1400 1625.0000 ;
        RECT 2473.7800 1624.5200 2476.7800 1625.0000 ;
        RECT 2473.7800 1619.0800 2476.7800 1619.5600 ;
        RECT 2473.7800 1629.9600 2476.7800 1630.4400 ;
        RECT 2485.5400 1629.9600 2487.1400 1630.4400 ;
        RECT 2575.5400 1602.7600 2577.1400 1603.2400 ;
        RECT 2575.5400 1608.2000 2577.1400 1608.6800 ;
        RECT 2575.5400 1613.6400 2577.1400 1614.1200 ;
        RECT 2575.5400 1591.8800 2577.1400 1592.3600 ;
        RECT 2575.5400 1597.3200 2577.1400 1597.8000 ;
        RECT 2530.5400 1602.7600 2532.1400 1603.2400 ;
        RECT 2530.5400 1608.2000 2532.1400 1608.6800 ;
        RECT 2530.5400 1613.6400 2532.1400 1614.1200 ;
        RECT 2530.5400 1591.8800 2532.1400 1592.3600 ;
        RECT 2530.5400 1597.3200 2532.1400 1597.8000 ;
        RECT 2575.5400 1575.5600 2577.1400 1576.0400 ;
        RECT 2575.5400 1581.0000 2577.1400 1581.4800 ;
        RECT 2575.5400 1586.4400 2577.1400 1586.9200 ;
        RECT 2575.5400 1564.6800 2577.1400 1565.1600 ;
        RECT 2575.5400 1570.1200 2577.1400 1570.6000 ;
        RECT 2530.5400 1575.5600 2532.1400 1576.0400 ;
        RECT 2530.5400 1581.0000 2532.1400 1581.4800 ;
        RECT 2530.5400 1586.4400 2532.1400 1586.9200 ;
        RECT 2530.5400 1564.6800 2532.1400 1565.1600 ;
        RECT 2530.5400 1570.1200 2532.1400 1570.6000 ;
        RECT 2485.5400 1602.7600 2487.1400 1603.2400 ;
        RECT 2485.5400 1608.2000 2487.1400 1608.6800 ;
        RECT 2485.5400 1613.6400 2487.1400 1614.1200 ;
        RECT 2473.7800 1602.7600 2476.7800 1603.2400 ;
        RECT 2473.7800 1608.2000 2476.7800 1608.6800 ;
        RECT 2473.7800 1613.6400 2476.7800 1614.1200 ;
        RECT 2485.5400 1591.8800 2487.1400 1592.3600 ;
        RECT 2485.5400 1597.3200 2487.1400 1597.8000 ;
        RECT 2473.7800 1591.8800 2476.7800 1592.3600 ;
        RECT 2473.7800 1597.3200 2476.7800 1597.8000 ;
        RECT 2485.5400 1575.5600 2487.1400 1576.0400 ;
        RECT 2485.5400 1581.0000 2487.1400 1581.4800 ;
        RECT 2485.5400 1586.4400 2487.1400 1586.9200 ;
        RECT 2473.7800 1575.5600 2476.7800 1576.0400 ;
        RECT 2473.7800 1581.0000 2476.7800 1581.4800 ;
        RECT 2473.7800 1586.4400 2476.7800 1586.9200 ;
        RECT 2485.5400 1564.6800 2487.1400 1565.1600 ;
        RECT 2485.5400 1570.1200 2487.1400 1570.6000 ;
        RECT 2473.7800 1564.6800 2476.7800 1565.1600 ;
        RECT 2473.7800 1570.1200 2476.7800 1570.6000 ;
        RECT 2677.8800 1548.3600 2680.8800 1548.8400 ;
        RECT 2677.8800 1553.8000 2680.8800 1554.2800 ;
        RECT 2677.8800 1559.2400 2680.8800 1559.7200 ;
        RECT 2665.5400 1548.3600 2667.1400 1548.8400 ;
        RECT 2665.5400 1553.8000 2667.1400 1554.2800 ;
        RECT 2665.5400 1559.2400 2667.1400 1559.7200 ;
        RECT 2677.8800 1537.4800 2680.8800 1537.9600 ;
        RECT 2677.8800 1542.9200 2680.8800 1543.4000 ;
        RECT 2665.5400 1537.4800 2667.1400 1537.9600 ;
        RECT 2665.5400 1542.9200 2667.1400 1543.4000 ;
        RECT 2677.8800 1521.1600 2680.8800 1521.6400 ;
        RECT 2677.8800 1526.6000 2680.8800 1527.0800 ;
        RECT 2677.8800 1532.0400 2680.8800 1532.5200 ;
        RECT 2665.5400 1521.1600 2667.1400 1521.6400 ;
        RECT 2665.5400 1526.6000 2667.1400 1527.0800 ;
        RECT 2665.5400 1532.0400 2667.1400 1532.5200 ;
        RECT 2677.8800 1510.2800 2680.8800 1510.7600 ;
        RECT 2677.8800 1515.7200 2680.8800 1516.2000 ;
        RECT 2665.5400 1510.2800 2667.1400 1510.7600 ;
        RECT 2665.5400 1515.7200 2667.1400 1516.2000 ;
        RECT 2620.5400 1548.3600 2622.1400 1548.8400 ;
        RECT 2620.5400 1553.8000 2622.1400 1554.2800 ;
        RECT 2620.5400 1559.2400 2622.1400 1559.7200 ;
        RECT 2620.5400 1537.4800 2622.1400 1537.9600 ;
        RECT 2620.5400 1542.9200 2622.1400 1543.4000 ;
        RECT 2620.5400 1521.1600 2622.1400 1521.6400 ;
        RECT 2620.5400 1526.6000 2622.1400 1527.0800 ;
        RECT 2620.5400 1532.0400 2622.1400 1532.5200 ;
        RECT 2620.5400 1510.2800 2622.1400 1510.7600 ;
        RECT 2620.5400 1515.7200 2622.1400 1516.2000 ;
        RECT 2677.8800 1493.9600 2680.8800 1494.4400 ;
        RECT 2677.8800 1499.4000 2680.8800 1499.8800 ;
        RECT 2677.8800 1504.8400 2680.8800 1505.3200 ;
        RECT 2665.5400 1493.9600 2667.1400 1494.4400 ;
        RECT 2665.5400 1499.4000 2667.1400 1499.8800 ;
        RECT 2665.5400 1504.8400 2667.1400 1505.3200 ;
        RECT 2677.8800 1483.0800 2680.8800 1483.5600 ;
        RECT 2677.8800 1488.5200 2680.8800 1489.0000 ;
        RECT 2665.5400 1483.0800 2667.1400 1483.5600 ;
        RECT 2665.5400 1488.5200 2667.1400 1489.0000 ;
        RECT 2677.8800 1466.7600 2680.8800 1467.2400 ;
        RECT 2677.8800 1472.2000 2680.8800 1472.6800 ;
        RECT 2677.8800 1477.6400 2680.8800 1478.1200 ;
        RECT 2665.5400 1466.7600 2667.1400 1467.2400 ;
        RECT 2665.5400 1472.2000 2667.1400 1472.6800 ;
        RECT 2665.5400 1477.6400 2667.1400 1478.1200 ;
        RECT 2677.8800 1461.3200 2680.8800 1461.8000 ;
        RECT 2665.5400 1461.3200 2667.1400 1461.8000 ;
        RECT 2620.5400 1493.9600 2622.1400 1494.4400 ;
        RECT 2620.5400 1499.4000 2622.1400 1499.8800 ;
        RECT 2620.5400 1504.8400 2622.1400 1505.3200 ;
        RECT 2620.5400 1483.0800 2622.1400 1483.5600 ;
        RECT 2620.5400 1488.5200 2622.1400 1489.0000 ;
        RECT 2620.5400 1466.7600 2622.1400 1467.2400 ;
        RECT 2620.5400 1472.2000 2622.1400 1472.6800 ;
        RECT 2620.5400 1477.6400 2622.1400 1478.1200 ;
        RECT 2620.5400 1461.3200 2622.1400 1461.8000 ;
        RECT 2575.5400 1548.3600 2577.1400 1548.8400 ;
        RECT 2575.5400 1553.8000 2577.1400 1554.2800 ;
        RECT 2575.5400 1559.2400 2577.1400 1559.7200 ;
        RECT 2575.5400 1537.4800 2577.1400 1537.9600 ;
        RECT 2575.5400 1542.9200 2577.1400 1543.4000 ;
        RECT 2530.5400 1548.3600 2532.1400 1548.8400 ;
        RECT 2530.5400 1553.8000 2532.1400 1554.2800 ;
        RECT 2530.5400 1559.2400 2532.1400 1559.7200 ;
        RECT 2530.5400 1537.4800 2532.1400 1537.9600 ;
        RECT 2530.5400 1542.9200 2532.1400 1543.4000 ;
        RECT 2575.5400 1521.1600 2577.1400 1521.6400 ;
        RECT 2575.5400 1526.6000 2577.1400 1527.0800 ;
        RECT 2575.5400 1532.0400 2577.1400 1532.5200 ;
        RECT 2575.5400 1510.2800 2577.1400 1510.7600 ;
        RECT 2575.5400 1515.7200 2577.1400 1516.2000 ;
        RECT 2530.5400 1521.1600 2532.1400 1521.6400 ;
        RECT 2530.5400 1526.6000 2532.1400 1527.0800 ;
        RECT 2530.5400 1532.0400 2532.1400 1532.5200 ;
        RECT 2530.5400 1510.2800 2532.1400 1510.7600 ;
        RECT 2530.5400 1515.7200 2532.1400 1516.2000 ;
        RECT 2485.5400 1548.3600 2487.1400 1548.8400 ;
        RECT 2485.5400 1553.8000 2487.1400 1554.2800 ;
        RECT 2485.5400 1559.2400 2487.1400 1559.7200 ;
        RECT 2473.7800 1548.3600 2476.7800 1548.8400 ;
        RECT 2473.7800 1553.8000 2476.7800 1554.2800 ;
        RECT 2473.7800 1559.2400 2476.7800 1559.7200 ;
        RECT 2485.5400 1537.4800 2487.1400 1537.9600 ;
        RECT 2485.5400 1542.9200 2487.1400 1543.4000 ;
        RECT 2473.7800 1537.4800 2476.7800 1537.9600 ;
        RECT 2473.7800 1542.9200 2476.7800 1543.4000 ;
        RECT 2485.5400 1521.1600 2487.1400 1521.6400 ;
        RECT 2485.5400 1526.6000 2487.1400 1527.0800 ;
        RECT 2485.5400 1532.0400 2487.1400 1532.5200 ;
        RECT 2473.7800 1521.1600 2476.7800 1521.6400 ;
        RECT 2473.7800 1526.6000 2476.7800 1527.0800 ;
        RECT 2473.7800 1532.0400 2476.7800 1532.5200 ;
        RECT 2485.5400 1510.2800 2487.1400 1510.7600 ;
        RECT 2485.5400 1515.7200 2487.1400 1516.2000 ;
        RECT 2473.7800 1510.2800 2476.7800 1510.7600 ;
        RECT 2473.7800 1515.7200 2476.7800 1516.2000 ;
        RECT 2575.5400 1493.9600 2577.1400 1494.4400 ;
        RECT 2575.5400 1499.4000 2577.1400 1499.8800 ;
        RECT 2575.5400 1504.8400 2577.1400 1505.3200 ;
        RECT 2575.5400 1483.0800 2577.1400 1483.5600 ;
        RECT 2575.5400 1488.5200 2577.1400 1489.0000 ;
        RECT 2530.5400 1493.9600 2532.1400 1494.4400 ;
        RECT 2530.5400 1499.4000 2532.1400 1499.8800 ;
        RECT 2530.5400 1504.8400 2532.1400 1505.3200 ;
        RECT 2530.5400 1483.0800 2532.1400 1483.5600 ;
        RECT 2530.5400 1488.5200 2532.1400 1489.0000 ;
        RECT 2575.5400 1466.7600 2577.1400 1467.2400 ;
        RECT 2575.5400 1472.2000 2577.1400 1472.6800 ;
        RECT 2575.5400 1477.6400 2577.1400 1478.1200 ;
        RECT 2575.5400 1461.3200 2577.1400 1461.8000 ;
        RECT 2530.5400 1466.7600 2532.1400 1467.2400 ;
        RECT 2530.5400 1472.2000 2532.1400 1472.6800 ;
        RECT 2530.5400 1477.6400 2532.1400 1478.1200 ;
        RECT 2530.5400 1461.3200 2532.1400 1461.8000 ;
        RECT 2485.5400 1493.9600 2487.1400 1494.4400 ;
        RECT 2485.5400 1499.4000 2487.1400 1499.8800 ;
        RECT 2485.5400 1504.8400 2487.1400 1505.3200 ;
        RECT 2473.7800 1493.9600 2476.7800 1494.4400 ;
        RECT 2473.7800 1499.4000 2476.7800 1499.8800 ;
        RECT 2473.7800 1504.8400 2476.7800 1505.3200 ;
        RECT 2485.5400 1483.0800 2487.1400 1483.5600 ;
        RECT 2485.5400 1488.5200 2487.1400 1489.0000 ;
        RECT 2473.7800 1483.0800 2476.7800 1483.5600 ;
        RECT 2473.7800 1488.5200 2476.7800 1489.0000 ;
        RECT 2485.5400 1466.7600 2487.1400 1467.2400 ;
        RECT 2485.5400 1472.2000 2487.1400 1472.6800 ;
        RECT 2485.5400 1477.6400 2487.1400 1478.1200 ;
        RECT 2473.7800 1466.7600 2476.7800 1467.2400 ;
        RECT 2473.7800 1472.2000 2476.7800 1472.6800 ;
        RECT 2473.7800 1477.6400 2476.7800 1478.1200 ;
        RECT 2473.7800 1461.3200 2476.7800 1461.8000 ;
        RECT 2485.5400 1461.3200 2487.1400 1461.8000 ;
        RECT 2473.7800 1666.2300 2680.8800 1669.2300 ;
        RECT 2473.7800 1453.1300 2680.8800 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 1223.4900 2667.1400 1439.5900 ;
        RECT 2620.5400 1223.4900 2622.1400 1439.5900 ;
        RECT 2575.5400 1223.4900 2577.1400 1439.5900 ;
        RECT 2530.5400 1223.4900 2532.1400 1439.5900 ;
        RECT 2485.5400 1223.4900 2487.1400 1439.5900 ;
        RECT 2677.8800 1223.4900 2680.8800 1439.5900 ;
        RECT 2473.7800 1223.4900 2476.7800 1439.5900 ;
      LAYER met3 ;
        RECT 2677.8800 1416.6400 2680.8800 1417.1200 ;
        RECT 2677.8800 1422.0800 2680.8800 1422.5600 ;
        RECT 2665.5400 1416.6400 2667.1400 1417.1200 ;
        RECT 2665.5400 1422.0800 2667.1400 1422.5600 ;
        RECT 2677.8800 1427.5200 2680.8800 1428.0000 ;
        RECT 2665.5400 1427.5200 2667.1400 1428.0000 ;
        RECT 2677.8800 1405.7600 2680.8800 1406.2400 ;
        RECT 2677.8800 1411.2000 2680.8800 1411.6800 ;
        RECT 2665.5400 1405.7600 2667.1400 1406.2400 ;
        RECT 2665.5400 1411.2000 2667.1400 1411.6800 ;
        RECT 2677.8800 1389.4400 2680.8800 1389.9200 ;
        RECT 2677.8800 1394.8800 2680.8800 1395.3600 ;
        RECT 2665.5400 1389.4400 2667.1400 1389.9200 ;
        RECT 2665.5400 1394.8800 2667.1400 1395.3600 ;
        RECT 2677.8800 1400.3200 2680.8800 1400.8000 ;
        RECT 2665.5400 1400.3200 2667.1400 1400.8000 ;
        RECT 2620.5400 1416.6400 2622.1400 1417.1200 ;
        RECT 2620.5400 1422.0800 2622.1400 1422.5600 ;
        RECT 2620.5400 1427.5200 2622.1400 1428.0000 ;
        RECT 2620.5400 1405.7600 2622.1400 1406.2400 ;
        RECT 2620.5400 1411.2000 2622.1400 1411.6800 ;
        RECT 2620.5400 1389.4400 2622.1400 1389.9200 ;
        RECT 2620.5400 1394.8800 2622.1400 1395.3600 ;
        RECT 2620.5400 1400.3200 2622.1400 1400.8000 ;
        RECT 2677.8800 1373.1200 2680.8800 1373.6000 ;
        RECT 2677.8800 1378.5600 2680.8800 1379.0400 ;
        RECT 2677.8800 1384.0000 2680.8800 1384.4800 ;
        RECT 2665.5400 1373.1200 2667.1400 1373.6000 ;
        RECT 2665.5400 1378.5600 2667.1400 1379.0400 ;
        RECT 2665.5400 1384.0000 2667.1400 1384.4800 ;
        RECT 2677.8800 1362.2400 2680.8800 1362.7200 ;
        RECT 2677.8800 1367.6800 2680.8800 1368.1600 ;
        RECT 2665.5400 1362.2400 2667.1400 1362.7200 ;
        RECT 2665.5400 1367.6800 2667.1400 1368.1600 ;
        RECT 2677.8800 1345.9200 2680.8800 1346.4000 ;
        RECT 2677.8800 1351.3600 2680.8800 1351.8400 ;
        RECT 2677.8800 1356.8000 2680.8800 1357.2800 ;
        RECT 2665.5400 1345.9200 2667.1400 1346.4000 ;
        RECT 2665.5400 1351.3600 2667.1400 1351.8400 ;
        RECT 2665.5400 1356.8000 2667.1400 1357.2800 ;
        RECT 2677.8800 1335.0400 2680.8800 1335.5200 ;
        RECT 2677.8800 1340.4800 2680.8800 1340.9600 ;
        RECT 2665.5400 1335.0400 2667.1400 1335.5200 ;
        RECT 2665.5400 1340.4800 2667.1400 1340.9600 ;
        RECT 2620.5400 1373.1200 2622.1400 1373.6000 ;
        RECT 2620.5400 1378.5600 2622.1400 1379.0400 ;
        RECT 2620.5400 1384.0000 2622.1400 1384.4800 ;
        RECT 2620.5400 1362.2400 2622.1400 1362.7200 ;
        RECT 2620.5400 1367.6800 2622.1400 1368.1600 ;
        RECT 2620.5400 1345.9200 2622.1400 1346.4000 ;
        RECT 2620.5400 1351.3600 2622.1400 1351.8400 ;
        RECT 2620.5400 1356.8000 2622.1400 1357.2800 ;
        RECT 2620.5400 1335.0400 2622.1400 1335.5200 ;
        RECT 2620.5400 1340.4800 2622.1400 1340.9600 ;
        RECT 2575.5400 1416.6400 2577.1400 1417.1200 ;
        RECT 2575.5400 1422.0800 2577.1400 1422.5600 ;
        RECT 2575.5400 1427.5200 2577.1400 1428.0000 ;
        RECT 2530.5400 1416.6400 2532.1400 1417.1200 ;
        RECT 2530.5400 1422.0800 2532.1400 1422.5600 ;
        RECT 2530.5400 1427.5200 2532.1400 1428.0000 ;
        RECT 2575.5400 1405.7600 2577.1400 1406.2400 ;
        RECT 2575.5400 1411.2000 2577.1400 1411.6800 ;
        RECT 2575.5400 1389.4400 2577.1400 1389.9200 ;
        RECT 2575.5400 1394.8800 2577.1400 1395.3600 ;
        RECT 2575.5400 1400.3200 2577.1400 1400.8000 ;
        RECT 2530.5400 1405.7600 2532.1400 1406.2400 ;
        RECT 2530.5400 1411.2000 2532.1400 1411.6800 ;
        RECT 2530.5400 1389.4400 2532.1400 1389.9200 ;
        RECT 2530.5400 1394.8800 2532.1400 1395.3600 ;
        RECT 2530.5400 1400.3200 2532.1400 1400.8000 ;
        RECT 2485.5400 1416.6400 2487.1400 1417.1200 ;
        RECT 2485.5400 1422.0800 2487.1400 1422.5600 ;
        RECT 2473.7800 1422.0800 2476.7800 1422.5600 ;
        RECT 2473.7800 1416.6400 2476.7800 1417.1200 ;
        RECT 2473.7800 1427.5200 2476.7800 1428.0000 ;
        RECT 2485.5400 1427.5200 2487.1400 1428.0000 ;
        RECT 2485.5400 1405.7600 2487.1400 1406.2400 ;
        RECT 2485.5400 1411.2000 2487.1400 1411.6800 ;
        RECT 2473.7800 1411.2000 2476.7800 1411.6800 ;
        RECT 2473.7800 1405.7600 2476.7800 1406.2400 ;
        RECT 2485.5400 1389.4400 2487.1400 1389.9200 ;
        RECT 2485.5400 1394.8800 2487.1400 1395.3600 ;
        RECT 2473.7800 1394.8800 2476.7800 1395.3600 ;
        RECT 2473.7800 1389.4400 2476.7800 1389.9200 ;
        RECT 2473.7800 1400.3200 2476.7800 1400.8000 ;
        RECT 2485.5400 1400.3200 2487.1400 1400.8000 ;
        RECT 2575.5400 1373.1200 2577.1400 1373.6000 ;
        RECT 2575.5400 1378.5600 2577.1400 1379.0400 ;
        RECT 2575.5400 1384.0000 2577.1400 1384.4800 ;
        RECT 2575.5400 1362.2400 2577.1400 1362.7200 ;
        RECT 2575.5400 1367.6800 2577.1400 1368.1600 ;
        RECT 2530.5400 1373.1200 2532.1400 1373.6000 ;
        RECT 2530.5400 1378.5600 2532.1400 1379.0400 ;
        RECT 2530.5400 1384.0000 2532.1400 1384.4800 ;
        RECT 2530.5400 1362.2400 2532.1400 1362.7200 ;
        RECT 2530.5400 1367.6800 2532.1400 1368.1600 ;
        RECT 2575.5400 1345.9200 2577.1400 1346.4000 ;
        RECT 2575.5400 1351.3600 2577.1400 1351.8400 ;
        RECT 2575.5400 1356.8000 2577.1400 1357.2800 ;
        RECT 2575.5400 1335.0400 2577.1400 1335.5200 ;
        RECT 2575.5400 1340.4800 2577.1400 1340.9600 ;
        RECT 2530.5400 1345.9200 2532.1400 1346.4000 ;
        RECT 2530.5400 1351.3600 2532.1400 1351.8400 ;
        RECT 2530.5400 1356.8000 2532.1400 1357.2800 ;
        RECT 2530.5400 1335.0400 2532.1400 1335.5200 ;
        RECT 2530.5400 1340.4800 2532.1400 1340.9600 ;
        RECT 2485.5400 1373.1200 2487.1400 1373.6000 ;
        RECT 2485.5400 1378.5600 2487.1400 1379.0400 ;
        RECT 2485.5400 1384.0000 2487.1400 1384.4800 ;
        RECT 2473.7800 1373.1200 2476.7800 1373.6000 ;
        RECT 2473.7800 1378.5600 2476.7800 1379.0400 ;
        RECT 2473.7800 1384.0000 2476.7800 1384.4800 ;
        RECT 2485.5400 1362.2400 2487.1400 1362.7200 ;
        RECT 2485.5400 1367.6800 2487.1400 1368.1600 ;
        RECT 2473.7800 1362.2400 2476.7800 1362.7200 ;
        RECT 2473.7800 1367.6800 2476.7800 1368.1600 ;
        RECT 2485.5400 1345.9200 2487.1400 1346.4000 ;
        RECT 2485.5400 1351.3600 2487.1400 1351.8400 ;
        RECT 2485.5400 1356.8000 2487.1400 1357.2800 ;
        RECT 2473.7800 1345.9200 2476.7800 1346.4000 ;
        RECT 2473.7800 1351.3600 2476.7800 1351.8400 ;
        RECT 2473.7800 1356.8000 2476.7800 1357.2800 ;
        RECT 2485.5400 1335.0400 2487.1400 1335.5200 ;
        RECT 2485.5400 1340.4800 2487.1400 1340.9600 ;
        RECT 2473.7800 1335.0400 2476.7800 1335.5200 ;
        RECT 2473.7800 1340.4800 2476.7800 1340.9600 ;
        RECT 2677.8800 1318.7200 2680.8800 1319.2000 ;
        RECT 2677.8800 1324.1600 2680.8800 1324.6400 ;
        RECT 2677.8800 1329.6000 2680.8800 1330.0800 ;
        RECT 2665.5400 1318.7200 2667.1400 1319.2000 ;
        RECT 2665.5400 1324.1600 2667.1400 1324.6400 ;
        RECT 2665.5400 1329.6000 2667.1400 1330.0800 ;
        RECT 2677.8800 1307.8400 2680.8800 1308.3200 ;
        RECT 2677.8800 1313.2800 2680.8800 1313.7600 ;
        RECT 2665.5400 1307.8400 2667.1400 1308.3200 ;
        RECT 2665.5400 1313.2800 2667.1400 1313.7600 ;
        RECT 2677.8800 1291.5200 2680.8800 1292.0000 ;
        RECT 2677.8800 1296.9600 2680.8800 1297.4400 ;
        RECT 2677.8800 1302.4000 2680.8800 1302.8800 ;
        RECT 2665.5400 1291.5200 2667.1400 1292.0000 ;
        RECT 2665.5400 1296.9600 2667.1400 1297.4400 ;
        RECT 2665.5400 1302.4000 2667.1400 1302.8800 ;
        RECT 2677.8800 1280.6400 2680.8800 1281.1200 ;
        RECT 2677.8800 1286.0800 2680.8800 1286.5600 ;
        RECT 2665.5400 1280.6400 2667.1400 1281.1200 ;
        RECT 2665.5400 1286.0800 2667.1400 1286.5600 ;
        RECT 2620.5400 1318.7200 2622.1400 1319.2000 ;
        RECT 2620.5400 1324.1600 2622.1400 1324.6400 ;
        RECT 2620.5400 1329.6000 2622.1400 1330.0800 ;
        RECT 2620.5400 1307.8400 2622.1400 1308.3200 ;
        RECT 2620.5400 1313.2800 2622.1400 1313.7600 ;
        RECT 2620.5400 1291.5200 2622.1400 1292.0000 ;
        RECT 2620.5400 1296.9600 2622.1400 1297.4400 ;
        RECT 2620.5400 1302.4000 2622.1400 1302.8800 ;
        RECT 2620.5400 1280.6400 2622.1400 1281.1200 ;
        RECT 2620.5400 1286.0800 2622.1400 1286.5600 ;
        RECT 2677.8800 1264.3200 2680.8800 1264.8000 ;
        RECT 2677.8800 1269.7600 2680.8800 1270.2400 ;
        RECT 2677.8800 1275.2000 2680.8800 1275.6800 ;
        RECT 2665.5400 1264.3200 2667.1400 1264.8000 ;
        RECT 2665.5400 1269.7600 2667.1400 1270.2400 ;
        RECT 2665.5400 1275.2000 2667.1400 1275.6800 ;
        RECT 2677.8800 1253.4400 2680.8800 1253.9200 ;
        RECT 2677.8800 1258.8800 2680.8800 1259.3600 ;
        RECT 2665.5400 1253.4400 2667.1400 1253.9200 ;
        RECT 2665.5400 1258.8800 2667.1400 1259.3600 ;
        RECT 2677.8800 1237.1200 2680.8800 1237.6000 ;
        RECT 2677.8800 1242.5600 2680.8800 1243.0400 ;
        RECT 2677.8800 1248.0000 2680.8800 1248.4800 ;
        RECT 2665.5400 1237.1200 2667.1400 1237.6000 ;
        RECT 2665.5400 1242.5600 2667.1400 1243.0400 ;
        RECT 2665.5400 1248.0000 2667.1400 1248.4800 ;
        RECT 2677.8800 1231.6800 2680.8800 1232.1600 ;
        RECT 2665.5400 1231.6800 2667.1400 1232.1600 ;
        RECT 2620.5400 1264.3200 2622.1400 1264.8000 ;
        RECT 2620.5400 1269.7600 2622.1400 1270.2400 ;
        RECT 2620.5400 1275.2000 2622.1400 1275.6800 ;
        RECT 2620.5400 1253.4400 2622.1400 1253.9200 ;
        RECT 2620.5400 1258.8800 2622.1400 1259.3600 ;
        RECT 2620.5400 1237.1200 2622.1400 1237.6000 ;
        RECT 2620.5400 1242.5600 2622.1400 1243.0400 ;
        RECT 2620.5400 1248.0000 2622.1400 1248.4800 ;
        RECT 2620.5400 1231.6800 2622.1400 1232.1600 ;
        RECT 2575.5400 1318.7200 2577.1400 1319.2000 ;
        RECT 2575.5400 1324.1600 2577.1400 1324.6400 ;
        RECT 2575.5400 1329.6000 2577.1400 1330.0800 ;
        RECT 2575.5400 1307.8400 2577.1400 1308.3200 ;
        RECT 2575.5400 1313.2800 2577.1400 1313.7600 ;
        RECT 2530.5400 1318.7200 2532.1400 1319.2000 ;
        RECT 2530.5400 1324.1600 2532.1400 1324.6400 ;
        RECT 2530.5400 1329.6000 2532.1400 1330.0800 ;
        RECT 2530.5400 1307.8400 2532.1400 1308.3200 ;
        RECT 2530.5400 1313.2800 2532.1400 1313.7600 ;
        RECT 2575.5400 1291.5200 2577.1400 1292.0000 ;
        RECT 2575.5400 1296.9600 2577.1400 1297.4400 ;
        RECT 2575.5400 1302.4000 2577.1400 1302.8800 ;
        RECT 2575.5400 1280.6400 2577.1400 1281.1200 ;
        RECT 2575.5400 1286.0800 2577.1400 1286.5600 ;
        RECT 2530.5400 1291.5200 2532.1400 1292.0000 ;
        RECT 2530.5400 1296.9600 2532.1400 1297.4400 ;
        RECT 2530.5400 1302.4000 2532.1400 1302.8800 ;
        RECT 2530.5400 1280.6400 2532.1400 1281.1200 ;
        RECT 2530.5400 1286.0800 2532.1400 1286.5600 ;
        RECT 2485.5400 1318.7200 2487.1400 1319.2000 ;
        RECT 2485.5400 1324.1600 2487.1400 1324.6400 ;
        RECT 2485.5400 1329.6000 2487.1400 1330.0800 ;
        RECT 2473.7800 1318.7200 2476.7800 1319.2000 ;
        RECT 2473.7800 1324.1600 2476.7800 1324.6400 ;
        RECT 2473.7800 1329.6000 2476.7800 1330.0800 ;
        RECT 2485.5400 1307.8400 2487.1400 1308.3200 ;
        RECT 2485.5400 1313.2800 2487.1400 1313.7600 ;
        RECT 2473.7800 1307.8400 2476.7800 1308.3200 ;
        RECT 2473.7800 1313.2800 2476.7800 1313.7600 ;
        RECT 2485.5400 1291.5200 2487.1400 1292.0000 ;
        RECT 2485.5400 1296.9600 2487.1400 1297.4400 ;
        RECT 2485.5400 1302.4000 2487.1400 1302.8800 ;
        RECT 2473.7800 1291.5200 2476.7800 1292.0000 ;
        RECT 2473.7800 1296.9600 2476.7800 1297.4400 ;
        RECT 2473.7800 1302.4000 2476.7800 1302.8800 ;
        RECT 2485.5400 1280.6400 2487.1400 1281.1200 ;
        RECT 2485.5400 1286.0800 2487.1400 1286.5600 ;
        RECT 2473.7800 1280.6400 2476.7800 1281.1200 ;
        RECT 2473.7800 1286.0800 2476.7800 1286.5600 ;
        RECT 2575.5400 1264.3200 2577.1400 1264.8000 ;
        RECT 2575.5400 1269.7600 2577.1400 1270.2400 ;
        RECT 2575.5400 1275.2000 2577.1400 1275.6800 ;
        RECT 2575.5400 1253.4400 2577.1400 1253.9200 ;
        RECT 2575.5400 1258.8800 2577.1400 1259.3600 ;
        RECT 2530.5400 1264.3200 2532.1400 1264.8000 ;
        RECT 2530.5400 1269.7600 2532.1400 1270.2400 ;
        RECT 2530.5400 1275.2000 2532.1400 1275.6800 ;
        RECT 2530.5400 1253.4400 2532.1400 1253.9200 ;
        RECT 2530.5400 1258.8800 2532.1400 1259.3600 ;
        RECT 2575.5400 1237.1200 2577.1400 1237.6000 ;
        RECT 2575.5400 1242.5600 2577.1400 1243.0400 ;
        RECT 2575.5400 1248.0000 2577.1400 1248.4800 ;
        RECT 2575.5400 1231.6800 2577.1400 1232.1600 ;
        RECT 2530.5400 1237.1200 2532.1400 1237.6000 ;
        RECT 2530.5400 1242.5600 2532.1400 1243.0400 ;
        RECT 2530.5400 1248.0000 2532.1400 1248.4800 ;
        RECT 2530.5400 1231.6800 2532.1400 1232.1600 ;
        RECT 2485.5400 1264.3200 2487.1400 1264.8000 ;
        RECT 2485.5400 1269.7600 2487.1400 1270.2400 ;
        RECT 2485.5400 1275.2000 2487.1400 1275.6800 ;
        RECT 2473.7800 1264.3200 2476.7800 1264.8000 ;
        RECT 2473.7800 1269.7600 2476.7800 1270.2400 ;
        RECT 2473.7800 1275.2000 2476.7800 1275.6800 ;
        RECT 2485.5400 1253.4400 2487.1400 1253.9200 ;
        RECT 2485.5400 1258.8800 2487.1400 1259.3600 ;
        RECT 2473.7800 1253.4400 2476.7800 1253.9200 ;
        RECT 2473.7800 1258.8800 2476.7800 1259.3600 ;
        RECT 2485.5400 1237.1200 2487.1400 1237.6000 ;
        RECT 2485.5400 1242.5600 2487.1400 1243.0400 ;
        RECT 2485.5400 1248.0000 2487.1400 1248.4800 ;
        RECT 2473.7800 1237.1200 2476.7800 1237.6000 ;
        RECT 2473.7800 1242.5600 2476.7800 1243.0400 ;
        RECT 2473.7800 1248.0000 2476.7800 1248.4800 ;
        RECT 2473.7800 1231.6800 2476.7800 1232.1600 ;
        RECT 2485.5400 1231.6800 2487.1400 1232.1600 ;
        RECT 2473.7800 1436.5900 2680.8800 1439.5900 ;
        RECT 2473.7800 1223.4900 2680.8800 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 993.8500 2667.1400 1209.9500 ;
        RECT 2620.5400 993.8500 2622.1400 1209.9500 ;
        RECT 2575.5400 993.8500 2577.1400 1209.9500 ;
        RECT 2530.5400 993.8500 2532.1400 1209.9500 ;
        RECT 2485.5400 993.8500 2487.1400 1209.9500 ;
        RECT 2677.8800 993.8500 2680.8800 1209.9500 ;
        RECT 2473.7800 993.8500 2476.7800 1209.9500 ;
      LAYER met3 ;
        RECT 2677.8800 1187.0000 2680.8800 1187.4800 ;
        RECT 2677.8800 1192.4400 2680.8800 1192.9200 ;
        RECT 2665.5400 1187.0000 2667.1400 1187.4800 ;
        RECT 2665.5400 1192.4400 2667.1400 1192.9200 ;
        RECT 2677.8800 1197.8800 2680.8800 1198.3600 ;
        RECT 2665.5400 1197.8800 2667.1400 1198.3600 ;
        RECT 2677.8800 1176.1200 2680.8800 1176.6000 ;
        RECT 2677.8800 1181.5600 2680.8800 1182.0400 ;
        RECT 2665.5400 1176.1200 2667.1400 1176.6000 ;
        RECT 2665.5400 1181.5600 2667.1400 1182.0400 ;
        RECT 2677.8800 1159.8000 2680.8800 1160.2800 ;
        RECT 2677.8800 1165.2400 2680.8800 1165.7200 ;
        RECT 2665.5400 1159.8000 2667.1400 1160.2800 ;
        RECT 2665.5400 1165.2400 2667.1400 1165.7200 ;
        RECT 2677.8800 1170.6800 2680.8800 1171.1600 ;
        RECT 2665.5400 1170.6800 2667.1400 1171.1600 ;
        RECT 2620.5400 1187.0000 2622.1400 1187.4800 ;
        RECT 2620.5400 1192.4400 2622.1400 1192.9200 ;
        RECT 2620.5400 1197.8800 2622.1400 1198.3600 ;
        RECT 2620.5400 1176.1200 2622.1400 1176.6000 ;
        RECT 2620.5400 1181.5600 2622.1400 1182.0400 ;
        RECT 2620.5400 1159.8000 2622.1400 1160.2800 ;
        RECT 2620.5400 1165.2400 2622.1400 1165.7200 ;
        RECT 2620.5400 1170.6800 2622.1400 1171.1600 ;
        RECT 2677.8800 1143.4800 2680.8800 1143.9600 ;
        RECT 2677.8800 1148.9200 2680.8800 1149.4000 ;
        RECT 2677.8800 1154.3600 2680.8800 1154.8400 ;
        RECT 2665.5400 1143.4800 2667.1400 1143.9600 ;
        RECT 2665.5400 1148.9200 2667.1400 1149.4000 ;
        RECT 2665.5400 1154.3600 2667.1400 1154.8400 ;
        RECT 2677.8800 1132.6000 2680.8800 1133.0800 ;
        RECT 2677.8800 1138.0400 2680.8800 1138.5200 ;
        RECT 2665.5400 1132.6000 2667.1400 1133.0800 ;
        RECT 2665.5400 1138.0400 2667.1400 1138.5200 ;
        RECT 2677.8800 1116.2800 2680.8800 1116.7600 ;
        RECT 2677.8800 1121.7200 2680.8800 1122.2000 ;
        RECT 2677.8800 1127.1600 2680.8800 1127.6400 ;
        RECT 2665.5400 1116.2800 2667.1400 1116.7600 ;
        RECT 2665.5400 1121.7200 2667.1400 1122.2000 ;
        RECT 2665.5400 1127.1600 2667.1400 1127.6400 ;
        RECT 2677.8800 1105.4000 2680.8800 1105.8800 ;
        RECT 2677.8800 1110.8400 2680.8800 1111.3200 ;
        RECT 2665.5400 1105.4000 2667.1400 1105.8800 ;
        RECT 2665.5400 1110.8400 2667.1400 1111.3200 ;
        RECT 2620.5400 1143.4800 2622.1400 1143.9600 ;
        RECT 2620.5400 1148.9200 2622.1400 1149.4000 ;
        RECT 2620.5400 1154.3600 2622.1400 1154.8400 ;
        RECT 2620.5400 1132.6000 2622.1400 1133.0800 ;
        RECT 2620.5400 1138.0400 2622.1400 1138.5200 ;
        RECT 2620.5400 1116.2800 2622.1400 1116.7600 ;
        RECT 2620.5400 1121.7200 2622.1400 1122.2000 ;
        RECT 2620.5400 1127.1600 2622.1400 1127.6400 ;
        RECT 2620.5400 1105.4000 2622.1400 1105.8800 ;
        RECT 2620.5400 1110.8400 2622.1400 1111.3200 ;
        RECT 2575.5400 1187.0000 2577.1400 1187.4800 ;
        RECT 2575.5400 1192.4400 2577.1400 1192.9200 ;
        RECT 2575.5400 1197.8800 2577.1400 1198.3600 ;
        RECT 2530.5400 1187.0000 2532.1400 1187.4800 ;
        RECT 2530.5400 1192.4400 2532.1400 1192.9200 ;
        RECT 2530.5400 1197.8800 2532.1400 1198.3600 ;
        RECT 2575.5400 1176.1200 2577.1400 1176.6000 ;
        RECT 2575.5400 1181.5600 2577.1400 1182.0400 ;
        RECT 2575.5400 1159.8000 2577.1400 1160.2800 ;
        RECT 2575.5400 1165.2400 2577.1400 1165.7200 ;
        RECT 2575.5400 1170.6800 2577.1400 1171.1600 ;
        RECT 2530.5400 1176.1200 2532.1400 1176.6000 ;
        RECT 2530.5400 1181.5600 2532.1400 1182.0400 ;
        RECT 2530.5400 1159.8000 2532.1400 1160.2800 ;
        RECT 2530.5400 1165.2400 2532.1400 1165.7200 ;
        RECT 2530.5400 1170.6800 2532.1400 1171.1600 ;
        RECT 2485.5400 1187.0000 2487.1400 1187.4800 ;
        RECT 2485.5400 1192.4400 2487.1400 1192.9200 ;
        RECT 2473.7800 1192.4400 2476.7800 1192.9200 ;
        RECT 2473.7800 1187.0000 2476.7800 1187.4800 ;
        RECT 2473.7800 1197.8800 2476.7800 1198.3600 ;
        RECT 2485.5400 1197.8800 2487.1400 1198.3600 ;
        RECT 2485.5400 1176.1200 2487.1400 1176.6000 ;
        RECT 2485.5400 1181.5600 2487.1400 1182.0400 ;
        RECT 2473.7800 1181.5600 2476.7800 1182.0400 ;
        RECT 2473.7800 1176.1200 2476.7800 1176.6000 ;
        RECT 2485.5400 1159.8000 2487.1400 1160.2800 ;
        RECT 2485.5400 1165.2400 2487.1400 1165.7200 ;
        RECT 2473.7800 1165.2400 2476.7800 1165.7200 ;
        RECT 2473.7800 1159.8000 2476.7800 1160.2800 ;
        RECT 2473.7800 1170.6800 2476.7800 1171.1600 ;
        RECT 2485.5400 1170.6800 2487.1400 1171.1600 ;
        RECT 2575.5400 1143.4800 2577.1400 1143.9600 ;
        RECT 2575.5400 1148.9200 2577.1400 1149.4000 ;
        RECT 2575.5400 1154.3600 2577.1400 1154.8400 ;
        RECT 2575.5400 1132.6000 2577.1400 1133.0800 ;
        RECT 2575.5400 1138.0400 2577.1400 1138.5200 ;
        RECT 2530.5400 1143.4800 2532.1400 1143.9600 ;
        RECT 2530.5400 1148.9200 2532.1400 1149.4000 ;
        RECT 2530.5400 1154.3600 2532.1400 1154.8400 ;
        RECT 2530.5400 1132.6000 2532.1400 1133.0800 ;
        RECT 2530.5400 1138.0400 2532.1400 1138.5200 ;
        RECT 2575.5400 1116.2800 2577.1400 1116.7600 ;
        RECT 2575.5400 1121.7200 2577.1400 1122.2000 ;
        RECT 2575.5400 1127.1600 2577.1400 1127.6400 ;
        RECT 2575.5400 1105.4000 2577.1400 1105.8800 ;
        RECT 2575.5400 1110.8400 2577.1400 1111.3200 ;
        RECT 2530.5400 1116.2800 2532.1400 1116.7600 ;
        RECT 2530.5400 1121.7200 2532.1400 1122.2000 ;
        RECT 2530.5400 1127.1600 2532.1400 1127.6400 ;
        RECT 2530.5400 1105.4000 2532.1400 1105.8800 ;
        RECT 2530.5400 1110.8400 2532.1400 1111.3200 ;
        RECT 2485.5400 1143.4800 2487.1400 1143.9600 ;
        RECT 2485.5400 1148.9200 2487.1400 1149.4000 ;
        RECT 2485.5400 1154.3600 2487.1400 1154.8400 ;
        RECT 2473.7800 1143.4800 2476.7800 1143.9600 ;
        RECT 2473.7800 1148.9200 2476.7800 1149.4000 ;
        RECT 2473.7800 1154.3600 2476.7800 1154.8400 ;
        RECT 2485.5400 1132.6000 2487.1400 1133.0800 ;
        RECT 2485.5400 1138.0400 2487.1400 1138.5200 ;
        RECT 2473.7800 1132.6000 2476.7800 1133.0800 ;
        RECT 2473.7800 1138.0400 2476.7800 1138.5200 ;
        RECT 2485.5400 1116.2800 2487.1400 1116.7600 ;
        RECT 2485.5400 1121.7200 2487.1400 1122.2000 ;
        RECT 2485.5400 1127.1600 2487.1400 1127.6400 ;
        RECT 2473.7800 1116.2800 2476.7800 1116.7600 ;
        RECT 2473.7800 1121.7200 2476.7800 1122.2000 ;
        RECT 2473.7800 1127.1600 2476.7800 1127.6400 ;
        RECT 2485.5400 1105.4000 2487.1400 1105.8800 ;
        RECT 2485.5400 1110.8400 2487.1400 1111.3200 ;
        RECT 2473.7800 1105.4000 2476.7800 1105.8800 ;
        RECT 2473.7800 1110.8400 2476.7800 1111.3200 ;
        RECT 2677.8800 1089.0800 2680.8800 1089.5600 ;
        RECT 2677.8800 1094.5200 2680.8800 1095.0000 ;
        RECT 2677.8800 1099.9600 2680.8800 1100.4400 ;
        RECT 2665.5400 1089.0800 2667.1400 1089.5600 ;
        RECT 2665.5400 1094.5200 2667.1400 1095.0000 ;
        RECT 2665.5400 1099.9600 2667.1400 1100.4400 ;
        RECT 2677.8800 1078.2000 2680.8800 1078.6800 ;
        RECT 2677.8800 1083.6400 2680.8800 1084.1200 ;
        RECT 2665.5400 1078.2000 2667.1400 1078.6800 ;
        RECT 2665.5400 1083.6400 2667.1400 1084.1200 ;
        RECT 2677.8800 1061.8800 2680.8800 1062.3600 ;
        RECT 2677.8800 1067.3200 2680.8800 1067.8000 ;
        RECT 2677.8800 1072.7600 2680.8800 1073.2400 ;
        RECT 2665.5400 1061.8800 2667.1400 1062.3600 ;
        RECT 2665.5400 1067.3200 2667.1400 1067.8000 ;
        RECT 2665.5400 1072.7600 2667.1400 1073.2400 ;
        RECT 2677.8800 1051.0000 2680.8800 1051.4800 ;
        RECT 2677.8800 1056.4400 2680.8800 1056.9200 ;
        RECT 2665.5400 1051.0000 2667.1400 1051.4800 ;
        RECT 2665.5400 1056.4400 2667.1400 1056.9200 ;
        RECT 2620.5400 1089.0800 2622.1400 1089.5600 ;
        RECT 2620.5400 1094.5200 2622.1400 1095.0000 ;
        RECT 2620.5400 1099.9600 2622.1400 1100.4400 ;
        RECT 2620.5400 1078.2000 2622.1400 1078.6800 ;
        RECT 2620.5400 1083.6400 2622.1400 1084.1200 ;
        RECT 2620.5400 1061.8800 2622.1400 1062.3600 ;
        RECT 2620.5400 1067.3200 2622.1400 1067.8000 ;
        RECT 2620.5400 1072.7600 2622.1400 1073.2400 ;
        RECT 2620.5400 1051.0000 2622.1400 1051.4800 ;
        RECT 2620.5400 1056.4400 2622.1400 1056.9200 ;
        RECT 2677.8800 1034.6800 2680.8800 1035.1600 ;
        RECT 2677.8800 1040.1200 2680.8800 1040.6000 ;
        RECT 2677.8800 1045.5600 2680.8800 1046.0400 ;
        RECT 2665.5400 1034.6800 2667.1400 1035.1600 ;
        RECT 2665.5400 1040.1200 2667.1400 1040.6000 ;
        RECT 2665.5400 1045.5600 2667.1400 1046.0400 ;
        RECT 2677.8800 1023.8000 2680.8800 1024.2800 ;
        RECT 2677.8800 1029.2400 2680.8800 1029.7200 ;
        RECT 2665.5400 1023.8000 2667.1400 1024.2800 ;
        RECT 2665.5400 1029.2400 2667.1400 1029.7200 ;
        RECT 2677.8800 1007.4800 2680.8800 1007.9600 ;
        RECT 2677.8800 1012.9200 2680.8800 1013.4000 ;
        RECT 2677.8800 1018.3600 2680.8800 1018.8400 ;
        RECT 2665.5400 1007.4800 2667.1400 1007.9600 ;
        RECT 2665.5400 1012.9200 2667.1400 1013.4000 ;
        RECT 2665.5400 1018.3600 2667.1400 1018.8400 ;
        RECT 2677.8800 1002.0400 2680.8800 1002.5200 ;
        RECT 2665.5400 1002.0400 2667.1400 1002.5200 ;
        RECT 2620.5400 1034.6800 2622.1400 1035.1600 ;
        RECT 2620.5400 1040.1200 2622.1400 1040.6000 ;
        RECT 2620.5400 1045.5600 2622.1400 1046.0400 ;
        RECT 2620.5400 1023.8000 2622.1400 1024.2800 ;
        RECT 2620.5400 1029.2400 2622.1400 1029.7200 ;
        RECT 2620.5400 1007.4800 2622.1400 1007.9600 ;
        RECT 2620.5400 1012.9200 2622.1400 1013.4000 ;
        RECT 2620.5400 1018.3600 2622.1400 1018.8400 ;
        RECT 2620.5400 1002.0400 2622.1400 1002.5200 ;
        RECT 2575.5400 1089.0800 2577.1400 1089.5600 ;
        RECT 2575.5400 1094.5200 2577.1400 1095.0000 ;
        RECT 2575.5400 1099.9600 2577.1400 1100.4400 ;
        RECT 2575.5400 1078.2000 2577.1400 1078.6800 ;
        RECT 2575.5400 1083.6400 2577.1400 1084.1200 ;
        RECT 2530.5400 1089.0800 2532.1400 1089.5600 ;
        RECT 2530.5400 1094.5200 2532.1400 1095.0000 ;
        RECT 2530.5400 1099.9600 2532.1400 1100.4400 ;
        RECT 2530.5400 1078.2000 2532.1400 1078.6800 ;
        RECT 2530.5400 1083.6400 2532.1400 1084.1200 ;
        RECT 2575.5400 1061.8800 2577.1400 1062.3600 ;
        RECT 2575.5400 1067.3200 2577.1400 1067.8000 ;
        RECT 2575.5400 1072.7600 2577.1400 1073.2400 ;
        RECT 2575.5400 1051.0000 2577.1400 1051.4800 ;
        RECT 2575.5400 1056.4400 2577.1400 1056.9200 ;
        RECT 2530.5400 1061.8800 2532.1400 1062.3600 ;
        RECT 2530.5400 1067.3200 2532.1400 1067.8000 ;
        RECT 2530.5400 1072.7600 2532.1400 1073.2400 ;
        RECT 2530.5400 1051.0000 2532.1400 1051.4800 ;
        RECT 2530.5400 1056.4400 2532.1400 1056.9200 ;
        RECT 2485.5400 1089.0800 2487.1400 1089.5600 ;
        RECT 2485.5400 1094.5200 2487.1400 1095.0000 ;
        RECT 2485.5400 1099.9600 2487.1400 1100.4400 ;
        RECT 2473.7800 1089.0800 2476.7800 1089.5600 ;
        RECT 2473.7800 1094.5200 2476.7800 1095.0000 ;
        RECT 2473.7800 1099.9600 2476.7800 1100.4400 ;
        RECT 2485.5400 1078.2000 2487.1400 1078.6800 ;
        RECT 2485.5400 1083.6400 2487.1400 1084.1200 ;
        RECT 2473.7800 1078.2000 2476.7800 1078.6800 ;
        RECT 2473.7800 1083.6400 2476.7800 1084.1200 ;
        RECT 2485.5400 1061.8800 2487.1400 1062.3600 ;
        RECT 2485.5400 1067.3200 2487.1400 1067.8000 ;
        RECT 2485.5400 1072.7600 2487.1400 1073.2400 ;
        RECT 2473.7800 1061.8800 2476.7800 1062.3600 ;
        RECT 2473.7800 1067.3200 2476.7800 1067.8000 ;
        RECT 2473.7800 1072.7600 2476.7800 1073.2400 ;
        RECT 2485.5400 1051.0000 2487.1400 1051.4800 ;
        RECT 2485.5400 1056.4400 2487.1400 1056.9200 ;
        RECT 2473.7800 1051.0000 2476.7800 1051.4800 ;
        RECT 2473.7800 1056.4400 2476.7800 1056.9200 ;
        RECT 2575.5400 1034.6800 2577.1400 1035.1600 ;
        RECT 2575.5400 1040.1200 2577.1400 1040.6000 ;
        RECT 2575.5400 1045.5600 2577.1400 1046.0400 ;
        RECT 2575.5400 1023.8000 2577.1400 1024.2800 ;
        RECT 2575.5400 1029.2400 2577.1400 1029.7200 ;
        RECT 2530.5400 1034.6800 2532.1400 1035.1600 ;
        RECT 2530.5400 1040.1200 2532.1400 1040.6000 ;
        RECT 2530.5400 1045.5600 2532.1400 1046.0400 ;
        RECT 2530.5400 1023.8000 2532.1400 1024.2800 ;
        RECT 2530.5400 1029.2400 2532.1400 1029.7200 ;
        RECT 2575.5400 1007.4800 2577.1400 1007.9600 ;
        RECT 2575.5400 1012.9200 2577.1400 1013.4000 ;
        RECT 2575.5400 1018.3600 2577.1400 1018.8400 ;
        RECT 2575.5400 1002.0400 2577.1400 1002.5200 ;
        RECT 2530.5400 1007.4800 2532.1400 1007.9600 ;
        RECT 2530.5400 1012.9200 2532.1400 1013.4000 ;
        RECT 2530.5400 1018.3600 2532.1400 1018.8400 ;
        RECT 2530.5400 1002.0400 2532.1400 1002.5200 ;
        RECT 2485.5400 1034.6800 2487.1400 1035.1600 ;
        RECT 2485.5400 1040.1200 2487.1400 1040.6000 ;
        RECT 2485.5400 1045.5600 2487.1400 1046.0400 ;
        RECT 2473.7800 1034.6800 2476.7800 1035.1600 ;
        RECT 2473.7800 1040.1200 2476.7800 1040.6000 ;
        RECT 2473.7800 1045.5600 2476.7800 1046.0400 ;
        RECT 2485.5400 1023.8000 2487.1400 1024.2800 ;
        RECT 2485.5400 1029.2400 2487.1400 1029.7200 ;
        RECT 2473.7800 1023.8000 2476.7800 1024.2800 ;
        RECT 2473.7800 1029.2400 2476.7800 1029.7200 ;
        RECT 2485.5400 1007.4800 2487.1400 1007.9600 ;
        RECT 2485.5400 1012.9200 2487.1400 1013.4000 ;
        RECT 2485.5400 1018.3600 2487.1400 1018.8400 ;
        RECT 2473.7800 1007.4800 2476.7800 1007.9600 ;
        RECT 2473.7800 1012.9200 2476.7800 1013.4000 ;
        RECT 2473.7800 1018.3600 2476.7800 1018.8400 ;
        RECT 2473.7800 1002.0400 2476.7800 1002.5200 ;
        RECT 2485.5400 1002.0400 2487.1400 1002.5200 ;
        RECT 2473.7800 1206.9500 2680.8800 1209.9500 ;
        RECT 2473.7800 993.8500 2680.8800 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2665.5400 764.2100 2667.1400 980.3100 ;
        RECT 2620.5400 764.2100 2622.1400 980.3100 ;
        RECT 2575.5400 764.2100 2577.1400 980.3100 ;
        RECT 2530.5400 764.2100 2532.1400 980.3100 ;
        RECT 2485.5400 764.2100 2487.1400 980.3100 ;
        RECT 2677.8800 764.2100 2680.8800 980.3100 ;
        RECT 2473.7800 764.2100 2476.7800 980.3100 ;
      LAYER met3 ;
        RECT 2677.8800 957.3600 2680.8800 957.8400 ;
        RECT 2677.8800 962.8000 2680.8800 963.2800 ;
        RECT 2665.5400 957.3600 2667.1400 957.8400 ;
        RECT 2665.5400 962.8000 2667.1400 963.2800 ;
        RECT 2677.8800 968.2400 2680.8800 968.7200 ;
        RECT 2665.5400 968.2400 2667.1400 968.7200 ;
        RECT 2677.8800 946.4800 2680.8800 946.9600 ;
        RECT 2677.8800 951.9200 2680.8800 952.4000 ;
        RECT 2665.5400 946.4800 2667.1400 946.9600 ;
        RECT 2665.5400 951.9200 2667.1400 952.4000 ;
        RECT 2677.8800 930.1600 2680.8800 930.6400 ;
        RECT 2677.8800 935.6000 2680.8800 936.0800 ;
        RECT 2665.5400 930.1600 2667.1400 930.6400 ;
        RECT 2665.5400 935.6000 2667.1400 936.0800 ;
        RECT 2677.8800 941.0400 2680.8800 941.5200 ;
        RECT 2665.5400 941.0400 2667.1400 941.5200 ;
        RECT 2620.5400 957.3600 2622.1400 957.8400 ;
        RECT 2620.5400 962.8000 2622.1400 963.2800 ;
        RECT 2620.5400 968.2400 2622.1400 968.7200 ;
        RECT 2620.5400 946.4800 2622.1400 946.9600 ;
        RECT 2620.5400 951.9200 2622.1400 952.4000 ;
        RECT 2620.5400 930.1600 2622.1400 930.6400 ;
        RECT 2620.5400 935.6000 2622.1400 936.0800 ;
        RECT 2620.5400 941.0400 2622.1400 941.5200 ;
        RECT 2677.8800 913.8400 2680.8800 914.3200 ;
        RECT 2677.8800 919.2800 2680.8800 919.7600 ;
        RECT 2677.8800 924.7200 2680.8800 925.2000 ;
        RECT 2665.5400 913.8400 2667.1400 914.3200 ;
        RECT 2665.5400 919.2800 2667.1400 919.7600 ;
        RECT 2665.5400 924.7200 2667.1400 925.2000 ;
        RECT 2677.8800 902.9600 2680.8800 903.4400 ;
        RECT 2677.8800 908.4000 2680.8800 908.8800 ;
        RECT 2665.5400 902.9600 2667.1400 903.4400 ;
        RECT 2665.5400 908.4000 2667.1400 908.8800 ;
        RECT 2677.8800 886.6400 2680.8800 887.1200 ;
        RECT 2677.8800 892.0800 2680.8800 892.5600 ;
        RECT 2677.8800 897.5200 2680.8800 898.0000 ;
        RECT 2665.5400 886.6400 2667.1400 887.1200 ;
        RECT 2665.5400 892.0800 2667.1400 892.5600 ;
        RECT 2665.5400 897.5200 2667.1400 898.0000 ;
        RECT 2677.8800 875.7600 2680.8800 876.2400 ;
        RECT 2677.8800 881.2000 2680.8800 881.6800 ;
        RECT 2665.5400 875.7600 2667.1400 876.2400 ;
        RECT 2665.5400 881.2000 2667.1400 881.6800 ;
        RECT 2620.5400 913.8400 2622.1400 914.3200 ;
        RECT 2620.5400 919.2800 2622.1400 919.7600 ;
        RECT 2620.5400 924.7200 2622.1400 925.2000 ;
        RECT 2620.5400 902.9600 2622.1400 903.4400 ;
        RECT 2620.5400 908.4000 2622.1400 908.8800 ;
        RECT 2620.5400 886.6400 2622.1400 887.1200 ;
        RECT 2620.5400 892.0800 2622.1400 892.5600 ;
        RECT 2620.5400 897.5200 2622.1400 898.0000 ;
        RECT 2620.5400 875.7600 2622.1400 876.2400 ;
        RECT 2620.5400 881.2000 2622.1400 881.6800 ;
        RECT 2575.5400 957.3600 2577.1400 957.8400 ;
        RECT 2575.5400 962.8000 2577.1400 963.2800 ;
        RECT 2575.5400 968.2400 2577.1400 968.7200 ;
        RECT 2530.5400 957.3600 2532.1400 957.8400 ;
        RECT 2530.5400 962.8000 2532.1400 963.2800 ;
        RECT 2530.5400 968.2400 2532.1400 968.7200 ;
        RECT 2575.5400 946.4800 2577.1400 946.9600 ;
        RECT 2575.5400 951.9200 2577.1400 952.4000 ;
        RECT 2575.5400 930.1600 2577.1400 930.6400 ;
        RECT 2575.5400 935.6000 2577.1400 936.0800 ;
        RECT 2575.5400 941.0400 2577.1400 941.5200 ;
        RECT 2530.5400 946.4800 2532.1400 946.9600 ;
        RECT 2530.5400 951.9200 2532.1400 952.4000 ;
        RECT 2530.5400 930.1600 2532.1400 930.6400 ;
        RECT 2530.5400 935.6000 2532.1400 936.0800 ;
        RECT 2530.5400 941.0400 2532.1400 941.5200 ;
        RECT 2485.5400 957.3600 2487.1400 957.8400 ;
        RECT 2485.5400 962.8000 2487.1400 963.2800 ;
        RECT 2473.7800 962.8000 2476.7800 963.2800 ;
        RECT 2473.7800 957.3600 2476.7800 957.8400 ;
        RECT 2473.7800 968.2400 2476.7800 968.7200 ;
        RECT 2485.5400 968.2400 2487.1400 968.7200 ;
        RECT 2485.5400 946.4800 2487.1400 946.9600 ;
        RECT 2485.5400 951.9200 2487.1400 952.4000 ;
        RECT 2473.7800 951.9200 2476.7800 952.4000 ;
        RECT 2473.7800 946.4800 2476.7800 946.9600 ;
        RECT 2485.5400 930.1600 2487.1400 930.6400 ;
        RECT 2485.5400 935.6000 2487.1400 936.0800 ;
        RECT 2473.7800 935.6000 2476.7800 936.0800 ;
        RECT 2473.7800 930.1600 2476.7800 930.6400 ;
        RECT 2473.7800 941.0400 2476.7800 941.5200 ;
        RECT 2485.5400 941.0400 2487.1400 941.5200 ;
        RECT 2575.5400 913.8400 2577.1400 914.3200 ;
        RECT 2575.5400 919.2800 2577.1400 919.7600 ;
        RECT 2575.5400 924.7200 2577.1400 925.2000 ;
        RECT 2575.5400 902.9600 2577.1400 903.4400 ;
        RECT 2575.5400 908.4000 2577.1400 908.8800 ;
        RECT 2530.5400 913.8400 2532.1400 914.3200 ;
        RECT 2530.5400 919.2800 2532.1400 919.7600 ;
        RECT 2530.5400 924.7200 2532.1400 925.2000 ;
        RECT 2530.5400 902.9600 2532.1400 903.4400 ;
        RECT 2530.5400 908.4000 2532.1400 908.8800 ;
        RECT 2575.5400 886.6400 2577.1400 887.1200 ;
        RECT 2575.5400 892.0800 2577.1400 892.5600 ;
        RECT 2575.5400 897.5200 2577.1400 898.0000 ;
        RECT 2575.5400 875.7600 2577.1400 876.2400 ;
        RECT 2575.5400 881.2000 2577.1400 881.6800 ;
        RECT 2530.5400 886.6400 2532.1400 887.1200 ;
        RECT 2530.5400 892.0800 2532.1400 892.5600 ;
        RECT 2530.5400 897.5200 2532.1400 898.0000 ;
        RECT 2530.5400 875.7600 2532.1400 876.2400 ;
        RECT 2530.5400 881.2000 2532.1400 881.6800 ;
        RECT 2485.5400 913.8400 2487.1400 914.3200 ;
        RECT 2485.5400 919.2800 2487.1400 919.7600 ;
        RECT 2485.5400 924.7200 2487.1400 925.2000 ;
        RECT 2473.7800 913.8400 2476.7800 914.3200 ;
        RECT 2473.7800 919.2800 2476.7800 919.7600 ;
        RECT 2473.7800 924.7200 2476.7800 925.2000 ;
        RECT 2485.5400 902.9600 2487.1400 903.4400 ;
        RECT 2485.5400 908.4000 2487.1400 908.8800 ;
        RECT 2473.7800 902.9600 2476.7800 903.4400 ;
        RECT 2473.7800 908.4000 2476.7800 908.8800 ;
        RECT 2485.5400 886.6400 2487.1400 887.1200 ;
        RECT 2485.5400 892.0800 2487.1400 892.5600 ;
        RECT 2485.5400 897.5200 2487.1400 898.0000 ;
        RECT 2473.7800 886.6400 2476.7800 887.1200 ;
        RECT 2473.7800 892.0800 2476.7800 892.5600 ;
        RECT 2473.7800 897.5200 2476.7800 898.0000 ;
        RECT 2485.5400 875.7600 2487.1400 876.2400 ;
        RECT 2485.5400 881.2000 2487.1400 881.6800 ;
        RECT 2473.7800 875.7600 2476.7800 876.2400 ;
        RECT 2473.7800 881.2000 2476.7800 881.6800 ;
        RECT 2677.8800 859.4400 2680.8800 859.9200 ;
        RECT 2677.8800 864.8800 2680.8800 865.3600 ;
        RECT 2677.8800 870.3200 2680.8800 870.8000 ;
        RECT 2665.5400 859.4400 2667.1400 859.9200 ;
        RECT 2665.5400 864.8800 2667.1400 865.3600 ;
        RECT 2665.5400 870.3200 2667.1400 870.8000 ;
        RECT 2677.8800 848.5600 2680.8800 849.0400 ;
        RECT 2677.8800 854.0000 2680.8800 854.4800 ;
        RECT 2665.5400 848.5600 2667.1400 849.0400 ;
        RECT 2665.5400 854.0000 2667.1400 854.4800 ;
        RECT 2677.8800 832.2400 2680.8800 832.7200 ;
        RECT 2677.8800 837.6800 2680.8800 838.1600 ;
        RECT 2677.8800 843.1200 2680.8800 843.6000 ;
        RECT 2665.5400 832.2400 2667.1400 832.7200 ;
        RECT 2665.5400 837.6800 2667.1400 838.1600 ;
        RECT 2665.5400 843.1200 2667.1400 843.6000 ;
        RECT 2677.8800 821.3600 2680.8800 821.8400 ;
        RECT 2677.8800 826.8000 2680.8800 827.2800 ;
        RECT 2665.5400 821.3600 2667.1400 821.8400 ;
        RECT 2665.5400 826.8000 2667.1400 827.2800 ;
        RECT 2620.5400 859.4400 2622.1400 859.9200 ;
        RECT 2620.5400 864.8800 2622.1400 865.3600 ;
        RECT 2620.5400 870.3200 2622.1400 870.8000 ;
        RECT 2620.5400 848.5600 2622.1400 849.0400 ;
        RECT 2620.5400 854.0000 2622.1400 854.4800 ;
        RECT 2620.5400 832.2400 2622.1400 832.7200 ;
        RECT 2620.5400 837.6800 2622.1400 838.1600 ;
        RECT 2620.5400 843.1200 2622.1400 843.6000 ;
        RECT 2620.5400 821.3600 2622.1400 821.8400 ;
        RECT 2620.5400 826.8000 2622.1400 827.2800 ;
        RECT 2677.8800 805.0400 2680.8800 805.5200 ;
        RECT 2677.8800 810.4800 2680.8800 810.9600 ;
        RECT 2677.8800 815.9200 2680.8800 816.4000 ;
        RECT 2665.5400 805.0400 2667.1400 805.5200 ;
        RECT 2665.5400 810.4800 2667.1400 810.9600 ;
        RECT 2665.5400 815.9200 2667.1400 816.4000 ;
        RECT 2677.8800 794.1600 2680.8800 794.6400 ;
        RECT 2677.8800 799.6000 2680.8800 800.0800 ;
        RECT 2665.5400 794.1600 2667.1400 794.6400 ;
        RECT 2665.5400 799.6000 2667.1400 800.0800 ;
        RECT 2677.8800 777.8400 2680.8800 778.3200 ;
        RECT 2677.8800 783.2800 2680.8800 783.7600 ;
        RECT 2677.8800 788.7200 2680.8800 789.2000 ;
        RECT 2665.5400 777.8400 2667.1400 778.3200 ;
        RECT 2665.5400 783.2800 2667.1400 783.7600 ;
        RECT 2665.5400 788.7200 2667.1400 789.2000 ;
        RECT 2677.8800 772.4000 2680.8800 772.8800 ;
        RECT 2665.5400 772.4000 2667.1400 772.8800 ;
        RECT 2620.5400 805.0400 2622.1400 805.5200 ;
        RECT 2620.5400 810.4800 2622.1400 810.9600 ;
        RECT 2620.5400 815.9200 2622.1400 816.4000 ;
        RECT 2620.5400 794.1600 2622.1400 794.6400 ;
        RECT 2620.5400 799.6000 2622.1400 800.0800 ;
        RECT 2620.5400 777.8400 2622.1400 778.3200 ;
        RECT 2620.5400 783.2800 2622.1400 783.7600 ;
        RECT 2620.5400 788.7200 2622.1400 789.2000 ;
        RECT 2620.5400 772.4000 2622.1400 772.8800 ;
        RECT 2575.5400 859.4400 2577.1400 859.9200 ;
        RECT 2575.5400 864.8800 2577.1400 865.3600 ;
        RECT 2575.5400 870.3200 2577.1400 870.8000 ;
        RECT 2575.5400 848.5600 2577.1400 849.0400 ;
        RECT 2575.5400 854.0000 2577.1400 854.4800 ;
        RECT 2530.5400 859.4400 2532.1400 859.9200 ;
        RECT 2530.5400 864.8800 2532.1400 865.3600 ;
        RECT 2530.5400 870.3200 2532.1400 870.8000 ;
        RECT 2530.5400 848.5600 2532.1400 849.0400 ;
        RECT 2530.5400 854.0000 2532.1400 854.4800 ;
        RECT 2575.5400 832.2400 2577.1400 832.7200 ;
        RECT 2575.5400 837.6800 2577.1400 838.1600 ;
        RECT 2575.5400 843.1200 2577.1400 843.6000 ;
        RECT 2575.5400 821.3600 2577.1400 821.8400 ;
        RECT 2575.5400 826.8000 2577.1400 827.2800 ;
        RECT 2530.5400 832.2400 2532.1400 832.7200 ;
        RECT 2530.5400 837.6800 2532.1400 838.1600 ;
        RECT 2530.5400 843.1200 2532.1400 843.6000 ;
        RECT 2530.5400 821.3600 2532.1400 821.8400 ;
        RECT 2530.5400 826.8000 2532.1400 827.2800 ;
        RECT 2485.5400 859.4400 2487.1400 859.9200 ;
        RECT 2485.5400 864.8800 2487.1400 865.3600 ;
        RECT 2485.5400 870.3200 2487.1400 870.8000 ;
        RECT 2473.7800 859.4400 2476.7800 859.9200 ;
        RECT 2473.7800 864.8800 2476.7800 865.3600 ;
        RECT 2473.7800 870.3200 2476.7800 870.8000 ;
        RECT 2485.5400 848.5600 2487.1400 849.0400 ;
        RECT 2485.5400 854.0000 2487.1400 854.4800 ;
        RECT 2473.7800 848.5600 2476.7800 849.0400 ;
        RECT 2473.7800 854.0000 2476.7800 854.4800 ;
        RECT 2485.5400 832.2400 2487.1400 832.7200 ;
        RECT 2485.5400 837.6800 2487.1400 838.1600 ;
        RECT 2485.5400 843.1200 2487.1400 843.6000 ;
        RECT 2473.7800 832.2400 2476.7800 832.7200 ;
        RECT 2473.7800 837.6800 2476.7800 838.1600 ;
        RECT 2473.7800 843.1200 2476.7800 843.6000 ;
        RECT 2485.5400 821.3600 2487.1400 821.8400 ;
        RECT 2485.5400 826.8000 2487.1400 827.2800 ;
        RECT 2473.7800 821.3600 2476.7800 821.8400 ;
        RECT 2473.7800 826.8000 2476.7800 827.2800 ;
        RECT 2575.5400 805.0400 2577.1400 805.5200 ;
        RECT 2575.5400 810.4800 2577.1400 810.9600 ;
        RECT 2575.5400 815.9200 2577.1400 816.4000 ;
        RECT 2575.5400 794.1600 2577.1400 794.6400 ;
        RECT 2575.5400 799.6000 2577.1400 800.0800 ;
        RECT 2530.5400 805.0400 2532.1400 805.5200 ;
        RECT 2530.5400 810.4800 2532.1400 810.9600 ;
        RECT 2530.5400 815.9200 2532.1400 816.4000 ;
        RECT 2530.5400 794.1600 2532.1400 794.6400 ;
        RECT 2530.5400 799.6000 2532.1400 800.0800 ;
        RECT 2575.5400 777.8400 2577.1400 778.3200 ;
        RECT 2575.5400 783.2800 2577.1400 783.7600 ;
        RECT 2575.5400 788.7200 2577.1400 789.2000 ;
        RECT 2575.5400 772.4000 2577.1400 772.8800 ;
        RECT 2530.5400 777.8400 2532.1400 778.3200 ;
        RECT 2530.5400 783.2800 2532.1400 783.7600 ;
        RECT 2530.5400 788.7200 2532.1400 789.2000 ;
        RECT 2530.5400 772.4000 2532.1400 772.8800 ;
        RECT 2485.5400 805.0400 2487.1400 805.5200 ;
        RECT 2485.5400 810.4800 2487.1400 810.9600 ;
        RECT 2485.5400 815.9200 2487.1400 816.4000 ;
        RECT 2473.7800 805.0400 2476.7800 805.5200 ;
        RECT 2473.7800 810.4800 2476.7800 810.9600 ;
        RECT 2473.7800 815.9200 2476.7800 816.4000 ;
        RECT 2485.5400 794.1600 2487.1400 794.6400 ;
        RECT 2485.5400 799.6000 2487.1400 800.0800 ;
        RECT 2473.7800 794.1600 2476.7800 794.6400 ;
        RECT 2473.7800 799.6000 2476.7800 800.0800 ;
        RECT 2485.5400 777.8400 2487.1400 778.3200 ;
        RECT 2485.5400 783.2800 2487.1400 783.7600 ;
        RECT 2485.5400 788.7200 2487.1400 789.2000 ;
        RECT 2473.7800 777.8400 2476.7800 778.3200 ;
        RECT 2473.7800 783.2800 2476.7800 783.7600 ;
        RECT 2473.7800 788.7200 2476.7800 789.2000 ;
        RECT 2473.7800 772.4000 2476.7800 772.8800 ;
        RECT 2485.5400 772.4000 2487.1400 772.8800 ;
        RECT 2473.7800 977.3100 2680.8800 980.3100 ;
        RECT 2473.7800 764.2100 2680.8800 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2788.1600 2830.6100 2790.1600 2857.5400 ;
        RECT 2695.0000 2830.6100 2697.0000 2857.5400 ;
      LAYER met3 ;
        RECT 2788.1600 2847.3200 2790.1600 2847.8000 ;
        RECT 2695.0000 2847.3200 2697.0000 2847.8000 ;
        RECT 2788.1600 2836.4400 2790.1600 2836.9200 ;
        RECT 2788.1600 2841.8800 2790.1600 2842.3600 ;
        RECT 2695.0000 2836.4400 2697.0000 2836.9200 ;
        RECT 2695.0000 2841.8800 2697.0000 2842.3600 ;
        RECT 2695.0000 2855.5400 2790.1600 2857.5400 ;
        RECT 2695.0000 2830.6100 2790.1600 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 536.0700 2697.0000 749.1700 ;
        RECT 2788.1600 536.0700 2789.6600 749.1700 ;
      LAYER met3 ;
        RECT 2788.1600 733.1600 2789.6600 733.6400 ;
        RECT 2788.1600 727.7200 2789.6600 728.2000 ;
        RECT 2788.1600 738.6000 2789.6600 739.0800 ;
        RECT 2788.1600 722.2800 2789.6600 722.7600 ;
        RECT 2788.1600 716.8400 2789.6600 717.3200 ;
        RECT 2788.1600 705.9600 2789.6600 706.4400 ;
        RECT 2788.1600 700.5200 2789.6600 701.0000 ;
        RECT 2788.1600 711.4000 2789.6600 711.8800 ;
        RECT 2788.1600 695.0800 2789.6600 695.5600 ;
        RECT 2788.1600 689.6400 2789.6600 690.1200 ;
        RECT 2788.1600 684.2000 2789.6600 684.6800 ;
        RECT 2788.1600 678.7600 2789.6600 679.2400 ;
        RECT 2788.1600 673.3200 2789.6600 673.8000 ;
        RECT 2788.1600 667.8800 2789.6600 668.3600 ;
        RECT 2788.1600 662.4400 2789.6600 662.9200 ;
        RECT 2788.1600 657.0000 2789.6600 657.4800 ;
        RECT 2788.1600 651.5600 2789.6600 652.0400 ;
        RECT 2788.1600 646.1200 2789.6600 646.6000 ;
        RECT 2695.5000 733.1600 2697.0000 733.6400 ;
        RECT 2695.5000 727.7200 2697.0000 728.2000 ;
        RECT 2695.5000 738.6000 2697.0000 739.0800 ;
        RECT 2695.5000 722.2800 2697.0000 722.7600 ;
        RECT 2695.5000 716.8400 2697.0000 717.3200 ;
        RECT 2695.5000 705.9600 2697.0000 706.4400 ;
        RECT 2695.5000 700.5200 2697.0000 701.0000 ;
        RECT 2695.5000 711.4000 2697.0000 711.8800 ;
        RECT 2695.5000 695.0800 2697.0000 695.5600 ;
        RECT 2695.5000 689.6400 2697.0000 690.1200 ;
        RECT 2695.5000 684.2000 2697.0000 684.6800 ;
        RECT 2695.5000 678.7600 2697.0000 679.2400 ;
        RECT 2695.5000 673.3200 2697.0000 673.8000 ;
        RECT 2695.5000 667.8800 2697.0000 668.3600 ;
        RECT 2695.5000 662.4400 2697.0000 662.9200 ;
        RECT 2695.5000 657.0000 2697.0000 657.4800 ;
        RECT 2695.5000 651.5600 2697.0000 652.0400 ;
        RECT 2695.5000 646.1200 2697.0000 646.6000 ;
        RECT 2788.1600 640.6800 2789.6600 641.1600 ;
        RECT 2788.1600 635.2400 2789.6600 635.7200 ;
        RECT 2788.1600 629.8000 2789.6600 630.2800 ;
        RECT 2788.1600 624.3600 2789.6600 624.8400 ;
        RECT 2788.1600 618.9200 2789.6600 619.4000 ;
        RECT 2788.1600 613.4800 2789.6600 613.9600 ;
        RECT 2788.1600 608.0400 2789.6600 608.5200 ;
        RECT 2788.1600 602.6000 2789.6600 603.0800 ;
        RECT 2788.1600 597.1600 2789.6600 597.6400 ;
        RECT 2788.1600 591.7200 2789.6600 592.2000 ;
        RECT 2788.1600 586.2800 2789.6600 586.7600 ;
        RECT 2788.1600 580.8400 2789.6600 581.3200 ;
        RECT 2788.1600 575.4000 2789.6600 575.8800 ;
        RECT 2788.1600 569.9600 2789.6600 570.4400 ;
        RECT 2788.1600 564.5200 2789.6600 565.0000 ;
        RECT 2788.1600 559.0800 2789.6600 559.5600 ;
        RECT 2788.1600 553.6400 2789.6600 554.1200 ;
        RECT 2788.1600 548.2000 2789.6600 548.6800 ;
        RECT 2788.1600 542.7600 2789.6600 543.2400 ;
        RECT 2695.5000 640.6800 2697.0000 641.1600 ;
        RECT 2695.5000 635.2400 2697.0000 635.7200 ;
        RECT 2695.5000 629.8000 2697.0000 630.2800 ;
        RECT 2695.5000 624.3600 2697.0000 624.8400 ;
        RECT 2695.5000 618.9200 2697.0000 619.4000 ;
        RECT 2695.5000 613.4800 2697.0000 613.9600 ;
        RECT 2695.5000 608.0400 2697.0000 608.5200 ;
        RECT 2695.5000 602.6000 2697.0000 603.0800 ;
        RECT 2695.5000 597.1600 2697.0000 597.6400 ;
        RECT 2695.5000 591.7200 2697.0000 592.2000 ;
        RECT 2695.5000 586.2800 2697.0000 586.7600 ;
        RECT 2695.5000 580.8400 2697.0000 581.3200 ;
        RECT 2695.5000 575.4000 2697.0000 575.8800 ;
        RECT 2695.5000 569.9600 2697.0000 570.4400 ;
        RECT 2695.5000 564.5200 2697.0000 565.0000 ;
        RECT 2695.5000 559.0800 2697.0000 559.5600 ;
        RECT 2695.5000 553.6400 2697.0000 554.1200 ;
        RECT 2695.5000 548.2000 2697.0000 548.6800 ;
        RECT 2695.5000 542.7600 2697.0000 543.2400 ;
        RECT 2695.5000 747.6700 2789.6600 749.1700 ;
        RECT 2695.5000 536.0700 2789.6600 537.5700 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 306.4300 2697.0000 519.5300 ;
        RECT 2788.1600 306.4300 2789.6600 519.5300 ;
      LAYER met3 ;
        RECT 2788.1600 503.5200 2789.6600 504.0000 ;
        RECT 2788.1600 498.0800 2789.6600 498.5600 ;
        RECT 2788.1600 508.9600 2789.6600 509.4400 ;
        RECT 2788.1600 492.6400 2789.6600 493.1200 ;
        RECT 2788.1600 487.2000 2789.6600 487.6800 ;
        RECT 2788.1600 476.3200 2789.6600 476.8000 ;
        RECT 2788.1600 470.8800 2789.6600 471.3600 ;
        RECT 2788.1600 481.7600 2789.6600 482.2400 ;
        RECT 2788.1600 465.4400 2789.6600 465.9200 ;
        RECT 2788.1600 460.0000 2789.6600 460.4800 ;
        RECT 2788.1600 454.5600 2789.6600 455.0400 ;
        RECT 2788.1600 449.1200 2789.6600 449.6000 ;
        RECT 2788.1600 443.6800 2789.6600 444.1600 ;
        RECT 2788.1600 438.2400 2789.6600 438.7200 ;
        RECT 2788.1600 432.8000 2789.6600 433.2800 ;
        RECT 2788.1600 427.3600 2789.6600 427.8400 ;
        RECT 2788.1600 421.9200 2789.6600 422.4000 ;
        RECT 2788.1600 416.4800 2789.6600 416.9600 ;
        RECT 2695.5000 503.5200 2697.0000 504.0000 ;
        RECT 2695.5000 498.0800 2697.0000 498.5600 ;
        RECT 2695.5000 508.9600 2697.0000 509.4400 ;
        RECT 2695.5000 492.6400 2697.0000 493.1200 ;
        RECT 2695.5000 487.2000 2697.0000 487.6800 ;
        RECT 2695.5000 476.3200 2697.0000 476.8000 ;
        RECT 2695.5000 470.8800 2697.0000 471.3600 ;
        RECT 2695.5000 481.7600 2697.0000 482.2400 ;
        RECT 2695.5000 465.4400 2697.0000 465.9200 ;
        RECT 2695.5000 460.0000 2697.0000 460.4800 ;
        RECT 2695.5000 454.5600 2697.0000 455.0400 ;
        RECT 2695.5000 449.1200 2697.0000 449.6000 ;
        RECT 2695.5000 443.6800 2697.0000 444.1600 ;
        RECT 2695.5000 438.2400 2697.0000 438.7200 ;
        RECT 2695.5000 432.8000 2697.0000 433.2800 ;
        RECT 2695.5000 427.3600 2697.0000 427.8400 ;
        RECT 2695.5000 421.9200 2697.0000 422.4000 ;
        RECT 2695.5000 416.4800 2697.0000 416.9600 ;
        RECT 2788.1600 411.0400 2789.6600 411.5200 ;
        RECT 2788.1600 405.6000 2789.6600 406.0800 ;
        RECT 2788.1600 400.1600 2789.6600 400.6400 ;
        RECT 2788.1600 394.7200 2789.6600 395.2000 ;
        RECT 2788.1600 389.2800 2789.6600 389.7600 ;
        RECT 2788.1600 383.8400 2789.6600 384.3200 ;
        RECT 2788.1600 378.4000 2789.6600 378.8800 ;
        RECT 2788.1600 372.9600 2789.6600 373.4400 ;
        RECT 2788.1600 367.5200 2789.6600 368.0000 ;
        RECT 2788.1600 362.0800 2789.6600 362.5600 ;
        RECT 2788.1600 356.6400 2789.6600 357.1200 ;
        RECT 2788.1600 351.2000 2789.6600 351.6800 ;
        RECT 2788.1600 345.7600 2789.6600 346.2400 ;
        RECT 2788.1600 340.3200 2789.6600 340.8000 ;
        RECT 2788.1600 334.8800 2789.6600 335.3600 ;
        RECT 2788.1600 329.4400 2789.6600 329.9200 ;
        RECT 2788.1600 324.0000 2789.6600 324.4800 ;
        RECT 2788.1600 318.5600 2789.6600 319.0400 ;
        RECT 2788.1600 313.1200 2789.6600 313.6000 ;
        RECT 2695.5000 411.0400 2697.0000 411.5200 ;
        RECT 2695.5000 405.6000 2697.0000 406.0800 ;
        RECT 2695.5000 400.1600 2697.0000 400.6400 ;
        RECT 2695.5000 394.7200 2697.0000 395.2000 ;
        RECT 2695.5000 389.2800 2697.0000 389.7600 ;
        RECT 2695.5000 383.8400 2697.0000 384.3200 ;
        RECT 2695.5000 378.4000 2697.0000 378.8800 ;
        RECT 2695.5000 372.9600 2697.0000 373.4400 ;
        RECT 2695.5000 367.5200 2697.0000 368.0000 ;
        RECT 2695.5000 362.0800 2697.0000 362.5600 ;
        RECT 2695.5000 356.6400 2697.0000 357.1200 ;
        RECT 2695.5000 351.2000 2697.0000 351.6800 ;
        RECT 2695.5000 345.7600 2697.0000 346.2400 ;
        RECT 2695.5000 340.3200 2697.0000 340.8000 ;
        RECT 2695.5000 334.8800 2697.0000 335.3600 ;
        RECT 2695.5000 329.4400 2697.0000 329.9200 ;
        RECT 2695.5000 324.0000 2697.0000 324.4800 ;
        RECT 2695.5000 318.5600 2697.0000 319.0400 ;
        RECT 2695.5000 313.1200 2697.0000 313.6000 ;
        RECT 2695.5000 518.0300 2789.6600 519.5300 ;
        RECT 2695.5000 306.4300 2789.6600 307.9300 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 76.7900 2697.0000 289.8900 ;
        RECT 2788.1600 76.7900 2789.6600 289.8900 ;
      LAYER met3 ;
        RECT 2788.1600 273.8800 2789.6600 274.3600 ;
        RECT 2788.1600 268.4400 2789.6600 268.9200 ;
        RECT 2788.1600 279.3200 2789.6600 279.8000 ;
        RECT 2788.1600 263.0000 2789.6600 263.4800 ;
        RECT 2788.1600 257.5600 2789.6600 258.0400 ;
        RECT 2788.1600 246.6800 2789.6600 247.1600 ;
        RECT 2788.1600 241.2400 2789.6600 241.7200 ;
        RECT 2788.1600 252.1200 2789.6600 252.6000 ;
        RECT 2788.1600 235.8000 2789.6600 236.2800 ;
        RECT 2788.1600 230.3600 2789.6600 230.8400 ;
        RECT 2788.1600 224.9200 2789.6600 225.4000 ;
        RECT 2788.1600 219.4800 2789.6600 219.9600 ;
        RECT 2788.1600 214.0400 2789.6600 214.5200 ;
        RECT 2788.1600 208.6000 2789.6600 209.0800 ;
        RECT 2788.1600 203.1600 2789.6600 203.6400 ;
        RECT 2788.1600 197.7200 2789.6600 198.2000 ;
        RECT 2788.1600 192.2800 2789.6600 192.7600 ;
        RECT 2788.1600 186.8400 2789.6600 187.3200 ;
        RECT 2695.5000 273.8800 2697.0000 274.3600 ;
        RECT 2695.5000 268.4400 2697.0000 268.9200 ;
        RECT 2695.5000 279.3200 2697.0000 279.8000 ;
        RECT 2695.5000 263.0000 2697.0000 263.4800 ;
        RECT 2695.5000 257.5600 2697.0000 258.0400 ;
        RECT 2695.5000 246.6800 2697.0000 247.1600 ;
        RECT 2695.5000 241.2400 2697.0000 241.7200 ;
        RECT 2695.5000 252.1200 2697.0000 252.6000 ;
        RECT 2695.5000 235.8000 2697.0000 236.2800 ;
        RECT 2695.5000 230.3600 2697.0000 230.8400 ;
        RECT 2695.5000 224.9200 2697.0000 225.4000 ;
        RECT 2695.5000 219.4800 2697.0000 219.9600 ;
        RECT 2695.5000 214.0400 2697.0000 214.5200 ;
        RECT 2695.5000 208.6000 2697.0000 209.0800 ;
        RECT 2695.5000 203.1600 2697.0000 203.6400 ;
        RECT 2695.5000 197.7200 2697.0000 198.2000 ;
        RECT 2695.5000 192.2800 2697.0000 192.7600 ;
        RECT 2695.5000 186.8400 2697.0000 187.3200 ;
        RECT 2788.1600 181.4000 2789.6600 181.8800 ;
        RECT 2788.1600 175.9600 2789.6600 176.4400 ;
        RECT 2788.1600 170.5200 2789.6600 171.0000 ;
        RECT 2788.1600 165.0800 2789.6600 165.5600 ;
        RECT 2788.1600 159.6400 2789.6600 160.1200 ;
        RECT 2788.1600 154.2000 2789.6600 154.6800 ;
        RECT 2788.1600 148.7600 2789.6600 149.2400 ;
        RECT 2788.1600 143.3200 2789.6600 143.8000 ;
        RECT 2788.1600 137.8800 2789.6600 138.3600 ;
        RECT 2788.1600 132.4400 2789.6600 132.9200 ;
        RECT 2788.1600 127.0000 2789.6600 127.4800 ;
        RECT 2788.1600 121.5600 2789.6600 122.0400 ;
        RECT 2788.1600 116.1200 2789.6600 116.6000 ;
        RECT 2788.1600 110.6800 2789.6600 111.1600 ;
        RECT 2788.1600 105.2400 2789.6600 105.7200 ;
        RECT 2788.1600 99.8000 2789.6600 100.2800 ;
        RECT 2788.1600 94.3600 2789.6600 94.8400 ;
        RECT 2788.1600 88.9200 2789.6600 89.4000 ;
        RECT 2788.1600 83.4800 2789.6600 83.9600 ;
        RECT 2695.5000 181.4000 2697.0000 181.8800 ;
        RECT 2695.5000 175.9600 2697.0000 176.4400 ;
        RECT 2695.5000 170.5200 2697.0000 171.0000 ;
        RECT 2695.5000 165.0800 2697.0000 165.5600 ;
        RECT 2695.5000 159.6400 2697.0000 160.1200 ;
        RECT 2695.5000 154.2000 2697.0000 154.6800 ;
        RECT 2695.5000 148.7600 2697.0000 149.2400 ;
        RECT 2695.5000 143.3200 2697.0000 143.8000 ;
        RECT 2695.5000 137.8800 2697.0000 138.3600 ;
        RECT 2695.5000 132.4400 2697.0000 132.9200 ;
        RECT 2695.5000 127.0000 2697.0000 127.4800 ;
        RECT 2695.5000 121.5600 2697.0000 122.0400 ;
        RECT 2695.5000 116.1200 2697.0000 116.6000 ;
        RECT 2695.5000 110.6800 2697.0000 111.1600 ;
        RECT 2695.5000 105.2400 2697.0000 105.7200 ;
        RECT 2695.5000 99.8000 2697.0000 100.2800 ;
        RECT 2695.5000 94.3600 2697.0000 94.8400 ;
        RECT 2695.5000 88.9200 2697.0000 89.4000 ;
        RECT 2695.5000 83.4800 2697.0000 83.9600 ;
        RECT 2695.5000 288.3900 2789.6600 289.8900 ;
        RECT 2695.5000 76.7900 2789.6600 78.2900 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'S_term_RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2788.1600 34.6700 2790.1600 61.6000 ;
        RECT 2695.0000 34.6700 2697.0000 61.6000 ;
      LAYER met3 ;
        RECT 2788.1600 51.3800 2790.1600 51.8600 ;
        RECT 2695.0000 51.3800 2697.0000 51.8600 ;
        RECT 2788.1600 40.5000 2790.1600 40.9800 ;
        RECT 2788.1600 45.9400 2790.1600 46.4200 ;
        RECT 2695.0000 40.5000 2697.0000 40.9800 ;
        RECT 2695.0000 45.9400 2697.0000 46.4200 ;
        RECT 2695.0000 59.6000 2790.1600 61.6000 ;
        RECT 2695.0000 34.6700 2790.1600 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 2602.8300 2697.0000 2815.9300 ;
        RECT 2788.1600 2602.8300 2789.6600 2815.9300 ;
      LAYER met3 ;
        RECT 2788.1600 2799.9200 2789.6600 2800.4000 ;
        RECT 2788.1600 2794.4800 2789.6600 2794.9600 ;
        RECT 2788.1600 2805.3600 2789.6600 2805.8400 ;
        RECT 2788.1600 2789.0400 2789.6600 2789.5200 ;
        RECT 2788.1600 2783.6000 2789.6600 2784.0800 ;
        RECT 2788.1600 2772.7200 2789.6600 2773.2000 ;
        RECT 2788.1600 2767.2800 2789.6600 2767.7600 ;
        RECT 2788.1600 2778.1600 2789.6600 2778.6400 ;
        RECT 2788.1600 2761.8400 2789.6600 2762.3200 ;
        RECT 2788.1600 2756.4000 2789.6600 2756.8800 ;
        RECT 2788.1600 2750.9600 2789.6600 2751.4400 ;
        RECT 2788.1600 2745.5200 2789.6600 2746.0000 ;
        RECT 2788.1600 2740.0800 2789.6600 2740.5600 ;
        RECT 2788.1600 2734.6400 2789.6600 2735.1200 ;
        RECT 2788.1600 2729.2000 2789.6600 2729.6800 ;
        RECT 2788.1600 2723.7600 2789.6600 2724.2400 ;
        RECT 2788.1600 2718.3200 2789.6600 2718.8000 ;
        RECT 2788.1600 2712.8800 2789.6600 2713.3600 ;
        RECT 2695.5000 2799.9200 2697.0000 2800.4000 ;
        RECT 2695.5000 2794.4800 2697.0000 2794.9600 ;
        RECT 2695.5000 2805.3600 2697.0000 2805.8400 ;
        RECT 2695.5000 2789.0400 2697.0000 2789.5200 ;
        RECT 2695.5000 2783.6000 2697.0000 2784.0800 ;
        RECT 2695.5000 2772.7200 2697.0000 2773.2000 ;
        RECT 2695.5000 2767.2800 2697.0000 2767.7600 ;
        RECT 2695.5000 2778.1600 2697.0000 2778.6400 ;
        RECT 2695.5000 2761.8400 2697.0000 2762.3200 ;
        RECT 2695.5000 2756.4000 2697.0000 2756.8800 ;
        RECT 2695.5000 2750.9600 2697.0000 2751.4400 ;
        RECT 2695.5000 2745.5200 2697.0000 2746.0000 ;
        RECT 2695.5000 2740.0800 2697.0000 2740.5600 ;
        RECT 2695.5000 2734.6400 2697.0000 2735.1200 ;
        RECT 2695.5000 2729.2000 2697.0000 2729.6800 ;
        RECT 2695.5000 2723.7600 2697.0000 2724.2400 ;
        RECT 2695.5000 2718.3200 2697.0000 2718.8000 ;
        RECT 2695.5000 2712.8800 2697.0000 2713.3600 ;
        RECT 2788.1600 2707.4400 2789.6600 2707.9200 ;
        RECT 2788.1600 2702.0000 2789.6600 2702.4800 ;
        RECT 2788.1600 2696.5600 2789.6600 2697.0400 ;
        RECT 2788.1600 2691.1200 2789.6600 2691.6000 ;
        RECT 2788.1600 2685.6800 2789.6600 2686.1600 ;
        RECT 2788.1600 2680.2400 2789.6600 2680.7200 ;
        RECT 2788.1600 2674.8000 2789.6600 2675.2800 ;
        RECT 2788.1600 2669.3600 2789.6600 2669.8400 ;
        RECT 2788.1600 2663.9200 2789.6600 2664.4000 ;
        RECT 2788.1600 2658.4800 2789.6600 2658.9600 ;
        RECT 2788.1600 2653.0400 2789.6600 2653.5200 ;
        RECT 2788.1600 2647.6000 2789.6600 2648.0800 ;
        RECT 2788.1600 2642.1600 2789.6600 2642.6400 ;
        RECT 2788.1600 2636.7200 2789.6600 2637.2000 ;
        RECT 2788.1600 2631.2800 2789.6600 2631.7600 ;
        RECT 2788.1600 2625.8400 2789.6600 2626.3200 ;
        RECT 2788.1600 2620.4000 2789.6600 2620.8800 ;
        RECT 2788.1600 2614.9600 2789.6600 2615.4400 ;
        RECT 2788.1600 2609.5200 2789.6600 2610.0000 ;
        RECT 2695.5000 2707.4400 2697.0000 2707.9200 ;
        RECT 2695.5000 2702.0000 2697.0000 2702.4800 ;
        RECT 2695.5000 2696.5600 2697.0000 2697.0400 ;
        RECT 2695.5000 2691.1200 2697.0000 2691.6000 ;
        RECT 2695.5000 2685.6800 2697.0000 2686.1600 ;
        RECT 2695.5000 2680.2400 2697.0000 2680.7200 ;
        RECT 2695.5000 2674.8000 2697.0000 2675.2800 ;
        RECT 2695.5000 2669.3600 2697.0000 2669.8400 ;
        RECT 2695.5000 2663.9200 2697.0000 2664.4000 ;
        RECT 2695.5000 2658.4800 2697.0000 2658.9600 ;
        RECT 2695.5000 2653.0400 2697.0000 2653.5200 ;
        RECT 2695.5000 2647.6000 2697.0000 2648.0800 ;
        RECT 2695.5000 2642.1600 2697.0000 2642.6400 ;
        RECT 2695.5000 2636.7200 2697.0000 2637.2000 ;
        RECT 2695.5000 2631.2800 2697.0000 2631.7600 ;
        RECT 2695.5000 2625.8400 2697.0000 2626.3200 ;
        RECT 2695.5000 2620.4000 2697.0000 2620.8800 ;
        RECT 2695.5000 2614.9600 2697.0000 2615.4400 ;
        RECT 2695.5000 2609.5200 2697.0000 2610.0000 ;
        RECT 2695.5000 2814.4300 2789.6600 2815.9300 ;
        RECT 2695.5000 2602.8300 2789.6600 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 2373.1900 2697.0000 2586.2900 ;
        RECT 2788.1600 2373.1900 2789.6600 2586.2900 ;
      LAYER met3 ;
        RECT 2788.1600 2570.2800 2789.6600 2570.7600 ;
        RECT 2788.1600 2564.8400 2789.6600 2565.3200 ;
        RECT 2788.1600 2575.7200 2789.6600 2576.2000 ;
        RECT 2788.1600 2559.4000 2789.6600 2559.8800 ;
        RECT 2788.1600 2553.9600 2789.6600 2554.4400 ;
        RECT 2788.1600 2543.0800 2789.6600 2543.5600 ;
        RECT 2788.1600 2537.6400 2789.6600 2538.1200 ;
        RECT 2788.1600 2548.5200 2789.6600 2549.0000 ;
        RECT 2788.1600 2532.2000 2789.6600 2532.6800 ;
        RECT 2788.1600 2526.7600 2789.6600 2527.2400 ;
        RECT 2788.1600 2521.3200 2789.6600 2521.8000 ;
        RECT 2788.1600 2515.8800 2789.6600 2516.3600 ;
        RECT 2788.1600 2510.4400 2789.6600 2510.9200 ;
        RECT 2788.1600 2505.0000 2789.6600 2505.4800 ;
        RECT 2788.1600 2499.5600 2789.6600 2500.0400 ;
        RECT 2788.1600 2494.1200 2789.6600 2494.6000 ;
        RECT 2788.1600 2488.6800 2789.6600 2489.1600 ;
        RECT 2788.1600 2483.2400 2789.6600 2483.7200 ;
        RECT 2695.5000 2570.2800 2697.0000 2570.7600 ;
        RECT 2695.5000 2564.8400 2697.0000 2565.3200 ;
        RECT 2695.5000 2575.7200 2697.0000 2576.2000 ;
        RECT 2695.5000 2559.4000 2697.0000 2559.8800 ;
        RECT 2695.5000 2553.9600 2697.0000 2554.4400 ;
        RECT 2695.5000 2543.0800 2697.0000 2543.5600 ;
        RECT 2695.5000 2537.6400 2697.0000 2538.1200 ;
        RECT 2695.5000 2548.5200 2697.0000 2549.0000 ;
        RECT 2695.5000 2532.2000 2697.0000 2532.6800 ;
        RECT 2695.5000 2526.7600 2697.0000 2527.2400 ;
        RECT 2695.5000 2521.3200 2697.0000 2521.8000 ;
        RECT 2695.5000 2515.8800 2697.0000 2516.3600 ;
        RECT 2695.5000 2510.4400 2697.0000 2510.9200 ;
        RECT 2695.5000 2505.0000 2697.0000 2505.4800 ;
        RECT 2695.5000 2499.5600 2697.0000 2500.0400 ;
        RECT 2695.5000 2494.1200 2697.0000 2494.6000 ;
        RECT 2695.5000 2488.6800 2697.0000 2489.1600 ;
        RECT 2695.5000 2483.2400 2697.0000 2483.7200 ;
        RECT 2788.1600 2477.8000 2789.6600 2478.2800 ;
        RECT 2788.1600 2472.3600 2789.6600 2472.8400 ;
        RECT 2788.1600 2466.9200 2789.6600 2467.4000 ;
        RECT 2788.1600 2461.4800 2789.6600 2461.9600 ;
        RECT 2788.1600 2456.0400 2789.6600 2456.5200 ;
        RECT 2788.1600 2450.6000 2789.6600 2451.0800 ;
        RECT 2788.1600 2445.1600 2789.6600 2445.6400 ;
        RECT 2788.1600 2439.7200 2789.6600 2440.2000 ;
        RECT 2788.1600 2434.2800 2789.6600 2434.7600 ;
        RECT 2788.1600 2428.8400 2789.6600 2429.3200 ;
        RECT 2788.1600 2423.4000 2789.6600 2423.8800 ;
        RECT 2788.1600 2417.9600 2789.6600 2418.4400 ;
        RECT 2788.1600 2412.5200 2789.6600 2413.0000 ;
        RECT 2788.1600 2407.0800 2789.6600 2407.5600 ;
        RECT 2788.1600 2401.6400 2789.6600 2402.1200 ;
        RECT 2788.1600 2396.2000 2789.6600 2396.6800 ;
        RECT 2788.1600 2390.7600 2789.6600 2391.2400 ;
        RECT 2788.1600 2385.3200 2789.6600 2385.8000 ;
        RECT 2788.1600 2379.8800 2789.6600 2380.3600 ;
        RECT 2695.5000 2477.8000 2697.0000 2478.2800 ;
        RECT 2695.5000 2472.3600 2697.0000 2472.8400 ;
        RECT 2695.5000 2466.9200 2697.0000 2467.4000 ;
        RECT 2695.5000 2461.4800 2697.0000 2461.9600 ;
        RECT 2695.5000 2456.0400 2697.0000 2456.5200 ;
        RECT 2695.5000 2450.6000 2697.0000 2451.0800 ;
        RECT 2695.5000 2445.1600 2697.0000 2445.6400 ;
        RECT 2695.5000 2439.7200 2697.0000 2440.2000 ;
        RECT 2695.5000 2434.2800 2697.0000 2434.7600 ;
        RECT 2695.5000 2428.8400 2697.0000 2429.3200 ;
        RECT 2695.5000 2423.4000 2697.0000 2423.8800 ;
        RECT 2695.5000 2417.9600 2697.0000 2418.4400 ;
        RECT 2695.5000 2412.5200 2697.0000 2413.0000 ;
        RECT 2695.5000 2407.0800 2697.0000 2407.5600 ;
        RECT 2695.5000 2401.6400 2697.0000 2402.1200 ;
        RECT 2695.5000 2396.2000 2697.0000 2396.6800 ;
        RECT 2695.5000 2390.7600 2697.0000 2391.2400 ;
        RECT 2695.5000 2385.3200 2697.0000 2385.8000 ;
        RECT 2695.5000 2379.8800 2697.0000 2380.3600 ;
        RECT 2695.5000 2584.7900 2789.6600 2586.2900 ;
        RECT 2695.5000 2373.1900 2789.6600 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 2143.5500 2697.0000 2356.6500 ;
        RECT 2788.1600 2143.5500 2789.6600 2356.6500 ;
      LAYER met3 ;
        RECT 2788.1600 2340.6400 2789.6600 2341.1200 ;
        RECT 2788.1600 2335.2000 2789.6600 2335.6800 ;
        RECT 2788.1600 2346.0800 2789.6600 2346.5600 ;
        RECT 2788.1600 2329.7600 2789.6600 2330.2400 ;
        RECT 2788.1600 2324.3200 2789.6600 2324.8000 ;
        RECT 2788.1600 2313.4400 2789.6600 2313.9200 ;
        RECT 2788.1600 2308.0000 2789.6600 2308.4800 ;
        RECT 2788.1600 2318.8800 2789.6600 2319.3600 ;
        RECT 2788.1600 2302.5600 2789.6600 2303.0400 ;
        RECT 2788.1600 2297.1200 2789.6600 2297.6000 ;
        RECT 2788.1600 2291.6800 2789.6600 2292.1600 ;
        RECT 2788.1600 2286.2400 2789.6600 2286.7200 ;
        RECT 2788.1600 2280.8000 2789.6600 2281.2800 ;
        RECT 2788.1600 2275.3600 2789.6600 2275.8400 ;
        RECT 2788.1600 2269.9200 2789.6600 2270.4000 ;
        RECT 2788.1600 2264.4800 2789.6600 2264.9600 ;
        RECT 2788.1600 2259.0400 2789.6600 2259.5200 ;
        RECT 2788.1600 2253.6000 2789.6600 2254.0800 ;
        RECT 2695.5000 2340.6400 2697.0000 2341.1200 ;
        RECT 2695.5000 2335.2000 2697.0000 2335.6800 ;
        RECT 2695.5000 2346.0800 2697.0000 2346.5600 ;
        RECT 2695.5000 2329.7600 2697.0000 2330.2400 ;
        RECT 2695.5000 2324.3200 2697.0000 2324.8000 ;
        RECT 2695.5000 2313.4400 2697.0000 2313.9200 ;
        RECT 2695.5000 2308.0000 2697.0000 2308.4800 ;
        RECT 2695.5000 2318.8800 2697.0000 2319.3600 ;
        RECT 2695.5000 2302.5600 2697.0000 2303.0400 ;
        RECT 2695.5000 2297.1200 2697.0000 2297.6000 ;
        RECT 2695.5000 2291.6800 2697.0000 2292.1600 ;
        RECT 2695.5000 2286.2400 2697.0000 2286.7200 ;
        RECT 2695.5000 2280.8000 2697.0000 2281.2800 ;
        RECT 2695.5000 2275.3600 2697.0000 2275.8400 ;
        RECT 2695.5000 2269.9200 2697.0000 2270.4000 ;
        RECT 2695.5000 2264.4800 2697.0000 2264.9600 ;
        RECT 2695.5000 2259.0400 2697.0000 2259.5200 ;
        RECT 2695.5000 2253.6000 2697.0000 2254.0800 ;
        RECT 2788.1600 2248.1600 2789.6600 2248.6400 ;
        RECT 2788.1600 2242.7200 2789.6600 2243.2000 ;
        RECT 2788.1600 2237.2800 2789.6600 2237.7600 ;
        RECT 2788.1600 2231.8400 2789.6600 2232.3200 ;
        RECT 2788.1600 2226.4000 2789.6600 2226.8800 ;
        RECT 2788.1600 2220.9600 2789.6600 2221.4400 ;
        RECT 2788.1600 2215.5200 2789.6600 2216.0000 ;
        RECT 2788.1600 2210.0800 2789.6600 2210.5600 ;
        RECT 2788.1600 2204.6400 2789.6600 2205.1200 ;
        RECT 2788.1600 2199.2000 2789.6600 2199.6800 ;
        RECT 2788.1600 2193.7600 2789.6600 2194.2400 ;
        RECT 2788.1600 2188.3200 2789.6600 2188.8000 ;
        RECT 2788.1600 2182.8800 2789.6600 2183.3600 ;
        RECT 2788.1600 2177.4400 2789.6600 2177.9200 ;
        RECT 2788.1600 2172.0000 2789.6600 2172.4800 ;
        RECT 2788.1600 2166.5600 2789.6600 2167.0400 ;
        RECT 2788.1600 2161.1200 2789.6600 2161.6000 ;
        RECT 2788.1600 2155.6800 2789.6600 2156.1600 ;
        RECT 2788.1600 2150.2400 2789.6600 2150.7200 ;
        RECT 2695.5000 2248.1600 2697.0000 2248.6400 ;
        RECT 2695.5000 2242.7200 2697.0000 2243.2000 ;
        RECT 2695.5000 2237.2800 2697.0000 2237.7600 ;
        RECT 2695.5000 2231.8400 2697.0000 2232.3200 ;
        RECT 2695.5000 2226.4000 2697.0000 2226.8800 ;
        RECT 2695.5000 2220.9600 2697.0000 2221.4400 ;
        RECT 2695.5000 2215.5200 2697.0000 2216.0000 ;
        RECT 2695.5000 2210.0800 2697.0000 2210.5600 ;
        RECT 2695.5000 2204.6400 2697.0000 2205.1200 ;
        RECT 2695.5000 2199.2000 2697.0000 2199.6800 ;
        RECT 2695.5000 2193.7600 2697.0000 2194.2400 ;
        RECT 2695.5000 2188.3200 2697.0000 2188.8000 ;
        RECT 2695.5000 2182.8800 2697.0000 2183.3600 ;
        RECT 2695.5000 2177.4400 2697.0000 2177.9200 ;
        RECT 2695.5000 2172.0000 2697.0000 2172.4800 ;
        RECT 2695.5000 2166.5600 2697.0000 2167.0400 ;
        RECT 2695.5000 2161.1200 2697.0000 2161.6000 ;
        RECT 2695.5000 2155.6800 2697.0000 2156.1600 ;
        RECT 2695.5000 2150.2400 2697.0000 2150.7200 ;
        RECT 2695.5000 2355.1500 2789.6600 2356.6500 ;
        RECT 2695.5000 2143.5500 2789.6600 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 1913.9100 2697.0000 2127.0100 ;
        RECT 2788.1600 1913.9100 2789.6600 2127.0100 ;
      LAYER met3 ;
        RECT 2788.1600 2111.0000 2789.6600 2111.4800 ;
        RECT 2788.1600 2105.5600 2789.6600 2106.0400 ;
        RECT 2788.1600 2116.4400 2789.6600 2116.9200 ;
        RECT 2788.1600 2100.1200 2789.6600 2100.6000 ;
        RECT 2788.1600 2094.6800 2789.6600 2095.1600 ;
        RECT 2788.1600 2083.8000 2789.6600 2084.2800 ;
        RECT 2788.1600 2078.3600 2789.6600 2078.8400 ;
        RECT 2788.1600 2089.2400 2789.6600 2089.7200 ;
        RECT 2788.1600 2072.9200 2789.6600 2073.4000 ;
        RECT 2788.1600 2067.4800 2789.6600 2067.9600 ;
        RECT 2788.1600 2062.0400 2789.6600 2062.5200 ;
        RECT 2788.1600 2056.6000 2789.6600 2057.0800 ;
        RECT 2788.1600 2051.1600 2789.6600 2051.6400 ;
        RECT 2788.1600 2045.7200 2789.6600 2046.2000 ;
        RECT 2788.1600 2040.2800 2789.6600 2040.7600 ;
        RECT 2788.1600 2034.8400 2789.6600 2035.3200 ;
        RECT 2788.1600 2029.4000 2789.6600 2029.8800 ;
        RECT 2788.1600 2023.9600 2789.6600 2024.4400 ;
        RECT 2695.5000 2111.0000 2697.0000 2111.4800 ;
        RECT 2695.5000 2105.5600 2697.0000 2106.0400 ;
        RECT 2695.5000 2116.4400 2697.0000 2116.9200 ;
        RECT 2695.5000 2100.1200 2697.0000 2100.6000 ;
        RECT 2695.5000 2094.6800 2697.0000 2095.1600 ;
        RECT 2695.5000 2083.8000 2697.0000 2084.2800 ;
        RECT 2695.5000 2078.3600 2697.0000 2078.8400 ;
        RECT 2695.5000 2089.2400 2697.0000 2089.7200 ;
        RECT 2695.5000 2072.9200 2697.0000 2073.4000 ;
        RECT 2695.5000 2067.4800 2697.0000 2067.9600 ;
        RECT 2695.5000 2062.0400 2697.0000 2062.5200 ;
        RECT 2695.5000 2056.6000 2697.0000 2057.0800 ;
        RECT 2695.5000 2051.1600 2697.0000 2051.6400 ;
        RECT 2695.5000 2045.7200 2697.0000 2046.2000 ;
        RECT 2695.5000 2040.2800 2697.0000 2040.7600 ;
        RECT 2695.5000 2034.8400 2697.0000 2035.3200 ;
        RECT 2695.5000 2029.4000 2697.0000 2029.8800 ;
        RECT 2695.5000 2023.9600 2697.0000 2024.4400 ;
        RECT 2788.1600 2018.5200 2789.6600 2019.0000 ;
        RECT 2788.1600 2013.0800 2789.6600 2013.5600 ;
        RECT 2788.1600 2007.6400 2789.6600 2008.1200 ;
        RECT 2788.1600 2002.2000 2789.6600 2002.6800 ;
        RECT 2788.1600 1996.7600 2789.6600 1997.2400 ;
        RECT 2788.1600 1991.3200 2789.6600 1991.8000 ;
        RECT 2788.1600 1985.8800 2789.6600 1986.3600 ;
        RECT 2788.1600 1980.4400 2789.6600 1980.9200 ;
        RECT 2788.1600 1975.0000 2789.6600 1975.4800 ;
        RECT 2788.1600 1969.5600 2789.6600 1970.0400 ;
        RECT 2788.1600 1964.1200 2789.6600 1964.6000 ;
        RECT 2788.1600 1958.6800 2789.6600 1959.1600 ;
        RECT 2788.1600 1953.2400 2789.6600 1953.7200 ;
        RECT 2788.1600 1947.8000 2789.6600 1948.2800 ;
        RECT 2788.1600 1942.3600 2789.6600 1942.8400 ;
        RECT 2788.1600 1936.9200 2789.6600 1937.4000 ;
        RECT 2788.1600 1931.4800 2789.6600 1931.9600 ;
        RECT 2788.1600 1926.0400 2789.6600 1926.5200 ;
        RECT 2788.1600 1920.6000 2789.6600 1921.0800 ;
        RECT 2695.5000 2018.5200 2697.0000 2019.0000 ;
        RECT 2695.5000 2013.0800 2697.0000 2013.5600 ;
        RECT 2695.5000 2007.6400 2697.0000 2008.1200 ;
        RECT 2695.5000 2002.2000 2697.0000 2002.6800 ;
        RECT 2695.5000 1996.7600 2697.0000 1997.2400 ;
        RECT 2695.5000 1991.3200 2697.0000 1991.8000 ;
        RECT 2695.5000 1985.8800 2697.0000 1986.3600 ;
        RECT 2695.5000 1980.4400 2697.0000 1980.9200 ;
        RECT 2695.5000 1975.0000 2697.0000 1975.4800 ;
        RECT 2695.5000 1969.5600 2697.0000 1970.0400 ;
        RECT 2695.5000 1964.1200 2697.0000 1964.6000 ;
        RECT 2695.5000 1958.6800 2697.0000 1959.1600 ;
        RECT 2695.5000 1953.2400 2697.0000 1953.7200 ;
        RECT 2695.5000 1947.8000 2697.0000 1948.2800 ;
        RECT 2695.5000 1942.3600 2697.0000 1942.8400 ;
        RECT 2695.5000 1936.9200 2697.0000 1937.4000 ;
        RECT 2695.5000 1931.4800 2697.0000 1931.9600 ;
        RECT 2695.5000 1926.0400 2697.0000 1926.5200 ;
        RECT 2695.5000 1920.6000 2697.0000 1921.0800 ;
        RECT 2695.5000 2125.5100 2789.6600 2127.0100 ;
        RECT 2695.5000 1913.9100 2789.6600 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 1684.2700 2697.0000 1897.3700 ;
        RECT 2788.1600 1684.2700 2789.6600 1897.3700 ;
      LAYER met3 ;
        RECT 2788.1600 1881.3600 2789.6600 1881.8400 ;
        RECT 2788.1600 1875.9200 2789.6600 1876.4000 ;
        RECT 2788.1600 1886.8000 2789.6600 1887.2800 ;
        RECT 2788.1600 1870.4800 2789.6600 1870.9600 ;
        RECT 2788.1600 1865.0400 2789.6600 1865.5200 ;
        RECT 2788.1600 1854.1600 2789.6600 1854.6400 ;
        RECT 2788.1600 1848.7200 2789.6600 1849.2000 ;
        RECT 2788.1600 1859.6000 2789.6600 1860.0800 ;
        RECT 2788.1600 1843.2800 2789.6600 1843.7600 ;
        RECT 2788.1600 1837.8400 2789.6600 1838.3200 ;
        RECT 2788.1600 1832.4000 2789.6600 1832.8800 ;
        RECT 2788.1600 1826.9600 2789.6600 1827.4400 ;
        RECT 2788.1600 1821.5200 2789.6600 1822.0000 ;
        RECT 2788.1600 1816.0800 2789.6600 1816.5600 ;
        RECT 2788.1600 1810.6400 2789.6600 1811.1200 ;
        RECT 2788.1600 1805.2000 2789.6600 1805.6800 ;
        RECT 2788.1600 1799.7600 2789.6600 1800.2400 ;
        RECT 2788.1600 1794.3200 2789.6600 1794.8000 ;
        RECT 2695.5000 1881.3600 2697.0000 1881.8400 ;
        RECT 2695.5000 1875.9200 2697.0000 1876.4000 ;
        RECT 2695.5000 1886.8000 2697.0000 1887.2800 ;
        RECT 2695.5000 1870.4800 2697.0000 1870.9600 ;
        RECT 2695.5000 1865.0400 2697.0000 1865.5200 ;
        RECT 2695.5000 1854.1600 2697.0000 1854.6400 ;
        RECT 2695.5000 1848.7200 2697.0000 1849.2000 ;
        RECT 2695.5000 1859.6000 2697.0000 1860.0800 ;
        RECT 2695.5000 1843.2800 2697.0000 1843.7600 ;
        RECT 2695.5000 1837.8400 2697.0000 1838.3200 ;
        RECT 2695.5000 1832.4000 2697.0000 1832.8800 ;
        RECT 2695.5000 1826.9600 2697.0000 1827.4400 ;
        RECT 2695.5000 1821.5200 2697.0000 1822.0000 ;
        RECT 2695.5000 1816.0800 2697.0000 1816.5600 ;
        RECT 2695.5000 1810.6400 2697.0000 1811.1200 ;
        RECT 2695.5000 1805.2000 2697.0000 1805.6800 ;
        RECT 2695.5000 1799.7600 2697.0000 1800.2400 ;
        RECT 2695.5000 1794.3200 2697.0000 1794.8000 ;
        RECT 2788.1600 1788.8800 2789.6600 1789.3600 ;
        RECT 2788.1600 1783.4400 2789.6600 1783.9200 ;
        RECT 2788.1600 1778.0000 2789.6600 1778.4800 ;
        RECT 2788.1600 1772.5600 2789.6600 1773.0400 ;
        RECT 2788.1600 1767.1200 2789.6600 1767.6000 ;
        RECT 2788.1600 1761.6800 2789.6600 1762.1600 ;
        RECT 2788.1600 1756.2400 2789.6600 1756.7200 ;
        RECT 2788.1600 1750.8000 2789.6600 1751.2800 ;
        RECT 2788.1600 1745.3600 2789.6600 1745.8400 ;
        RECT 2788.1600 1739.9200 2789.6600 1740.4000 ;
        RECT 2788.1600 1734.4800 2789.6600 1734.9600 ;
        RECT 2788.1600 1729.0400 2789.6600 1729.5200 ;
        RECT 2788.1600 1723.6000 2789.6600 1724.0800 ;
        RECT 2788.1600 1718.1600 2789.6600 1718.6400 ;
        RECT 2788.1600 1712.7200 2789.6600 1713.2000 ;
        RECT 2788.1600 1707.2800 2789.6600 1707.7600 ;
        RECT 2788.1600 1701.8400 2789.6600 1702.3200 ;
        RECT 2788.1600 1696.4000 2789.6600 1696.8800 ;
        RECT 2788.1600 1690.9600 2789.6600 1691.4400 ;
        RECT 2695.5000 1788.8800 2697.0000 1789.3600 ;
        RECT 2695.5000 1783.4400 2697.0000 1783.9200 ;
        RECT 2695.5000 1778.0000 2697.0000 1778.4800 ;
        RECT 2695.5000 1772.5600 2697.0000 1773.0400 ;
        RECT 2695.5000 1767.1200 2697.0000 1767.6000 ;
        RECT 2695.5000 1761.6800 2697.0000 1762.1600 ;
        RECT 2695.5000 1756.2400 2697.0000 1756.7200 ;
        RECT 2695.5000 1750.8000 2697.0000 1751.2800 ;
        RECT 2695.5000 1745.3600 2697.0000 1745.8400 ;
        RECT 2695.5000 1739.9200 2697.0000 1740.4000 ;
        RECT 2695.5000 1734.4800 2697.0000 1734.9600 ;
        RECT 2695.5000 1729.0400 2697.0000 1729.5200 ;
        RECT 2695.5000 1723.6000 2697.0000 1724.0800 ;
        RECT 2695.5000 1718.1600 2697.0000 1718.6400 ;
        RECT 2695.5000 1712.7200 2697.0000 1713.2000 ;
        RECT 2695.5000 1707.2800 2697.0000 1707.7600 ;
        RECT 2695.5000 1701.8400 2697.0000 1702.3200 ;
        RECT 2695.5000 1696.4000 2697.0000 1696.8800 ;
        RECT 2695.5000 1690.9600 2697.0000 1691.4400 ;
        RECT 2695.5000 1895.8700 2789.6600 1897.3700 ;
        RECT 2695.5000 1684.2700 2789.6600 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 1454.6300 2697.0000 1667.7300 ;
        RECT 2788.1600 1454.6300 2789.6600 1667.7300 ;
      LAYER met3 ;
        RECT 2788.1600 1651.7200 2789.6600 1652.2000 ;
        RECT 2788.1600 1646.2800 2789.6600 1646.7600 ;
        RECT 2788.1600 1657.1600 2789.6600 1657.6400 ;
        RECT 2788.1600 1640.8400 2789.6600 1641.3200 ;
        RECT 2788.1600 1635.4000 2789.6600 1635.8800 ;
        RECT 2788.1600 1624.5200 2789.6600 1625.0000 ;
        RECT 2788.1600 1619.0800 2789.6600 1619.5600 ;
        RECT 2788.1600 1629.9600 2789.6600 1630.4400 ;
        RECT 2788.1600 1613.6400 2789.6600 1614.1200 ;
        RECT 2788.1600 1608.2000 2789.6600 1608.6800 ;
        RECT 2788.1600 1602.7600 2789.6600 1603.2400 ;
        RECT 2788.1600 1597.3200 2789.6600 1597.8000 ;
        RECT 2788.1600 1591.8800 2789.6600 1592.3600 ;
        RECT 2788.1600 1586.4400 2789.6600 1586.9200 ;
        RECT 2788.1600 1581.0000 2789.6600 1581.4800 ;
        RECT 2788.1600 1575.5600 2789.6600 1576.0400 ;
        RECT 2788.1600 1570.1200 2789.6600 1570.6000 ;
        RECT 2788.1600 1564.6800 2789.6600 1565.1600 ;
        RECT 2695.5000 1651.7200 2697.0000 1652.2000 ;
        RECT 2695.5000 1646.2800 2697.0000 1646.7600 ;
        RECT 2695.5000 1657.1600 2697.0000 1657.6400 ;
        RECT 2695.5000 1640.8400 2697.0000 1641.3200 ;
        RECT 2695.5000 1635.4000 2697.0000 1635.8800 ;
        RECT 2695.5000 1624.5200 2697.0000 1625.0000 ;
        RECT 2695.5000 1619.0800 2697.0000 1619.5600 ;
        RECT 2695.5000 1629.9600 2697.0000 1630.4400 ;
        RECT 2695.5000 1613.6400 2697.0000 1614.1200 ;
        RECT 2695.5000 1608.2000 2697.0000 1608.6800 ;
        RECT 2695.5000 1602.7600 2697.0000 1603.2400 ;
        RECT 2695.5000 1597.3200 2697.0000 1597.8000 ;
        RECT 2695.5000 1591.8800 2697.0000 1592.3600 ;
        RECT 2695.5000 1586.4400 2697.0000 1586.9200 ;
        RECT 2695.5000 1581.0000 2697.0000 1581.4800 ;
        RECT 2695.5000 1575.5600 2697.0000 1576.0400 ;
        RECT 2695.5000 1570.1200 2697.0000 1570.6000 ;
        RECT 2695.5000 1564.6800 2697.0000 1565.1600 ;
        RECT 2788.1600 1559.2400 2789.6600 1559.7200 ;
        RECT 2788.1600 1553.8000 2789.6600 1554.2800 ;
        RECT 2788.1600 1548.3600 2789.6600 1548.8400 ;
        RECT 2788.1600 1542.9200 2789.6600 1543.4000 ;
        RECT 2788.1600 1537.4800 2789.6600 1537.9600 ;
        RECT 2788.1600 1532.0400 2789.6600 1532.5200 ;
        RECT 2788.1600 1526.6000 2789.6600 1527.0800 ;
        RECT 2788.1600 1521.1600 2789.6600 1521.6400 ;
        RECT 2788.1600 1515.7200 2789.6600 1516.2000 ;
        RECT 2788.1600 1510.2800 2789.6600 1510.7600 ;
        RECT 2788.1600 1504.8400 2789.6600 1505.3200 ;
        RECT 2788.1600 1499.4000 2789.6600 1499.8800 ;
        RECT 2788.1600 1493.9600 2789.6600 1494.4400 ;
        RECT 2788.1600 1488.5200 2789.6600 1489.0000 ;
        RECT 2788.1600 1483.0800 2789.6600 1483.5600 ;
        RECT 2788.1600 1477.6400 2789.6600 1478.1200 ;
        RECT 2788.1600 1472.2000 2789.6600 1472.6800 ;
        RECT 2788.1600 1466.7600 2789.6600 1467.2400 ;
        RECT 2788.1600 1461.3200 2789.6600 1461.8000 ;
        RECT 2695.5000 1559.2400 2697.0000 1559.7200 ;
        RECT 2695.5000 1553.8000 2697.0000 1554.2800 ;
        RECT 2695.5000 1548.3600 2697.0000 1548.8400 ;
        RECT 2695.5000 1542.9200 2697.0000 1543.4000 ;
        RECT 2695.5000 1537.4800 2697.0000 1537.9600 ;
        RECT 2695.5000 1532.0400 2697.0000 1532.5200 ;
        RECT 2695.5000 1526.6000 2697.0000 1527.0800 ;
        RECT 2695.5000 1521.1600 2697.0000 1521.6400 ;
        RECT 2695.5000 1515.7200 2697.0000 1516.2000 ;
        RECT 2695.5000 1510.2800 2697.0000 1510.7600 ;
        RECT 2695.5000 1504.8400 2697.0000 1505.3200 ;
        RECT 2695.5000 1499.4000 2697.0000 1499.8800 ;
        RECT 2695.5000 1493.9600 2697.0000 1494.4400 ;
        RECT 2695.5000 1488.5200 2697.0000 1489.0000 ;
        RECT 2695.5000 1483.0800 2697.0000 1483.5600 ;
        RECT 2695.5000 1477.6400 2697.0000 1478.1200 ;
        RECT 2695.5000 1472.2000 2697.0000 1472.6800 ;
        RECT 2695.5000 1466.7600 2697.0000 1467.2400 ;
        RECT 2695.5000 1461.3200 2697.0000 1461.8000 ;
        RECT 2695.5000 1666.2300 2789.6600 1667.7300 ;
        RECT 2695.5000 1454.6300 2789.6600 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 1224.9900 2697.0000 1438.0900 ;
        RECT 2788.1600 1224.9900 2789.6600 1438.0900 ;
      LAYER met3 ;
        RECT 2788.1600 1422.0800 2789.6600 1422.5600 ;
        RECT 2788.1600 1416.6400 2789.6600 1417.1200 ;
        RECT 2788.1600 1427.5200 2789.6600 1428.0000 ;
        RECT 2788.1600 1411.2000 2789.6600 1411.6800 ;
        RECT 2788.1600 1405.7600 2789.6600 1406.2400 ;
        RECT 2788.1600 1394.8800 2789.6600 1395.3600 ;
        RECT 2788.1600 1389.4400 2789.6600 1389.9200 ;
        RECT 2788.1600 1400.3200 2789.6600 1400.8000 ;
        RECT 2788.1600 1384.0000 2789.6600 1384.4800 ;
        RECT 2788.1600 1378.5600 2789.6600 1379.0400 ;
        RECT 2788.1600 1373.1200 2789.6600 1373.6000 ;
        RECT 2788.1600 1367.6800 2789.6600 1368.1600 ;
        RECT 2788.1600 1362.2400 2789.6600 1362.7200 ;
        RECT 2788.1600 1356.8000 2789.6600 1357.2800 ;
        RECT 2788.1600 1351.3600 2789.6600 1351.8400 ;
        RECT 2788.1600 1345.9200 2789.6600 1346.4000 ;
        RECT 2788.1600 1340.4800 2789.6600 1340.9600 ;
        RECT 2788.1600 1335.0400 2789.6600 1335.5200 ;
        RECT 2695.5000 1422.0800 2697.0000 1422.5600 ;
        RECT 2695.5000 1416.6400 2697.0000 1417.1200 ;
        RECT 2695.5000 1427.5200 2697.0000 1428.0000 ;
        RECT 2695.5000 1411.2000 2697.0000 1411.6800 ;
        RECT 2695.5000 1405.7600 2697.0000 1406.2400 ;
        RECT 2695.5000 1394.8800 2697.0000 1395.3600 ;
        RECT 2695.5000 1389.4400 2697.0000 1389.9200 ;
        RECT 2695.5000 1400.3200 2697.0000 1400.8000 ;
        RECT 2695.5000 1384.0000 2697.0000 1384.4800 ;
        RECT 2695.5000 1378.5600 2697.0000 1379.0400 ;
        RECT 2695.5000 1373.1200 2697.0000 1373.6000 ;
        RECT 2695.5000 1367.6800 2697.0000 1368.1600 ;
        RECT 2695.5000 1362.2400 2697.0000 1362.7200 ;
        RECT 2695.5000 1356.8000 2697.0000 1357.2800 ;
        RECT 2695.5000 1351.3600 2697.0000 1351.8400 ;
        RECT 2695.5000 1345.9200 2697.0000 1346.4000 ;
        RECT 2695.5000 1340.4800 2697.0000 1340.9600 ;
        RECT 2695.5000 1335.0400 2697.0000 1335.5200 ;
        RECT 2788.1600 1329.6000 2789.6600 1330.0800 ;
        RECT 2788.1600 1324.1600 2789.6600 1324.6400 ;
        RECT 2788.1600 1318.7200 2789.6600 1319.2000 ;
        RECT 2788.1600 1313.2800 2789.6600 1313.7600 ;
        RECT 2788.1600 1307.8400 2789.6600 1308.3200 ;
        RECT 2788.1600 1302.4000 2789.6600 1302.8800 ;
        RECT 2788.1600 1296.9600 2789.6600 1297.4400 ;
        RECT 2788.1600 1291.5200 2789.6600 1292.0000 ;
        RECT 2788.1600 1286.0800 2789.6600 1286.5600 ;
        RECT 2788.1600 1280.6400 2789.6600 1281.1200 ;
        RECT 2788.1600 1275.2000 2789.6600 1275.6800 ;
        RECT 2788.1600 1269.7600 2789.6600 1270.2400 ;
        RECT 2788.1600 1264.3200 2789.6600 1264.8000 ;
        RECT 2788.1600 1258.8800 2789.6600 1259.3600 ;
        RECT 2788.1600 1253.4400 2789.6600 1253.9200 ;
        RECT 2788.1600 1248.0000 2789.6600 1248.4800 ;
        RECT 2788.1600 1242.5600 2789.6600 1243.0400 ;
        RECT 2788.1600 1237.1200 2789.6600 1237.6000 ;
        RECT 2788.1600 1231.6800 2789.6600 1232.1600 ;
        RECT 2695.5000 1329.6000 2697.0000 1330.0800 ;
        RECT 2695.5000 1324.1600 2697.0000 1324.6400 ;
        RECT 2695.5000 1318.7200 2697.0000 1319.2000 ;
        RECT 2695.5000 1313.2800 2697.0000 1313.7600 ;
        RECT 2695.5000 1307.8400 2697.0000 1308.3200 ;
        RECT 2695.5000 1302.4000 2697.0000 1302.8800 ;
        RECT 2695.5000 1296.9600 2697.0000 1297.4400 ;
        RECT 2695.5000 1291.5200 2697.0000 1292.0000 ;
        RECT 2695.5000 1286.0800 2697.0000 1286.5600 ;
        RECT 2695.5000 1280.6400 2697.0000 1281.1200 ;
        RECT 2695.5000 1275.2000 2697.0000 1275.6800 ;
        RECT 2695.5000 1269.7600 2697.0000 1270.2400 ;
        RECT 2695.5000 1264.3200 2697.0000 1264.8000 ;
        RECT 2695.5000 1258.8800 2697.0000 1259.3600 ;
        RECT 2695.5000 1253.4400 2697.0000 1253.9200 ;
        RECT 2695.5000 1248.0000 2697.0000 1248.4800 ;
        RECT 2695.5000 1242.5600 2697.0000 1243.0400 ;
        RECT 2695.5000 1237.1200 2697.0000 1237.6000 ;
        RECT 2695.5000 1231.6800 2697.0000 1232.1600 ;
        RECT 2695.5000 1436.5900 2789.6600 1438.0900 ;
        RECT 2695.5000 1224.9900 2789.6600 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 995.3500 2697.0000 1208.4500 ;
        RECT 2788.1600 995.3500 2789.6600 1208.4500 ;
      LAYER met3 ;
        RECT 2788.1600 1192.4400 2789.6600 1192.9200 ;
        RECT 2788.1600 1187.0000 2789.6600 1187.4800 ;
        RECT 2788.1600 1197.8800 2789.6600 1198.3600 ;
        RECT 2788.1600 1181.5600 2789.6600 1182.0400 ;
        RECT 2788.1600 1176.1200 2789.6600 1176.6000 ;
        RECT 2788.1600 1165.2400 2789.6600 1165.7200 ;
        RECT 2788.1600 1159.8000 2789.6600 1160.2800 ;
        RECT 2788.1600 1170.6800 2789.6600 1171.1600 ;
        RECT 2788.1600 1154.3600 2789.6600 1154.8400 ;
        RECT 2788.1600 1148.9200 2789.6600 1149.4000 ;
        RECT 2788.1600 1143.4800 2789.6600 1143.9600 ;
        RECT 2788.1600 1138.0400 2789.6600 1138.5200 ;
        RECT 2788.1600 1132.6000 2789.6600 1133.0800 ;
        RECT 2788.1600 1127.1600 2789.6600 1127.6400 ;
        RECT 2788.1600 1121.7200 2789.6600 1122.2000 ;
        RECT 2788.1600 1116.2800 2789.6600 1116.7600 ;
        RECT 2788.1600 1110.8400 2789.6600 1111.3200 ;
        RECT 2788.1600 1105.4000 2789.6600 1105.8800 ;
        RECT 2695.5000 1192.4400 2697.0000 1192.9200 ;
        RECT 2695.5000 1187.0000 2697.0000 1187.4800 ;
        RECT 2695.5000 1197.8800 2697.0000 1198.3600 ;
        RECT 2695.5000 1181.5600 2697.0000 1182.0400 ;
        RECT 2695.5000 1176.1200 2697.0000 1176.6000 ;
        RECT 2695.5000 1165.2400 2697.0000 1165.7200 ;
        RECT 2695.5000 1159.8000 2697.0000 1160.2800 ;
        RECT 2695.5000 1170.6800 2697.0000 1171.1600 ;
        RECT 2695.5000 1154.3600 2697.0000 1154.8400 ;
        RECT 2695.5000 1148.9200 2697.0000 1149.4000 ;
        RECT 2695.5000 1143.4800 2697.0000 1143.9600 ;
        RECT 2695.5000 1138.0400 2697.0000 1138.5200 ;
        RECT 2695.5000 1132.6000 2697.0000 1133.0800 ;
        RECT 2695.5000 1127.1600 2697.0000 1127.6400 ;
        RECT 2695.5000 1121.7200 2697.0000 1122.2000 ;
        RECT 2695.5000 1116.2800 2697.0000 1116.7600 ;
        RECT 2695.5000 1110.8400 2697.0000 1111.3200 ;
        RECT 2695.5000 1105.4000 2697.0000 1105.8800 ;
        RECT 2788.1600 1099.9600 2789.6600 1100.4400 ;
        RECT 2788.1600 1094.5200 2789.6600 1095.0000 ;
        RECT 2788.1600 1089.0800 2789.6600 1089.5600 ;
        RECT 2788.1600 1083.6400 2789.6600 1084.1200 ;
        RECT 2788.1600 1078.2000 2789.6600 1078.6800 ;
        RECT 2788.1600 1072.7600 2789.6600 1073.2400 ;
        RECT 2788.1600 1067.3200 2789.6600 1067.8000 ;
        RECT 2788.1600 1061.8800 2789.6600 1062.3600 ;
        RECT 2788.1600 1056.4400 2789.6600 1056.9200 ;
        RECT 2788.1600 1051.0000 2789.6600 1051.4800 ;
        RECT 2788.1600 1045.5600 2789.6600 1046.0400 ;
        RECT 2788.1600 1040.1200 2789.6600 1040.6000 ;
        RECT 2788.1600 1034.6800 2789.6600 1035.1600 ;
        RECT 2788.1600 1029.2400 2789.6600 1029.7200 ;
        RECT 2788.1600 1023.8000 2789.6600 1024.2800 ;
        RECT 2788.1600 1018.3600 2789.6600 1018.8400 ;
        RECT 2788.1600 1012.9200 2789.6600 1013.4000 ;
        RECT 2788.1600 1007.4800 2789.6600 1007.9600 ;
        RECT 2788.1600 1002.0400 2789.6600 1002.5200 ;
        RECT 2695.5000 1099.9600 2697.0000 1100.4400 ;
        RECT 2695.5000 1094.5200 2697.0000 1095.0000 ;
        RECT 2695.5000 1089.0800 2697.0000 1089.5600 ;
        RECT 2695.5000 1083.6400 2697.0000 1084.1200 ;
        RECT 2695.5000 1078.2000 2697.0000 1078.6800 ;
        RECT 2695.5000 1072.7600 2697.0000 1073.2400 ;
        RECT 2695.5000 1067.3200 2697.0000 1067.8000 ;
        RECT 2695.5000 1061.8800 2697.0000 1062.3600 ;
        RECT 2695.5000 1056.4400 2697.0000 1056.9200 ;
        RECT 2695.5000 1051.0000 2697.0000 1051.4800 ;
        RECT 2695.5000 1045.5600 2697.0000 1046.0400 ;
        RECT 2695.5000 1040.1200 2697.0000 1040.6000 ;
        RECT 2695.5000 1034.6800 2697.0000 1035.1600 ;
        RECT 2695.5000 1029.2400 2697.0000 1029.7200 ;
        RECT 2695.5000 1023.8000 2697.0000 1024.2800 ;
        RECT 2695.5000 1018.3600 2697.0000 1018.8400 ;
        RECT 2695.5000 1012.9200 2697.0000 1013.4000 ;
        RECT 2695.5000 1007.4800 2697.0000 1007.9600 ;
        RECT 2695.5000 1002.0400 2697.0000 1002.5200 ;
        RECT 2695.5000 1206.9500 2789.6600 1208.4500 ;
        RECT 2695.5000 995.3500 2789.6600 996.8500 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'RAM_IO'
    PORT
      LAYER met4 ;
        RECT 2695.5000 765.7100 2697.0000 978.8100 ;
        RECT 2788.1600 765.7100 2789.6600 978.8100 ;
      LAYER met3 ;
        RECT 2788.1600 962.8000 2789.6600 963.2800 ;
        RECT 2788.1600 957.3600 2789.6600 957.8400 ;
        RECT 2788.1600 968.2400 2789.6600 968.7200 ;
        RECT 2788.1600 951.9200 2789.6600 952.4000 ;
        RECT 2788.1600 946.4800 2789.6600 946.9600 ;
        RECT 2788.1600 935.6000 2789.6600 936.0800 ;
        RECT 2788.1600 930.1600 2789.6600 930.6400 ;
        RECT 2788.1600 941.0400 2789.6600 941.5200 ;
        RECT 2788.1600 924.7200 2789.6600 925.2000 ;
        RECT 2788.1600 919.2800 2789.6600 919.7600 ;
        RECT 2788.1600 913.8400 2789.6600 914.3200 ;
        RECT 2788.1600 908.4000 2789.6600 908.8800 ;
        RECT 2788.1600 902.9600 2789.6600 903.4400 ;
        RECT 2788.1600 897.5200 2789.6600 898.0000 ;
        RECT 2788.1600 892.0800 2789.6600 892.5600 ;
        RECT 2788.1600 886.6400 2789.6600 887.1200 ;
        RECT 2788.1600 881.2000 2789.6600 881.6800 ;
        RECT 2788.1600 875.7600 2789.6600 876.2400 ;
        RECT 2695.5000 962.8000 2697.0000 963.2800 ;
        RECT 2695.5000 957.3600 2697.0000 957.8400 ;
        RECT 2695.5000 968.2400 2697.0000 968.7200 ;
        RECT 2695.5000 951.9200 2697.0000 952.4000 ;
        RECT 2695.5000 946.4800 2697.0000 946.9600 ;
        RECT 2695.5000 935.6000 2697.0000 936.0800 ;
        RECT 2695.5000 930.1600 2697.0000 930.6400 ;
        RECT 2695.5000 941.0400 2697.0000 941.5200 ;
        RECT 2695.5000 924.7200 2697.0000 925.2000 ;
        RECT 2695.5000 919.2800 2697.0000 919.7600 ;
        RECT 2695.5000 913.8400 2697.0000 914.3200 ;
        RECT 2695.5000 908.4000 2697.0000 908.8800 ;
        RECT 2695.5000 902.9600 2697.0000 903.4400 ;
        RECT 2695.5000 897.5200 2697.0000 898.0000 ;
        RECT 2695.5000 892.0800 2697.0000 892.5600 ;
        RECT 2695.5000 886.6400 2697.0000 887.1200 ;
        RECT 2695.5000 881.2000 2697.0000 881.6800 ;
        RECT 2695.5000 875.7600 2697.0000 876.2400 ;
        RECT 2788.1600 870.3200 2789.6600 870.8000 ;
        RECT 2788.1600 864.8800 2789.6600 865.3600 ;
        RECT 2788.1600 859.4400 2789.6600 859.9200 ;
        RECT 2788.1600 854.0000 2789.6600 854.4800 ;
        RECT 2788.1600 848.5600 2789.6600 849.0400 ;
        RECT 2788.1600 843.1200 2789.6600 843.6000 ;
        RECT 2788.1600 837.6800 2789.6600 838.1600 ;
        RECT 2788.1600 832.2400 2789.6600 832.7200 ;
        RECT 2788.1600 826.8000 2789.6600 827.2800 ;
        RECT 2788.1600 821.3600 2789.6600 821.8400 ;
        RECT 2788.1600 815.9200 2789.6600 816.4000 ;
        RECT 2788.1600 810.4800 2789.6600 810.9600 ;
        RECT 2788.1600 805.0400 2789.6600 805.5200 ;
        RECT 2788.1600 799.6000 2789.6600 800.0800 ;
        RECT 2788.1600 794.1600 2789.6600 794.6400 ;
        RECT 2788.1600 788.7200 2789.6600 789.2000 ;
        RECT 2788.1600 783.2800 2789.6600 783.7600 ;
        RECT 2788.1600 777.8400 2789.6600 778.3200 ;
        RECT 2788.1600 772.4000 2789.6600 772.8800 ;
        RECT 2695.5000 870.3200 2697.0000 870.8000 ;
        RECT 2695.5000 864.8800 2697.0000 865.3600 ;
        RECT 2695.5000 859.4400 2697.0000 859.9200 ;
        RECT 2695.5000 854.0000 2697.0000 854.4800 ;
        RECT 2695.5000 848.5600 2697.0000 849.0400 ;
        RECT 2695.5000 843.1200 2697.0000 843.6000 ;
        RECT 2695.5000 837.6800 2697.0000 838.1600 ;
        RECT 2695.5000 832.2400 2697.0000 832.7200 ;
        RECT 2695.5000 826.8000 2697.0000 827.2800 ;
        RECT 2695.5000 821.3600 2697.0000 821.8400 ;
        RECT 2695.5000 815.9200 2697.0000 816.4000 ;
        RECT 2695.5000 810.4800 2697.0000 810.9600 ;
        RECT 2695.5000 805.0400 2697.0000 805.5200 ;
        RECT 2695.5000 799.6000 2697.0000 800.0800 ;
        RECT 2695.5000 794.1600 2697.0000 794.6400 ;
        RECT 2695.5000 788.7200 2697.0000 789.2000 ;
        RECT 2695.5000 783.2800 2697.0000 783.7600 ;
        RECT 2695.5000 777.8400 2697.0000 778.3200 ;
        RECT 2695.5000 772.4000 2697.0000 772.8800 ;
        RECT 2695.5000 977.3100 2789.6600 978.8100 ;
        RECT 2695.5000 765.7100 2789.6600 767.2100 ;
    END
# end of P/G pin shape extracted from block 'RAM_IO'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 242.6800 2830.6100 244.6800 2857.5400 ;
        RECT 445.7800 2830.6100 447.7800 2857.5400 ;
      LAYER met3 ;
        RECT 445.7800 2847.3200 447.7800 2847.8000 ;
        RECT 242.6800 2847.3200 244.6800 2847.8000 ;
        RECT 445.7800 2841.8800 447.7800 2842.3600 ;
        RECT 445.7800 2836.4400 447.7800 2836.9200 ;
        RECT 242.6800 2841.8800 244.6800 2842.3600 ;
        RECT 242.6800 2836.4400 244.6800 2836.9200 ;
        RECT 242.6800 2855.5400 447.7800 2857.5400 ;
        RECT 242.6800 2830.6100 447.7800 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 534.5700 435.0400 750.6700 ;
        RECT 388.4400 534.5700 390.0400 750.6700 ;
        RECT 343.4400 534.5700 345.0400 750.6700 ;
        RECT 298.4400 534.5700 300.0400 750.6700 ;
        RECT 253.4400 534.5700 255.0400 750.6700 ;
        RECT 445.7800 534.5700 448.7800 750.6700 ;
        RECT 241.6800 534.5700 244.6800 750.6700 ;
      LAYER met3 ;
        RECT 445.7800 727.7200 448.7800 728.2000 ;
        RECT 445.7800 733.1600 448.7800 733.6400 ;
        RECT 433.4400 727.7200 435.0400 728.2000 ;
        RECT 433.4400 733.1600 435.0400 733.6400 ;
        RECT 445.7800 738.6000 448.7800 739.0800 ;
        RECT 433.4400 738.6000 435.0400 739.0800 ;
        RECT 445.7800 716.8400 448.7800 717.3200 ;
        RECT 445.7800 722.2800 448.7800 722.7600 ;
        RECT 433.4400 716.8400 435.0400 717.3200 ;
        RECT 433.4400 722.2800 435.0400 722.7600 ;
        RECT 445.7800 700.5200 448.7800 701.0000 ;
        RECT 445.7800 705.9600 448.7800 706.4400 ;
        RECT 433.4400 700.5200 435.0400 701.0000 ;
        RECT 433.4400 705.9600 435.0400 706.4400 ;
        RECT 445.7800 711.4000 448.7800 711.8800 ;
        RECT 433.4400 711.4000 435.0400 711.8800 ;
        RECT 388.4400 727.7200 390.0400 728.2000 ;
        RECT 388.4400 733.1600 390.0400 733.6400 ;
        RECT 388.4400 738.6000 390.0400 739.0800 ;
        RECT 388.4400 716.8400 390.0400 717.3200 ;
        RECT 388.4400 722.2800 390.0400 722.7600 ;
        RECT 388.4400 700.5200 390.0400 701.0000 ;
        RECT 388.4400 705.9600 390.0400 706.4400 ;
        RECT 388.4400 711.4000 390.0400 711.8800 ;
        RECT 445.7800 684.2000 448.7800 684.6800 ;
        RECT 445.7800 689.6400 448.7800 690.1200 ;
        RECT 445.7800 695.0800 448.7800 695.5600 ;
        RECT 433.4400 684.2000 435.0400 684.6800 ;
        RECT 433.4400 689.6400 435.0400 690.1200 ;
        RECT 433.4400 695.0800 435.0400 695.5600 ;
        RECT 445.7800 673.3200 448.7800 673.8000 ;
        RECT 445.7800 678.7600 448.7800 679.2400 ;
        RECT 433.4400 673.3200 435.0400 673.8000 ;
        RECT 433.4400 678.7600 435.0400 679.2400 ;
        RECT 445.7800 657.0000 448.7800 657.4800 ;
        RECT 445.7800 662.4400 448.7800 662.9200 ;
        RECT 445.7800 667.8800 448.7800 668.3600 ;
        RECT 433.4400 657.0000 435.0400 657.4800 ;
        RECT 433.4400 662.4400 435.0400 662.9200 ;
        RECT 433.4400 667.8800 435.0400 668.3600 ;
        RECT 445.7800 646.1200 448.7800 646.6000 ;
        RECT 445.7800 651.5600 448.7800 652.0400 ;
        RECT 433.4400 646.1200 435.0400 646.6000 ;
        RECT 433.4400 651.5600 435.0400 652.0400 ;
        RECT 388.4400 684.2000 390.0400 684.6800 ;
        RECT 388.4400 689.6400 390.0400 690.1200 ;
        RECT 388.4400 695.0800 390.0400 695.5600 ;
        RECT 388.4400 673.3200 390.0400 673.8000 ;
        RECT 388.4400 678.7600 390.0400 679.2400 ;
        RECT 388.4400 657.0000 390.0400 657.4800 ;
        RECT 388.4400 662.4400 390.0400 662.9200 ;
        RECT 388.4400 667.8800 390.0400 668.3600 ;
        RECT 388.4400 646.1200 390.0400 646.6000 ;
        RECT 388.4400 651.5600 390.0400 652.0400 ;
        RECT 343.4400 727.7200 345.0400 728.2000 ;
        RECT 343.4400 733.1600 345.0400 733.6400 ;
        RECT 343.4400 738.6000 345.0400 739.0800 ;
        RECT 298.4400 727.7200 300.0400 728.2000 ;
        RECT 298.4400 733.1600 300.0400 733.6400 ;
        RECT 298.4400 738.6000 300.0400 739.0800 ;
        RECT 343.4400 716.8400 345.0400 717.3200 ;
        RECT 343.4400 722.2800 345.0400 722.7600 ;
        RECT 343.4400 700.5200 345.0400 701.0000 ;
        RECT 343.4400 705.9600 345.0400 706.4400 ;
        RECT 343.4400 711.4000 345.0400 711.8800 ;
        RECT 298.4400 716.8400 300.0400 717.3200 ;
        RECT 298.4400 722.2800 300.0400 722.7600 ;
        RECT 298.4400 700.5200 300.0400 701.0000 ;
        RECT 298.4400 705.9600 300.0400 706.4400 ;
        RECT 298.4400 711.4000 300.0400 711.8800 ;
        RECT 253.4400 727.7200 255.0400 728.2000 ;
        RECT 253.4400 733.1600 255.0400 733.6400 ;
        RECT 241.6800 733.1600 244.6800 733.6400 ;
        RECT 241.6800 727.7200 244.6800 728.2000 ;
        RECT 241.6800 738.6000 244.6800 739.0800 ;
        RECT 253.4400 738.6000 255.0400 739.0800 ;
        RECT 253.4400 716.8400 255.0400 717.3200 ;
        RECT 253.4400 722.2800 255.0400 722.7600 ;
        RECT 241.6800 722.2800 244.6800 722.7600 ;
        RECT 241.6800 716.8400 244.6800 717.3200 ;
        RECT 253.4400 700.5200 255.0400 701.0000 ;
        RECT 253.4400 705.9600 255.0400 706.4400 ;
        RECT 241.6800 705.9600 244.6800 706.4400 ;
        RECT 241.6800 700.5200 244.6800 701.0000 ;
        RECT 241.6800 711.4000 244.6800 711.8800 ;
        RECT 253.4400 711.4000 255.0400 711.8800 ;
        RECT 343.4400 684.2000 345.0400 684.6800 ;
        RECT 343.4400 689.6400 345.0400 690.1200 ;
        RECT 343.4400 695.0800 345.0400 695.5600 ;
        RECT 343.4400 673.3200 345.0400 673.8000 ;
        RECT 343.4400 678.7600 345.0400 679.2400 ;
        RECT 298.4400 684.2000 300.0400 684.6800 ;
        RECT 298.4400 689.6400 300.0400 690.1200 ;
        RECT 298.4400 695.0800 300.0400 695.5600 ;
        RECT 298.4400 673.3200 300.0400 673.8000 ;
        RECT 298.4400 678.7600 300.0400 679.2400 ;
        RECT 343.4400 657.0000 345.0400 657.4800 ;
        RECT 343.4400 662.4400 345.0400 662.9200 ;
        RECT 343.4400 667.8800 345.0400 668.3600 ;
        RECT 343.4400 646.1200 345.0400 646.6000 ;
        RECT 343.4400 651.5600 345.0400 652.0400 ;
        RECT 298.4400 657.0000 300.0400 657.4800 ;
        RECT 298.4400 662.4400 300.0400 662.9200 ;
        RECT 298.4400 667.8800 300.0400 668.3600 ;
        RECT 298.4400 646.1200 300.0400 646.6000 ;
        RECT 298.4400 651.5600 300.0400 652.0400 ;
        RECT 253.4400 684.2000 255.0400 684.6800 ;
        RECT 253.4400 689.6400 255.0400 690.1200 ;
        RECT 253.4400 695.0800 255.0400 695.5600 ;
        RECT 241.6800 684.2000 244.6800 684.6800 ;
        RECT 241.6800 689.6400 244.6800 690.1200 ;
        RECT 241.6800 695.0800 244.6800 695.5600 ;
        RECT 253.4400 673.3200 255.0400 673.8000 ;
        RECT 253.4400 678.7600 255.0400 679.2400 ;
        RECT 241.6800 673.3200 244.6800 673.8000 ;
        RECT 241.6800 678.7600 244.6800 679.2400 ;
        RECT 253.4400 657.0000 255.0400 657.4800 ;
        RECT 253.4400 662.4400 255.0400 662.9200 ;
        RECT 253.4400 667.8800 255.0400 668.3600 ;
        RECT 241.6800 657.0000 244.6800 657.4800 ;
        RECT 241.6800 662.4400 244.6800 662.9200 ;
        RECT 241.6800 667.8800 244.6800 668.3600 ;
        RECT 253.4400 646.1200 255.0400 646.6000 ;
        RECT 253.4400 651.5600 255.0400 652.0400 ;
        RECT 241.6800 646.1200 244.6800 646.6000 ;
        RECT 241.6800 651.5600 244.6800 652.0400 ;
        RECT 445.7800 629.8000 448.7800 630.2800 ;
        RECT 445.7800 635.2400 448.7800 635.7200 ;
        RECT 445.7800 640.6800 448.7800 641.1600 ;
        RECT 433.4400 629.8000 435.0400 630.2800 ;
        RECT 433.4400 635.2400 435.0400 635.7200 ;
        RECT 433.4400 640.6800 435.0400 641.1600 ;
        RECT 445.7800 618.9200 448.7800 619.4000 ;
        RECT 445.7800 624.3600 448.7800 624.8400 ;
        RECT 433.4400 618.9200 435.0400 619.4000 ;
        RECT 433.4400 624.3600 435.0400 624.8400 ;
        RECT 445.7800 602.6000 448.7800 603.0800 ;
        RECT 445.7800 608.0400 448.7800 608.5200 ;
        RECT 445.7800 613.4800 448.7800 613.9600 ;
        RECT 433.4400 602.6000 435.0400 603.0800 ;
        RECT 433.4400 608.0400 435.0400 608.5200 ;
        RECT 433.4400 613.4800 435.0400 613.9600 ;
        RECT 445.7800 591.7200 448.7800 592.2000 ;
        RECT 445.7800 597.1600 448.7800 597.6400 ;
        RECT 433.4400 591.7200 435.0400 592.2000 ;
        RECT 433.4400 597.1600 435.0400 597.6400 ;
        RECT 388.4400 629.8000 390.0400 630.2800 ;
        RECT 388.4400 635.2400 390.0400 635.7200 ;
        RECT 388.4400 640.6800 390.0400 641.1600 ;
        RECT 388.4400 618.9200 390.0400 619.4000 ;
        RECT 388.4400 624.3600 390.0400 624.8400 ;
        RECT 388.4400 602.6000 390.0400 603.0800 ;
        RECT 388.4400 608.0400 390.0400 608.5200 ;
        RECT 388.4400 613.4800 390.0400 613.9600 ;
        RECT 388.4400 591.7200 390.0400 592.2000 ;
        RECT 388.4400 597.1600 390.0400 597.6400 ;
        RECT 445.7800 575.4000 448.7800 575.8800 ;
        RECT 445.7800 580.8400 448.7800 581.3200 ;
        RECT 445.7800 586.2800 448.7800 586.7600 ;
        RECT 433.4400 575.4000 435.0400 575.8800 ;
        RECT 433.4400 580.8400 435.0400 581.3200 ;
        RECT 433.4400 586.2800 435.0400 586.7600 ;
        RECT 445.7800 564.5200 448.7800 565.0000 ;
        RECT 445.7800 569.9600 448.7800 570.4400 ;
        RECT 433.4400 564.5200 435.0400 565.0000 ;
        RECT 433.4400 569.9600 435.0400 570.4400 ;
        RECT 445.7800 548.2000 448.7800 548.6800 ;
        RECT 445.7800 553.6400 448.7800 554.1200 ;
        RECT 445.7800 559.0800 448.7800 559.5600 ;
        RECT 433.4400 548.2000 435.0400 548.6800 ;
        RECT 433.4400 553.6400 435.0400 554.1200 ;
        RECT 433.4400 559.0800 435.0400 559.5600 ;
        RECT 445.7800 542.7600 448.7800 543.2400 ;
        RECT 433.4400 542.7600 435.0400 543.2400 ;
        RECT 388.4400 575.4000 390.0400 575.8800 ;
        RECT 388.4400 580.8400 390.0400 581.3200 ;
        RECT 388.4400 586.2800 390.0400 586.7600 ;
        RECT 388.4400 564.5200 390.0400 565.0000 ;
        RECT 388.4400 569.9600 390.0400 570.4400 ;
        RECT 388.4400 548.2000 390.0400 548.6800 ;
        RECT 388.4400 553.6400 390.0400 554.1200 ;
        RECT 388.4400 559.0800 390.0400 559.5600 ;
        RECT 388.4400 542.7600 390.0400 543.2400 ;
        RECT 343.4400 629.8000 345.0400 630.2800 ;
        RECT 343.4400 635.2400 345.0400 635.7200 ;
        RECT 343.4400 640.6800 345.0400 641.1600 ;
        RECT 343.4400 618.9200 345.0400 619.4000 ;
        RECT 343.4400 624.3600 345.0400 624.8400 ;
        RECT 298.4400 629.8000 300.0400 630.2800 ;
        RECT 298.4400 635.2400 300.0400 635.7200 ;
        RECT 298.4400 640.6800 300.0400 641.1600 ;
        RECT 298.4400 618.9200 300.0400 619.4000 ;
        RECT 298.4400 624.3600 300.0400 624.8400 ;
        RECT 343.4400 602.6000 345.0400 603.0800 ;
        RECT 343.4400 608.0400 345.0400 608.5200 ;
        RECT 343.4400 613.4800 345.0400 613.9600 ;
        RECT 343.4400 591.7200 345.0400 592.2000 ;
        RECT 343.4400 597.1600 345.0400 597.6400 ;
        RECT 298.4400 602.6000 300.0400 603.0800 ;
        RECT 298.4400 608.0400 300.0400 608.5200 ;
        RECT 298.4400 613.4800 300.0400 613.9600 ;
        RECT 298.4400 591.7200 300.0400 592.2000 ;
        RECT 298.4400 597.1600 300.0400 597.6400 ;
        RECT 253.4400 629.8000 255.0400 630.2800 ;
        RECT 253.4400 635.2400 255.0400 635.7200 ;
        RECT 253.4400 640.6800 255.0400 641.1600 ;
        RECT 241.6800 629.8000 244.6800 630.2800 ;
        RECT 241.6800 635.2400 244.6800 635.7200 ;
        RECT 241.6800 640.6800 244.6800 641.1600 ;
        RECT 253.4400 618.9200 255.0400 619.4000 ;
        RECT 253.4400 624.3600 255.0400 624.8400 ;
        RECT 241.6800 618.9200 244.6800 619.4000 ;
        RECT 241.6800 624.3600 244.6800 624.8400 ;
        RECT 253.4400 602.6000 255.0400 603.0800 ;
        RECT 253.4400 608.0400 255.0400 608.5200 ;
        RECT 253.4400 613.4800 255.0400 613.9600 ;
        RECT 241.6800 602.6000 244.6800 603.0800 ;
        RECT 241.6800 608.0400 244.6800 608.5200 ;
        RECT 241.6800 613.4800 244.6800 613.9600 ;
        RECT 253.4400 591.7200 255.0400 592.2000 ;
        RECT 253.4400 597.1600 255.0400 597.6400 ;
        RECT 241.6800 591.7200 244.6800 592.2000 ;
        RECT 241.6800 597.1600 244.6800 597.6400 ;
        RECT 343.4400 575.4000 345.0400 575.8800 ;
        RECT 343.4400 580.8400 345.0400 581.3200 ;
        RECT 343.4400 586.2800 345.0400 586.7600 ;
        RECT 343.4400 564.5200 345.0400 565.0000 ;
        RECT 343.4400 569.9600 345.0400 570.4400 ;
        RECT 298.4400 575.4000 300.0400 575.8800 ;
        RECT 298.4400 580.8400 300.0400 581.3200 ;
        RECT 298.4400 586.2800 300.0400 586.7600 ;
        RECT 298.4400 564.5200 300.0400 565.0000 ;
        RECT 298.4400 569.9600 300.0400 570.4400 ;
        RECT 343.4400 548.2000 345.0400 548.6800 ;
        RECT 343.4400 553.6400 345.0400 554.1200 ;
        RECT 343.4400 559.0800 345.0400 559.5600 ;
        RECT 343.4400 542.7600 345.0400 543.2400 ;
        RECT 298.4400 548.2000 300.0400 548.6800 ;
        RECT 298.4400 553.6400 300.0400 554.1200 ;
        RECT 298.4400 559.0800 300.0400 559.5600 ;
        RECT 298.4400 542.7600 300.0400 543.2400 ;
        RECT 253.4400 575.4000 255.0400 575.8800 ;
        RECT 253.4400 580.8400 255.0400 581.3200 ;
        RECT 253.4400 586.2800 255.0400 586.7600 ;
        RECT 241.6800 575.4000 244.6800 575.8800 ;
        RECT 241.6800 580.8400 244.6800 581.3200 ;
        RECT 241.6800 586.2800 244.6800 586.7600 ;
        RECT 253.4400 564.5200 255.0400 565.0000 ;
        RECT 253.4400 569.9600 255.0400 570.4400 ;
        RECT 241.6800 564.5200 244.6800 565.0000 ;
        RECT 241.6800 569.9600 244.6800 570.4400 ;
        RECT 253.4400 548.2000 255.0400 548.6800 ;
        RECT 253.4400 553.6400 255.0400 554.1200 ;
        RECT 253.4400 559.0800 255.0400 559.5600 ;
        RECT 241.6800 548.2000 244.6800 548.6800 ;
        RECT 241.6800 553.6400 244.6800 554.1200 ;
        RECT 241.6800 559.0800 244.6800 559.5600 ;
        RECT 241.6800 542.7600 244.6800 543.2400 ;
        RECT 253.4400 542.7600 255.0400 543.2400 ;
        RECT 241.6800 747.6700 448.7800 750.6700 ;
        RECT 241.6800 534.5700 448.7800 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 304.9300 435.0400 521.0300 ;
        RECT 388.4400 304.9300 390.0400 521.0300 ;
        RECT 343.4400 304.9300 345.0400 521.0300 ;
        RECT 298.4400 304.9300 300.0400 521.0300 ;
        RECT 253.4400 304.9300 255.0400 521.0300 ;
        RECT 445.7800 304.9300 448.7800 521.0300 ;
        RECT 241.6800 304.9300 244.6800 521.0300 ;
      LAYER met3 ;
        RECT 445.7800 498.0800 448.7800 498.5600 ;
        RECT 445.7800 503.5200 448.7800 504.0000 ;
        RECT 433.4400 498.0800 435.0400 498.5600 ;
        RECT 433.4400 503.5200 435.0400 504.0000 ;
        RECT 445.7800 508.9600 448.7800 509.4400 ;
        RECT 433.4400 508.9600 435.0400 509.4400 ;
        RECT 445.7800 487.2000 448.7800 487.6800 ;
        RECT 445.7800 492.6400 448.7800 493.1200 ;
        RECT 433.4400 487.2000 435.0400 487.6800 ;
        RECT 433.4400 492.6400 435.0400 493.1200 ;
        RECT 445.7800 470.8800 448.7800 471.3600 ;
        RECT 445.7800 476.3200 448.7800 476.8000 ;
        RECT 433.4400 470.8800 435.0400 471.3600 ;
        RECT 433.4400 476.3200 435.0400 476.8000 ;
        RECT 445.7800 481.7600 448.7800 482.2400 ;
        RECT 433.4400 481.7600 435.0400 482.2400 ;
        RECT 388.4400 498.0800 390.0400 498.5600 ;
        RECT 388.4400 503.5200 390.0400 504.0000 ;
        RECT 388.4400 508.9600 390.0400 509.4400 ;
        RECT 388.4400 487.2000 390.0400 487.6800 ;
        RECT 388.4400 492.6400 390.0400 493.1200 ;
        RECT 388.4400 470.8800 390.0400 471.3600 ;
        RECT 388.4400 476.3200 390.0400 476.8000 ;
        RECT 388.4400 481.7600 390.0400 482.2400 ;
        RECT 445.7800 454.5600 448.7800 455.0400 ;
        RECT 445.7800 460.0000 448.7800 460.4800 ;
        RECT 445.7800 465.4400 448.7800 465.9200 ;
        RECT 433.4400 454.5600 435.0400 455.0400 ;
        RECT 433.4400 460.0000 435.0400 460.4800 ;
        RECT 433.4400 465.4400 435.0400 465.9200 ;
        RECT 445.7800 443.6800 448.7800 444.1600 ;
        RECT 445.7800 449.1200 448.7800 449.6000 ;
        RECT 433.4400 443.6800 435.0400 444.1600 ;
        RECT 433.4400 449.1200 435.0400 449.6000 ;
        RECT 445.7800 427.3600 448.7800 427.8400 ;
        RECT 445.7800 432.8000 448.7800 433.2800 ;
        RECT 445.7800 438.2400 448.7800 438.7200 ;
        RECT 433.4400 427.3600 435.0400 427.8400 ;
        RECT 433.4400 432.8000 435.0400 433.2800 ;
        RECT 433.4400 438.2400 435.0400 438.7200 ;
        RECT 445.7800 416.4800 448.7800 416.9600 ;
        RECT 445.7800 421.9200 448.7800 422.4000 ;
        RECT 433.4400 416.4800 435.0400 416.9600 ;
        RECT 433.4400 421.9200 435.0400 422.4000 ;
        RECT 388.4400 454.5600 390.0400 455.0400 ;
        RECT 388.4400 460.0000 390.0400 460.4800 ;
        RECT 388.4400 465.4400 390.0400 465.9200 ;
        RECT 388.4400 443.6800 390.0400 444.1600 ;
        RECT 388.4400 449.1200 390.0400 449.6000 ;
        RECT 388.4400 427.3600 390.0400 427.8400 ;
        RECT 388.4400 432.8000 390.0400 433.2800 ;
        RECT 388.4400 438.2400 390.0400 438.7200 ;
        RECT 388.4400 416.4800 390.0400 416.9600 ;
        RECT 388.4400 421.9200 390.0400 422.4000 ;
        RECT 343.4400 498.0800 345.0400 498.5600 ;
        RECT 343.4400 503.5200 345.0400 504.0000 ;
        RECT 343.4400 508.9600 345.0400 509.4400 ;
        RECT 298.4400 498.0800 300.0400 498.5600 ;
        RECT 298.4400 503.5200 300.0400 504.0000 ;
        RECT 298.4400 508.9600 300.0400 509.4400 ;
        RECT 343.4400 487.2000 345.0400 487.6800 ;
        RECT 343.4400 492.6400 345.0400 493.1200 ;
        RECT 343.4400 470.8800 345.0400 471.3600 ;
        RECT 343.4400 476.3200 345.0400 476.8000 ;
        RECT 343.4400 481.7600 345.0400 482.2400 ;
        RECT 298.4400 487.2000 300.0400 487.6800 ;
        RECT 298.4400 492.6400 300.0400 493.1200 ;
        RECT 298.4400 470.8800 300.0400 471.3600 ;
        RECT 298.4400 476.3200 300.0400 476.8000 ;
        RECT 298.4400 481.7600 300.0400 482.2400 ;
        RECT 253.4400 498.0800 255.0400 498.5600 ;
        RECT 253.4400 503.5200 255.0400 504.0000 ;
        RECT 241.6800 503.5200 244.6800 504.0000 ;
        RECT 241.6800 498.0800 244.6800 498.5600 ;
        RECT 241.6800 508.9600 244.6800 509.4400 ;
        RECT 253.4400 508.9600 255.0400 509.4400 ;
        RECT 253.4400 487.2000 255.0400 487.6800 ;
        RECT 253.4400 492.6400 255.0400 493.1200 ;
        RECT 241.6800 492.6400 244.6800 493.1200 ;
        RECT 241.6800 487.2000 244.6800 487.6800 ;
        RECT 253.4400 470.8800 255.0400 471.3600 ;
        RECT 253.4400 476.3200 255.0400 476.8000 ;
        RECT 241.6800 476.3200 244.6800 476.8000 ;
        RECT 241.6800 470.8800 244.6800 471.3600 ;
        RECT 241.6800 481.7600 244.6800 482.2400 ;
        RECT 253.4400 481.7600 255.0400 482.2400 ;
        RECT 343.4400 454.5600 345.0400 455.0400 ;
        RECT 343.4400 460.0000 345.0400 460.4800 ;
        RECT 343.4400 465.4400 345.0400 465.9200 ;
        RECT 343.4400 443.6800 345.0400 444.1600 ;
        RECT 343.4400 449.1200 345.0400 449.6000 ;
        RECT 298.4400 454.5600 300.0400 455.0400 ;
        RECT 298.4400 460.0000 300.0400 460.4800 ;
        RECT 298.4400 465.4400 300.0400 465.9200 ;
        RECT 298.4400 443.6800 300.0400 444.1600 ;
        RECT 298.4400 449.1200 300.0400 449.6000 ;
        RECT 343.4400 427.3600 345.0400 427.8400 ;
        RECT 343.4400 432.8000 345.0400 433.2800 ;
        RECT 343.4400 438.2400 345.0400 438.7200 ;
        RECT 343.4400 416.4800 345.0400 416.9600 ;
        RECT 343.4400 421.9200 345.0400 422.4000 ;
        RECT 298.4400 427.3600 300.0400 427.8400 ;
        RECT 298.4400 432.8000 300.0400 433.2800 ;
        RECT 298.4400 438.2400 300.0400 438.7200 ;
        RECT 298.4400 416.4800 300.0400 416.9600 ;
        RECT 298.4400 421.9200 300.0400 422.4000 ;
        RECT 253.4400 454.5600 255.0400 455.0400 ;
        RECT 253.4400 460.0000 255.0400 460.4800 ;
        RECT 253.4400 465.4400 255.0400 465.9200 ;
        RECT 241.6800 454.5600 244.6800 455.0400 ;
        RECT 241.6800 460.0000 244.6800 460.4800 ;
        RECT 241.6800 465.4400 244.6800 465.9200 ;
        RECT 253.4400 443.6800 255.0400 444.1600 ;
        RECT 253.4400 449.1200 255.0400 449.6000 ;
        RECT 241.6800 443.6800 244.6800 444.1600 ;
        RECT 241.6800 449.1200 244.6800 449.6000 ;
        RECT 253.4400 427.3600 255.0400 427.8400 ;
        RECT 253.4400 432.8000 255.0400 433.2800 ;
        RECT 253.4400 438.2400 255.0400 438.7200 ;
        RECT 241.6800 427.3600 244.6800 427.8400 ;
        RECT 241.6800 432.8000 244.6800 433.2800 ;
        RECT 241.6800 438.2400 244.6800 438.7200 ;
        RECT 253.4400 416.4800 255.0400 416.9600 ;
        RECT 253.4400 421.9200 255.0400 422.4000 ;
        RECT 241.6800 416.4800 244.6800 416.9600 ;
        RECT 241.6800 421.9200 244.6800 422.4000 ;
        RECT 445.7800 400.1600 448.7800 400.6400 ;
        RECT 445.7800 405.6000 448.7800 406.0800 ;
        RECT 445.7800 411.0400 448.7800 411.5200 ;
        RECT 433.4400 400.1600 435.0400 400.6400 ;
        RECT 433.4400 405.6000 435.0400 406.0800 ;
        RECT 433.4400 411.0400 435.0400 411.5200 ;
        RECT 445.7800 389.2800 448.7800 389.7600 ;
        RECT 445.7800 394.7200 448.7800 395.2000 ;
        RECT 433.4400 389.2800 435.0400 389.7600 ;
        RECT 433.4400 394.7200 435.0400 395.2000 ;
        RECT 445.7800 372.9600 448.7800 373.4400 ;
        RECT 445.7800 378.4000 448.7800 378.8800 ;
        RECT 445.7800 383.8400 448.7800 384.3200 ;
        RECT 433.4400 372.9600 435.0400 373.4400 ;
        RECT 433.4400 378.4000 435.0400 378.8800 ;
        RECT 433.4400 383.8400 435.0400 384.3200 ;
        RECT 445.7800 362.0800 448.7800 362.5600 ;
        RECT 445.7800 367.5200 448.7800 368.0000 ;
        RECT 433.4400 362.0800 435.0400 362.5600 ;
        RECT 433.4400 367.5200 435.0400 368.0000 ;
        RECT 388.4400 400.1600 390.0400 400.6400 ;
        RECT 388.4400 405.6000 390.0400 406.0800 ;
        RECT 388.4400 411.0400 390.0400 411.5200 ;
        RECT 388.4400 389.2800 390.0400 389.7600 ;
        RECT 388.4400 394.7200 390.0400 395.2000 ;
        RECT 388.4400 372.9600 390.0400 373.4400 ;
        RECT 388.4400 378.4000 390.0400 378.8800 ;
        RECT 388.4400 383.8400 390.0400 384.3200 ;
        RECT 388.4400 362.0800 390.0400 362.5600 ;
        RECT 388.4400 367.5200 390.0400 368.0000 ;
        RECT 445.7800 345.7600 448.7800 346.2400 ;
        RECT 445.7800 351.2000 448.7800 351.6800 ;
        RECT 445.7800 356.6400 448.7800 357.1200 ;
        RECT 433.4400 345.7600 435.0400 346.2400 ;
        RECT 433.4400 351.2000 435.0400 351.6800 ;
        RECT 433.4400 356.6400 435.0400 357.1200 ;
        RECT 445.7800 334.8800 448.7800 335.3600 ;
        RECT 445.7800 340.3200 448.7800 340.8000 ;
        RECT 433.4400 334.8800 435.0400 335.3600 ;
        RECT 433.4400 340.3200 435.0400 340.8000 ;
        RECT 445.7800 318.5600 448.7800 319.0400 ;
        RECT 445.7800 324.0000 448.7800 324.4800 ;
        RECT 445.7800 329.4400 448.7800 329.9200 ;
        RECT 433.4400 318.5600 435.0400 319.0400 ;
        RECT 433.4400 324.0000 435.0400 324.4800 ;
        RECT 433.4400 329.4400 435.0400 329.9200 ;
        RECT 445.7800 313.1200 448.7800 313.6000 ;
        RECT 433.4400 313.1200 435.0400 313.6000 ;
        RECT 388.4400 345.7600 390.0400 346.2400 ;
        RECT 388.4400 351.2000 390.0400 351.6800 ;
        RECT 388.4400 356.6400 390.0400 357.1200 ;
        RECT 388.4400 334.8800 390.0400 335.3600 ;
        RECT 388.4400 340.3200 390.0400 340.8000 ;
        RECT 388.4400 318.5600 390.0400 319.0400 ;
        RECT 388.4400 324.0000 390.0400 324.4800 ;
        RECT 388.4400 329.4400 390.0400 329.9200 ;
        RECT 388.4400 313.1200 390.0400 313.6000 ;
        RECT 343.4400 400.1600 345.0400 400.6400 ;
        RECT 343.4400 405.6000 345.0400 406.0800 ;
        RECT 343.4400 411.0400 345.0400 411.5200 ;
        RECT 343.4400 389.2800 345.0400 389.7600 ;
        RECT 343.4400 394.7200 345.0400 395.2000 ;
        RECT 298.4400 400.1600 300.0400 400.6400 ;
        RECT 298.4400 405.6000 300.0400 406.0800 ;
        RECT 298.4400 411.0400 300.0400 411.5200 ;
        RECT 298.4400 389.2800 300.0400 389.7600 ;
        RECT 298.4400 394.7200 300.0400 395.2000 ;
        RECT 343.4400 372.9600 345.0400 373.4400 ;
        RECT 343.4400 378.4000 345.0400 378.8800 ;
        RECT 343.4400 383.8400 345.0400 384.3200 ;
        RECT 343.4400 362.0800 345.0400 362.5600 ;
        RECT 343.4400 367.5200 345.0400 368.0000 ;
        RECT 298.4400 372.9600 300.0400 373.4400 ;
        RECT 298.4400 378.4000 300.0400 378.8800 ;
        RECT 298.4400 383.8400 300.0400 384.3200 ;
        RECT 298.4400 362.0800 300.0400 362.5600 ;
        RECT 298.4400 367.5200 300.0400 368.0000 ;
        RECT 253.4400 400.1600 255.0400 400.6400 ;
        RECT 253.4400 405.6000 255.0400 406.0800 ;
        RECT 253.4400 411.0400 255.0400 411.5200 ;
        RECT 241.6800 400.1600 244.6800 400.6400 ;
        RECT 241.6800 405.6000 244.6800 406.0800 ;
        RECT 241.6800 411.0400 244.6800 411.5200 ;
        RECT 253.4400 389.2800 255.0400 389.7600 ;
        RECT 253.4400 394.7200 255.0400 395.2000 ;
        RECT 241.6800 389.2800 244.6800 389.7600 ;
        RECT 241.6800 394.7200 244.6800 395.2000 ;
        RECT 253.4400 372.9600 255.0400 373.4400 ;
        RECT 253.4400 378.4000 255.0400 378.8800 ;
        RECT 253.4400 383.8400 255.0400 384.3200 ;
        RECT 241.6800 372.9600 244.6800 373.4400 ;
        RECT 241.6800 378.4000 244.6800 378.8800 ;
        RECT 241.6800 383.8400 244.6800 384.3200 ;
        RECT 253.4400 362.0800 255.0400 362.5600 ;
        RECT 253.4400 367.5200 255.0400 368.0000 ;
        RECT 241.6800 362.0800 244.6800 362.5600 ;
        RECT 241.6800 367.5200 244.6800 368.0000 ;
        RECT 343.4400 345.7600 345.0400 346.2400 ;
        RECT 343.4400 351.2000 345.0400 351.6800 ;
        RECT 343.4400 356.6400 345.0400 357.1200 ;
        RECT 343.4400 334.8800 345.0400 335.3600 ;
        RECT 343.4400 340.3200 345.0400 340.8000 ;
        RECT 298.4400 345.7600 300.0400 346.2400 ;
        RECT 298.4400 351.2000 300.0400 351.6800 ;
        RECT 298.4400 356.6400 300.0400 357.1200 ;
        RECT 298.4400 334.8800 300.0400 335.3600 ;
        RECT 298.4400 340.3200 300.0400 340.8000 ;
        RECT 343.4400 318.5600 345.0400 319.0400 ;
        RECT 343.4400 324.0000 345.0400 324.4800 ;
        RECT 343.4400 329.4400 345.0400 329.9200 ;
        RECT 343.4400 313.1200 345.0400 313.6000 ;
        RECT 298.4400 318.5600 300.0400 319.0400 ;
        RECT 298.4400 324.0000 300.0400 324.4800 ;
        RECT 298.4400 329.4400 300.0400 329.9200 ;
        RECT 298.4400 313.1200 300.0400 313.6000 ;
        RECT 253.4400 345.7600 255.0400 346.2400 ;
        RECT 253.4400 351.2000 255.0400 351.6800 ;
        RECT 253.4400 356.6400 255.0400 357.1200 ;
        RECT 241.6800 345.7600 244.6800 346.2400 ;
        RECT 241.6800 351.2000 244.6800 351.6800 ;
        RECT 241.6800 356.6400 244.6800 357.1200 ;
        RECT 253.4400 334.8800 255.0400 335.3600 ;
        RECT 253.4400 340.3200 255.0400 340.8000 ;
        RECT 241.6800 334.8800 244.6800 335.3600 ;
        RECT 241.6800 340.3200 244.6800 340.8000 ;
        RECT 253.4400 318.5600 255.0400 319.0400 ;
        RECT 253.4400 324.0000 255.0400 324.4800 ;
        RECT 253.4400 329.4400 255.0400 329.9200 ;
        RECT 241.6800 318.5600 244.6800 319.0400 ;
        RECT 241.6800 324.0000 244.6800 324.4800 ;
        RECT 241.6800 329.4400 244.6800 329.9200 ;
        RECT 241.6800 313.1200 244.6800 313.6000 ;
        RECT 253.4400 313.1200 255.0400 313.6000 ;
        RECT 241.6800 518.0300 448.7800 521.0300 ;
        RECT 241.6800 304.9300 448.7800 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 75.2900 435.0400 291.3900 ;
        RECT 388.4400 75.2900 390.0400 291.3900 ;
        RECT 343.4400 75.2900 345.0400 291.3900 ;
        RECT 298.4400 75.2900 300.0400 291.3900 ;
        RECT 253.4400 75.2900 255.0400 291.3900 ;
        RECT 445.7800 75.2900 448.7800 291.3900 ;
        RECT 241.6800 75.2900 244.6800 291.3900 ;
      LAYER met3 ;
        RECT 445.7800 268.4400 448.7800 268.9200 ;
        RECT 445.7800 273.8800 448.7800 274.3600 ;
        RECT 433.4400 268.4400 435.0400 268.9200 ;
        RECT 433.4400 273.8800 435.0400 274.3600 ;
        RECT 445.7800 279.3200 448.7800 279.8000 ;
        RECT 433.4400 279.3200 435.0400 279.8000 ;
        RECT 445.7800 257.5600 448.7800 258.0400 ;
        RECT 445.7800 263.0000 448.7800 263.4800 ;
        RECT 433.4400 257.5600 435.0400 258.0400 ;
        RECT 433.4400 263.0000 435.0400 263.4800 ;
        RECT 445.7800 241.2400 448.7800 241.7200 ;
        RECT 445.7800 246.6800 448.7800 247.1600 ;
        RECT 433.4400 241.2400 435.0400 241.7200 ;
        RECT 433.4400 246.6800 435.0400 247.1600 ;
        RECT 445.7800 252.1200 448.7800 252.6000 ;
        RECT 433.4400 252.1200 435.0400 252.6000 ;
        RECT 388.4400 268.4400 390.0400 268.9200 ;
        RECT 388.4400 273.8800 390.0400 274.3600 ;
        RECT 388.4400 279.3200 390.0400 279.8000 ;
        RECT 388.4400 257.5600 390.0400 258.0400 ;
        RECT 388.4400 263.0000 390.0400 263.4800 ;
        RECT 388.4400 241.2400 390.0400 241.7200 ;
        RECT 388.4400 246.6800 390.0400 247.1600 ;
        RECT 388.4400 252.1200 390.0400 252.6000 ;
        RECT 445.7800 224.9200 448.7800 225.4000 ;
        RECT 445.7800 230.3600 448.7800 230.8400 ;
        RECT 445.7800 235.8000 448.7800 236.2800 ;
        RECT 433.4400 224.9200 435.0400 225.4000 ;
        RECT 433.4400 230.3600 435.0400 230.8400 ;
        RECT 433.4400 235.8000 435.0400 236.2800 ;
        RECT 445.7800 214.0400 448.7800 214.5200 ;
        RECT 445.7800 219.4800 448.7800 219.9600 ;
        RECT 433.4400 214.0400 435.0400 214.5200 ;
        RECT 433.4400 219.4800 435.0400 219.9600 ;
        RECT 445.7800 197.7200 448.7800 198.2000 ;
        RECT 445.7800 203.1600 448.7800 203.6400 ;
        RECT 445.7800 208.6000 448.7800 209.0800 ;
        RECT 433.4400 197.7200 435.0400 198.2000 ;
        RECT 433.4400 203.1600 435.0400 203.6400 ;
        RECT 433.4400 208.6000 435.0400 209.0800 ;
        RECT 445.7800 186.8400 448.7800 187.3200 ;
        RECT 445.7800 192.2800 448.7800 192.7600 ;
        RECT 433.4400 186.8400 435.0400 187.3200 ;
        RECT 433.4400 192.2800 435.0400 192.7600 ;
        RECT 388.4400 224.9200 390.0400 225.4000 ;
        RECT 388.4400 230.3600 390.0400 230.8400 ;
        RECT 388.4400 235.8000 390.0400 236.2800 ;
        RECT 388.4400 214.0400 390.0400 214.5200 ;
        RECT 388.4400 219.4800 390.0400 219.9600 ;
        RECT 388.4400 197.7200 390.0400 198.2000 ;
        RECT 388.4400 203.1600 390.0400 203.6400 ;
        RECT 388.4400 208.6000 390.0400 209.0800 ;
        RECT 388.4400 186.8400 390.0400 187.3200 ;
        RECT 388.4400 192.2800 390.0400 192.7600 ;
        RECT 343.4400 268.4400 345.0400 268.9200 ;
        RECT 343.4400 273.8800 345.0400 274.3600 ;
        RECT 343.4400 279.3200 345.0400 279.8000 ;
        RECT 298.4400 268.4400 300.0400 268.9200 ;
        RECT 298.4400 273.8800 300.0400 274.3600 ;
        RECT 298.4400 279.3200 300.0400 279.8000 ;
        RECT 343.4400 257.5600 345.0400 258.0400 ;
        RECT 343.4400 263.0000 345.0400 263.4800 ;
        RECT 343.4400 241.2400 345.0400 241.7200 ;
        RECT 343.4400 246.6800 345.0400 247.1600 ;
        RECT 343.4400 252.1200 345.0400 252.6000 ;
        RECT 298.4400 257.5600 300.0400 258.0400 ;
        RECT 298.4400 263.0000 300.0400 263.4800 ;
        RECT 298.4400 241.2400 300.0400 241.7200 ;
        RECT 298.4400 246.6800 300.0400 247.1600 ;
        RECT 298.4400 252.1200 300.0400 252.6000 ;
        RECT 253.4400 268.4400 255.0400 268.9200 ;
        RECT 253.4400 273.8800 255.0400 274.3600 ;
        RECT 241.6800 273.8800 244.6800 274.3600 ;
        RECT 241.6800 268.4400 244.6800 268.9200 ;
        RECT 241.6800 279.3200 244.6800 279.8000 ;
        RECT 253.4400 279.3200 255.0400 279.8000 ;
        RECT 253.4400 257.5600 255.0400 258.0400 ;
        RECT 253.4400 263.0000 255.0400 263.4800 ;
        RECT 241.6800 263.0000 244.6800 263.4800 ;
        RECT 241.6800 257.5600 244.6800 258.0400 ;
        RECT 253.4400 241.2400 255.0400 241.7200 ;
        RECT 253.4400 246.6800 255.0400 247.1600 ;
        RECT 241.6800 246.6800 244.6800 247.1600 ;
        RECT 241.6800 241.2400 244.6800 241.7200 ;
        RECT 241.6800 252.1200 244.6800 252.6000 ;
        RECT 253.4400 252.1200 255.0400 252.6000 ;
        RECT 343.4400 224.9200 345.0400 225.4000 ;
        RECT 343.4400 230.3600 345.0400 230.8400 ;
        RECT 343.4400 235.8000 345.0400 236.2800 ;
        RECT 343.4400 214.0400 345.0400 214.5200 ;
        RECT 343.4400 219.4800 345.0400 219.9600 ;
        RECT 298.4400 224.9200 300.0400 225.4000 ;
        RECT 298.4400 230.3600 300.0400 230.8400 ;
        RECT 298.4400 235.8000 300.0400 236.2800 ;
        RECT 298.4400 214.0400 300.0400 214.5200 ;
        RECT 298.4400 219.4800 300.0400 219.9600 ;
        RECT 343.4400 197.7200 345.0400 198.2000 ;
        RECT 343.4400 203.1600 345.0400 203.6400 ;
        RECT 343.4400 208.6000 345.0400 209.0800 ;
        RECT 343.4400 186.8400 345.0400 187.3200 ;
        RECT 343.4400 192.2800 345.0400 192.7600 ;
        RECT 298.4400 197.7200 300.0400 198.2000 ;
        RECT 298.4400 203.1600 300.0400 203.6400 ;
        RECT 298.4400 208.6000 300.0400 209.0800 ;
        RECT 298.4400 186.8400 300.0400 187.3200 ;
        RECT 298.4400 192.2800 300.0400 192.7600 ;
        RECT 253.4400 224.9200 255.0400 225.4000 ;
        RECT 253.4400 230.3600 255.0400 230.8400 ;
        RECT 253.4400 235.8000 255.0400 236.2800 ;
        RECT 241.6800 224.9200 244.6800 225.4000 ;
        RECT 241.6800 230.3600 244.6800 230.8400 ;
        RECT 241.6800 235.8000 244.6800 236.2800 ;
        RECT 253.4400 214.0400 255.0400 214.5200 ;
        RECT 253.4400 219.4800 255.0400 219.9600 ;
        RECT 241.6800 214.0400 244.6800 214.5200 ;
        RECT 241.6800 219.4800 244.6800 219.9600 ;
        RECT 253.4400 197.7200 255.0400 198.2000 ;
        RECT 253.4400 203.1600 255.0400 203.6400 ;
        RECT 253.4400 208.6000 255.0400 209.0800 ;
        RECT 241.6800 197.7200 244.6800 198.2000 ;
        RECT 241.6800 203.1600 244.6800 203.6400 ;
        RECT 241.6800 208.6000 244.6800 209.0800 ;
        RECT 253.4400 186.8400 255.0400 187.3200 ;
        RECT 253.4400 192.2800 255.0400 192.7600 ;
        RECT 241.6800 186.8400 244.6800 187.3200 ;
        RECT 241.6800 192.2800 244.6800 192.7600 ;
        RECT 445.7800 170.5200 448.7800 171.0000 ;
        RECT 445.7800 175.9600 448.7800 176.4400 ;
        RECT 445.7800 181.4000 448.7800 181.8800 ;
        RECT 433.4400 170.5200 435.0400 171.0000 ;
        RECT 433.4400 175.9600 435.0400 176.4400 ;
        RECT 433.4400 181.4000 435.0400 181.8800 ;
        RECT 445.7800 159.6400 448.7800 160.1200 ;
        RECT 445.7800 165.0800 448.7800 165.5600 ;
        RECT 433.4400 159.6400 435.0400 160.1200 ;
        RECT 433.4400 165.0800 435.0400 165.5600 ;
        RECT 445.7800 143.3200 448.7800 143.8000 ;
        RECT 445.7800 148.7600 448.7800 149.2400 ;
        RECT 445.7800 154.2000 448.7800 154.6800 ;
        RECT 433.4400 143.3200 435.0400 143.8000 ;
        RECT 433.4400 148.7600 435.0400 149.2400 ;
        RECT 433.4400 154.2000 435.0400 154.6800 ;
        RECT 445.7800 132.4400 448.7800 132.9200 ;
        RECT 445.7800 137.8800 448.7800 138.3600 ;
        RECT 433.4400 132.4400 435.0400 132.9200 ;
        RECT 433.4400 137.8800 435.0400 138.3600 ;
        RECT 388.4400 170.5200 390.0400 171.0000 ;
        RECT 388.4400 175.9600 390.0400 176.4400 ;
        RECT 388.4400 181.4000 390.0400 181.8800 ;
        RECT 388.4400 159.6400 390.0400 160.1200 ;
        RECT 388.4400 165.0800 390.0400 165.5600 ;
        RECT 388.4400 143.3200 390.0400 143.8000 ;
        RECT 388.4400 148.7600 390.0400 149.2400 ;
        RECT 388.4400 154.2000 390.0400 154.6800 ;
        RECT 388.4400 132.4400 390.0400 132.9200 ;
        RECT 388.4400 137.8800 390.0400 138.3600 ;
        RECT 445.7800 116.1200 448.7800 116.6000 ;
        RECT 445.7800 121.5600 448.7800 122.0400 ;
        RECT 445.7800 127.0000 448.7800 127.4800 ;
        RECT 433.4400 116.1200 435.0400 116.6000 ;
        RECT 433.4400 121.5600 435.0400 122.0400 ;
        RECT 433.4400 127.0000 435.0400 127.4800 ;
        RECT 445.7800 105.2400 448.7800 105.7200 ;
        RECT 445.7800 110.6800 448.7800 111.1600 ;
        RECT 433.4400 105.2400 435.0400 105.7200 ;
        RECT 433.4400 110.6800 435.0400 111.1600 ;
        RECT 445.7800 88.9200 448.7800 89.4000 ;
        RECT 445.7800 94.3600 448.7800 94.8400 ;
        RECT 445.7800 99.8000 448.7800 100.2800 ;
        RECT 433.4400 88.9200 435.0400 89.4000 ;
        RECT 433.4400 94.3600 435.0400 94.8400 ;
        RECT 433.4400 99.8000 435.0400 100.2800 ;
        RECT 445.7800 83.4800 448.7800 83.9600 ;
        RECT 433.4400 83.4800 435.0400 83.9600 ;
        RECT 388.4400 116.1200 390.0400 116.6000 ;
        RECT 388.4400 121.5600 390.0400 122.0400 ;
        RECT 388.4400 127.0000 390.0400 127.4800 ;
        RECT 388.4400 105.2400 390.0400 105.7200 ;
        RECT 388.4400 110.6800 390.0400 111.1600 ;
        RECT 388.4400 88.9200 390.0400 89.4000 ;
        RECT 388.4400 94.3600 390.0400 94.8400 ;
        RECT 388.4400 99.8000 390.0400 100.2800 ;
        RECT 388.4400 83.4800 390.0400 83.9600 ;
        RECT 343.4400 170.5200 345.0400 171.0000 ;
        RECT 343.4400 175.9600 345.0400 176.4400 ;
        RECT 343.4400 181.4000 345.0400 181.8800 ;
        RECT 343.4400 159.6400 345.0400 160.1200 ;
        RECT 343.4400 165.0800 345.0400 165.5600 ;
        RECT 298.4400 170.5200 300.0400 171.0000 ;
        RECT 298.4400 175.9600 300.0400 176.4400 ;
        RECT 298.4400 181.4000 300.0400 181.8800 ;
        RECT 298.4400 159.6400 300.0400 160.1200 ;
        RECT 298.4400 165.0800 300.0400 165.5600 ;
        RECT 343.4400 143.3200 345.0400 143.8000 ;
        RECT 343.4400 148.7600 345.0400 149.2400 ;
        RECT 343.4400 154.2000 345.0400 154.6800 ;
        RECT 343.4400 132.4400 345.0400 132.9200 ;
        RECT 343.4400 137.8800 345.0400 138.3600 ;
        RECT 298.4400 143.3200 300.0400 143.8000 ;
        RECT 298.4400 148.7600 300.0400 149.2400 ;
        RECT 298.4400 154.2000 300.0400 154.6800 ;
        RECT 298.4400 132.4400 300.0400 132.9200 ;
        RECT 298.4400 137.8800 300.0400 138.3600 ;
        RECT 253.4400 170.5200 255.0400 171.0000 ;
        RECT 253.4400 175.9600 255.0400 176.4400 ;
        RECT 253.4400 181.4000 255.0400 181.8800 ;
        RECT 241.6800 170.5200 244.6800 171.0000 ;
        RECT 241.6800 175.9600 244.6800 176.4400 ;
        RECT 241.6800 181.4000 244.6800 181.8800 ;
        RECT 253.4400 159.6400 255.0400 160.1200 ;
        RECT 253.4400 165.0800 255.0400 165.5600 ;
        RECT 241.6800 159.6400 244.6800 160.1200 ;
        RECT 241.6800 165.0800 244.6800 165.5600 ;
        RECT 253.4400 143.3200 255.0400 143.8000 ;
        RECT 253.4400 148.7600 255.0400 149.2400 ;
        RECT 253.4400 154.2000 255.0400 154.6800 ;
        RECT 241.6800 143.3200 244.6800 143.8000 ;
        RECT 241.6800 148.7600 244.6800 149.2400 ;
        RECT 241.6800 154.2000 244.6800 154.6800 ;
        RECT 253.4400 132.4400 255.0400 132.9200 ;
        RECT 253.4400 137.8800 255.0400 138.3600 ;
        RECT 241.6800 132.4400 244.6800 132.9200 ;
        RECT 241.6800 137.8800 244.6800 138.3600 ;
        RECT 343.4400 116.1200 345.0400 116.6000 ;
        RECT 343.4400 121.5600 345.0400 122.0400 ;
        RECT 343.4400 127.0000 345.0400 127.4800 ;
        RECT 343.4400 105.2400 345.0400 105.7200 ;
        RECT 343.4400 110.6800 345.0400 111.1600 ;
        RECT 298.4400 116.1200 300.0400 116.6000 ;
        RECT 298.4400 121.5600 300.0400 122.0400 ;
        RECT 298.4400 127.0000 300.0400 127.4800 ;
        RECT 298.4400 105.2400 300.0400 105.7200 ;
        RECT 298.4400 110.6800 300.0400 111.1600 ;
        RECT 343.4400 88.9200 345.0400 89.4000 ;
        RECT 343.4400 94.3600 345.0400 94.8400 ;
        RECT 343.4400 99.8000 345.0400 100.2800 ;
        RECT 343.4400 83.4800 345.0400 83.9600 ;
        RECT 298.4400 88.9200 300.0400 89.4000 ;
        RECT 298.4400 94.3600 300.0400 94.8400 ;
        RECT 298.4400 99.8000 300.0400 100.2800 ;
        RECT 298.4400 83.4800 300.0400 83.9600 ;
        RECT 253.4400 116.1200 255.0400 116.6000 ;
        RECT 253.4400 121.5600 255.0400 122.0400 ;
        RECT 253.4400 127.0000 255.0400 127.4800 ;
        RECT 241.6800 116.1200 244.6800 116.6000 ;
        RECT 241.6800 121.5600 244.6800 122.0400 ;
        RECT 241.6800 127.0000 244.6800 127.4800 ;
        RECT 253.4400 105.2400 255.0400 105.7200 ;
        RECT 253.4400 110.6800 255.0400 111.1600 ;
        RECT 241.6800 105.2400 244.6800 105.7200 ;
        RECT 241.6800 110.6800 244.6800 111.1600 ;
        RECT 253.4400 88.9200 255.0400 89.4000 ;
        RECT 253.4400 94.3600 255.0400 94.8400 ;
        RECT 253.4400 99.8000 255.0400 100.2800 ;
        RECT 241.6800 88.9200 244.6800 89.4000 ;
        RECT 241.6800 94.3600 244.6800 94.8400 ;
        RECT 241.6800 99.8000 244.6800 100.2800 ;
        RECT 241.6800 83.4800 244.6800 83.9600 ;
        RECT 253.4400 83.4800 255.0400 83.9600 ;
        RECT 241.6800 288.3900 448.7800 291.3900 ;
        RECT 241.6800 75.2900 448.7800 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 242.6800 34.6700 244.6800 61.6000 ;
        RECT 445.7800 34.6700 447.7800 61.6000 ;
      LAYER met3 ;
        RECT 445.7800 51.3800 447.7800 51.8600 ;
        RECT 242.6800 51.3800 244.6800 51.8600 ;
        RECT 445.7800 45.9400 447.7800 46.4200 ;
        RECT 445.7800 40.5000 447.7800 40.9800 ;
        RECT 242.6800 45.9400 244.6800 46.4200 ;
        RECT 242.6800 40.5000 244.6800 40.9800 ;
        RECT 242.6800 59.6000 447.7800 61.6000 ;
        RECT 242.6800 34.6700 447.7800 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 2601.3300 435.0400 2817.4300 ;
        RECT 388.4400 2601.3300 390.0400 2817.4300 ;
        RECT 343.4400 2601.3300 345.0400 2817.4300 ;
        RECT 298.4400 2601.3300 300.0400 2817.4300 ;
        RECT 253.4400 2601.3300 255.0400 2817.4300 ;
        RECT 445.7800 2601.3300 448.7800 2817.4300 ;
        RECT 241.6800 2601.3300 244.6800 2817.4300 ;
      LAYER met3 ;
        RECT 445.7800 2794.4800 448.7800 2794.9600 ;
        RECT 445.7800 2799.9200 448.7800 2800.4000 ;
        RECT 433.4400 2794.4800 435.0400 2794.9600 ;
        RECT 433.4400 2799.9200 435.0400 2800.4000 ;
        RECT 445.7800 2805.3600 448.7800 2805.8400 ;
        RECT 433.4400 2805.3600 435.0400 2805.8400 ;
        RECT 445.7800 2783.6000 448.7800 2784.0800 ;
        RECT 445.7800 2789.0400 448.7800 2789.5200 ;
        RECT 433.4400 2783.6000 435.0400 2784.0800 ;
        RECT 433.4400 2789.0400 435.0400 2789.5200 ;
        RECT 445.7800 2767.2800 448.7800 2767.7600 ;
        RECT 445.7800 2772.7200 448.7800 2773.2000 ;
        RECT 433.4400 2767.2800 435.0400 2767.7600 ;
        RECT 433.4400 2772.7200 435.0400 2773.2000 ;
        RECT 445.7800 2778.1600 448.7800 2778.6400 ;
        RECT 433.4400 2778.1600 435.0400 2778.6400 ;
        RECT 388.4400 2794.4800 390.0400 2794.9600 ;
        RECT 388.4400 2799.9200 390.0400 2800.4000 ;
        RECT 388.4400 2805.3600 390.0400 2805.8400 ;
        RECT 388.4400 2783.6000 390.0400 2784.0800 ;
        RECT 388.4400 2789.0400 390.0400 2789.5200 ;
        RECT 388.4400 2767.2800 390.0400 2767.7600 ;
        RECT 388.4400 2772.7200 390.0400 2773.2000 ;
        RECT 388.4400 2778.1600 390.0400 2778.6400 ;
        RECT 445.7800 2750.9600 448.7800 2751.4400 ;
        RECT 445.7800 2756.4000 448.7800 2756.8800 ;
        RECT 445.7800 2761.8400 448.7800 2762.3200 ;
        RECT 433.4400 2750.9600 435.0400 2751.4400 ;
        RECT 433.4400 2756.4000 435.0400 2756.8800 ;
        RECT 433.4400 2761.8400 435.0400 2762.3200 ;
        RECT 445.7800 2740.0800 448.7800 2740.5600 ;
        RECT 445.7800 2745.5200 448.7800 2746.0000 ;
        RECT 433.4400 2740.0800 435.0400 2740.5600 ;
        RECT 433.4400 2745.5200 435.0400 2746.0000 ;
        RECT 445.7800 2723.7600 448.7800 2724.2400 ;
        RECT 445.7800 2729.2000 448.7800 2729.6800 ;
        RECT 445.7800 2734.6400 448.7800 2735.1200 ;
        RECT 433.4400 2723.7600 435.0400 2724.2400 ;
        RECT 433.4400 2729.2000 435.0400 2729.6800 ;
        RECT 433.4400 2734.6400 435.0400 2735.1200 ;
        RECT 445.7800 2712.8800 448.7800 2713.3600 ;
        RECT 445.7800 2718.3200 448.7800 2718.8000 ;
        RECT 433.4400 2712.8800 435.0400 2713.3600 ;
        RECT 433.4400 2718.3200 435.0400 2718.8000 ;
        RECT 388.4400 2750.9600 390.0400 2751.4400 ;
        RECT 388.4400 2756.4000 390.0400 2756.8800 ;
        RECT 388.4400 2761.8400 390.0400 2762.3200 ;
        RECT 388.4400 2740.0800 390.0400 2740.5600 ;
        RECT 388.4400 2745.5200 390.0400 2746.0000 ;
        RECT 388.4400 2723.7600 390.0400 2724.2400 ;
        RECT 388.4400 2729.2000 390.0400 2729.6800 ;
        RECT 388.4400 2734.6400 390.0400 2735.1200 ;
        RECT 388.4400 2712.8800 390.0400 2713.3600 ;
        RECT 388.4400 2718.3200 390.0400 2718.8000 ;
        RECT 343.4400 2794.4800 345.0400 2794.9600 ;
        RECT 343.4400 2799.9200 345.0400 2800.4000 ;
        RECT 343.4400 2805.3600 345.0400 2805.8400 ;
        RECT 298.4400 2794.4800 300.0400 2794.9600 ;
        RECT 298.4400 2799.9200 300.0400 2800.4000 ;
        RECT 298.4400 2805.3600 300.0400 2805.8400 ;
        RECT 343.4400 2783.6000 345.0400 2784.0800 ;
        RECT 343.4400 2789.0400 345.0400 2789.5200 ;
        RECT 343.4400 2767.2800 345.0400 2767.7600 ;
        RECT 343.4400 2772.7200 345.0400 2773.2000 ;
        RECT 343.4400 2778.1600 345.0400 2778.6400 ;
        RECT 298.4400 2783.6000 300.0400 2784.0800 ;
        RECT 298.4400 2789.0400 300.0400 2789.5200 ;
        RECT 298.4400 2767.2800 300.0400 2767.7600 ;
        RECT 298.4400 2772.7200 300.0400 2773.2000 ;
        RECT 298.4400 2778.1600 300.0400 2778.6400 ;
        RECT 253.4400 2794.4800 255.0400 2794.9600 ;
        RECT 253.4400 2799.9200 255.0400 2800.4000 ;
        RECT 241.6800 2799.9200 244.6800 2800.4000 ;
        RECT 241.6800 2794.4800 244.6800 2794.9600 ;
        RECT 241.6800 2805.3600 244.6800 2805.8400 ;
        RECT 253.4400 2805.3600 255.0400 2805.8400 ;
        RECT 253.4400 2783.6000 255.0400 2784.0800 ;
        RECT 253.4400 2789.0400 255.0400 2789.5200 ;
        RECT 241.6800 2789.0400 244.6800 2789.5200 ;
        RECT 241.6800 2783.6000 244.6800 2784.0800 ;
        RECT 253.4400 2767.2800 255.0400 2767.7600 ;
        RECT 253.4400 2772.7200 255.0400 2773.2000 ;
        RECT 241.6800 2772.7200 244.6800 2773.2000 ;
        RECT 241.6800 2767.2800 244.6800 2767.7600 ;
        RECT 241.6800 2778.1600 244.6800 2778.6400 ;
        RECT 253.4400 2778.1600 255.0400 2778.6400 ;
        RECT 343.4400 2750.9600 345.0400 2751.4400 ;
        RECT 343.4400 2756.4000 345.0400 2756.8800 ;
        RECT 343.4400 2761.8400 345.0400 2762.3200 ;
        RECT 343.4400 2740.0800 345.0400 2740.5600 ;
        RECT 343.4400 2745.5200 345.0400 2746.0000 ;
        RECT 298.4400 2750.9600 300.0400 2751.4400 ;
        RECT 298.4400 2756.4000 300.0400 2756.8800 ;
        RECT 298.4400 2761.8400 300.0400 2762.3200 ;
        RECT 298.4400 2740.0800 300.0400 2740.5600 ;
        RECT 298.4400 2745.5200 300.0400 2746.0000 ;
        RECT 343.4400 2723.7600 345.0400 2724.2400 ;
        RECT 343.4400 2729.2000 345.0400 2729.6800 ;
        RECT 343.4400 2734.6400 345.0400 2735.1200 ;
        RECT 343.4400 2712.8800 345.0400 2713.3600 ;
        RECT 343.4400 2718.3200 345.0400 2718.8000 ;
        RECT 298.4400 2723.7600 300.0400 2724.2400 ;
        RECT 298.4400 2729.2000 300.0400 2729.6800 ;
        RECT 298.4400 2734.6400 300.0400 2735.1200 ;
        RECT 298.4400 2712.8800 300.0400 2713.3600 ;
        RECT 298.4400 2718.3200 300.0400 2718.8000 ;
        RECT 253.4400 2750.9600 255.0400 2751.4400 ;
        RECT 253.4400 2756.4000 255.0400 2756.8800 ;
        RECT 253.4400 2761.8400 255.0400 2762.3200 ;
        RECT 241.6800 2750.9600 244.6800 2751.4400 ;
        RECT 241.6800 2756.4000 244.6800 2756.8800 ;
        RECT 241.6800 2761.8400 244.6800 2762.3200 ;
        RECT 253.4400 2740.0800 255.0400 2740.5600 ;
        RECT 253.4400 2745.5200 255.0400 2746.0000 ;
        RECT 241.6800 2740.0800 244.6800 2740.5600 ;
        RECT 241.6800 2745.5200 244.6800 2746.0000 ;
        RECT 253.4400 2723.7600 255.0400 2724.2400 ;
        RECT 253.4400 2729.2000 255.0400 2729.6800 ;
        RECT 253.4400 2734.6400 255.0400 2735.1200 ;
        RECT 241.6800 2723.7600 244.6800 2724.2400 ;
        RECT 241.6800 2729.2000 244.6800 2729.6800 ;
        RECT 241.6800 2734.6400 244.6800 2735.1200 ;
        RECT 253.4400 2712.8800 255.0400 2713.3600 ;
        RECT 253.4400 2718.3200 255.0400 2718.8000 ;
        RECT 241.6800 2712.8800 244.6800 2713.3600 ;
        RECT 241.6800 2718.3200 244.6800 2718.8000 ;
        RECT 445.7800 2696.5600 448.7800 2697.0400 ;
        RECT 445.7800 2702.0000 448.7800 2702.4800 ;
        RECT 445.7800 2707.4400 448.7800 2707.9200 ;
        RECT 433.4400 2696.5600 435.0400 2697.0400 ;
        RECT 433.4400 2702.0000 435.0400 2702.4800 ;
        RECT 433.4400 2707.4400 435.0400 2707.9200 ;
        RECT 445.7800 2685.6800 448.7800 2686.1600 ;
        RECT 445.7800 2691.1200 448.7800 2691.6000 ;
        RECT 433.4400 2685.6800 435.0400 2686.1600 ;
        RECT 433.4400 2691.1200 435.0400 2691.6000 ;
        RECT 445.7800 2669.3600 448.7800 2669.8400 ;
        RECT 445.7800 2674.8000 448.7800 2675.2800 ;
        RECT 445.7800 2680.2400 448.7800 2680.7200 ;
        RECT 433.4400 2669.3600 435.0400 2669.8400 ;
        RECT 433.4400 2674.8000 435.0400 2675.2800 ;
        RECT 433.4400 2680.2400 435.0400 2680.7200 ;
        RECT 445.7800 2658.4800 448.7800 2658.9600 ;
        RECT 445.7800 2663.9200 448.7800 2664.4000 ;
        RECT 433.4400 2658.4800 435.0400 2658.9600 ;
        RECT 433.4400 2663.9200 435.0400 2664.4000 ;
        RECT 388.4400 2696.5600 390.0400 2697.0400 ;
        RECT 388.4400 2702.0000 390.0400 2702.4800 ;
        RECT 388.4400 2707.4400 390.0400 2707.9200 ;
        RECT 388.4400 2685.6800 390.0400 2686.1600 ;
        RECT 388.4400 2691.1200 390.0400 2691.6000 ;
        RECT 388.4400 2669.3600 390.0400 2669.8400 ;
        RECT 388.4400 2674.8000 390.0400 2675.2800 ;
        RECT 388.4400 2680.2400 390.0400 2680.7200 ;
        RECT 388.4400 2658.4800 390.0400 2658.9600 ;
        RECT 388.4400 2663.9200 390.0400 2664.4000 ;
        RECT 445.7800 2642.1600 448.7800 2642.6400 ;
        RECT 445.7800 2647.6000 448.7800 2648.0800 ;
        RECT 445.7800 2653.0400 448.7800 2653.5200 ;
        RECT 433.4400 2642.1600 435.0400 2642.6400 ;
        RECT 433.4400 2647.6000 435.0400 2648.0800 ;
        RECT 433.4400 2653.0400 435.0400 2653.5200 ;
        RECT 445.7800 2631.2800 448.7800 2631.7600 ;
        RECT 445.7800 2636.7200 448.7800 2637.2000 ;
        RECT 433.4400 2631.2800 435.0400 2631.7600 ;
        RECT 433.4400 2636.7200 435.0400 2637.2000 ;
        RECT 445.7800 2614.9600 448.7800 2615.4400 ;
        RECT 445.7800 2620.4000 448.7800 2620.8800 ;
        RECT 445.7800 2625.8400 448.7800 2626.3200 ;
        RECT 433.4400 2614.9600 435.0400 2615.4400 ;
        RECT 433.4400 2620.4000 435.0400 2620.8800 ;
        RECT 433.4400 2625.8400 435.0400 2626.3200 ;
        RECT 445.7800 2609.5200 448.7800 2610.0000 ;
        RECT 433.4400 2609.5200 435.0400 2610.0000 ;
        RECT 388.4400 2642.1600 390.0400 2642.6400 ;
        RECT 388.4400 2647.6000 390.0400 2648.0800 ;
        RECT 388.4400 2653.0400 390.0400 2653.5200 ;
        RECT 388.4400 2631.2800 390.0400 2631.7600 ;
        RECT 388.4400 2636.7200 390.0400 2637.2000 ;
        RECT 388.4400 2614.9600 390.0400 2615.4400 ;
        RECT 388.4400 2620.4000 390.0400 2620.8800 ;
        RECT 388.4400 2625.8400 390.0400 2626.3200 ;
        RECT 388.4400 2609.5200 390.0400 2610.0000 ;
        RECT 343.4400 2696.5600 345.0400 2697.0400 ;
        RECT 343.4400 2702.0000 345.0400 2702.4800 ;
        RECT 343.4400 2707.4400 345.0400 2707.9200 ;
        RECT 343.4400 2685.6800 345.0400 2686.1600 ;
        RECT 343.4400 2691.1200 345.0400 2691.6000 ;
        RECT 298.4400 2696.5600 300.0400 2697.0400 ;
        RECT 298.4400 2702.0000 300.0400 2702.4800 ;
        RECT 298.4400 2707.4400 300.0400 2707.9200 ;
        RECT 298.4400 2685.6800 300.0400 2686.1600 ;
        RECT 298.4400 2691.1200 300.0400 2691.6000 ;
        RECT 343.4400 2669.3600 345.0400 2669.8400 ;
        RECT 343.4400 2674.8000 345.0400 2675.2800 ;
        RECT 343.4400 2680.2400 345.0400 2680.7200 ;
        RECT 343.4400 2658.4800 345.0400 2658.9600 ;
        RECT 343.4400 2663.9200 345.0400 2664.4000 ;
        RECT 298.4400 2669.3600 300.0400 2669.8400 ;
        RECT 298.4400 2674.8000 300.0400 2675.2800 ;
        RECT 298.4400 2680.2400 300.0400 2680.7200 ;
        RECT 298.4400 2658.4800 300.0400 2658.9600 ;
        RECT 298.4400 2663.9200 300.0400 2664.4000 ;
        RECT 253.4400 2696.5600 255.0400 2697.0400 ;
        RECT 253.4400 2702.0000 255.0400 2702.4800 ;
        RECT 253.4400 2707.4400 255.0400 2707.9200 ;
        RECT 241.6800 2696.5600 244.6800 2697.0400 ;
        RECT 241.6800 2702.0000 244.6800 2702.4800 ;
        RECT 241.6800 2707.4400 244.6800 2707.9200 ;
        RECT 253.4400 2685.6800 255.0400 2686.1600 ;
        RECT 253.4400 2691.1200 255.0400 2691.6000 ;
        RECT 241.6800 2685.6800 244.6800 2686.1600 ;
        RECT 241.6800 2691.1200 244.6800 2691.6000 ;
        RECT 253.4400 2669.3600 255.0400 2669.8400 ;
        RECT 253.4400 2674.8000 255.0400 2675.2800 ;
        RECT 253.4400 2680.2400 255.0400 2680.7200 ;
        RECT 241.6800 2669.3600 244.6800 2669.8400 ;
        RECT 241.6800 2674.8000 244.6800 2675.2800 ;
        RECT 241.6800 2680.2400 244.6800 2680.7200 ;
        RECT 253.4400 2658.4800 255.0400 2658.9600 ;
        RECT 253.4400 2663.9200 255.0400 2664.4000 ;
        RECT 241.6800 2658.4800 244.6800 2658.9600 ;
        RECT 241.6800 2663.9200 244.6800 2664.4000 ;
        RECT 343.4400 2642.1600 345.0400 2642.6400 ;
        RECT 343.4400 2647.6000 345.0400 2648.0800 ;
        RECT 343.4400 2653.0400 345.0400 2653.5200 ;
        RECT 343.4400 2631.2800 345.0400 2631.7600 ;
        RECT 343.4400 2636.7200 345.0400 2637.2000 ;
        RECT 298.4400 2642.1600 300.0400 2642.6400 ;
        RECT 298.4400 2647.6000 300.0400 2648.0800 ;
        RECT 298.4400 2653.0400 300.0400 2653.5200 ;
        RECT 298.4400 2631.2800 300.0400 2631.7600 ;
        RECT 298.4400 2636.7200 300.0400 2637.2000 ;
        RECT 343.4400 2614.9600 345.0400 2615.4400 ;
        RECT 343.4400 2620.4000 345.0400 2620.8800 ;
        RECT 343.4400 2625.8400 345.0400 2626.3200 ;
        RECT 343.4400 2609.5200 345.0400 2610.0000 ;
        RECT 298.4400 2614.9600 300.0400 2615.4400 ;
        RECT 298.4400 2620.4000 300.0400 2620.8800 ;
        RECT 298.4400 2625.8400 300.0400 2626.3200 ;
        RECT 298.4400 2609.5200 300.0400 2610.0000 ;
        RECT 253.4400 2642.1600 255.0400 2642.6400 ;
        RECT 253.4400 2647.6000 255.0400 2648.0800 ;
        RECT 253.4400 2653.0400 255.0400 2653.5200 ;
        RECT 241.6800 2642.1600 244.6800 2642.6400 ;
        RECT 241.6800 2647.6000 244.6800 2648.0800 ;
        RECT 241.6800 2653.0400 244.6800 2653.5200 ;
        RECT 253.4400 2631.2800 255.0400 2631.7600 ;
        RECT 253.4400 2636.7200 255.0400 2637.2000 ;
        RECT 241.6800 2631.2800 244.6800 2631.7600 ;
        RECT 241.6800 2636.7200 244.6800 2637.2000 ;
        RECT 253.4400 2614.9600 255.0400 2615.4400 ;
        RECT 253.4400 2620.4000 255.0400 2620.8800 ;
        RECT 253.4400 2625.8400 255.0400 2626.3200 ;
        RECT 241.6800 2614.9600 244.6800 2615.4400 ;
        RECT 241.6800 2620.4000 244.6800 2620.8800 ;
        RECT 241.6800 2625.8400 244.6800 2626.3200 ;
        RECT 241.6800 2609.5200 244.6800 2610.0000 ;
        RECT 253.4400 2609.5200 255.0400 2610.0000 ;
        RECT 241.6800 2814.4300 448.7800 2817.4300 ;
        RECT 241.6800 2601.3300 448.7800 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 2371.6900 435.0400 2587.7900 ;
        RECT 388.4400 2371.6900 390.0400 2587.7900 ;
        RECT 343.4400 2371.6900 345.0400 2587.7900 ;
        RECT 298.4400 2371.6900 300.0400 2587.7900 ;
        RECT 253.4400 2371.6900 255.0400 2587.7900 ;
        RECT 445.7800 2371.6900 448.7800 2587.7900 ;
        RECT 241.6800 2371.6900 244.6800 2587.7900 ;
      LAYER met3 ;
        RECT 445.7800 2564.8400 448.7800 2565.3200 ;
        RECT 445.7800 2570.2800 448.7800 2570.7600 ;
        RECT 433.4400 2564.8400 435.0400 2565.3200 ;
        RECT 433.4400 2570.2800 435.0400 2570.7600 ;
        RECT 445.7800 2575.7200 448.7800 2576.2000 ;
        RECT 433.4400 2575.7200 435.0400 2576.2000 ;
        RECT 445.7800 2553.9600 448.7800 2554.4400 ;
        RECT 445.7800 2559.4000 448.7800 2559.8800 ;
        RECT 433.4400 2553.9600 435.0400 2554.4400 ;
        RECT 433.4400 2559.4000 435.0400 2559.8800 ;
        RECT 445.7800 2537.6400 448.7800 2538.1200 ;
        RECT 445.7800 2543.0800 448.7800 2543.5600 ;
        RECT 433.4400 2537.6400 435.0400 2538.1200 ;
        RECT 433.4400 2543.0800 435.0400 2543.5600 ;
        RECT 445.7800 2548.5200 448.7800 2549.0000 ;
        RECT 433.4400 2548.5200 435.0400 2549.0000 ;
        RECT 388.4400 2564.8400 390.0400 2565.3200 ;
        RECT 388.4400 2570.2800 390.0400 2570.7600 ;
        RECT 388.4400 2575.7200 390.0400 2576.2000 ;
        RECT 388.4400 2553.9600 390.0400 2554.4400 ;
        RECT 388.4400 2559.4000 390.0400 2559.8800 ;
        RECT 388.4400 2537.6400 390.0400 2538.1200 ;
        RECT 388.4400 2543.0800 390.0400 2543.5600 ;
        RECT 388.4400 2548.5200 390.0400 2549.0000 ;
        RECT 445.7800 2521.3200 448.7800 2521.8000 ;
        RECT 445.7800 2526.7600 448.7800 2527.2400 ;
        RECT 445.7800 2532.2000 448.7800 2532.6800 ;
        RECT 433.4400 2521.3200 435.0400 2521.8000 ;
        RECT 433.4400 2526.7600 435.0400 2527.2400 ;
        RECT 433.4400 2532.2000 435.0400 2532.6800 ;
        RECT 445.7800 2510.4400 448.7800 2510.9200 ;
        RECT 445.7800 2515.8800 448.7800 2516.3600 ;
        RECT 433.4400 2510.4400 435.0400 2510.9200 ;
        RECT 433.4400 2515.8800 435.0400 2516.3600 ;
        RECT 445.7800 2494.1200 448.7800 2494.6000 ;
        RECT 445.7800 2499.5600 448.7800 2500.0400 ;
        RECT 445.7800 2505.0000 448.7800 2505.4800 ;
        RECT 433.4400 2494.1200 435.0400 2494.6000 ;
        RECT 433.4400 2499.5600 435.0400 2500.0400 ;
        RECT 433.4400 2505.0000 435.0400 2505.4800 ;
        RECT 445.7800 2483.2400 448.7800 2483.7200 ;
        RECT 445.7800 2488.6800 448.7800 2489.1600 ;
        RECT 433.4400 2483.2400 435.0400 2483.7200 ;
        RECT 433.4400 2488.6800 435.0400 2489.1600 ;
        RECT 388.4400 2521.3200 390.0400 2521.8000 ;
        RECT 388.4400 2526.7600 390.0400 2527.2400 ;
        RECT 388.4400 2532.2000 390.0400 2532.6800 ;
        RECT 388.4400 2510.4400 390.0400 2510.9200 ;
        RECT 388.4400 2515.8800 390.0400 2516.3600 ;
        RECT 388.4400 2494.1200 390.0400 2494.6000 ;
        RECT 388.4400 2499.5600 390.0400 2500.0400 ;
        RECT 388.4400 2505.0000 390.0400 2505.4800 ;
        RECT 388.4400 2483.2400 390.0400 2483.7200 ;
        RECT 388.4400 2488.6800 390.0400 2489.1600 ;
        RECT 343.4400 2564.8400 345.0400 2565.3200 ;
        RECT 343.4400 2570.2800 345.0400 2570.7600 ;
        RECT 343.4400 2575.7200 345.0400 2576.2000 ;
        RECT 298.4400 2564.8400 300.0400 2565.3200 ;
        RECT 298.4400 2570.2800 300.0400 2570.7600 ;
        RECT 298.4400 2575.7200 300.0400 2576.2000 ;
        RECT 343.4400 2553.9600 345.0400 2554.4400 ;
        RECT 343.4400 2559.4000 345.0400 2559.8800 ;
        RECT 343.4400 2537.6400 345.0400 2538.1200 ;
        RECT 343.4400 2543.0800 345.0400 2543.5600 ;
        RECT 343.4400 2548.5200 345.0400 2549.0000 ;
        RECT 298.4400 2553.9600 300.0400 2554.4400 ;
        RECT 298.4400 2559.4000 300.0400 2559.8800 ;
        RECT 298.4400 2537.6400 300.0400 2538.1200 ;
        RECT 298.4400 2543.0800 300.0400 2543.5600 ;
        RECT 298.4400 2548.5200 300.0400 2549.0000 ;
        RECT 253.4400 2564.8400 255.0400 2565.3200 ;
        RECT 253.4400 2570.2800 255.0400 2570.7600 ;
        RECT 241.6800 2570.2800 244.6800 2570.7600 ;
        RECT 241.6800 2564.8400 244.6800 2565.3200 ;
        RECT 241.6800 2575.7200 244.6800 2576.2000 ;
        RECT 253.4400 2575.7200 255.0400 2576.2000 ;
        RECT 253.4400 2553.9600 255.0400 2554.4400 ;
        RECT 253.4400 2559.4000 255.0400 2559.8800 ;
        RECT 241.6800 2559.4000 244.6800 2559.8800 ;
        RECT 241.6800 2553.9600 244.6800 2554.4400 ;
        RECT 253.4400 2537.6400 255.0400 2538.1200 ;
        RECT 253.4400 2543.0800 255.0400 2543.5600 ;
        RECT 241.6800 2543.0800 244.6800 2543.5600 ;
        RECT 241.6800 2537.6400 244.6800 2538.1200 ;
        RECT 241.6800 2548.5200 244.6800 2549.0000 ;
        RECT 253.4400 2548.5200 255.0400 2549.0000 ;
        RECT 343.4400 2521.3200 345.0400 2521.8000 ;
        RECT 343.4400 2526.7600 345.0400 2527.2400 ;
        RECT 343.4400 2532.2000 345.0400 2532.6800 ;
        RECT 343.4400 2510.4400 345.0400 2510.9200 ;
        RECT 343.4400 2515.8800 345.0400 2516.3600 ;
        RECT 298.4400 2521.3200 300.0400 2521.8000 ;
        RECT 298.4400 2526.7600 300.0400 2527.2400 ;
        RECT 298.4400 2532.2000 300.0400 2532.6800 ;
        RECT 298.4400 2510.4400 300.0400 2510.9200 ;
        RECT 298.4400 2515.8800 300.0400 2516.3600 ;
        RECT 343.4400 2494.1200 345.0400 2494.6000 ;
        RECT 343.4400 2499.5600 345.0400 2500.0400 ;
        RECT 343.4400 2505.0000 345.0400 2505.4800 ;
        RECT 343.4400 2483.2400 345.0400 2483.7200 ;
        RECT 343.4400 2488.6800 345.0400 2489.1600 ;
        RECT 298.4400 2494.1200 300.0400 2494.6000 ;
        RECT 298.4400 2499.5600 300.0400 2500.0400 ;
        RECT 298.4400 2505.0000 300.0400 2505.4800 ;
        RECT 298.4400 2483.2400 300.0400 2483.7200 ;
        RECT 298.4400 2488.6800 300.0400 2489.1600 ;
        RECT 253.4400 2521.3200 255.0400 2521.8000 ;
        RECT 253.4400 2526.7600 255.0400 2527.2400 ;
        RECT 253.4400 2532.2000 255.0400 2532.6800 ;
        RECT 241.6800 2521.3200 244.6800 2521.8000 ;
        RECT 241.6800 2526.7600 244.6800 2527.2400 ;
        RECT 241.6800 2532.2000 244.6800 2532.6800 ;
        RECT 253.4400 2510.4400 255.0400 2510.9200 ;
        RECT 253.4400 2515.8800 255.0400 2516.3600 ;
        RECT 241.6800 2510.4400 244.6800 2510.9200 ;
        RECT 241.6800 2515.8800 244.6800 2516.3600 ;
        RECT 253.4400 2494.1200 255.0400 2494.6000 ;
        RECT 253.4400 2499.5600 255.0400 2500.0400 ;
        RECT 253.4400 2505.0000 255.0400 2505.4800 ;
        RECT 241.6800 2494.1200 244.6800 2494.6000 ;
        RECT 241.6800 2499.5600 244.6800 2500.0400 ;
        RECT 241.6800 2505.0000 244.6800 2505.4800 ;
        RECT 253.4400 2483.2400 255.0400 2483.7200 ;
        RECT 253.4400 2488.6800 255.0400 2489.1600 ;
        RECT 241.6800 2483.2400 244.6800 2483.7200 ;
        RECT 241.6800 2488.6800 244.6800 2489.1600 ;
        RECT 445.7800 2466.9200 448.7800 2467.4000 ;
        RECT 445.7800 2472.3600 448.7800 2472.8400 ;
        RECT 445.7800 2477.8000 448.7800 2478.2800 ;
        RECT 433.4400 2466.9200 435.0400 2467.4000 ;
        RECT 433.4400 2472.3600 435.0400 2472.8400 ;
        RECT 433.4400 2477.8000 435.0400 2478.2800 ;
        RECT 445.7800 2456.0400 448.7800 2456.5200 ;
        RECT 445.7800 2461.4800 448.7800 2461.9600 ;
        RECT 433.4400 2456.0400 435.0400 2456.5200 ;
        RECT 433.4400 2461.4800 435.0400 2461.9600 ;
        RECT 445.7800 2439.7200 448.7800 2440.2000 ;
        RECT 445.7800 2445.1600 448.7800 2445.6400 ;
        RECT 445.7800 2450.6000 448.7800 2451.0800 ;
        RECT 433.4400 2439.7200 435.0400 2440.2000 ;
        RECT 433.4400 2445.1600 435.0400 2445.6400 ;
        RECT 433.4400 2450.6000 435.0400 2451.0800 ;
        RECT 445.7800 2428.8400 448.7800 2429.3200 ;
        RECT 445.7800 2434.2800 448.7800 2434.7600 ;
        RECT 433.4400 2428.8400 435.0400 2429.3200 ;
        RECT 433.4400 2434.2800 435.0400 2434.7600 ;
        RECT 388.4400 2466.9200 390.0400 2467.4000 ;
        RECT 388.4400 2472.3600 390.0400 2472.8400 ;
        RECT 388.4400 2477.8000 390.0400 2478.2800 ;
        RECT 388.4400 2456.0400 390.0400 2456.5200 ;
        RECT 388.4400 2461.4800 390.0400 2461.9600 ;
        RECT 388.4400 2439.7200 390.0400 2440.2000 ;
        RECT 388.4400 2445.1600 390.0400 2445.6400 ;
        RECT 388.4400 2450.6000 390.0400 2451.0800 ;
        RECT 388.4400 2428.8400 390.0400 2429.3200 ;
        RECT 388.4400 2434.2800 390.0400 2434.7600 ;
        RECT 445.7800 2412.5200 448.7800 2413.0000 ;
        RECT 445.7800 2417.9600 448.7800 2418.4400 ;
        RECT 445.7800 2423.4000 448.7800 2423.8800 ;
        RECT 433.4400 2412.5200 435.0400 2413.0000 ;
        RECT 433.4400 2417.9600 435.0400 2418.4400 ;
        RECT 433.4400 2423.4000 435.0400 2423.8800 ;
        RECT 445.7800 2401.6400 448.7800 2402.1200 ;
        RECT 445.7800 2407.0800 448.7800 2407.5600 ;
        RECT 433.4400 2401.6400 435.0400 2402.1200 ;
        RECT 433.4400 2407.0800 435.0400 2407.5600 ;
        RECT 445.7800 2385.3200 448.7800 2385.8000 ;
        RECT 445.7800 2390.7600 448.7800 2391.2400 ;
        RECT 445.7800 2396.2000 448.7800 2396.6800 ;
        RECT 433.4400 2385.3200 435.0400 2385.8000 ;
        RECT 433.4400 2390.7600 435.0400 2391.2400 ;
        RECT 433.4400 2396.2000 435.0400 2396.6800 ;
        RECT 445.7800 2379.8800 448.7800 2380.3600 ;
        RECT 433.4400 2379.8800 435.0400 2380.3600 ;
        RECT 388.4400 2412.5200 390.0400 2413.0000 ;
        RECT 388.4400 2417.9600 390.0400 2418.4400 ;
        RECT 388.4400 2423.4000 390.0400 2423.8800 ;
        RECT 388.4400 2401.6400 390.0400 2402.1200 ;
        RECT 388.4400 2407.0800 390.0400 2407.5600 ;
        RECT 388.4400 2385.3200 390.0400 2385.8000 ;
        RECT 388.4400 2390.7600 390.0400 2391.2400 ;
        RECT 388.4400 2396.2000 390.0400 2396.6800 ;
        RECT 388.4400 2379.8800 390.0400 2380.3600 ;
        RECT 343.4400 2466.9200 345.0400 2467.4000 ;
        RECT 343.4400 2472.3600 345.0400 2472.8400 ;
        RECT 343.4400 2477.8000 345.0400 2478.2800 ;
        RECT 343.4400 2456.0400 345.0400 2456.5200 ;
        RECT 343.4400 2461.4800 345.0400 2461.9600 ;
        RECT 298.4400 2466.9200 300.0400 2467.4000 ;
        RECT 298.4400 2472.3600 300.0400 2472.8400 ;
        RECT 298.4400 2477.8000 300.0400 2478.2800 ;
        RECT 298.4400 2456.0400 300.0400 2456.5200 ;
        RECT 298.4400 2461.4800 300.0400 2461.9600 ;
        RECT 343.4400 2439.7200 345.0400 2440.2000 ;
        RECT 343.4400 2445.1600 345.0400 2445.6400 ;
        RECT 343.4400 2450.6000 345.0400 2451.0800 ;
        RECT 343.4400 2428.8400 345.0400 2429.3200 ;
        RECT 343.4400 2434.2800 345.0400 2434.7600 ;
        RECT 298.4400 2439.7200 300.0400 2440.2000 ;
        RECT 298.4400 2445.1600 300.0400 2445.6400 ;
        RECT 298.4400 2450.6000 300.0400 2451.0800 ;
        RECT 298.4400 2428.8400 300.0400 2429.3200 ;
        RECT 298.4400 2434.2800 300.0400 2434.7600 ;
        RECT 253.4400 2466.9200 255.0400 2467.4000 ;
        RECT 253.4400 2472.3600 255.0400 2472.8400 ;
        RECT 253.4400 2477.8000 255.0400 2478.2800 ;
        RECT 241.6800 2466.9200 244.6800 2467.4000 ;
        RECT 241.6800 2472.3600 244.6800 2472.8400 ;
        RECT 241.6800 2477.8000 244.6800 2478.2800 ;
        RECT 253.4400 2456.0400 255.0400 2456.5200 ;
        RECT 253.4400 2461.4800 255.0400 2461.9600 ;
        RECT 241.6800 2456.0400 244.6800 2456.5200 ;
        RECT 241.6800 2461.4800 244.6800 2461.9600 ;
        RECT 253.4400 2439.7200 255.0400 2440.2000 ;
        RECT 253.4400 2445.1600 255.0400 2445.6400 ;
        RECT 253.4400 2450.6000 255.0400 2451.0800 ;
        RECT 241.6800 2439.7200 244.6800 2440.2000 ;
        RECT 241.6800 2445.1600 244.6800 2445.6400 ;
        RECT 241.6800 2450.6000 244.6800 2451.0800 ;
        RECT 253.4400 2428.8400 255.0400 2429.3200 ;
        RECT 253.4400 2434.2800 255.0400 2434.7600 ;
        RECT 241.6800 2428.8400 244.6800 2429.3200 ;
        RECT 241.6800 2434.2800 244.6800 2434.7600 ;
        RECT 343.4400 2412.5200 345.0400 2413.0000 ;
        RECT 343.4400 2417.9600 345.0400 2418.4400 ;
        RECT 343.4400 2423.4000 345.0400 2423.8800 ;
        RECT 343.4400 2401.6400 345.0400 2402.1200 ;
        RECT 343.4400 2407.0800 345.0400 2407.5600 ;
        RECT 298.4400 2412.5200 300.0400 2413.0000 ;
        RECT 298.4400 2417.9600 300.0400 2418.4400 ;
        RECT 298.4400 2423.4000 300.0400 2423.8800 ;
        RECT 298.4400 2401.6400 300.0400 2402.1200 ;
        RECT 298.4400 2407.0800 300.0400 2407.5600 ;
        RECT 343.4400 2385.3200 345.0400 2385.8000 ;
        RECT 343.4400 2390.7600 345.0400 2391.2400 ;
        RECT 343.4400 2396.2000 345.0400 2396.6800 ;
        RECT 343.4400 2379.8800 345.0400 2380.3600 ;
        RECT 298.4400 2385.3200 300.0400 2385.8000 ;
        RECT 298.4400 2390.7600 300.0400 2391.2400 ;
        RECT 298.4400 2396.2000 300.0400 2396.6800 ;
        RECT 298.4400 2379.8800 300.0400 2380.3600 ;
        RECT 253.4400 2412.5200 255.0400 2413.0000 ;
        RECT 253.4400 2417.9600 255.0400 2418.4400 ;
        RECT 253.4400 2423.4000 255.0400 2423.8800 ;
        RECT 241.6800 2412.5200 244.6800 2413.0000 ;
        RECT 241.6800 2417.9600 244.6800 2418.4400 ;
        RECT 241.6800 2423.4000 244.6800 2423.8800 ;
        RECT 253.4400 2401.6400 255.0400 2402.1200 ;
        RECT 253.4400 2407.0800 255.0400 2407.5600 ;
        RECT 241.6800 2401.6400 244.6800 2402.1200 ;
        RECT 241.6800 2407.0800 244.6800 2407.5600 ;
        RECT 253.4400 2385.3200 255.0400 2385.8000 ;
        RECT 253.4400 2390.7600 255.0400 2391.2400 ;
        RECT 253.4400 2396.2000 255.0400 2396.6800 ;
        RECT 241.6800 2385.3200 244.6800 2385.8000 ;
        RECT 241.6800 2390.7600 244.6800 2391.2400 ;
        RECT 241.6800 2396.2000 244.6800 2396.6800 ;
        RECT 241.6800 2379.8800 244.6800 2380.3600 ;
        RECT 253.4400 2379.8800 255.0400 2380.3600 ;
        RECT 241.6800 2584.7900 448.7800 2587.7900 ;
        RECT 241.6800 2371.6900 448.7800 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 2142.0500 435.0400 2358.1500 ;
        RECT 388.4400 2142.0500 390.0400 2358.1500 ;
        RECT 343.4400 2142.0500 345.0400 2358.1500 ;
        RECT 298.4400 2142.0500 300.0400 2358.1500 ;
        RECT 253.4400 2142.0500 255.0400 2358.1500 ;
        RECT 445.7800 2142.0500 448.7800 2358.1500 ;
        RECT 241.6800 2142.0500 244.6800 2358.1500 ;
      LAYER met3 ;
        RECT 445.7800 2335.2000 448.7800 2335.6800 ;
        RECT 445.7800 2340.6400 448.7800 2341.1200 ;
        RECT 433.4400 2335.2000 435.0400 2335.6800 ;
        RECT 433.4400 2340.6400 435.0400 2341.1200 ;
        RECT 445.7800 2346.0800 448.7800 2346.5600 ;
        RECT 433.4400 2346.0800 435.0400 2346.5600 ;
        RECT 445.7800 2324.3200 448.7800 2324.8000 ;
        RECT 445.7800 2329.7600 448.7800 2330.2400 ;
        RECT 433.4400 2324.3200 435.0400 2324.8000 ;
        RECT 433.4400 2329.7600 435.0400 2330.2400 ;
        RECT 445.7800 2308.0000 448.7800 2308.4800 ;
        RECT 445.7800 2313.4400 448.7800 2313.9200 ;
        RECT 433.4400 2308.0000 435.0400 2308.4800 ;
        RECT 433.4400 2313.4400 435.0400 2313.9200 ;
        RECT 445.7800 2318.8800 448.7800 2319.3600 ;
        RECT 433.4400 2318.8800 435.0400 2319.3600 ;
        RECT 388.4400 2335.2000 390.0400 2335.6800 ;
        RECT 388.4400 2340.6400 390.0400 2341.1200 ;
        RECT 388.4400 2346.0800 390.0400 2346.5600 ;
        RECT 388.4400 2324.3200 390.0400 2324.8000 ;
        RECT 388.4400 2329.7600 390.0400 2330.2400 ;
        RECT 388.4400 2308.0000 390.0400 2308.4800 ;
        RECT 388.4400 2313.4400 390.0400 2313.9200 ;
        RECT 388.4400 2318.8800 390.0400 2319.3600 ;
        RECT 445.7800 2291.6800 448.7800 2292.1600 ;
        RECT 445.7800 2297.1200 448.7800 2297.6000 ;
        RECT 445.7800 2302.5600 448.7800 2303.0400 ;
        RECT 433.4400 2291.6800 435.0400 2292.1600 ;
        RECT 433.4400 2297.1200 435.0400 2297.6000 ;
        RECT 433.4400 2302.5600 435.0400 2303.0400 ;
        RECT 445.7800 2280.8000 448.7800 2281.2800 ;
        RECT 445.7800 2286.2400 448.7800 2286.7200 ;
        RECT 433.4400 2280.8000 435.0400 2281.2800 ;
        RECT 433.4400 2286.2400 435.0400 2286.7200 ;
        RECT 445.7800 2264.4800 448.7800 2264.9600 ;
        RECT 445.7800 2269.9200 448.7800 2270.4000 ;
        RECT 445.7800 2275.3600 448.7800 2275.8400 ;
        RECT 433.4400 2264.4800 435.0400 2264.9600 ;
        RECT 433.4400 2269.9200 435.0400 2270.4000 ;
        RECT 433.4400 2275.3600 435.0400 2275.8400 ;
        RECT 445.7800 2253.6000 448.7800 2254.0800 ;
        RECT 445.7800 2259.0400 448.7800 2259.5200 ;
        RECT 433.4400 2253.6000 435.0400 2254.0800 ;
        RECT 433.4400 2259.0400 435.0400 2259.5200 ;
        RECT 388.4400 2291.6800 390.0400 2292.1600 ;
        RECT 388.4400 2297.1200 390.0400 2297.6000 ;
        RECT 388.4400 2302.5600 390.0400 2303.0400 ;
        RECT 388.4400 2280.8000 390.0400 2281.2800 ;
        RECT 388.4400 2286.2400 390.0400 2286.7200 ;
        RECT 388.4400 2264.4800 390.0400 2264.9600 ;
        RECT 388.4400 2269.9200 390.0400 2270.4000 ;
        RECT 388.4400 2275.3600 390.0400 2275.8400 ;
        RECT 388.4400 2253.6000 390.0400 2254.0800 ;
        RECT 388.4400 2259.0400 390.0400 2259.5200 ;
        RECT 343.4400 2335.2000 345.0400 2335.6800 ;
        RECT 343.4400 2340.6400 345.0400 2341.1200 ;
        RECT 343.4400 2346.0800 345.0400 2346.5600 ;
        RECT 298.4400 2335.2000 300.0400 2335.6800 ;
        RECT 298.4400 2340.6400 300.0400 2341.1200 ;
        RECT 298.4400 2346.0800 300.0400 2346.5600 ;
        RECT 343.4400 2324.3200 345.0400 2324.8000 ;
        RECT 343.4400 2329.7600 345.0400 2330.2400 ;
        RECT 343.4400 2308.0000 345.0400 2308.4800 ;
        RECT 343.4400 2313.4400 345.0400 2313.9200 ;
        RECT 343.4400 2318.8800 345.0400 2319.3600 ;
        RECT 298.4400 2324.3200 300.0400 2324.8000 ;
        RECT 298.4400 2329.7600 300.0400 2330.2400 ;
        RECT 298.4400 2308.0000 300.0400 2308.4800 ;
        RECT 298.4400 2313.4400 300.0400 2313.9200 ;
        RECT 298.4400 2318.8800 300.0400 2319.3600 ;
        RECT 253.4400 2335.2000 255.0400 2335.6800 ;
        RECT 253.4400 2340.6400 255.0400 2341.1200 ;
        RECT 241.6800 2340.6400 244.6800 2341.1200 ;
        RECT 241.6800 2335.2000 244.6800 2335.6800 ;
        RECT 241.6800 2346.0800 244.6800 2346.5600 ;
        RECT 253.4400 2346.0800 255.0400 2346.5600 ;
        RECT 253.4400 2324.3200 255.0400 2324.8000 ;
        RECT 253.4400 2329.7600 255.0400 2330.2400 ;
        RECT 241.6800 2329.7600 244.6800 2330.2400 ;
        RECT 241.6800 2324.3200 244.6800 2324.8000 ;
        RECT 253.4400 2308.0000 255.0400 2308.4800 ;
        RECT 253.4400 2313.4400 255.0400 2313.9200 ;
        RECT 241.6800 2313.4400 244.6800 2313.9200 ;
        RECT 241.6800 2308.0000 244.6800 2308.4800 ;
        RECT 241.6800 2318.8800 244.6800 2319.3600 ;
        RECT 253.4400 2318.8800 255.0400 2319.3600 ;
        RECT 343.4400 2291.6800 345.0400 2292.1600 ;
        RECT 343.4400 2297.1200 345.0400 2297.6000 ;
        RECT 343.4400 2302.5600 345.0400 2303.0400 ;
        RECT 343.4400 2280.8000 345.0400 2281.2800 ;
        RECT 343.4400 2286.2400 345.0400 2286.7200 ;
        RECT 298.4400 2291.6800 300.0400 2292.1600 ;
        RECT 298.4400 2297.1200 300.0400 2297.6000 ;
        RECT 298.4400 2302.5600 300.0400 2303.0400 ;
        RECT 298.4400 2280.8000 300.0400 2281.2800 ;
        RECT 298.4400 2286.2400 300.0400 2286.7200 ;
        RECT 343.4400 2264.4800 345.0400 2264.9600 ;
        RECT 343.4400 2269.9200 345.0400 2270.4000 ;
        RECT 343.4400 2275.3600 345.0400 2275.8400 ;
        RECT 343.4400 2253.6000 345.0400 2254.0800 ;
        RECT 343.4400 2259.0400 345.0400 2259.5200 ;
        RECT 298.4400 2264.4800 300.0400 2264.9600 ;
        RECT 298.4400 2269.9200 300.0400 2270.4000 ;
        RECT 298.4400 2275.3600 300.0400 2275.8400 ;
        RECT 298.4400 2253.6000 300.0400 2254.0800 ;
        RECT 298.4400 2259.0400 300.0400 2259.5200 ;
        RECT 253.4400 2291.6800 255.0400 2292.1600 ;
        RECT 253.4400 2297.1200 255.0400 2297.6000 ;
        RECT 253.4400 2302.5600 255.0400 2303.0400 ;
        RECT 241.6800 2291.6800 244.6800 2292.1600 ;
        RECT 241.6800 2297.1200 244.6800 2297.6000 ;
        RECT 241.6800 2302.5600 244.6800 2303.0400 ;
        RECT 253.4400 2280.8000 255.0400 2281.2800 ;
        RECT 253.4400 2286.2400 255.0400 2286.7200 ;
        RECT 241.6800 2280.8000 244.6800 2281.2800 ;
        RECT 241.6800 2286.2400 244.6800 2286.7200 ;
        RECT 253.4400 2264.4800 255.0400 2264.9600 ;
        RECT 253.4400 2269.9200 255.0400 2270.4000 ;
        RECT 253.4400 2275.3600 255.0400 2275.8400 ;
        RECT 241.6800 2264.4800 244.6800 2264.9600 ;
        RECT 241.6800 2269.9200 244.6800 2270.4000 ;
        RECT 241.6800 2275.3600 244.6800 2275.8400 ;
        RECT 253.4400 2253.6000 255.0400 2254.0800 ;
        RECT 253.4400 2259.0400 255.0400 2259.5200 ;
        RECT 241.6800 2253.6000 244.6800 2254.0800 ;
        RECT 241.6800 2259.0400 244.6800 2259.5200 ;
        RECT 445.7800 2237.2800 448.7800 2237.7600 ;
        RECT 445.7800 2242.7200 448.7800 2243.2000 ;
        RECT 445.7800 2248.1600 448.7800 2248.6400 ;
        RECT 433.4400 2237.2800 435.0400 2237.7600 ;
        RECT 433.4400 2242.7200 435.0400 2243.2000 ;
        RECT 433.4400 2248.1600 435.0400 2248.6400 ;
        RECT 445.7800 2226.4000 448.7800 2226.8800 ;
        RECT 445.7800 2231.8400 448.7800 2232.3200 ;
        RECT 433.4400 2226.4000 435.0400 2226.8800 ;
        RECT 433.4400 2231.8400 435.0400 2232.3200 ;
        RECT 445.7800 2210.0800 448.7800 2210.5600 ;
        RECT 445.7800 2215.5200 448.7800 2216.0000 ;
        RECT 445.7800 2220.9600 448.7800 2221.4400 ;
        RECT 433.4400 2210.0800 435.0400 2210.5600 ;
        RECT 433.4400 2215.5200 435.0400 2216.0000 ;
        RECT 433.4400 2220.9600 435.0400 2221.4400 ;
        RECT 445.7800 2199.2000 448.7800 2199.6800 ;
        RECT 445.7800 2204.6400 448.7800 2205.1200 ;
        RECT 433.4400 2199.2000 435.0400 2199.6800 ;
        RECT 433.4400 2204.6400 435.0400 2205.1200 ;
        RECT 388.4400 2237.2800 390.0400 2237.7600 ;
        RECT 388.4400 2242.7200 390.0400 2243.2000 ;
        RECT 388.4400 2248.1600 390.0400 2248.6400 ;
        RECT 388.4400 2226.4000 390.0400 2226.8800 ;
        RECT 388.4400 2231.8400 390.0400 2232.3200 ;
        RECT 388.4400 2210.0800 390.0400 2210.5600 ;
        RECT 388.4400 2215.5200 390.0400 2216.0000 ;
        RECT 388.4400 2220.9600 390.0400 2221.4400 ;
        RECT 388.4400 2199.2000 390.0400 2199.6800 ;
        RECT 388.4400 2204.6400 390.0400 2205.1200 ;
        RECT 445.7800 2182.8800 448.7800 2183.3600 ;
        RECT 445.7800 2188.3200 448.7800 2188.8000 ;
        RECT 445.7800 2193.7600 448.7800 2194.2400 ;
        RECT 433.4400 2182.8800 435.0400 2183.3600 ;
        RECT 433.4400 2188.3200 435.0400 2188.8000 ;
        RECT 433.4400 2193.7600 435.0400 2194.2400 ;
        RECT 445.7800 2172.0000 448.7800 2172.4800 ;
        RECT 445.7800 2177.4400 448.7800 2177.9200 ;
        RECT 433.4400 2172.0000 435.0400 2172.4800 ;
        RECT 433.4400 2177.4400 435.0400 2177.9200 ;
        RECT 445.7800 2155.6800 448.7800 2156.1600 ;
        RECT 445.7800 2161.1200 448.7800 2161.6000 ;
        RECT 445.7800 2166.5600 448.7800 2167.0400 ;
        RECT 433.4400 2155.6800 435.0400 2156.1600 ;
        RECT 433.4400 2161.1200 435.0400 2161.6000 ;
        RECT 433.4400 2166.5600 435.0400 2167.0400 ;
        RECT 445.7800 2150.2400 448.7800 2150.7200 ;
        RECT 433.4400 2150.2400 435.0400 2150.7200 ;
        RECT 388.4400 2182.8800 390.0400 2183.3600 ;
        RECT 388.4400 2188.3200 390.0400 2188.8000 ;
        RECT 388.4400 2193.7600 390.0400 2194.2400 ;
        RECT 388.4400 2172.0000 390.0400 2172.4800 ;
        RECT 388.4400 2177.4400 390.0400 2177.9200 ;
        RECT 388.4400 2155.6800 390.0400 2156.1600 ;
        RECT 388.4400 2161.1200 390.0400 2161.6000 ;
        RECT 388.4400 2166.5600 390.0400 2167.0400 ;
        RECT 388.4400 2150.2400 390.0400 2150.7200 ;
        RECT 343.4400 2237.2800 345.0400 2237.7600 ;
        RECT 343.4400 2242.7200 345.0400 2243.2000 ;
        RECT 343.4400 2248.1600 345.0400 2248.6400 ;
        RECT 343.4400 2226.4000 345.0400 2226.8800 ;
        RECT 343.4400 2231.8400 345.0400 2232.3200 ;
        RECT 298.4400 2237.2800 300.0400 2237.7600 ;
        RECT 298.4400 2242.7200 300.0400 2243.2000 ;
        RECT 298.4400 2248.1600 300.0400 2248.6400 ;
        RECT 298.4400 2226.4000 300.0400 2226.8800 ;
        RECT 298.4400 2231.8400 300.0400 2232.3200 ;
        RECT 343.4400 2210.0800 345.0400 2210.5600 ;
        RECT 343.4400 2215.5200 345.0400 2216.0000 ;
        RECT 343.4400 2220.9600 345.0400 2221.4400 ;
        RECT 343.4400 2199.2000 345.0400 2199.6800 ;
        RECT 343.4400 2204.6400 345.0400 2205.1200 ;
        RECT 298.4400 2210.0800 300.0400 2210.5600 ;
        RECT 298.4400 2215.5200 300.0400 2216.0000 ;
        RECT 298.4400 2220.9600 300.0400 2221.4400 ;
        RECT 298.4400 2199.2000 300.0400 2199.6800 ;
        RECT 298.4400 2204.6400 300.0400 2205.1200 ;
        RECT 253.4400 2237.2800 255.0400 2237.7600 ;
        RECT 253.4400 2242.7200 255.0400 2243.2000 ;
        RECT 253.4400 2248.1600 255.0400 2248.6400 ;
        RECT 241.6800 2237.2800 244.6800 2237.7600 ;
        RECT 241.6800 2242.7200 244.6800 2243.2000 ;
        RECT 241.6800 2248.1600 244.6800 2248.6400 ;
        RECT 253.4400 2226.4000 255.0400 2226.8800 ;
        RECT 253.4400 2231.8400 255.0400 2232.3200 ;
        RECT 241.6800 2226.4000 244.6800 2226.8800 ;
        RECT 241.6800 2231.8400 244.6800 2232.3200 ;
        RECT 253.4400 2210.0800 255.0400 2210.5600 ;
        RECT 253.4400 2215.5200 255.0400 2216.0000 ;
        RECT 253.4400 2220.9600 255.0400 2221.4400 ;
        RECT 241.6800 2210.0800 244.6800 2210.5600 ;
        RECT 241.6800 2215.5200 244.6800 2216.0000 ;
        RECT 241.6800 2220.9600 244.6800 2221.4400 ;
        RECT 253.4400 2199.2000 255.0400 2199.6800 ;
        RECT 253.4400 2204.6400 255.0400 2205.1200 ;
        RECT 241.6800 2199.2000 244.6800 2199.6800 ;
        RECT 241.6800 2204.6400 244.6800 2205.1200 ;
        RECT 343.4400 2182.8800 345.0400 2183.3600 ;
        RECT 343.4400 2188.3200 345.0400 2188.8000 ;
        RECT 343.4400 2193.7600 345.0400 2194.2400 ;
        RECT 343.4400 2172.0000 345.0400 2172.4800 ;
        RECT 343.4400 2177.4400 345.0400 2177.9200 ;
        RECT 298.4400 2182.8800 300.0400 2183.3600 ;
        RECT 298.4400 2188.3200 300.0400 2188.8000 ;
        RECT 298.4400 2193.7600 300.0400 2194.2400 ;
        RECT 298.4400 2172.0000 300.0400 2172.4800 ;
        RECT 298.4400 2177.4400 300.0400 2177.9200 ;
        RECT 343.4400 2155.6800 345.0400 2156.1600 ;
        RECT 343.4400 2161.1200 345.0400 2161.6000 ;
        RECT 343.4400 2166.5600 345.0400 2167.0400 ;
        RECT 343.4400 2150.2400 345.0400 2150.7200 ;
        RECT 298.4400 2155.6800 300.0400 2156.1600 ;
        RECT 298.4400 2161.1200 300.0400 2161.6000 ;
        RECT 298.4400 2166.5600 300.0400 2167.0400 ;
        RECT 298.4400 2150.2400 300.0400 2150.7200 ;
        RECT 253.4400 2182.8800 255.0400 2183.3600 ;
        RECT 253.4400 2188.3200 255.0400 2188.8000 ;
        RECT 253.4400 2193.7600 255.0400 2194.2400 ;
        RECT 241.6800 2182.8800 244.6800 2183.3600 ;
        RECT 241.6800 2188.3200 244.6800 2188.8000 ;
        RECT 241.6800 2193.7600 244.6800 2194.2400 ;
        RECT 253.4400 2172.0000 255.0400 2172.4800 ;
        RECT 253.4400 2177.4400 255.0400 2177.9200 ;
        RECT 241.6800 2172.0000 244.6800 2172.4800 ;
        RECT 241.6800 2177.4400 244.6800 2177.9200 ;
        RECT 253.4400 2155.6800 255.0400 2156.1600 ;
        RECT 253.4400 2161.1200 255.0400 2161.6000 ;
        RECT 253.4400 2166.5600 255.0400 2167.0400 ;
        RECT 241.6800 2155.6800 244.6800 2156.1600 ;
        RECT 241.6800 2161.1200 244.6800 2161.6000 ;
        RECT 241.6800 2166.5600 244.6800 2167.0400 ;
        RECT 241.6800 2150.2400 244.6800 2150.7200 ;
        RECT 253.4400 2150.2400 255.0400 2150.7200 ;
        RECT 241.6800 2355.1500 448.7800 2358.1500 ;
        RECT 241.6800 2142.0500 448.7800 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 1912.4100 435.0400 2128.5100 ;
        RECT 388.4400 1912.4100 390.0400 2128.5100 ;
        RECT 343.4400 1912.4100 345.0400 2128.5100 ;
        RECT 298.4400 1912.4100 300.0400 2128.5100 ;
        RECT 253.4400 1912.4100 255.0400 2128.5100 ;
        RECT 445.7800 1912.4100 448.7800 2128.5100 ;
        RECT 241.6800 1912.4100 244.6800 2128.5100 ;
      LAYER met3 ;
        RECT 445.7800 2105.5600 448.7800 2106.0400 ;
        RECT 445.7800 2111.0000 448.7800 2111.4800 ;
        RECT 433.4400 2105.5600 435.0400 2106.0400 ;
        RECT 433.4400 2111.0000 435.0400 2111.4800 ;
        RECT 445.7800 2116.4400 448.7800 2116.9200 ;
        RECT 433.4400 2116.4400 435.0400 2116.9200 ;
        RECT 445.7800 2094.6800 448.7800 2095.1600 ;
        RECT 445.7800 2100.1200 448.7800 2100.6000 ;
        RECT 433.4400 2094.6800 435.0400 2095.1600 ;
        RECT 433.4400 2100.1200 435.0400 2100.6000 ;
        RECT 445.7800 2078.3600 448.7800 2078.8400 ;
        RECT 445.7800 2083.8000 448.7800 2084.2800 ;
        RECT 433.4400 2078.3600 435.0400 2078.8400 ;
        RECT 433.4400 2083.8000 435.0400 2084.2800 ;
        RECT 445.7800 2089.2400 448.7800 2089.7200 ;
        RECT 433.4400 2089.2400 435.0400 2089.7200 ;
        RECT 388.4400 2105.5600 390.0400 2106.0400 ;
        RECT 388.4400 2111.0000 390.0400 2111.4800 ;
        RECT 388.4400 2116.4400 390.0400 2116.9200 ;
        RECT 388.4400 2094.6800 390.0400 2095.1600 ;
        RECT 388.4400 2100.1200 390.0400 2100.6000 ;
        RECT 388.4400 2078.3600 390.0400 2078.8400 ;
        RECT 388.4400 2083.8000 390.0400 2084.2800 ;
        RECT 388.4400 2089.2400 390.0400 2089.7200 ;
        RECT 445.7800 2062.0400 448.7800 2062.5200 ;
        RECT 445.7800 2067.4800 448.7800 2067.9600 ;
        RECT 445.7800 2072.9200 448.7800 2073.4000 ;
        RECT 433.4400 2062.0400 435.0400 2062.5200 ;
        RECT 433.4400 2067.4800 435.0400 2067.9600 ;
        RECT 433.4400 2072.9200 435.0400 2073.4000 ;
        RECT 445.7800 2051.1600 448.7800 2051.6400 ;
        RECT 445.7800 2056.6000 448.7800 2057.0800 ;
        RECT 433.4400 2051.1600 435.0400 2051.6400 ;
        RECT 433.4400 2056.6000 435.0400 2057.0800 ;
        RECT 445.7800 2034.8400 448.7800 2035.3200 ;
        RECT 445.7800 2040.2800 448.7800 2040.7600 ;
        RECT 445.7800 2045.7200 448.7800 2046.2000 ;
        RECT 433.4400 2034.8400 435.0400 2035.3200 ;
        RECT 433.4400 2040.2800 435.0400 2040.7600 ;
        RECT 433.4400 2045.7200 435.0400 2046.2000 ;
        RECT 445.7800 2023.9600 448.7800 2024.4400 ;
        RECT 445.7800 2029.4000 448.7800 2029.8800 ;
        RECT 433.4400 2023.9600 435.0400 2024.4400 ;
        RECT 433.4400 2029.4000 435.0400 2029.8800 ;
        RECT 388.4400 2062.0400 390.0400 2062.5200 ;
        RECT 388.4400 2067.4800 390.0400 2067.9600 ;
        RECT 388.4400 2072.9200 390.0400 2073.4000 ;
        RECT 388.4400 2051.1600 390.0400 2051.6400 ;
        RECT 388.4400 2056.6000 390.0400 2057.0800 ;
        RECT 388.4400 2034.8400 390.0400 2035.3200 ;
        RECT 388.4400 2040.2800 390.0400 2040.7600 ;
        RECT 388.4400 2045.7200 390.0400 2046.2000 ;
        RECT 388.4400 2023.9600 390.0400 2024.4400 ;
        RECT 388.4400 2029.4000 390.0400 2029.8800 ;
        RECT 343.4400 2105.5600 345.0400 2106.0400 ;
        RECT 343.4400 2111.0000 345.0400 2111.4800 ;
        RECT 343.4400 2116.4400 345.0400 2116.9200 ;
        RECT 298.4400 2105.5600 300.0400 2106.0400 ;
        RECT 298.4400 2111.0000 300.0400 2111.4800 ;
        RECT 298.4400 2116.4400 300.0400 2116.9200 ;
        RECT 343.4400 2094.6800 345.0400 2095.1600 ;
        RECT 343.4400 2100.1200 345.0400 2100.6000 ;
        RECT 343.4400 2078.3600 345.0400 2078.8400 ;
        RECT 343.4400 2083.8000 345.0400 2084.2800 ;
        RECT 343.4400 2089.2400 345.0400 2089.7200 ;
        RECT 298.4400 2094.6800 300.0400 2095.1600 ;
        RECT 298.4400 2100.1200 300.0400 2100.6000 ;
        RECT 298.4400 2078.3600 300.0400 2078.8400 ;
        RECT 298.4400 2083.8000 300.0400 2084.2800 ;
        RECT 298.4400 2089.2400 300.0400 2089.7200 ;
        RECT 253.4400 2105.5600 255.0400 2106.0400 ;
        RECT 253.4400 2111.0000 255.0400 2111.4800 ;
        RECT 241.6800 2111.0000 244.6800 2111.4800 ;
        RECT 241.6800 2105.5600 244.6800 2106.0400 ;
        RECT 241.6800 2116.4400 244.6800 2116.9200 ;
        RECT 253.4400 2116.4400 255.0400 2116.9200 ;
        RECT 253.4400 2094.6800 255.0400 2095.1600 ;
        RECT 253.4400 2100.1200 255.0400 2100.6000 ;
        RECT 241.6800 2100.1200 244.6800 2100.6000 ;
        RECT 241.6800 2094.6800 244.6800 2095.1600 ;
        RECT 253.4400 2078.3600 255.0400 2078.8400 ;
        RECT 253.4400 2083.8000 255.0400 2084.2800 ;
        RECT 241.6800 2083.8000 244.6800 2084.2800 ;
        RECT 241.6800 2078.3600 244.6800 2078.8400 ;
        RECT 241.6800 2089.2400 244.6800 2089.7200 ;
        RECT 253.4400 2089.2400 255.0400 2089.7200 ;
        RECT 343.4400 2062.0400 345.0400 2062.5200 ;
        RECT 343.4400 2067.4800 345.0400 2067.9600 ;
        RECT 343.4400 2072.9200 345.0400 2073.4000 ;
        RECT 343.4400 2051.1600 345.0400 2051.6400 ;
        RECT 343.4400 2056.6000 345.0400 2057.0800 ;
        RECT 298.4400 2062.0400 300.0400 2062.5200 ;
        RECT 298.4400 2067.4800 300.0400 2067.9600 ;
        RECT 298.4400 2072.9200 300.0400 2073.4000 ;
        RECT 298.4400 2051.1600 300.0400 2051.6400 ;
        RECT 298.4400 2056.6000 300.0400 2057.0800 ;
        RECT 343.4400 2034.8400 345.0400 2035.3200 ;
        RECT 343.4400 2040.2800 345.0400 2040.7600 ;
        RECT 343.4400 2045.7200 345.0400 2046.2000 ;
        RECT 343.4400 2023.9600 345.0400 2024.4400 ;
        RECT 343.4400 2029.4000 345.0400 2029.8800 ;
        RECT 298.4400 2034.8400 300.0400 2035.3200 ;
        RECT 298.4400 2040.2800 300.0400 2040.7600 ;
        RECT 298.4400 2045.7200 300.0400 2046.2000 ;
        RECT 298.4400 2023.9600 300.0400 2024.4400 ;
        RECT 298.4400 2029.4000 300.0400 2029.8800 ;
        RECT 253.4400 2062.0400 255.0400 2062.5200 ;
        RECT 253.4400 2067.4800 255.0400 2067.9600 ;
        RECT 253.4400 2072.9200 255.0400 2073.4000 ;
        RECT 241.6800 2062.0400 244.6800 2062.5200 ;
        RECT 241.6800 2067.4800 244.6800 2067.9600 ;
        RECT 241.6800 2072.9200 244.6800 2073.4000 ;
        RECT 253.4400 2051.1600 255.0400 2051.6400 ;
        RECT 253.4400 2056.6000 255.0400 2057.0800 ;
        RECT 241.6800 2051.1600 244.6800 2051.6400 ;
        RECT 241.6800 2056.6000 244.6800 2057.0800 ;
        RECT 253.4400 2034.8400 255.0400 2035.3200 ;
        RECT 253.4400 2040.2800 255.0400 2040.7600 ;
        RECT 253.4400 2045.7200 255.0400 2046.2000 ;
        RECT 241.6800 2034.8400 244.6800 2035.3200 ;
        RECT 241.6800 2040.2800 244.6800 2040.7600 ;
        RECT 241.6800 2045.7200 244.6800 2046.2000 ;
        RECT 253.4400 2023.9600 255.0400 2024.4400 ;
        RECT 253.4400 2029.4000 255.0400 2029.8800 ;
        RECT 241.6800 2023.9600 244.6800 2024.4400 ;
        RECT 241.6800 2029.4000 244.6800 2029.8800 ;
        RECT 445.7800 2007.6400 448.7800 2008.1200 ;
        RECT 445.7800 2013.0800 448.7800 2013.5600 ;
        RECT 445.7800 2018.5200 448.7800 2019.0000 ;
        RECT 433.4400 2007.6400 435.0400 2008.1200 ;
        RECT 433.4400 2013.0800 435.0400 2013.5600 ;
        RECT 433.4400 2018.5200 435.0400 2019.0000 ;
        RECT 445.7800 1996.7600 448.7800 1997.2400 ;
        RECT 445.7800 2002.2000 448.7800 2002.6800 ;
        RECT 433.4400 1996.7600 435.0400 1997.2400 ;
        RECT 433.4400 2002.2000 435.0400 2002.6800 ;
        RECT 445.7800 1980.4400 448.7800 1980.9200 ;
        RECT 445.7800 1985.8800 448.7800 1986.3600 ;
        RECT 445.7800 1991.3200 448.7800 1991.8000 ;
        RECT 433.4400 1980.4400 435.0400 1980.9200 ;
        RECT 433.4400 1985.8800 435.0400 1986.3600 ;
        RECT 433.4400 1991.3200 435.0400 1991.8000 ;
        RECT 445.7800 1969.5600 448.7800 1970.0400 ;
        RECT 445.7800 1975.0000 448.7800 1975.4800 ;
        RECT 433.4400 1969.5600 435.0400 1970.0400 ;
        RECT 433.4400 1975.0000 435.0400 1975.4800 ;
        RECT 388.4400 2007.6400 390.0400 2008.1200 ;
        RECT 388.4400 2013.0800 390.0400 2013.5600 ;
        RECT 388.4400 2018.5200 390.0400 2019.0000 ;
        RECT 388.4400 1996.7600 390.0400 1997.2400 ;
        RECT 388.4400 2002.2000 390.0400 2002.6800 ;
        RECT 388.4400 1980.4400 390.0400 1980.9200 ;
        RECT 388.4400 1985.8800 390.0400 1986.3600 ;
        RECT 388.4400 1991.3200 390.0400 1991.8000 ;
        RECT 388.4400 1969.5600 390.0400 1970.0400 ;
        RECT 388.4400 1975.0000 390.0400 1975.4800 ;
        RECT 445.7800 1953.2400 448.7800 1953.7200 ;
        RECT 445.7800 1958.6800 448.7800 1959.1600 ;
        RECT 445.7800 1964.1200 448.7800 1964.6000 ;
        RECT 433.4400 1953.2400 435.0400 1953.7200 ;
        RECT 433.4400 1958.6800 435.0400 1959.1600 ;
        RECT 433.4400 1964.1200 435.0400 1964.6000 ;
        RECT 445.7800 1942.3600 448.7800 1942.8400 ;
        RECT 445.7800 1947.8000 448.7800 1948.2800 ;
        RECT 433.4400 1942.3600 435.0400 1942.8400 ;
        RECT 433.4400 1947.8000 435.0400 1948.2800 ;
        RECT 445.7800 1926.0400 448.7800 1926.5200 ;
        RECT 445.7800 1931.4800 448.7800 1931.9600 ;
        RECT 445.7800 1936.9200 448.7800 1937.4000 ;
        RECT 433.4400 1926.0400 435.0400 1926.5200 ;
        RECT 433.4400 1931.4800 435.0400 1931.9600 ;
        RECT 433.4400 1936.9200 435.0400 1937.4000 ;
        RECT 445.7800 1920.6000 448.7800 1921.0800 ;
        RECT 433.4400 1920.6000 435.0400 1921.0800 ;
        RECT 388.4400 1953.2400 390.0400 1953.7200 ;
        RECT 388.4400 1958.6800 390.0400 1959.1600 ;
        RECT 388.4400 1964.1200 390.0400 1964.6000 ;
        RECT 388.4400 1942.3600 390.0400 1942.8400 ;
        RECT 388.4400 1947.8000 390.0400 1948.2800 ;
        RECT 388.4400 1926.0400 390.0400 1926.5200 ;
        RECT 388.4400 1931.4800 390.0400 1931.9600 ;
        RECT 388.4400 1936.9200 390.0400 1937.4000 ;
        RECT 388.4400 1920.6000 390.0400 1921.0800 ;
        RECT 343.4400 2007.6400 345.0400 2008.1200 ;
        RECT 343.4400 2013.0800 345.0400 2013.5600 ;
        RECT 343.4400 2018.5200 345.0400 2019.0000 ;
        RECT 343.4400 1996.7600 345.0400 1997.2400 ;
        RECT 343.4400 2002.2000 345.0400 2002.6800 ;
        RECT 298.4400 2007.6400 300.0400 2008.1200 ;
        RECT 298.4400 2013.0800 300.0400 2013.5600 ;
        RECT 298.4400 2018.5200 300.0400 2019.0000 ;
        RECT 298.4400 1996.7600 300.0400 1997.2400 ;
        RECT 298.4400 2002.2000 300.0400 2002.6800 ;
        RECT 343.4400 1980.4400 345.0400 1980.9200 ;
        RECT 343.4400 1985.8800 345.0400 1986.3600 ;
        RECT 343.4400 1991.3200 345.0400 1991.8000 ;
        RECT 343.4400 1969.5600 345.0400 1970.0400 ;
        RECT 343.4400 1975.0000 345.0400 1975.4800 ;
        RECT 298.4400 1980.4400 300.0400 1980.9200 ;
        RECT 298.4400 1985.8800 300.0400 1986.3600 ;
        RECT 298.4400 1991.3200 300.0400 1991.8000 ;
        RECT 298.4400 1969.5600 300.0400 1970.0400 ;
        RECT 298.4400 1975.0000 300.0400 1975.4800 ;
        RECT 253.4400 2007.6400 255.0400 2008.1200 ;
        RECT 253.4400 2013.0800 255.0400 2013.5600 ;
        RECT 253.4400 2018.5200 255.0400 2019.0000 ;
        RECT 241.6800 2007.6400 244.6800 2008.1200 ;
        RECT 241.6800 2013.0800 244.6800 2013.5600 ;
        RECT 241.6800 2018.5200 244.6800 2019.0000 ;
        RECT 253.4400 1996.7600 255.0400 1997.2400 ;
        RECT 253.4400 2002.2000 255.0400 2002.6800 ;
        RECT 241.6800 1996.7600 244.6800 1997.2400 ;
        RECT 241.6800 2002.2000 244.6800 2002.6800 ;
        RECT 253.4400 1980.4400 255.0400 1980.9200 ;
        RECT 253.4400 1985.8800 255.0400 1986.3600 ;
        RECT 253.4400 1991.3200 255.0400 1991.8000 ;
        RECT 241.6800 1980.4400 244.6800 1980.9200 ;
        RECT 241.6800 1985.8800 244.6800 1986.3600 ;
        RECT 241.6800 1991.3200 244.6800 1991.8000 ;
        RECT 253.4400 1969.5600 255.0400 1970.0400 ;
        RECT 253.4400 1975.0000 255.0400 1975.4800 ;
        RECT 241.6800 1969.5600 244.6800 1970.0400 ;
        RECT 241.6800 1975.0000 244.6800 1975.4800 ;
        RECT 343.4400 1953.2400 345.0400 1953.7200 ;
        RECT 343.4400 1958.6800 345.0400 1959.1600 ;
        RECT 343.4400 1964.1200 345.0400 1964.6000 ;
        RECT 343.4400 1942.3600 345.0400 1942.8400 ;
        RECT 343.4400 1947.8000 345.0400 1948.2800 ;
        RECT 298.4400 1953.2400 300.0400 1953.7200 ;
        RECT 298.4400 1958.6800 300.0400 1959.1600 ;
        RECT 298.4400 1964.1200 300.0400 1964.6000 ;
        RECT 298.4400 1942.3600 300.0400 1942.8400 ;
        RECT 298.4400 1947.8000 300.0400 1948.2800 ;
        RECT 343.4400 1926.0400 345.0400 1926.5200 ;
        RECT 343.4400 1931.4800 345.0400 1931.9600 ;
        RECT 343.4400 1936.9200 345.0400 1937.4000 ;
        RECT 343.4400 1920.6000 345.0400 1921.0800 ;
        RECT 298.4400 1926.0400 300.0400 1926.5200 ;
        RECT 298.4400 1931.4800 300.0400 1931.9600 ;
        RECT 298.4400 1936.9200 300.0400 1937.4000 ;
        RECT 298.4400 1920.6000 300.0400 1921.0800 ;
        RECT 253.4400 1953.2400 255.0400 1953.7200 ;
        RECT 253.4400 1958.6800 255.0400 1959.1600 ;
        RECT 253.4400 1964.1200 255.0400 1964.6000 ;
        RECT 241.6800 1953.2400 244.6800 1953.7200 ;
        RECT 241.6800 1958.6800 244.6800 1959.1600 ;
        RECT 241.6800 1964.1200 244.6800 1964.6000 ;
        RECT 253.4400 1942.3600 255.0400 1942.8400 ;
        RECT 253.4400 1947.8000 255.0400 1948.2800 ;
        RECT 241.6800 1942.3600 244.6800 1942.8400 ;
        RECT 241.6800 1947.8000 244.6800 1948.2800 ;
        RECT 253.4400 1926.0400 255.0400 1926.5200 ;
        RECT 253.4400 1931.4800 255.0400 1931.9600 ;
        RECT 253.4400 1936.9200 255.0400 1937.4000 ;
        RECT 241.6800 1926.0400 244.6800 1926.5200 ;
        RECT 241.6800 1931.4800 244.6800 1931.9600 ;
        RECT 241.6800 1936.9200 244.6800 1937.4000 ;
        RECT 241.6800 1920.6000 244.6800 1921.0800 ;
        RECT 253.4400 1920.6000 255.0400 1921.0800 ;
        RECT 241.6800 2125.5100 448.7800 2128.5100 ;
        RECT 241.6800 1912.4100 448.7800 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 1682.7700 435.0400 1898.8700 ;
        RECT 388.4400 1682.7700 390.0400 1898.8700 ;
        RECT 343.4400 1682.7700 345.0400 1898.8700 ;
        RECT 298.4400 1682.7700 300.0400 1898.8700 ;
        RECT 253.4400 1682.7700 255.0400 1898.8700 ;
        RECT 445.7800 1682.7700 448.7800 1898.8700 ;
        RECT 241.6800 1682.7700 244.6800 1898.8700 ;
      LAYER met3 ;
        RECT 445.7800 1875.9200 448.7800 1876.4000 ;
        RECT 445.7800 1881.3600 448.7800 1881.8400 ;
        RECT 433.4400 1875.9200 435.0400 1876.4000 ;
        RECT 433.4400 1881.3600 435.0400 1881.8400 ;
        RECT 445.7800 1886.8000 448.7800 1887.2800 ;
        RECT 433.4400 1886.8000 435.0400 1887.2800 ;
        RECT 445.7800 1865.0400 448.7800 1865.5200 ;
        RECT 445.7800 1870.4800 448.7800 1870.9600 ;
        RECT 433.4400 1865.0400 435.0400 1865.5200 ;
        RECT 433.4400 1870.4800 435.0400 1870.9600 ;
        RECT 445.7800 1848.7200 448.7800 1849.2000 ;
        RECT 445.7800 1854.1600 448.7800 1854.6400 ;
        RECT 433.4400 1848.7200 435.0400 1849.2000 ;
        RECT 433.4400 1854.1600 435.0400 1854.6400 ;
        RECT 445.7800 1859.6000 448.7800 1860.0800 ;
        RECT 433.4400 1859.6000 435.0400 1860.0800 ;
        RECT 388.4400 1875.9200 390.0400 1876.4000 ;
        RECT 388.4400 1881.3600 390.0400 1881.8400 ;
        RECT 388.4400 1886.8000 390.0400 1887.2800 ;
        RECT 388.4400 1865.0400 390.0400 1865.5200 ;
        RECT 388.4400 1870.4800 390.0400 1870.9600 ;
        RECT 388.4400 1848.7200 390.0400 1849.2000 ;
        RECT 388.4400 1854.1600 390.0400 1854.6400 ;
        RECT 388.4400 1859.6000 390.0400 1860.0800 ;
        RECT 445.7800 1832.4000 448.7800 1832.8800 ;
        RECT 445.7800 1837.8400 448.7800 1838.3200 ;
        RECT 445.7800 1843.2800 448.7800 1843.7600 ;
        RECT 433.4400 1832.4000 435.0400 1832.8800 ;
        RECT 433.4400 1837.8400 435.0400 1838.3200 ;
        RECT 433.4400 1843.2800 435.0400 1843.7600 ;
        RECT 445.7800 1821.5200 448.7800 1822.0000 ;
        RECT 445.7800 1826.9600 448.7800 1827.4400 ;
        RECT 433.4400 1821.5200 435.0400 1822.0000 ;
        RECT 433.4400 1826.9600 435.0400 1827.4400 ;
        RECT 445.7800 1805.2000 448.7800 1805.6800 ;
        RECT 445.7800 1810.6400 448.7800 1811.1200 ;
        RECT 445.7800 1816.0800 448.7800 1816.5600 ;
        RECT 433.4400 1805.2000 435.0400 1805.6800 ;
        RECT 433.4400 1810.6400 435.0400 1811.1200 ;
        RECT 433.4400 1816.0800 435.0400 1816.5600 ;
        RECT 445.7800 1794.3200 448.7800 1794.8000 ;
        RECT 445.7800 1799.7600 448.7800 1800.2400 ;
        RECT 433.4400 1794.3200 435.0400 1794.8000 ;
        RECT 433.4400 1799.7600 435.0400 1800.2400 ;
        RECT 388.4400 1832.4000 390.0400 1832.8800 ;
        RECT 388.4400 1837.8400 390.0400 1838.3200 ;
        RECT 388.4400 1843.2800 390.0400 1843.7600 ;
        RECT 388.4400 1821.5200 390.0400 1822.0000 ;
        RECT 388.4400 1826.9600 390.0400 1827.4400 ;
        RECT 388.4400 1805.2000 390.0400 1805.6800 ;
        RECT 388.4400 1810.6400 390.0400 1811.1200 ;
        RECT 388.4400 1816.0800 390.0400 1816.5600 ;
        RECT 388.4400 1794.3200 390.0400 1794.8000 ;
        RECT 388.4400 1799.7600 390.0400 1800.2400 ;
        RECT 343.4400 1875.9200 345.0400 1876.4000 ;
        RECT 343.4400 1881.3600 345.0400 1881.8400 ;
        RECT 343.4400 1886.8000 345.0400 1887.2800 ;
        RECT 298.4400 1875.9200 300.0400 1876.4000 ;
        RECT 298.4400 1881.3600 300.0400 1881.8400 ;
        RECT 298.4400 1886.8000 300.0400 1887.2800 ;
        RECT 343.4400 1865.0400 345.0400 1865.5200 ;
        RECT 343.4400 1870.4800 345.0400 1870.9600 ;
        RECT 343.4400 1848.7200 345.0400 1849.2000 ;
        RECT 343.4400 1854.1600 345.0400 1854.6400 ;
        RECT 343.4400 1859.6000 345.0400 1860.0800 ;
        RECT 298.4400 1865.0400 300.0400 1865.5200 ;
        RECT 298.4400 1870.4800 300.0400 1870.9600 ;
        RECT 298.4400 1848.7200 300.0400 1849.2000 ;
        RECT 298.4400 1854.1600 300.0400 1854.6400 ;
        RECT 298.4400 1859.6000 300.0400 1860.0800 ;
        RECT 253.4400 1875.9200 255.0400 1876.4000 ;
        RECT 253.4400 1881.3600 255.0400 1881.8400 ;
        RECT 241.6800 1881.3600 244.6800 1881.8400 ;
        RECT 241.6800 1875.9200 244.6800 1876.4000 ;
        RECT 241.6800 1886.8000 244.6800 1887.2800 ;
        RECT 253.4400 1886.8000 255.0400 1887.2800 ;
        RECT 253.4400 1865.0400 255.0400 1865.5200 ;
        RECT 253.4400 1870.4800 255.0400 1870.9600 ;
        RECT 241.6800 1870.4800 244.6800 1870.9600 ;
        RECT 241.6800 1865.0400 244.6800 1865.5200 ;
        RECT 253.4400 1848.7200 255.0400 1849.2000 ;
        RECT 253.4400 1854.1600 255.0400 1854.6400 ;
        RECT 241.6800 1854.1600 244.6800 1854.6400 ;
        RECT 241.6800 1848.7200 244.6800 1849.2000 ;
        RECT 241.6800 1859.6000 244.6800 1860.0800 ;
        RECT 253.4400 1859.6000 255.0400 1860.0800 ;
        RECT 343.4400 1832.4000 345.0400 1832.8800 ;
        RECT 343.4400 1837.8400 345.0400 1838.3200 ;
        RECT 343.4400 1843.2800 345.0400 1843.7600 ;
        RECT 343.4400 1821.5200 345.0400 1822.0000 ;
        RECT 343.4400 1826.9600 345.0400 1827.4400 ;
        RECT 298.4400 1832.4000 300.0400 1832.8800 ;
        RECT 298.4400 1837.8400 300.0400 1838.3200 ;
        RECT 298.4400 1843.2800 300.0400 1843.7600 ;
        RECT 298.4400 1821.5200 300.0400 1822.0000 ;
        RECT 298.4400 1826.9600 300.0400 1827.4400 ;
        RECT 343.4400 1805.2000 345.0400 1805.6800 ;
        RECT 343.4400 1810.6400 345.0400 1811.1200 ;
        RECT 343.4400 1816.0800 345.0400 1816.5600 ;
        RECT 343.4400 1794.3200 345.0400 1794.8000 ;
        RECT 343.4400 1799.7600 345.0400 1800.2400 ;
        RECT 298.4400 1805.2000 300.0400 1805.6800 ;
        RECT 298.4400 1810.6400 300.0400 1811.1200 ;
        RECT 298.4400 1816.0800 300.0400 1816.5600 ;
        RECT 298.4400 1794.3200 300.0400 1794.8000 ;
        RECT 298.4400 1799.7600 300.0400 1800.2400 ;
        RECT 253.4400 1832.4000 255.0400 1832.8800 ;
        RECT 253.4400 1837.8400 255.0400 1838.3200 ;
        RECT 253.4400 1843.2800 255.0400 1843.7600 ;
        RECT 241.6800 1832.4000 244.6800 1832.8800 ;
        RECT 241.6800 1837.8400 244.6800 1838.3200 ;
        RECT 241.6800 1843.2800 244.6800 1843.7600 ;
        RECT 253.4400 1821.5200 255.0400 1822.0000 ;
        RECT 253.4400 1826.9600 255.0400 1827.4400 ;
        RECT 241.6800 1821.5200 244.6800 1822.0000 ;
        RECT 241.6800 1826.9600 244.6800 1827.4400 ;
        RECT 253.4400 1805.2000 255.0400 1805.6800 ;
        RECT 253.4400 1810.6400 255.0400 1811.1200 ;
        RECT 253.4400 1816.0800 255.0400 1816.5600 ;
        RECT 241.6800 1805.2000 244.6800 1805.6800 ;
        RECT 241.6800 1810.6400 244.6800 1811.1200 ;
        RECT 241.6800 1816.0800 244.6800 1816.5600 ;
        RECT 253.4400 1794.3200 255.0400 1794.8000 ;
        RECT 253.4400 1799.7600 255.0400 1800.2400 ;
        RECT 241.6800 1794.3200 244.6800 1794.8000 ;
        RECT 241.6800 1799.7600 244.6800 1800.2400 ;
        RECT 445.7800 1778.0000 448.7800 1778.4800 ;
        RECT 445.7800 1783.4400 448.7800 1783.9200 ;
        RECT 445.7800 1788.8800 448.7800 1789.3600 ;
        RECT 433.4400 1778.0000 435.0400 1778.4800 ;
        RECT 433.4400 1783.4400 435.0400 1783.9200 ;
        RECT 433.4400 1788.8800 435.0400 1789.3600 ;
        RECT 445.7800 1767.1200 448.7800 1767.6000 ;
        RECT 445.7800 1772.5600 448.7800 1773.0400 ;
        RECT 433.4400 1767.1200 435.0400 1767.6000 ;
        RECT 433.4400 1772.5600 435.0400 1773.0400 ;
        RECT 445.7800 1750.8000 448.7800 1751.2800 ;
        RECT 445.7800 1756.2400 448.7800 1756.7200 ;
        RECT 445.7800 1761.6800 448.7800 1762.1600 ;
        RECT 433.4400 1750.8000 435.0400 1751.2800 ;
        RECT 433.4400 1756.2400 435.0400 1756.7200 ;
        RECT 433.4400 1761.6800 435.0400 1762.1600 ;
        RECT 445.7800 1739.9200 448.7800 1740.4000 ;
        RECT 445.7800 1745.3600 448.7800 1745.8400 ;
        RECT 433.4400 1739.9200 435.0400 1740.4000 ;
        RECT 433.4400 1745.3600 435.0400 1745.8400 ;
        RECT 388.4400 1778.0000 390.0400 1778.4800 ;
        RECT 388.4400 1783.4400 390.0400 1783.9200 ;
        RECT 388.4400 1788.8800 390.0400 1789.3600 ;
        RECT 388.4400 1767.1200 390.0400 1767.6000 ;
        RECT 388.4400 1772.5600 390.0400 1773.0400 ;
        RECT 388.4400 1750.8000 390.0400 1751.2800 ;
        RECT 388.4400 1756.2400 390.0400 1756.7200 ;
        RECT 388.4400 1761.6800 390.0400 1762.1600 ;
        RECT 388.4400 1739.9200 390.0400 1740.4000 ;
        RECT 388.4400 1745.3600 390.0400 1745.8400 ;
        RECT 445.7800 1723.6000 448.7800 1724.0800 ;
        RECT 445.7800 1729.0400 448.7800 1729.5200 ;
        RECT 445.7800 1734.4800 448.7800 1734.9600 ;
        RECT 433.4400 1723.6000 435.0400 1724.0800 ;
        RECT 433.4400 1729.0400 435.0400 1729.5200 ;
        RECT 433.4400 1734.4800 435.0400 1734.9600 ;
        RECT 445.7800 1712.7200 448.7800 1713.2000 ;
        RECT 445.7800 1718.1600 448.7800 1718.6400 ;
        RECT 433.4400 1712.7200 435.0400 1713.2000 ;
        RECT 433.4400 1718.1600 435.0400 1718.6400 ;
        RECT 445.7800 1696.4000 448.7800 1696.8800 ;
        RECT 445.7800 1701.8400 448.7800 1702.3200 ;
        RECT 445.7800 1707.2800 448.7800 1707.7600 ;
        RECT 433.4400 1696.4000 435.0400 1696.8800 ;
        RECT 433.4400 1701.8400 435.0400 1702.3200 ;
        RECT 433.4400 1707.2800 435.0400 1707.7600 ;
        RECT 445.7800 1690.9600 448.7800 1691.4400 ;
        RECT 433.4400 1690.9600 435.0400 1691.4400 ;
        RECT 388.4400 1723.6000 390.0400 1724.0800 ;
        RECT 388.4400 1729.0400 390.0400 1729.5200 ;
        RECT 388.4400 1734.4800 390.0400 1734.9600 ;
        RECT 388.4400 1712.7200 390.0400 1713.2000 ;
        RECT 388.4400 1718.1600 390.0400 1718.6400 ;
        RECT 388.4400 1696.4000 390.0400 1696.8800 ;
        RECT 388.4400 1701.8400 390.0400 1702.3200 ;
        RECT 388.4400 1707.2800 390.0400 1707.7600 ;
        RECT 388.4400 1690.9600 390.0400 1691.4400 ;
        RECT 343.4400 1778.0000 345.0400 1778.4800 ;
        RECT 343.4400 1783.4400 345.0400 1783.9200 ;
        RECT 343.4400 1788.8800 345.0400 1789.3600 ;
        RECT 343.4400 1767.1200 345.0400 1767.6000 ;
        RECT 343.4400 1772.5600 345.0400 1773.0400 ;
        RECT 298.4400 1778.0000 300.0400 1778.4800 ;
        RECT 298.4400 1783.4400 300.0400 1783.9200 ;
        RECT 298.4400 1788.8800 300.0400 1789.3600 ;
        RECT 298.4400 1767.1200 300.0400 1767.6000 ;
        RECT 298.4400 1772.5600 300.0400 1773.0400 ;
        RECT 343.4400 1750.8000 345.0400 1751.2800 ;
        RECT 343.4400 1756.2400 345.0400 1756.7200 ;
        RECT 343.4400 1761.6800 345.0400 1762.1600 ;
        RECT 343.4400 1739.9200 345.0400 1740.4000 ;
        RECT 343.4400 1745.3600 345.0400 1745.8400 ;
        RECT 298.4400 1750.8000 300.0400 1751.2800 ;
        RECT 298.4400 1756.2400 300.0400 1756.7200 ;
        RECT 298.4400 1761.6800 300.0400 1762.1600 ;
        RECT 298.4400 1739.9200 300.0400 1740.4000 ;
        RECT 298.4400 1745.3600 300.0400 1745.8400 ;
        RECT 253.4400 1778.0000 255.0400 1778.4800 ;
        RECT 253.4400 1783.4400 255.0400 1783.9200 ;
        RECT 253.4400 1788.8800 255.0400 1789.3600 ;
        RECT 241.6800 1778.0000 244.6800 1778.4800 ;
        RECT 241.6800 1783.4400 244.6800 1783.9200 ;
        RECT 241.6800 1788.8800 244.6800 1789.3600 ;
        RECT 253.4400 1767.1200 255.0400 1767.6000 ;
        RECT 253.4400 1772.5600 255.0400 1773.0400 ;
        RECT 241.6800 1767.1200 244.6800 1767.6000 ;
        RECT 241.6800 1772.5600 244.6800 1773.0400 ;
        RECT 253.4400 1750.8000 255.0400 1751.2800 ;
        RECT 253.4400 1756.2400 255.0400 1756.7200 ;
        RECT 253.4400 1761.6800 255.0400 1762.1600 ;
        RECT 241.6800 1750.8000 244.6800 1751.2800 ;
        RECT 241.6800 1756.2400 244.6800 1756.7200 ;
        RECT 241.6800 1761.6800 244.6800 1762.1600 ;
        RECT 253.4400 1739.9200 255.0400 1740.4000 ;
        RECT 253.4400 1745.3600 255.0400 1745.8400 ;
        RECT 241.6800 1739.9200 244.6800 1740.4000 ;
        RECT 241.6800 1745.3600 244.6800 1745.8400 ;
        RECT 343.4400 1723.6000 345.0400 1724.0800 ;
        RECT 343.4400 1729.0400 345.0400 1729.5200 ;
        RECT 343.4400 1734.4800 345.0400 1734.9600 ;
        RECT 343.4400 1712.7200 345.0400 1713.2000 ;
        RECT 343.4400 1718.1600 345.0400 1718.6400 ;
        RECT 298.4400 1723.6000 300.0400 1724.0800 ;
        RECT 298.4400 1729.0400 300.0400 1729.5200 ;
        RECT 298.4400 1734.4800 300.0400 1734.9600 ;
        RECT 298.4400 1712.7200 300.0400 1713.2000 ;
        RECT 298.4400 1718.1600 300.0400 1718.6400 ;
        RECT 343.4400 1696.4000 345.0400 1696.8800 ;
        RECT 343.4400 1701.8400 345.0400 1702.3200 ;
        RECT 343.4400 1707.2800 345.0400 1707.7600 ;
        RECT 343.4400 1690.9600 345.0400 1691.4400 ;
        RECT 298.4400 1696.4000 300.0400 1696.8800 ;
        RECT 298.4400 1701.8400 300.0400 1702.3200 ;
        RECT 298.4400 1707.2800 300.0400 1707.7600 ;
        RECT 298.4400 1690.9600 300.0400 1691.4400 ;
        RECT 253.4400 1723.6000 255.0400 1724.0800 ;
        RECT 253.4400 1729.0400 255.0400 1729.5200 ;
        RECT 253.4400 1734.4800 255.0400 1734.9600 ;
        RECT 241.6800 1723.6000 244.6800 1724.0800 ;
        RECT 241.6800 1729.0400 244.6800 1729.5200 ;
        RECT 241.6800 1734.4800 244.6800 1734.9600 ;
        RECT 253.4400 1712.7200 255.0400 1713.2000 ;
        RECT 253.4400 1718.1600 255.0400 1718.6400 ;
        RECT 241.6800 1712.7200 244.6800 1713.2000 ;
        RECT 241.6800 1718.1600 244.6800 1718.6400 ;
        RECT 253.4400 1696.4000 255.0400 1696.8800 ;
        RECT 253.4400 1701.8400 255.0400 1702.3200 ;
        RECT 253.4400 1707.2800 255.0400 1707.7600 ;
        RECT 241.6800 1696.4000 244.6800 1696.8800 ;
        RECT 241.6800 1701.8400 244.6800 1702.3200 ;
        RECT 241.6800 1707.2800 244.6800 1707.7600 ;
        RECT 241.6800 1690.9600 244.6800 1691.4400 ;
        RECT 253.4400 1690.9600 255.0400 1691.4400 ;
        RECT 241.6800 1895.8700 448.7800 1898.8700 ;
        RECT 241.6800 1682.7700 448.7800 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 1453.1300 435.0400 1669.2300 ;
        RECT 388.4400 1453.1300 390.0400 1669.2300 ;
        RECT 343.4400 1453.1300 345.0400 1669.2300 ;
        RECT 298.4400 1453.1300 300.0400 1669.2300 ;
        RECT 253.4400 1453.1300 255.0400 1669.2300 ;
        RECT 445.7800 1453.1300 448.7800 1669.2300 ;
        RECT 241.6800 1453.1300 244.6800 1669.2300 ;
      LAYER met3 ;
        RECT 445.7800 1646.2800 448.7800 1646.7600 ;
        RECT 445.7800 1651.7200 448.7800 1652.2000 ;
        RECT 433.4400 1646.2800 435.0400 1646.7600 ;
        RECT 433.4400 1651.7200 435.0400 1652.2000 ;
        RECT 445.7800 1657.1600 448.7800 1657.6400 ;
        RECT 433.4400 1657.1600 435.0400 1657.6400 ;
        RECT 445.7800 1635.4000 448.7800 1635.8800 ;
        RECT 445.7800 1640.8400 448.7800 1641.3200 ;
        RECT 433.4400 1635.4000 435.0400 1635.8800 ;
        RECT 433.4400 1640.8400 435.0400 1641.3200 ;
        RECT 445.7800 1619.0800 448.7800 1619.5600 ;
        RECT 445.7800 1624.5200 448.7800 1625.0000 ;
        RECT 433.4400 1619.0800 435.0400 1619.5600 ;
        RECT 433.4400 1624.5200 435.0400 1625.0000 ;
        RECT 445.7800 1629.9600 448.7800 1630.4400 ;
        RECT 433.4400 1629.9600 435.0400 1630.4400 ;
        RECT 388.4400 1646.2800 390.0400 1646.7600 ;
        RECT 388.4400 1651.7200 390.0400 1652.2000 ;
        RECT 388.4400 1657.1600 390.0400 1657.6400 ;
        RECT 388.4400 1635.4000 390.0400 1635.8800 ;
        RECT 388.4400 1640.8400 390.0400 1641.3200 ;
        RECT 388.4400 1619.0800 390.0400 1619.5600 ;
        RECT 388.4400 1624.5200 390.0400 1625.0000 ;
        RECT 388.4400 1629.9600 390.0400 1630.4400 ;
        RECT 445.7800 1602.7600 448.7800 1603.2400 ;
        RECT 445.7800 1608.2000 448.7800 1608.6800 ;
        RECT 445.7800 1613.6400 448.7800 1614.1200 ;
        RECT 433.4400 1602.7600 435.0400 1603.2400 ;
        RECT 433.4400 1608.2000 435.0400 1608.6800 ;
        RECT 433.4400 1613.6400 435.0400 1614.1200 ;
        RECT 445.7800 1591.8800 448.7800 1592.3600 ;
        RECT 445.7800 1597.3200 448.7800 1597.8000 ;
        RECT 433.4400 1591.8800 435.0400 1592.3600 ;
        RECT 433.4400 1597.3200 435.0400 1597.8000 ;
        RECT 445.7800 1575.5600 448.7800 1576.0400 ;
        RECT 445.7800 1581.0000 448.7800 1581.4800 ;
        RECT 445.7800 1586.4400 448.7800 1586.9200 ;
        RECT 433.4400 1575.5600 435.0400 1576.0400 ;
        RECT 433.4400 1581.0000 435.0400 1581.4800 ;
        RECT 433.4400 1586.4400 435.0400 1586.9200 ;
        RECT 445.7800 1564.6800 448.7800 1565.1600 ;
        RECT 445.7800 1570.1200 448.7800 1570.6000 ;
        RECT 433.4400 1564.6800 435.0400 1565.1600 ;
        RECT 433.4400 1570.1200 435.0400 1570.6000 ;
        RECT 388.4400 1602.7600 390.0400 1603.2400 ;
        RECT 388.4400 1608.2000 390.0400 1608.6800 ;
        RECT 388.4400 1613.6400 390.0400 1614.1200 ;
        RECT 388.4400 1591.8800 390.0400 1592.3600 ;
        RECT 388.4400 1597.3200 390.0400 1597.8000 ;
        RECT 388.4400 1575.5600 390.0400 1576.0400 ;
        RECT 388.4400 1581.0000 390.0400 1581.4800 ;
        RECT 388.4400 1586.4400 390.0400 1586.9200 ;
        RECT 388.4400 1564.6800 390.0400 1565.1600 ;
        RECT 388.4400 1570.1200 390.0400 1570.6000 ;
        RECT 343.4400 1646.2800 345.0400 1646.7600 ;
        RECT 343.4400 1651.7200 345.0400 1652.2000 ;
        RECT 343.4400 1657.1600 345.0400 1657.6400 ;
        RECT 298.4400 1646.2800 300.0400 1646.7600 ;
        RECT 298.4400 1651.7200 300.0400 1652.2000 ;
        RECT 298.4400 1657.1600 300.0400 1657.6400 ;
        RECT 343.4400 1635.4000 345.0400 1635.8800 ;
        RECT 343.4400 1640.8400 345.0400 1641.3200 ;
        RECT 343.4400 1619.0800 345.0400 1619.5600 ;
        RECT 343.4400 1624.5200 345.0400 1625.0000 ;
        RECT 343.4400 1629.9600 345.0400 1630.4400 ;
        RECT 298.4400 1635.4000 300.0400 1635.8800 ;
        RECT 298.4400 1640.8400 300.0400 1641.3200 ;
        RECT 298.4400 1619.0800 300.0400 1619.5600 ;
        RECT 298.4400 1624.5200 300.0400 1625.0000 ;
        RECT 298.4400 1629.9600 300.0400 1630.4400 ;
        RECT 253.4400 1646.2800 255.0400 1646.7600 ;
        RECT 253.4400 1651.7200 255.0400 1652.2000 ;
        RECT 241.6800 1651.7200 244.6800 1652.2000 ;
        RECT 241.6800 1646.2800 244.6800 1646.7600 ;
        RECT 241.6800 1657.1600 244.6800 1657.6400 ;
        RECT 253.4400 1657.1600 255.0400 1657.6400 ;
        RECT 253.4400 1635.4000 255.0400 1635.8800 ;
        RECT 253.4400 1640.8400 255.0400 1641.3200 ;
        RECT 241.6800 1640.8400 244.6800 1641.3200 ;
        RECT 241.6800 1635.4000 244.6800 1635.8800 ;
        RECT 253.4400 1619.0800 255.0400 1619.5600 ;
        RECT 253.4400 1624.5200 255.0400 1625.0000 ;
        RECT 241.6800 1624.5200 244.6800 1625.0000 ;
        RECT 241.6800 1619.0800 244.6800 1619.5600 ;
        RECT 241.6800 1629.9600 244.6800 1630.4400 ;
        RECT 253.4400 1629.9600 255.0400 1630.4400 ;
        RECT 343.4400 1602.7600 345.0400 1603.2400 ;
        RECT 343.4400 1608.2000 345.0400 1608.6800 ;
        RECT 343.4400 1613.6400 345.0400 1614.1200 ;
        RECT 343.4400 1591.8800 345.0400 1592.3600 ;
        RECT 343.4400 1597.3200 345.0400 1597.8000 ;
        RECT 298.4400 1602.7600 300.0400 1603.2400 ;
        RECT 298.4400 1608.2000 300.0400 1608.6800 ;
        RECT 298.4400 1613.6400 300.0400 1614.1200 ;
        RECT 298.4400 1591.8800 300.0400 1592.3600 ;
        RECT 298.4400 1597.3200 300.0400 1597.8000 ;
        RECT 343.4400 1575.5600 345.0400 1576.0400 ;
        RECT 343.4400 1581.0000 345.0400 1581.4800 ;
        RECT 343.4400 1586.4400 345.0400 1586.9200 ;
        RECT 343.4400 1564.6800 345.0400 1565.1600 ;
        RECT 343.4400 1570.1200 345.0400 1570.6000 ;
        RECT 298.4400 1575.5600 300.0400 1576.0400 ;
        RECT 298.4400 1581.0000 300.0400 1581.4800 ;
        RECT 298.4400 1586.4400 300.0400 1586.9200 ;
        RECT 298.4400 1564.6800 300.0400 1565.1600 ;
        RECT 298.4400 1570.1200 300.0400 1570.6000 ;
        RECT 253.4400 1602.7600 255.0400 1603.2400 ;
        RECT 253.4400 1608.2000 255.0400 1608.6800 ;
        RECT 253.4400 1613.6400 255.0400 1614.1200 ;
        RECT 241.6800 1602.7600 244.6800 1603.2400 ;
        RECT 241.6800 1608.2000 244.6800 1608.6800 ;
        RECT 241.6800 1613.6400 244.6800 1614.1200 ;
        RECT 253.4400 1591.8800 255.0400 1592.3600 ;
        RECT 253.4400 1597.3200 255.0400 1597.8000 ;
        RECT 241.6800 1591.8800 244.6800 1592.3600 ;
        RECT 241.6800 1597.3200 244.6800 1597.8000 ;
        RECT 253.4400 1575.5600 255.0400 1576.0400 ;
        RECT 253.4400 1581.0000 255.0400 1581.4800 ;
        RECT 253.4400 1586.4400 255.0400 1586.9200 ;
        RECT 241.6800 1575.5600 244.6800 1576.0400 ;
        RECT 241.6800 1581.0000 244.6800 1581.4800 ;
        RECT 241.6800 1586.4400 244.6800 1586.9200 ;
        RECT 253.4400 1564.6800 255.0400 1565.1600 ;
        RECT 253.4400 1570.1200 255.0400 1570.6000 ;
        RECT 241.6800 1564.6800 244.6800 1565.1600 ;
        RECT 241.6800 1570.1200 244.6800 1570.6000 ;
        RECT 445.7800 1548.3600 448.7800 1548.8400 ;
        RECT 445.7800 1553.8000 448.7800 1554.2800 ;
        RECT 445.7800 1559.2400 448.7800 1559.7200 ;
        RECT 433.4400 1548.3600 435.0400 1548.8400 ;
        RECT 433.4400 1553.8000 435.0400 1554.2800 ;
        RECT 433.4400 1559.2400 435.0400 1559.7200 ;
        RECT 445.7800 1537.4800 448.7800 1537.9600 ;
        RECT 445.7800 1542.9200 448.7800 1543.4000 ;
        RECT 433.4400 1537.4800 435.0400 1537.9600 ;
        RECT 433.4400 1542.9200 435.0400 1543.4000 ;
        RECT 445.7800 1521.1600 448.7800 1521.6400 ;
        RECT 445.7800 1526.6000 448.7800 1527.0800 ;
        RECT 445.7800 1532.0400 448.7800 1532.5200 ;
        RECT 433.4400 1521.1600 435.0400 1521.6400 ;
        RECT 433.4400 1526.6000 435.0400 1527.0800 ;
        RECT 433.4400 1532.0400 435.0400 1532.5200 ;
        RECT 445.7800 1510.2800 448.7800 1510.7600 ;
        RECT 445.7800 1515.7200 448.7800 1516.2000 ;
        RECT 433.4400 1510.2800 435.0400 1510.7600 ;
        RECT 433.4400 1515.7200 435.0400 1516.2000 ;
        RECT 388.4400 1548.3600 390.0400 1548.8400 ;
        RECT 388.4400 1553.8000 390.0400 1554.2800 ;
        RECT 388.4400 1559.2400 390.0400 1559.7200 ;
        RECT 388.4400 1537.4800 390.0400 1537.9600 ;
        RECT 388.4400 1542.9200 390.0400 1543.4000 ;
        RECT 388.4400 1521.1600 390.0400 1521.6400 ;
        RECT 388.4400 1526.6000 390.0400 1527.0800 ;
        RECT 388.4400 1532.0400 390.0400 1532.5200 ;
        RECT 388.4400 1510.2800 390.0400 1510.7600 ;
        RECT 388.4400 1515.7200 390.0400 1516.2000 ;
        RECT 445.7800 1493.9600 448.7800 1494.4400 ;
        RECT 445.7800 1499.4000 448.7800 1499.8800 ;
        RECT 445.7800 1504.8400 448.7800 1505.3200 ;
        RECT 433.4400 1493.9600 435.0400 1494.4400 ;
        RECT 433.4400 1499.4000 435.0400 1499.8800 ;
        RECT 433.4400 1504.8400 435.0400 1505.3200 ;
        RECT 445.7800 1483.0800 448.7800 1483.5600 ;
        RECT 445.7800 1488.5200 448.7800 1489.0000 ;
        RECT 433.4400 1483.0800 435.0400 1483.5600 ;
        RECT 433.4400 1488.5200 435.0400 1489.0000 ;
        RECT 445.7800 1466.7600 448.7800 1467.2400 ;
        RECT 445.7800 1472.2000 448.7800 1472.6800 ;
        RECT 445.7800 1477.6400 448.7800 1478.1200 ;
        RECT 433.4400 1466.7600 435.0400 1467.2400 ;
        RECT 433.4400 1472.2000 435.0400 1472.6800 ;
        RECT 433.4400 1477.6400 435.0400 1478.1200 ;
        RECT 445.7800 1461.3200 448.7800 1461.8000 ;
        RECT 433.4400 1461.3200 435.0400 1461.8000 ;
        RECT 388.4400 1493.9600 390.0400 1494.4400 ;
        RECT 388.4400 1499.4000 390.0400 1499.8800 ;
        RECT 388.4400 1504.8400 390.0400 1505.3200 ;
        RECT 388.4400 1483.0800 390.0400 1483.5600 ;
        RECT 388.4400 1488.5200 390.0400 1489.0000 ;
        RECT 388.4400 1466.7600 390.0400 1467.2400 ;
        RECT 388.4400 1472.2000 390.0400 1472.6800 ;
        RECT 388.4400 1477.6400 390.0400 1478.1200 ;
        RECT 388.4400 1461.3200 390.0400 1461.8000 ;
        RECT 343.4400 1548.3600 345.0400 1548.8400 ;
        RECT 343.4400 1553.8000 345.0400 1554.2800 ;
        RECT 343.4400 1559.2400 345.0400 1559.7200 ;
        RECT 343.4400 1537.4800 345.0400 1537.9600 ;
        RECT 343.4400 1542.9200 345.0400 1543.4000 ;
        RECT 298.4400 1548.3600 300.0400 1548.8400 ;
        RECT 298.4400 1553.8000 300.0400 1554.2800 ;
        RECT 298.4400 1559.2400 300.0400 1559.7200 ;
        RECT 298.4400 1537.4800 300.0400 1537.9600 ;
        RECT 298.4400 1542.9200 300.0400 1543.4000 ;
        RECT 343.4400 1521.1600 345.0400 1521.6400 ;
        RECT 343.4400 1526.6000 345.0400 1527.0800 ;
        RECT 343.4400 1532.0400 345.0400 1532.5200 ;
        RECT 343.4400 1510.2800 345.0400 1510.7600 ;
        RECT 343.4400 1515.7200 345.0400 1516.2000 ;
        RECT 298.4400 1521.1600 300.0400 1521.6400 ;
        RECT 298.4400 1526.6000 300.0400 1527.0800 ;
        RECT 298.4400 1532.0400 300.0400 1532.5200 ;
        RECT 298.4400 1510.2800 300.0400 1510.7600 ;
        RECT 298.4400 1515.7200 300.0400 1516.2000 ;
        RECT 253.4400 1548.3600 255.0400 1548.8400 ;
        RECT 253.4400 1553.8000 255.0400 1554.2800 ;
        RECT 253.4400 1559.2400 255.0400 1559.7200 ;
        RECT 241.6800 1548.3600 244.6800 1548.8400 ;
        RECT 241.6800 1553.8000 244.6800 1554.2800 ;
        RECT 241.6800 1559.2400 244.6800 1559.7200 ;
        RECT 253.4400 1537.4800 255.0400 1537.9600 ;
        RECT 253.4400 1542.9200 255.0400 1543.4000 ;
        RECT 241.6800 1537.4800 244.6800 1537.9600 ;
        RECT 241.6800 1542.9200 244.6800 1543.4000 ;
        RECT 253.4400 1521.1600 255.0400 1521.6400 ;
        RECT 253.4400 1526.6000 255.0400 1527.0800 ;
        RECT 253.4400 1532.0400 255.0400 1532.5200 ;
        RECT 241.6800 1521.1600 244.6800 1521.6400 ;
        RECT 241.6800 1526.6000 244.6800 1527.0800 ;
        RECT 241.6800 1532.0400 244.6800 1532.5200 ;
        RECT 253.4400 1510.2800 255.0400 1510.7600 ;
        RECT 253.4400 1515.7200 255.0400 1516.2000 ;
        RECT 241.6800 1510.2800 244.6800 1510.7600 ;
        RECT 241.6800 1515.7200 244.6800 1516.2000 ;
        RECT 343.4400 1493.9600 345.0400 1494.4400 ;
        RECT 343.4400 1499.4000 345.0400 1499.8800 ;
        RECT 343.4400 1504.8400 345.0400 1505.3200 ;
        RECT 343.4400 1483.0800 345.0400 1483.5600 ;
        RECT 343.4400 1488.5200 345.0400 1489.0000 ;
        RECT 298.4400 1493.9600 300.0400 1494.4400 ;
        RECT 298.4400 1499.4000 300.0400 1499.8800 ;
        RECT 298.4400 1504.8400 300.0400 1505.3200 ;
        RECT 298.4400 1483.0800 300.0400 1483.5600 ;
        RECT 298.4400 1488.5200 300.0400 1489.0000 ;
        RECT 343.4400 1466.7600 345.0400 1467.2400 ;
        RECT 343.4400 1472.2000 345.0400 1472.6800 ;
        RECT 343.4400 1477.6400 345.0400 1478.1200 ;
        RECT 343.4400 1461.3200 345.0400 1461.8000 ;
        RECT 298.4400 1466.7600 300.0400 1467.2400 ;
        RECT 298.4400 1472.2000 300.0400 1472.6800 ;
        RECT 298.4400 1477.6400 300.0400 1478.1200 ;
        RECT 298.4400 1461.3200 300.0400 1461.8000 ;
        RECT 253.4400 1493.9600 255.0400 1494.4400 ;
        RECT 253.4400 1499.4000 255.0400 1499.8800 ;
        RECT 253.4400 1504.8400 255.0400 1505.3200 ;
        RECT 241.6800 1493.9600 244.6800 1494.4400 ;
        RECT 241.6800 1499.4000 244.6800 1499.8800 ;
        RECT 241.6800 1504.8400 244.6800 1505.3200 ;
        RECT 253.4400 1483.0800 255.0400 1483.5600 ;
        RECT 253.4400 1488.5200 255.0400 1489.0000 ;
        RECT 241.6800 1483.0800 244.6800 1483.5600 ;
        RECT 241.6800 1488.5200 244.6800 1489.0000 ;
        RECT 253.4400 1466.7600 255.0400 1467.2400 ;
        RECT 253.4400 1472.2000 255.0400 1472.6800 ;
        RECT 253.4400 1477.6400 255.0400 1478.1200 ;
        RECT 241.6800 1466.7600 244.6800 1467.2400 ;
        RECT 241.6800 1472.2000 244.6800 1472.6800 ;
        RECT 241.6800 1477.6400 244.6800 1478.1200 ;
        RECT 241.6800 1461.3200 244.6800 1461.8000 ;
        RECT 253.4400 1461.3200 255.0400 1461.8000 ;
        RECT 241.6800 1666.2300 448.7800 1669.2300 ;
        RECT 241.6800 1453.1300 448.7800 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 1223.4900 435.0400 1439.5900 ;
        RECT 388.4400 1223.4900 390.0400 1439.5900 ;
        RECT 343.4400 1223.4900 345.0400 1439.5900 ;
        RECT 298.4400 1223.4900 300.0400 1439.5900 ;
        RECT 253.4400 1223.4900 255.0400 1439.5900 ;
        RECT 445.7800 1223.4900 448.7800 1439.5900 ;
        RECT 241.6800 1223.4900 244.6800 1439.5900 ;
      LAYER met3 ;
        RECT 445.7800 1416.6400 448.7800 1417.1200 ;
        RECT 445.7800 1422.0800 448.7800 1422.5600 ;
        RECT 433.4400 1416.6400 435.0400 1417.1200 ;
        RECT 433.4400 1422.0800 435.0400 1422.5600 ;
        RECT 445.7800 1427.5200 448.7800 1428.0000 ;
        RECT 433.4400 1427.5200 435.0400 1428.0000 ;
        RECT 445.7800 1405.7600 448.7800 1406.2400 ;
        RECT 445.7800 1411.2000 448.7800 1411.6800 ;
        RECT 433.4400 1405.7600 435.0400 1406.2400 ;
        RECT 433.4400 1411.2000 435.0400 1411.6800 ;
        RECT 445.7800 1389.4400 448.7800 1389.9200 ;
        RECT 445.7800 1394.8800 448.7800 1395.3600 ;
        RECT 433.4400 1389.4400 435.0400 1389.9200 ;
        RECT 433.4400 1394.8800 435.0400 1395.3600 ;
        RECT 445.7800 1400.3200 448.7800 1400.8000 ;
        RECT 433.4400 1400.3200 435.0400 1400.8000 ;
        RECT 388.4400 1416.6400 390.0400 1417.1200 ;
        RECT 388.4400 1422.0800 390.0400 1422.5600 ;
        RECT 388.4400 1427.5200 390.0400 1428.0000 ;
        RECT 388.4400 1405.7600 390.0400 1406.2400 ;
        RECT 388.4400 1411.2000 390.0400 1411.6800 ;
        RECT 388.4400 1389.4400 390.0400 1389.9200 ;
        RECT 388.4400 1394.8800 390.0400 1395.3600 ;
        RECT 388.4400 1400.3200 390.0400 1400.8000 ;
        RECT 445.7800 1373.1200 448.7800 1373.6000 ;
        RECT 445.7800 1378.5600 448.7800 1379.0400 ;
        RECT 445.7800 1384.0000 448.7800 1384.4800 ;
        RECT 433.4400 1373.1200 435.0400 1373.6000 ;
        RECT 433.4400 1378.5600 435.0400 1379.0400 ;
        RECT 433.4400 1384.0000 435.0400 1384.4800 ;
        RECT 445.7800 1362.2400 448.7800 1362.7200 ;
        RECT 445.7800 1367.6800 448.7800 1368.1600 ;
        RECT 433.4400 1362.2400 435.0400 1362.7200 ;
        RECT 433.4400 1367.6800 435.0400 1368.1600 ;
        RECT 445.7800 1345.9200 448.7800 1346.4000 ;
        RECT 445.7800 1351.3600 448.7800 1351.8400 ;
        RECT 445.7800 1356.8000 448.7800 1357.2800 ;
        RECT 433.4400 1345.9200 435.0400 1346.4000 ;
        RECT 433.4400 1351.3600 435.0400 1351.8400 ;
        RECT 433.4400 1356.8000 435.0400 1357.2800 ;
        RECT 445.7800 1335.0400 448.7800 1335.5200 ;
        RECT 445.7800 1340.4800 448.7800 1340.9600 ;
        RECT 433.4400 1335.0400 435.0400 1335.5200 ;
        RECT 433.4400 1340.4800 435.0400 1340.9600 ;
        RECT 388.4400 1373.1200 390.0400 1373.6000 ;
        RECT 388.4400 1378.5600 390.0400 1379.0400 ;
        RECT 388.4400 1384.0000 390.0400 1384.4800 ;
        RECT 388.4400 1362.2400 390.0400 1362.7200 ;
        RECT 388.4400 1367.6800 390.0400 1368.1600 ;
        RECT 388.4400 1345.9200 390.0400 1346.4000 ;
        RECT 388.4400 1351.3600 390.0400 1351.8400 ;
        RECT 388.4400 1356.8000 390.0400 1357.2800 ;
        RECT 388.4400 1335.0400 390.0400 1335.5200 ;
        RECT 388.4400 1340.4800 390.0400 1340.9600 ;
        RECT 343.4400 1416.6400 345.0400 1417.1200 ;
        RECT 343.4400 1422.0800 345.0400 1422.5600 ;
        RECT 343.4400 1427.5200 345.0400 1428.0000 ;
        RECT 298.4400 1416.6400 300.0400 1417.1200 ;
        RECT 298.4400 1422.0800 300.0400 1422.5600 ;
        RECT 298.4400 1427.5200 300.0400 1428.0000 ;
        RECT 343.4400 1405.7600 345.0400 1406.2400 ;
        RECT 343.4400 1411.2000 345.0400 1411.6800 ;
        RECT 343.4400 1389.4400 345.0400 1389.9200 ;
        RECT 343.4400 1394.8800 345.0400 1395.3600 ;
        RECT 343.4400 1400.3200 345.0400 1400.8000 ;
        RECT 298.4400 1405.7600 300.0400 1406.2400 ;
        RECT 298.4400 1411.2000 300.0400 1411.6800 ;
        RECT 298.4400 1389.4400 300.0400 1389.9200 ;
        RECT 298.4400 1394.8800 300.0400 1395.3600 ;
        RECT 298.4400 1400.3200 300.0400 1400.8000 ;
        RECT 253.4400 1416.6400 255.0400 1417.1200 ;
        RECT 253.4400 1422.0800 255.0400 1422.5600 ;
        RECT 241.6800 1422.0800 244.6800 1422.5600 ;
        RECT 241.6800 1416.6400 244.6800 1417.1200 ;
        RECT 241.6800 1427.5200 244.6800 1428.0000 ;
        RECT 253.4400 1427.5200 255.0400 1428.0000 ;
        RECT 253.4400 1405.7600 255.0400 1406.2400 ;
        RECT 253.4400 1411.2000 255.0400 1411.6800 ;
        RECT 241.6800 1411.2000 244.6800 1411.6800 ;
        RECT 241.6800 1405.7600 244.6800 1406.2400 ;
        RECT 253.4400 1389.4400 255.0400 1389.9200 ;
        RECT 253.4400 1394.8800 255.0400 1395.3600 ;
        RECT 241.6800 1394.8800 244.6800 1395.3600 ;
        RECT 241.6800 1389.4400 244.6800 1389.9200 ;
        RECT 241.6800 1400.3200 244.6800 1400.8000 ;
        RECT 253.4400 1400.3200 255.0400 1400.8000 ;
        RECT 343.4400 1373.1200 345.0400 1373.6000 ;
        RECT 343.4400 1378.5600 345.0400 1379.0400 ;
        RECT 343.4400 1384.0000 345.0400 1384.4800 ;
        RECT 343.4400 1362.2400 345.0400 1362.7200 ;
        RECT 343.4400 1367.6800 345.0400 1368.1600 ;
        RECT 298.4400 1373.1200 300.0400 1373.6000 ;
        RECT 298.4400 1378.5600 300.0400 1379.0400 ;
        RECT 298.4400 1384.0000 300.0400 1384.4800 ;
        RECT 298.4400 1362.2400 300.0400 1362.7200 ;
        RECT 298.4400 1367.6800 300.0400 1368.1600 ;
        RECT 343.4400 1345.9200 345.0400 1346.4000 ;
        RECT 343.4400 1351.3600 345.0400 1351.8400 ;
        RECT 343.4400 1356.8000 345.0400 1357.2800 ;
        RECT 343.4400 1335.0400 345.0400 1335.5200 ;
        RECT 343.4400 1340.4800 345.0400 1340.9600 ;
        RECT 298.4400 1345.9200 300.0400 1346.4000 ;
        RECT 298.4400 1351.3600 300.0400 1351.8400 ;
        RECT 298.4400 1356.8000 300.0400 1357.2800 ;
        RECT 298.4400 1335.0400 300.0400 1335.5200 ;
        RECT 298.4400 1340.4800 300.0400 1340.9600 ;
        RECT 253.4400 1373.1200 255.0400 1373.6000 ;
        RECT 253.4400 1378.5600 255.0400 1379.0400 ;
        RECT 253.4400 1384.0000 255.0400 1384.4800 ;
        RECT 241.6800 1373.1200 244.6800 1373.6000 ;
        RECT 241.6800 1378.5600 244.6800 1379.0400 ;
        RECT 241.6800 1384.0000 244.6800 1384.4800 ;
        RECT 253.4400 1362.2400 255.0400 1362.7200 ;
        RECT 253.4400 1367.6800 255.0400 1368.1600 ;
        RECT 241.6800 1362.2400 244.6800 1362.7200 ;
        RECT 241.6800 1367.6800 244.6800 1368.1600 ;
        RECT 253.4400 1345.9200 255.0400 1346.4000 ;
        RECT 253.4400 1351.3600 255.0400 1351.8400 ;
        RECT 253.4400 1356.8000 255.0400 1357.2800 ;
        RECT 241.6800 1345.9200 244.6800 1346.4000 ;
        RECT 241.6800 1351.3600 244.6800 1351.8400 ;
        RECT 241.6800 1356.8000 244.6800 1357.2800 ;
        RECT 253.4400 1335.0400 255.0400 1335.5200 ;
        RECT 253.4400 1340.4800 255.0400 1340.9600 ;
        RECT 241.6800 1335.0400 244.6800 1335.5200 ;
        RECT 241.6800 1340.4800 244.6800 1340.9600 ;
        RECT 445.7800 1318.7200 448.7800 1319.2000 ;
        RECT 445.7800 1324.1600 448.7800 1324.6400 ;
        RECT 445.7800 1329.6000 448.7800 1330.0800 ;
        RECT 433.4400 1318.7200 435.0400 1319.2000 ;
        RECT 433.4400 1324.1600 435.0400 1324.6400 ;
        RECT 433.4400 1329.6000 435.0400 1330.0800 ;
        RECT 445.7800 1307.8400 448.7800 1308.3200 ;
        RECT 445.7800 1313.2800 448.7800 1313.7600 ;
        RECT 433.4400 1307.8400 435.0400 1308.3200 ;
        RECT 433.4400 1313.2800 435.0400 1313.7600 ;
        RECT 445.7800 1291.5200 448.7800 1292.0000 ;
        RECT 445.7800 1296.9600 448.7800 1297.4400 ;
        RECT 445.7800 1302.4000 448.7800 1302.8800 ;
        RECT 433.4400 1291.5200 435.0400 1292.0000 ;
        RECT 433.4400 1296.9600 435.0400 1297.4400 ;
        RECT 433.4400 1302.4000 435.0400 1302.8800 ;
        RECT 445.7800 1280.6400 448.7800 1281.1200 ;
        RECT 445.7800 1286.0800 448.7800 1286.5600 ;
        RECT 433.4400 1280.6400 435.0400 1281.1200 ;
        RECT 433.4400 1286.0800 435.0400 1286.5600 ;
        RECT 388.4400 1318.7200 390.0400 1319.2000 ;
        RECT 388.4400 1324.1600 390.0400 1324.6400 ;
        RECT 388.4400 1329.6000 390.0400 1330.0800 ;
        RECT 388.4400 1307.8400 390.0400 1308.3200 ;
        RECT 388.4400 1313.2800 390.0400 1313.7600 ;
        RECT 388.4400 1291.5200 390.0400 1292.0000 ;
        RECT 388.4400 1296.9600 390.0400 1297.4400 ;
        RECT 388.4400 1302.4000 390.0400 1302.8800 ;
        RECT 388.4400 1280.6400 390.0400 1281.1200 ;
        RECT 388.4400 1286.0800 390.0400 1286.5600 ;
        RECT 445.7800 1264.3200 448.7800 1264.8000 ;
        RECT 445.7800 1269.7600 448.7800 1270.2400 ;
        RECT 445.7800 1275.2000 448.7800 1275.6800 ;
        RECT 433.4400 1264.3200 435.0400 1264.8000 ;
        RECT 433.4400 1269.7600 435.0400 1270.2400 ;
        RECT 433.4400 1275.2000 435.0400 1275.6800 ;
        RECT 445.7800 1253.4400 448.7800 1253.9200 ;
        RECT 445.7800 1258.8800 448.7800 1259.3600 ;
        RECT 433.4400 1253.4400 435.0400 1253.9200 ;
        RECT 433.4400 1258.8800 435.0400 1259.3600 ;
        RECT 445.7800 1237.1200 448.7800 1237.6000 ;
        RECT 445.7800 1242.5600 448.7800 1243.0400 ;
        RECT 445.7800 1248.0000 448.7800 1248.4800 ;
        RECT 433.4400 1237.1200 435.0400 1237.6000 ;
        RECT 433.4400 1242.5600 435.0400 1243.0400 ;
        RECT 433.4400 1248.0000 435.0400 1248.4800 ;
        RECT 445.7800 1231.6800 448.7800 1232.1600 ;
        RECT 433.4400 1231.6800 435.0400 1232.1600 ;
        RECT 388.4400 1264.3200 390.0400 1264.8000 ;
        RECT 388.4400 1269.7600 390.0400 1270.2400 ;
        RECT 388.4400 1275.2000 390.0400 1275.6800 ;
        RECT 388.4400 1253.4400 390.0400 1253.9200 ;
        RECT 388.4400 1258.8800 390.0400 1259.3600 ;
        RECT 388.4400 1237.1200 390.0400 1237.6000 ;
        RECT 388.4400 1242.5600 390.0400 1243.0400 ;
        RECT 388.4400 1248.0000 390.0400 1248.4800 ;
        RECT 388.4400 1231.6800 390.0400 1232.1600 ;
        RECT 343.4400 1318.7200 345.0400 1319.2000 ;
        RECT 343.4400 1324.1600 345.0400 1324.6400 ;
        RECT 343.4400 1329.6000 345.0400 1330.0800 ;
        RECT 343.4400 1307.8400 345.0400 1308.3200 ;
        RECT 343.4400 1313.2800 345.0400 1313.7600 ;
        RECT 298.4400 1318.7200 300.0400 1319.2000 ;
        RECT 298.4400 1324.1600 300.0400 1324.6400 ;
        RECT 298.4400 1329.6000 300.0400 1330.0800 ;
        RECT 298.4400 1307.8400 300.0400 1308.3200 ;
        RECT 298.4400 1313.2800 300.0400 1313.7600 ;
        RECT 343.4400 1291.5200 345.0400 1292.0000 ;
        RECT 343.4400 1296.9600 345.0400 1297.4400 ;
        RECT 343.4400 1302.4000 345.0400 1302.8800 ;
        RECT 343.4400 1280.6400 345.0400 1281.1200 ;
        RECT 343.4400 1286.0800 345.0400 1286.5600 ;
        RECT 298.4400 1291.5200 300.0400 1292.0000 ;
        RECT 298.4400 1296.9600 300.0400 1297.4400 ;
        RECT 298.4400 1302.4000 300.0400 1302.8800 ;
        RECT 298.4400 1280.6400 300.0400 1281.1200 ;
        RECT 298.4400 1286.0800 300.0400 1286.5600 ;
        RECT 253.4400 1318.7200 255.0400 1319.2000 ;
        RECT 253.4400 1324.1600 255.0400 1324.6400 ;
        RECT 253.4400 1329.6000 255.0400 1330.0800 ;
        RECT 241.6800 1318.7200 244.6800 1319.2000 ;
        RECT 241.6800 1324.1600 244.6800 1324.6400 ;
        RECT 241.6800 1329.6000 244.6800 1330.0800 ;
        RECT 253.4400 1307.8400 255.0400 1308.3200 ;
        RECT 253.4400 1313.2800 255.0400 1313.7600 ;
        RECT 241.6800 1307.8400 244.6800 1308.3200 ;
        RECT 241.6800 1313.2800 244.6800 1313.7600 ;
        RECT 253.4400 1291.5200 255.0400 1292.0000 ;
        RECT 253.4400 1296.9600 255.0400 1297.4400 ;
        RECT 253.4400 1302.4000 255.0400 1302.8800 ;
        RECT 241.6800 1291.5200 244.6800 1292.0000 ;
        RECT 241.6800 1296.9600 244.6800 1297.4400 ;
        RECT 241.6800 1302.4000 244.6800 1302.8800 ;
        RECT 253.4400 1280.6400 255.0400 1281.1200 ;
        RECT 253.4400 1286.0800 255.0400 1286.5600 ;
        RECT 241.6800 1280.6400 244.6800 1281.1200 ;
        RECT 241.6800 1286.0800 244.6800 1286.5600 ;
        RECT 343.4400 1264.3200 345.0400 1264.8000 ;
        RECT 343.4400 1269.7600 345.0400 1270.2400 ;
        RECT 343.4400 1275.2000 345.0400 1275.6800 ;
        RECT 343.4400 1253.4400 345.0400 1253.9200 ;
        RECT 343.4400 1258.8800 345.0400 1259.3600 ;
        RECT 298.4400 1264.3200 300.0400 1264.8000 ;
        RECT 298.4400 1269.7600 300.0400 1270.2400 ;
        RECT 298.4400 1275.2000 300.0400 1275.6800 ;
        RECT 298.4400 1253.4400 300.0400 1253.9200 ;
        RECT 298.4400 1258.8800 300.0400 1259.3600 ;
        RECT 343.4400 1237.1200 345.0400 1237.6000 ;
        RECT 343.4400 1242.5600 345.0400 1243.0400 ;
        RECT 343.4400 1248.0000 345.0400 1248.4800 ;
        RECT 343.4400 1231.6800 345.0400 1232.1600 ;
        RECT 298.4400 1237.1200 300.0400 1237.6000 ;
        RECT 298.4400 1242.5600 300.0400 1243.0400 ;
        RECT 298.4400 1248.0000 300.0400 1248.4800 ;
        RECT 298.4400 1231.6800 300.0400 1232.1600 ;
        RECT 253.4400 1264.3200 255.0400 1264.8000 ;
        RECT 253.4400 1269.7600 255.0400 1270.2400 ;
        RECT 253.4400 1275.2000 255.0400 1275.6800 ;
        RECT 241.6800 1264.3200 244.6800 1264.8000 ;
        RECT 241.6800 1269.7600 244.6800 1270.2400 ;
        RECT 241.6800 1275.2000 244.6800 1275.6800 ;
        RECT 253.4400 1253.4400 255.0400 1253.9200 ;
        RECT 253.4400 1258.8800 255.0400 1259.3600 ;
        RECT 241.6800 1253.4400 244.6800 1253.9200 ;
        RECT 241.6800 1258.8800 244.6800 1259.3600 ;
        RECT 253.4400 1237.1200 255.0400 1237.6000 ;
        RECT 253.4400 1242.5600 255.0400 1243.0400 ;
        RECT 253.4400 1248.0000 255.0400 1248.4800 ;
        RECT 241.6800 1237.1200 244.6800 1237.6000 ;
        RECT 241.6800 1242.5600 244.6800 1243.0400 ;
        RECT 241.6800 1248.0000 244.6800 1248.4800 ;
        RECT 241.6800 1231.6800 244.6800 1232.1600 ;
        RECT 253.4400 1231.6800 255.0400 1232.1600 ;
        RECT 241.6800 1436.5900 448.7800 1439.5900 ;
        RECT 241.6800 1223.4900 448.7800 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 993.8500 435.0400 1209.9500 ;
        RECT 388.4400 993.8500 390.0400 1209.9500 ;
        RECT 343.4400 993.8500 345.0400 1209.9500 ;
        RECT 298.4400 993.8500 300.0400 1209.9500 ;
        RECT 253.4400 993.8500 255.0400 1209.9500 ;
        RECT 445.7800 993.8500 448.7800 1209.9500 ;
        RECT 241.6800 993.8500 244.6800 1209.9500 ;
      LAYER met3 ;
        RECT 445.7800 1187.0000 448.7800 1187.4800 ;
        RECT 445.7800 1192.4400 448.7800 1192.9200 ;
        RECT 433.4400 1187.0000 435.0400 1187.4800 ;
        RECT 433.4400 1192.4400 435.0400 1192.9200 ;
        RECT 445.7800 1197.8800 448.7800 1198.3600 ;
        RECT 433.4400 1197.8800 435.0400 1198.3600 ;
        RECT 445.7800 1176.1200 448.7800 1176.6000 ;
        RECT 445.7800 1181.5600 448.7800 1182.0400 ;
        RECT 433.4400 1176.1200 435.0400 1176.6000 ;
        RECT 433.4400 1181.5600 435.0400 1182.0400 ;
        RECT 445.7800 1159.8000 448.7800 1160.2800 ;
        RECT 445.7800 1165.2400 448.7800 1165.7200 ;
        RECT 433.4400 1159.8000 435.0400 1160.2800 ;
        RECT 433.4400 1165.2400 435.0400 1165.7200 ;
        RECT 445.7800 1170.6800 448.7800 1171.1600 ;
        RECT 433.4400 1170.6800 435.0400 1171.1600 ;
        RECT 388.4400 1187.0000 390.0400 1187.4800 ;
        RECT 388.4400 1192.4400 390.0400 1192.9200 ;
        RECT 388.4400 1197.8800 390.0400 1198.3600 ;
        RECT 388.4400 1176.1200 390.0400 1176.6000 ;
        RECT 388.4400 1181.5600 390.0400 1182.0400 ;
        RECT 388.4400 1159.8000 390.0400 1160.2800 ;
        RECT 388.4400 1165.2400 390.0400 1165.7200 ;
        RECT 388.4400 1170.6800 390.0400 1171.1600 ;
        RECT 445.7800 1143.4800 448.7800 1143.9600 ;
        RECT 445.7800 1148.9200 448.7800 1149.4000 ;
        RECT 445.7800 1154.3600 448.7800 1154.8400 ;
        RECT 433.4400 1143.4800 435.0400 1143.9600 ;
        RECT 433.4400 1148.9200 435.0400 1149.4000 ;
        RECT 433.4400 1154.3600 435.0400 1154.8400 ;
        RECT 445.7800 1132.6000 448.7800 1133.0800 ;
        RECT 445.7800 1138.0400 448.7800 1138.5200 ;
        RECT 433.4400 1132.6000 435.0400 1133.0800 ;
        RECT 433.4400 1138.0400 435.0400 1138.5200 ;
        RECT 445.7800 1116.2800 448.7800 1116.7600 ;
        RECT 445.7800 1121.7200 448.7800 1122.2000 ;
        RECT 445.7800 1127.1600 448.7800 1127.6400 ;
        RECT 433.4400 1116.2800 435.0400 1116.7600 ;
        RECT 433.4400 1121.7200 435.0400 1122.2000 ;
        RECT 433.4400 1127.1600 435.0400 1127.6400 ;
        RECT 445.7800 1105.4000 448.7800 1105.8800 ;
        RECT 445.7800 1110.8400 448.7800 1111.3200 ;
        RECT 433.4400 1105.4000 435.0400 1105.8800 ;
        RECT 433.4400 1110.8400 435.0400 1111.3200 ;
        RECT 388.4400 1143.4800 390.0400 1143.9600 ;
        RECT 388.4400 1148.9200 390.0400 1149.4000 ;
        RECT 388.4400 1154.3600 390.0400 1154.8400 ;
        RECT 388.4400 1132.6000 390.0400 1133.0800 ;
        RECT 388.4400 1138.0400 390.0400 1138.5200 ;
        RECT 388.4400 1116.2800 390.0400 1116.7600 ;
        RECT 388.4400 1121.7200 390.0400 1122.2000 ;
        RECT 388.4400 1127.1600 390.0400 1127.6400 ;
        RECT 388.4400 1105.4000 390.0400 1105.8800 ;
        RECT 388.4400 1110.8400 390.0400 1111.3200 ;
        RECT 343.4400 1187.0000 345.0400 1187.4800 ;
        RECT 343.4400 1192.4400 345.0400 1192.9200 ;
        RECT 343.4400 1197.8800 345.0400 1198.3600 ;
        RECT 298.4400 1187.0000 300.0400 1187.4800 ;
        RECT 298.4400 1192.4400 300.0400 1192.9200 ;
        RECT 298.4400 1197.8800 300.0400 1198.3600 ;
        RECT 343.4400 1176.1200 345.0400 1176.6000 ;
        RECT 343.4400 1181.5600 345.0400 1182.0400 ;
        RECT 343.4400 1159.8000 345.0400 1160.2800 ;
        RECT 343.4400 1165.2400 345.0400 1165.7200 ;
        RECT 343.4400 1170.6800 345.0400 1171.1600 ;
        RECT 298.4400 1176.1200 300.0400 1176.6000 ;
        RECT 298.4400 1181.5600 300.0400 1182.0400 ;
        RECT 298.4400 1159.8000 300.0400 1160.2800 ;
        RECT 298.4400 1165.2400 300.0400 1165.7200 ;
        RECT 298.4400 1170.6800 300.0400 1171.1600 ;
        RECT 253.4400 1187.0000 255.0400 1187.4800 ;
        RECT 253.4400 1192.4400 255.0400 1192.9200 ;
        RECT 241.6800 1192.4400 244.6800 1192.9200 ;
        RECT 241.6800 1187.0000 244.6800 1187.4800 ;
        RECT 241.6800 1197.8800 244.6800 1198.3600 ;
        RECT 253.4400 1197.8800 255.0400 1198.3600 ;
        RECT 253.4400 1176.1200 255.0400 1176.6000 ;
        RECT 253.4400 1181.5600 255.0400 1182.0400 ;
        RECT 241.6800 1181.5600 244.6800 1182.0400 ;
        RECT 241.6800 1176.1200 244.6800 1176.6000 ;
        RECT 253.4400 1159.8000 255.0400 1160.2800 ;
        RECT 253.4400 1165.2400 255.0400 1165.7200 ;
        RECT 241.6800 1165.2400 244.6800 1165.7200 ;
        RECT 241.6800 1159.8000 244.6800 1160.2800 ;
        RECT 241.6800 1170.6800 244.6800 1171.1600 ;
        RECT 253.4400 1170.6800 255.0400 1171.1600 ;
        RECT 343.4400 1143.4800 345.0400 1143.9600 ;
        RECT 343.4400 1148.9200 345.0400 1149.4000 ;
        RECT 343.4400 1154.3600 345.0400 1154.8400 ;
        RECT 343.4400 1132.6000 345.0400 1133.0800 ;
        RECT 343.4400 1138.0400 345.0400 1138.5200 ;
        RECT 298.4400 1143.4800 300.0400 1143.9600 ;
        RECT 298.4400 1148.9200 300.0400 1149.4000 ;
        RECT 298.4400 1154.3600 300.0400 1154.8400 ;
        RECT 298.4400 1132.6000 300.0400 1133.0800 ;
        RECT 298.4400 1138.0400 300.0400 1138.5200 ;
        RECT 343.4400 1116.2800 345.0400 1116.7600 ;
        RECT 343.4400 1121.7200 345.0400 1122.2000 ;
        RECT 343.4400 1127.1600 345.0400 1127.6400 ;
        RECT 343.4400 1105.4000 345.0400 1105.8800 ;
        RECT 343.4400 1110.8400 345.0400 1111.3200 ;
        RECT 298.4400 1116.2800 300.0400 1116.7600 ;
        RECT 298.4400 1121.7200 300.0400 1122.2000 ;
        RECT 298.4400 1127.1600 300.0400 1127.6400 ;
        RECT 298.4400 1105.4000 300.0400 1105.8800 ;
        RECT 298.4400 1110.8400 300.0400 1111.3200 ;
        RECT 253.4400 1143.4800 255.0400 1143.9600 ;
        RECT 253.4400 1148.9200 255.0400 1149.4000 ;
        RECT 253.4400 1154.3600 255.0400 1154.8400 ;
        RECT 241.6800 1143.4800 244.6800 1143.9600 ;
        RECT 241.6800 1148.9200 244.6800 1149.4000 ;
        RECT 241.6800 1154.3600 244.6800 1154.8400 ;
        RECT 253.4400 1132.6000 255.0400 1133.0800 ;
        RECT 253.4400 1138.0400 255.0400 1138.5200 ;
        RECT 241.6800 1132.6000 244.6800 1133.0800 ;
        RECT 241.6800 1138.0400 244.6800 1138.5200 ;
        RECT 253.4400 1116.2800 255.0400 1116.7600 ;
        RECT 253.4400 1121.7200 255.0400 1122.2000 ;
        RECT 253.4400 1127.1600 255.0400 1127.6400 ;
        RECT 241.6800 1116.2800 244.6800 1116.7600 ;
        RECT 241.6800 1121.7200 244.6800 1122.2000 ;
        RECT 241.6800 1127.1600 244.6800 1127.6400 ;
        RECT 253.4400 1105.4000 255.0400 1105.8800 ;
        RECT 253.4400 1110.8400 255.0400 1111.3200 ;
        RECT 241.6800 1105.4000 244.6800 1105.8800 ;
        RECT 241.6800 1110.8400 244.6800 1111.3200 ;
        RECT 445.7800 1089.0800 448.7800 1089.5600 ;
        RECT 445.7800 1094.5200 448.7800 1095.0000 ;
        RECT 445.7800 1099.9600 448.7800 1100.4400 ;
        RECT 433.4400 1089.0800 435.0400 1089.5600 ;
        RECT 433.4400 1094.5200 435.0400 1095.0000 ;
        RECT 433.4400 1099.9600 435.0400 1100.4400 ;
        RECT 445.7800 1078.2000 448.7800 1078.6800 ;
        RECT 445.7800 1083.6400 448.7800 1084.1200 ;
        RECT 433.4400 1078.2000 435.0400 1078.6800 ;
        RECT 433.4400 1083.6400 435.0400 1084.1200 ;
        RECT 445.7800 1061.8800 448.7800 1062.3600 ;
        RECT 445.7800 1067.3200 448.7800 1067.8000 ;
        RECT 445.7800 1072.7600 448.7800 1073.2400 ;
        RECT 433.4400 1061.8800 435.0400 1062.3600 ;
        RECT 433.4400 1067.3200 435.0400 1067.8000 ;
        RECT 433.4400 1072.7600 435.0400 1073.2400 ;
        RECT 445.7800 1051.0000 448.7800 1051.4800 ;
        RECT 445.7800 1056.4400 448.7800 1056.9200 ;
        RECT 433.4400 1051.0000 435.0400 1051.4800 ;
        RECT 433.4400 1056.4400 435.0400 1056.9200 ;
        RECT 388.4400 1089.0800 390.0400 1089.5600 ;
        RECT 388.4400 1094.5200 390.0400 1095.0000 ;
        RECT 388.4400 1099.9600 390.0400 1100.4400 ;
        RECT 388.4400 1078.2000 390.0400 1078.6800 ;
        RECT 388.4400 1083.6400 390.0400 1084.1200 ;
        RECT 388.4400 1061.8800 390.0400 1062.3600 ;
        RECT 388.4400 1067.3200 390.0400 1067.8000 ;
        RECT 388.4400 1072.7600 390.0400 1073.2400 ;
        RECT 388.4400 1051.0000 390.0400 1051.4800 ;
        RECT 388.4400 1056.4400 390.0400 1056.9200 ;
        RECT 445.7800 1034.6800 448.7800 1035.1600 ;
        RECT 445.7800 1040.1200 448.7800 1040.6000 ;
        RECT 445.7800 1045.5600 448.7800 1046.0400 ;
        RECT 433.4400 1034.6800 435.0400 1035.1600 ;
        RECT 433.4400 1040.1200 435.0400 1040.6000 ;
        RECT 433.4400 1045.5600 435.0400 1046.0400 ;
        RECT 445.7800 1023.8000 448.7800 1024.2800 ;
        RECT 445.7800 1029.2400 448.7800 1029.7200 ;
        RECT 433.4400 1023.8000 435.0400 1024.2800 ;
        RECT 433.4400 1029.2400 435.0400 1029.7200 ;
        RECT 445.7800 1007.4800 448.7800 1007.9600 ;
        RECT 445.7800 1012.9200 448.7800 1013.4000 ;
        RECT 445.7800 1018.3600 448.7800 1018.8400 ;
        RECT 433.4400 1007.4800 435.0400 1007.9600 ;
        RECT 433.4400 1012.9200 435.0400 1013.4000 ;
        RECT 433.4400 1018.3600 435.0400 1018.8400 ;
        RECT 445.7800 1002.0400 448.7800 1002.5200 ;
        RECT 433.4400 1002.0400 435.0400 1002.5200 ;
        RECT 388.4400 1034.6800 390.0400 1035.1600 ;
        RECT 388.4400 1040.1200 390.0400 1040.6000 ;
        RECT 388.4400 1045.5600 390.0400 1046.0400 ;
        RECT 388.4400 1023.8000 390.0400 1024.2800 ;
        RECT 388.4400 1029.2400 390.0400 1029.7200 ;
        RECT 388.4400 1007.4800 390.0400 1007.9600 ;
        RECT 388.4400 1012.9200 390.0400 1013.4000 ;
        RECT 388.4400 1018.3600 390.0400 1018.8400 ;
        RECT 388.4400 1002.0400 390.0400 1002.5200 ;
        RECT 343.4400 1089.0800 345.0400 1089.5600 ;
        RECT 343.4400 1094.5200 345.0400 1095.0000 ;
        RECT 343.4400 1099.9600 345.0400 1100.4400 ;
        RECT 343.4400 1078.2000 345.0400 1078.6800 ;
        RECT 343.4400 1083.6400 345.0400 1084.1200 ;
        RECT 298.4400 1089.0800 300.0400 1089.5600 ;
        RECT 298.4400 1094.5200 300.0400 1095.0000 ;
        RECT 298.4400 1099.9600 300.0400 1100.4400 ;
        RECT 298.4400 1078.2000 300.0400 1078.6800 ;
        RECT 298.4400 1083.6400 300.0400 1084.1200 ;
        RECT 343.4400 1061.8800 345.0400 1062.3600 ;
        RECT 343.4400 1067.3200 345.0400 1067.8000 ;
        RECT 343.4400 1072.7600 345.0400 1073.2400 ;
        RECT 343.4400 1051.0000 345.0400 1051.4800 ;
        RECT 343.4400 1056.4400 345.0400 1056.9200 ;
        RECT 298.4400 1061.8800 300.0400 1062.3600 ;
        RECT 298.4400 1067.3200 300.0400 1067.8000 ;
        RECT 298.4400 1072.7600 300.0400 1073.2400 ;
        RECT 298.4400 1051.0000 300.0400 1051.4800 ;
        RECT 298.4400 1056.4400 300.0400 1056.9200 ;
        RECT 253.4400 1089.0800 255.0400 1089.5600 ;
        RECT 253.4400 1094.5200 255.0400 1095.0000 ;
        RECT 253.4400 1099.9600 255.0400 1100.4400 ;
        RECT 241.6800 1089.0800 244.6800 1089.5600 ;
        RECT 241.6800 1094.5200 244.6800 1095.0000 ;
        RECT 241.6800 1099.9600 244.6800 1100.4400 ;
        RECT 253.4400 1078.2000 255.0400 1078.6800 ;
        RECT 253.4400 1083.6400 255.0400 1084.1200 ;
        RECT 241.6800 1078.2000 244.6800 1078.6800 ;
        RECT 241.6800 1083.6400 244.6800 1084.1200 ;
        RECT 253.4400 1061.8800 255.0400 1062.3600 ;
        RECT 253.4400 1067.3200 255.0400 1067.8000 ;
        RECT 253.4400 1072.7600 255.0400 1073.2400 ;
        RECT 241.6800 1061.8800 244.6800 1062.3600 ;
        RECT 241.6800 1067.3200 244.6800 1067.8000 ;
        RECT 241.6800 1072.7600 244.6800 1073.2400 ;
        RECT 253.4400 1051.0000 255.0400 1051.4800 ;
        RECT 253.4400 1056.4400 255.0400 1056.9200 ;
        RECT 241.6800 1051.0000 244.6800 1051.4800 ;
        RECT 241.6800 1056.4400 244.6800 1056.9200 ;
        RECT 343.4400 1034.6800 345.0400 1035.1600 ;
        RECT 343.4400 1040.1200 345.0400 1040.6000 ;
        RECT 343.4400 1045.5600 345.0400 1046.0400 ;
        RECT 343.4400 1023.8000 345.0400 1024.2800 ;
        RECT 343.4400 1029.2400 345.0400 1029.7200 ;
        RECT 298.4400 1034.6800 300.0400 1035.1600 ;
        RECT 298.4400 1040.1200 300.0400 1040.6000 ;
        RECT 298.4400 1045.5600 300.0400 1046.0400 ;
        RECT 298.4400 1023.8000 300.0400 1024.2800 ;
        RECT 298.4400 1029.2400 300.0400 1029.7200 ;
        RECT 343.4400 1007.4800 345.0400 1007.9600 ;
        RECT 343.4400 1012.9200 345.0400 1013.4000 ;
        RECT 343.4400 1018.3600 345.0400 1018.8400 ;
        RECT 343.4400 1002.0400 345.0400 1002.5200 ;
        RECT 298.4400 1007.4800 300.0400 1007.9600 ;
        RECT 298.4400 1012.9200 300.0400 1013.4000 ;
        RECT 298.4400 1018.3600 300.0400 1018.8400 ;
        RECT 298.4400 1002.0400 300.0400 1002.5200 ;
        RECT 253.4400 1034.6800 255.0400 1035.1600 ;
        RECT 253.4400 1040.1200 255.0400 1040.6000 ;
        RECT 253.4400 1045.5600 255.0400 1046.0400 ;
        RECT 241.6800 1034.6800 244.6800 1035.1600 ;
        RECT 241.6800 1040.1200 244.6800 1040.6000 ;
        RECT 241.6800 1045.5600 244.6800 1046.0400 ;
        RECT 253.4400 1023.8000 255.0400 1024.2800 ;
        RECT 253.4400 1029.2400 255.0400 1029.7200 ;
        RECT 241.6800 1023.8000 244.6800 1024.2800 ;
        RECT 241.6800 1029.2400 244.6800 1029.7200 ;
        RECT 253.4400 1007.4800 255.0400 1007.9600 ;
        RECT 253.4400 1012.9200 255.0400 1013.4000 ;
        RECT 253.4400 1018.3600 255.0400 1018.8400 ;
        RECT 241.6800 1007.4800 244.6800 1007.9600 ;
        RECT 241.6800 1012.9200 244.6800 1013.4000 ;
        RECT 241.6800 1018.3600 244.6800 1018.8400 ;
        RECT 241.6800 1002.0400 244.6800 1002.5200 ;
        RECT 253.4400 1002.0400 255.0400 1002.5200 ;
        RECT 241.6800 1206.9500 448.7800 1209.9500 ;
        RECT 241.6800 993.8500 448.7800 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 433.4400 764.2100 435.0400 980.3100 ;
        RECT 388.4400 764.2100 390.0400 980.3100 ;
        RECT 343.4400 764.2100 345.0400 980.3100 ;
        RECT 298.4400 764.2100 300.0400 980.3100 ;
        RECT 253.4400 764.2100 255.0400 980.3100 ;
        RECT 445.7800 764.2100 448.7800 980.3100 ;
        RECT 241.6800 764.2100 244.6800 980.3100 ;
      LAYER met3 ;
        RECT 445.7800 957.3600 448.7800 957.8400 ;
        RECT 445.7800 962.8000 448.7800 963.2800 ;
        RECT 433.4400 957.3600 435.0400 957.8400 ;
        RECT 433.4400 962.8000 435.0400 963.2800 ;
        RECT 445.7800 968.2400 448.7800 968.7200 ;
        RECT 433.4400 968.2400 435.0400 968.7200 ;
        RECT 445.7800 946.4800 448.7800 946.9600 ;
        RECT 445.7800 951.9200 448.7800 952.4000 ;
        RECT 433.4400 946.4800 435.0400 946.9600 ;
        RECT 433.4400 951.9200 435.0400 952.4000 ;
        RECT 445.7800 930.1600 448.7800 930.6400 ;
        RECT 445.7800 935.6000 448.7800 936.0800 ;
        RECT 433.4400 930.1600 435.0400 930.6400 ;
        RECT 433.4400 935.6000 435.0400 936.0800 ;
        RECT 445.7800 941.0400 448.7800 941.5200 ;
        RECT 433.4400 941.0400 435.0400 941.5200 ;
        RECT 388.4400 957.3600 390.0400 957.8400 ;
        RECT 388.4400 962.8000 390.0400 963.2800 ;
        RECT 388.4400 968.2400 390.0400 968.7200 ;
        RECT 388.4400 946.4800 390.0400 946.9600 ;
        RECT 388.4400 951.9200 390.0400 952.4000 ;
        RECT 388.4400 930.1600 390.0400 930.6400 ;
        RECT 388.4400 935.6000 390.0400 936.0800 ;
        RECT 388.4400 941.0400 390.0400 941.5200 ;
        RECT 445.7800 913.8400 448.7800 914.3200 ;
        RECT 445.7800 919.2800 448.7800 919.7600 ;
        RECT 445.7800 924.7200 448.7800 925.2000 ;
        RECT 433.4400 913.8400 435.0400 914.3200 ;
        RECT 433.4400 919.2800 435.0400 919.7600 ;
        RECT 433.4400 924.7200 435.0400 925.2000 ;
        RECT 445.7800 902.9600 448.7800 903.4400 ;
        RECT 445.7800 908.4000 448.7800 908.8800 ;
        RECT 433.4400 902.9600 435.0400 903.4400 ;
        RECT 433.4400 908.4000 435.0400 908.8800 ;
        RECT 445.7800 886.6400 448.7800 887.1200 ;
        RECT 445.7800 892.0800 448.7800 892.5600 ;
        RECT 445.7800 897.5200 448.7800 898.0000 ;
        RECT 433.4400 886.6400 435.0400 887.1200 ;
        RECT 433.4400 892.0800 435.0400 892.5600 ;
        RECT 433.4400 897.5200 435.0400 898.0000 ;
        RECT 445.7800 875.7600 448.7800 876.2400 ;
        RECT 445.7800 881.2000 448.7800 881.6800 ;
        RECT 433.4400 875.7600 435.0400 876.2400 ;
        RECT 433.4400 881.2000 435.0400 881.6800 ;
        RECT 388.4400 913.8400 390.0400 914.3200 ;
        RECT 388.4400 919.2800 390.0400 919.7600 ;
        RECT 388.4400 924.7200 390.0400 925.2000 ;
        RECT 388.4400 902.9600 390.0400 903.4400 ;
        RECT 388.4400 908.4000 390.0400 908.8800 ;
        RECT 388.4400 886.6400 390.0400 887.1200 ;
        RECT 388.4400 892.0800 390.0400 892.5600 ;
        RECT 388.4400 897.5200 390.0400 898.0000 ;
        RECT 388.4400 875.7600 390.0400 876.2400 ;
        RECT 388.4400 881.2000 390.0400 881.6800 ;
        RECT 343.4400 957.3600 345.0400 957.8400 ;
        RECT 343.4400 962.8000 345.0400 963.2800 ;
        RECT 343.4400 968.2400 345.0400 968.7200 ;
        RECT 298.4400 957.3600 300.0400 957.8400 ;
        RECT 298.4400 962.8000 300.0400 963.2800 ;
        RECT 298.4400 968.2400 300.0400 968.7200 ;
        RECT 343.4400 946.4800 345.0400 946.9600 ;
        RECT 343.4400 951.9200 345.0400 952.4000 ;
        RECT 343.4400 930.1600 345.0400 930.6400 ;
        RECT 343.4400 935.6000 345.0400 936.0800 ;
        RECT 343.4400 941.0400 345.0400 941.5200 ;
        RECT 298.4400 946.4800 300.0400 946.9600 ;
        RECT 298.4400 951.9200 300.0400 952.4000 ;
        RECT 298.4400 930.1600 300.0400 930.6400 ;
        RECT 298.4400 935.6000 300.0400 936.0800 ;
        RECT 298.4400 941.0400 300.0400 941.5200 ;
        RECT 253.4400 957.3600 255.0400 957.8400 ;
        RECT 253.4400 962.8000 255.0400 963.2800 ;
        RECT 241.6800 962.8000 244.6800 963.2800 ;
        RECT 241.6800 957.3600 244.6800 957.8400 ;
        RECT 241.6800 968.2400 244.6800 968.7200 ;
        RECT 253.4400 968.2400 255.0400 968.7200 ;
        RECT 253.4400 946.4800 255.0400 946.9600 ;
        RECT 253.4400 951.9200 255.0400 952.4000 ;
        RECT 241.6800 951.9200 244.6800 952.4000 ;
        RECT 241.6800 946.4800 244.6800 946.9600 ;
        RECT 253.4400 930.1600 255.0400 930.6400 ;
        RECT 253.4400 935.6000 255.0400 936.0800 ;
        RECT 241.6800 935.6000 244.6800 936.0800 ;
        RECT 241.6800 930.1600 244.6800 930.6400 ;
        RECT 241.6800 941.0400 244.6800 941.5200 ;
        RECT 253.4400 941.0400 255.0400 941.5200 ;
        RECT 343.4400 913.8400 345.0400 914.3200 ;
        RECT 343.4400 919.2800 345.0400 919.7600 ;
        RECT 343.4400 924.7200 345.0400 925.2000 ;
        RECT 343.4400 902.9600 345.0400 903.4400 ;
        RECT 343.4400 908.4000 345.0400 908.8800 ;
        RECT 298.4400 913.8400 300.0400 914.3200 ;
        RECT 298.4400 919.2800 300.0400 919.7600 ;
        RECT 298.4400 924.7200 300.0400 925.2000 ;
        RECT 298.4400 902.9600 300.0400 903.4400 ;
        RECT 298.4400 908.4000 300.0400 908.8800 ;
        RECT 343.4400 886.6400 345.0400 887.1200 ;
        RECT 343.4400 892.0800 345.0400 892.5600 ;
        RECT 343.4400 897.5200 345.0400 898.0000 ;
        RECT 343.4400 875.7600 345.0400 876.2400 ;
        RECT 343.4400 881.2000 345.0400 881.6800 ;
        RECT 298.4400 886.6400 300.0400 887.1200 ;
        RECT 298.4400 892.0800 300.0400 892.5600 ;
        RECT 298.4400 897.5200 300.0400 898.0000 ;
        RECT 298.4400 875.7600 300.0400 876.2400 ;
        RECT 298.4400 881.2000 300.0400 881.6800 ;
        RECT 253.4400 913.8400 255.0400 914.3200 ;
        RECT 253.4400 919.2800 255.0400 919.7600 ;
        RECT 253.4400 924.7200 255.0400 925.2000 ;
        RECT 241.6800 913.8400 244.6800 914.3200 ;
        RECT 241.6800 919.2800 244.6800 919.7600 ;
        RECT 241.6800 924.7200 244.6800 925.2000 ;
        RECT 253.4400 902.9600 255.0400 903.4400 ;
        RECT 253.4400 908.4000 255.0400 908.8800 ;
        RECT 241.6800 902.9600 244.6800 903.4400 ;
        RECT 241.6800 908.4000 244.6800 908.8800 ;
        RECT 253.4400 886.6400 255.0400 887.1200 ;
        RECT 253.4400 892.0800 255.0400 892.5600 ;
        RECT 253.4400 897.5200 255.0400 898.0000 ;
        RECT 241.6800 886.6400 244.6800 887.1200 ;
        RECT 241.6800 892.0800 244.6800 892.5600 ;
        RECT 241.6800 897.5200 244.6800 898.0000 ;
        RECT 253.4400 875.7600 255.0400 876.2400 ;
        RECT 253.4400 881.2000 255.0400 881.6800 ;
        RECT 241.6800 875.7600 244.6800 876.2400 ;
        RECT 241.6800 881.2000 244.6800 881.6800 ;
        RECT 445.7800 859.4400 448.7800 859.9200 ;
        RECT 445.7800 864.8800 448.7800 865.3600 ;
        RECT 445.7800 870.3200 448.7800 870.8000 ;
        RECT 433.4400 859.4400 435.0400 859.9200 ;
        RECT 433.4400 864.8800 435.0400 865.3600 ;
        RECT 433.4400 870.3200 435.0400 870.8000 ;
        RECT 445.7800 848.5600 448.7800 849.0400 ;
        RECT 445.7800 854.0000 448.7800 854.4800 ;
        RECT 433.4400 848.5600 435.0400 849.0400 ;
        RECT 433.4400 854.0000 435.0400 854.4800 ;
        RECT 445.7800 832.2400 448.7800 832.7200 ;
        RECT 445.7800 837.6800 448.7800 838.1600 ;
        RECT 445.7800 843.1200 448.7800 843.6000 ;
        RECT 433.4400 832.2400 435.0400 832.7200 ;
        RECT 433.4400 837.6800 435.0400 838.1600 ;
        RECT 433.4400 843.1200 435.0400 843.6000 ;
        RECT 445.7800 821.3600 448.7800 821.8400 ;
        RECT 445.7800 826.8000 448.7800 827.2800 ;
        RECT 433.4400 821.3600 435.0400 821.8400 ;
        RECT 433.4400 826.8000 435.0400 827.2800 ;
        RECT 388.4400 859.4400 390.0400 859.9200 ;
        RECT 388.4400 864.8800 390.0400 865.3600 ;
        RECT 388.4400 870.3200 390.0400 870.8000 ;
        RECT 388.4400 848.5600 390.0400 849.0400 ;
        RECT 388.4400 854.0000 390.0400 854.4800 ;
        RECT 388.4400 832.2400 390.0400 832.7200 ;
        RECT 388.4400 837.6800 390.0400 838.1600 ;
        RECT 388.4400 843.1200 390.0400 843.6000 ;
        RECT 388.4400 821.3600 390.0400 821.8400 ;
        RECT 388.4400 826.8000 390.0400 827.2800 ;
        RECT 445.7800 805.0400 448.7800 805.5200 ;
        RECT 445.7800 810.4800 448.7800 810.9600 ;
        RECT 445.7800 815.9200 448.7800 816.4000 ;
        RECT 433.4400 805.0400 435.0400 805.5200 ;
        RECT 433.4400 810.4800 435.0400 810.9600 ;
        RECT 433.4400 815.9200 435.0400 816.4000 ;
        RECT 445.7800 794.1600 448.7800 794.6400 ;
        RECT 445.7800 799.6000 448.7800 800.0800 ;
        RECT 433.4400 794.1600 435.0400 794.6400 ;
        RECT 433.4400 799.6000 435.0400 800.0800 ;
        RECT 445.7800 777.8400 448.7800 778.3200 ;
        RECT 445.7800 783.2800 448.7800 783.7600 ;
        RECT 445.7800 788.7200 448.7800 789.2000 ;
        RECT 433.4400 777.8400 435.0400 778.3200 ;
        RECT 433.4400 783.2800 435.0400 783.7600 ;
        RECT 433.4400 788.7200 435.0400 789.2000 ;
        RECT 445.7800 772.4000 448.7800 772.8800 ;
        RECT 433.4400 772.4000 435.0400 772.8800 ;
        RECT 388.4400 805.0400 390.0400 805.5200 ;
        RECT 388.4400 810.4800 390.0400 810.9600 ;
        RECT 388.4400 815.9200 390.0400 816.4000 ;
        RECT 388.4400 794.1600 390.0400 794.6400 ;
        RECT 388.4400 799.6000 390.0400 800.0800 ;
        RECT 388.4400 777.8400 390.0400 778.3200 ;
        RECT 388.4400 783.2800 390.0400 783.7600 ;
        RECT 388.4400 788.7200 390.0400 789.2000 ;
        RECT 388.4400 772.4000 390.0400 772.8800 ;
        RECT 343.4400 859.4400 345.0400 859.9200 ;
        RECT 343.4400 864.8800 345.0400 865.3600 ;
        RECT 343.4400 870.3200 345.0400 870.8000 ;
        RECT 343.4400 848.5600 345.0400 849.0400 ;
        RECT 343.4400 854.0000 345.0400 854.4800 ;
        RECT 298.4400 859.4400 300.0400 859.9200 ;
        RECT 298.4400 864.8800 300.0400 865.3600 ;
        RECT 298.4400 870.3200 300.0400 870.8000 ;
        RECT 298.4400 848.5600 300.0400 849.0400 ;
        RECT 298.4400 854.0000 300.0400 854.4800 ;
        RECT 343.4400 832.2400 345.0400 832.7200 ;
        RECT 343.4400 837.6800 345.0400 838.1600 ;
        RECT 343.4400 843.1200 345.0400 843.6000 ;
        RECT 343.4400 821.3600 345.0400 821.8400 ;
        RECT 343.4400 826.8000 345.0400 827.2800 ;
        RECT 298.4400 832.2400 300.0400 832.7200 ;
        RECT 298.4400 837.6800 300.0400 838.1600 ;
        RECT 298.4400 843.1200 300.0400 843.6000 ;
        RECT 298.4400 821.3600 300.0400 821.8400 ;
        RECT 298.4400 826.8000 300.0400 827.2800 ;
        RECT 253.4400 859.4400 255.0400 859.9200 ;
        RECT 253.4400 864.8800 255.0400 865.3600 ;
        RECT 253.4400 870.3200 255.0400 870.8000 ;
        RECT 241.6800 859.4400 244.6800 859.9200 ;
        RECT 241.6800 864.8800 244.6800 865.3600 ;
        RECT 241.6800 870.3200 244.6800 870.8000 ;
        RECT 253.4400 848.5600 255.0400 849.0400 ;
        RECT 253.4400 854.0000 255.0400 854.4800 ;
        RECT 241.6800 848.5600 244.6800 849.0400 ;
        RECT 241.6800 854.0000 244.6800 854.4800 ;
        RECT 253.4400 832.2400 255.0400 832.7200 ;
        RECT 253.4400 837.6800 255.0400 838.1600 ;
        RECT 253.4400 843.1200 255.0400 843.6000 ;
        RECT 241.6800 832.2400 244.6800 832.7200 ;
        RECT 241.6800 837.6800 244.6800 838.1600 ;
        RECT 241.6800 843.1200 244.6800 843.6000 ;
        RECT 253.4400 821.3600 255.0400 821.8400 ;
        RECT 253.4400 826.8000 255.0400 827.2800 ;
        RECT 241.6800 821.3600 244.6800 821.8400 ;
        RECT 241.6800 826.8000 244.6800 827.2800 ;
        RECT 343.4400 805.0400 345.0400 805.5200 ;
        RECT 343.4400 810.4800 345.0400 810.9600 ;
        RECT 343.4400 815.9200 345.0400 816.4000 ;
        RECT 343.4400 794.1600 345.0400 794.6400 ;
        RECT 343.4400 799.6000 345.0400 800.0800 ;
        RECT 298.4400 805.0400 300.0400 805.5200 ;
        RECT 298.4400 810.4800 300.0400 810.9600 ;
        RECT 298.4400 815.9200 300.0400 816.4000 ;
        RECT 298.4400 794.1600 300.0400 794.6400 ;
        RECT 298.4400 799.6000 300.0400 800.0800 ;
        RECT 343.4400 777.8400 345.0400 778.3200 ;
        RECT 343.4400 783.2800 345.0400 783.7600 ;
        RECT 343.4400 788.7200 345.0400 789.2000 ;
        RECT 343.4400 772.4000 345.0400 772.8800 ;
        RECT 298.4400 777.8400 300.0400 778.3200 ;
        RECT 298.4400 783.2800 300.0400 783.7600 ;
        RECT 298.4400 788.7200 300.0400 789.2000 ;
        RECT 298.4400 772.4000 300.0400 772.8800 ;
        RECT 253.4400 805.0400 255.0400 805.5200 ;
        RECT 253.4400 810.4800 255.0400 810.9600 ;
        RECT 253.4400 815.9200 255.0400 816.4000 ;
        RECT 241.6800 805.0400 244.6800 805.5200 ;
        RECT 241.6800 810.4800 244.6800 810.9600 ;
        RECT 241.6800 815.9200 244.6800 816.4000 ;
        RECT 253.4400 794.1600 255.0400 794.6400 ;
        RECT 253.4400 799.6000 255.0400 800.0800 ;
        RECT 241.6800 794.1600 244.6800 794.6400 ;
        RECT 241.6800 799.6000 244.6800 800.0800 ;
        RECT 253.4400 777.8400 255.0400 778.3200 ;
        RECT 253.4400 783.2800 255.0400 783.7600 ;
        RECT 253.4400 788.7200 255.0400 789.2000 ;
        RECT 241.6800 777.8400 244.6800 778.3200 ;
        RECT 241.6800 783.2800 244.6800 783.7600 ;
        RECT 241.6800 788.7200 244.6800 789.2000 ;
        RECT 241.6800 772.4000 244.6800 772.8800 ;
        RECT 253.4400 772.4000 255.0400 772.8800 ;
        RECT 241.6800 977.3100 448.7800 980.3100 ;
        RECT 241.6800 764.2100 448.7800 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 462.9000 2830.6100 464.9000 2857.5400 ;
        RECT 666.0000 2830.6100 668.0000 2857.5400 ;
      LAYER met3 ;
        RECT 666.0000 2847.3200 668.0000 2847.8000 ;
        RECT 462.9000 2847.3200 464.9000 2847.8000 ;
        RECT 666.0000 2841.8800 668.0000 2842.3600 ;
        RECT 666.0000 2836.4400 668.0000 2836.9200 ;
        RECT 462.9000 2841.8800 464.9000 2842.3600 ;
        RECT 462.9000 2836.4400 464.9000 2836.9200 ;
        RECT 462.9000 2855.5400 668.0000 2857.5400 ;
        RECT 462.9000 2830.6100 668.0000 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 534.5700 655.2600 750.6700 ;
        RECT 608.6600 534.5700 610.2600 750.6700 ;
        RECT 563.6600 534.5700 565.2600 750.6700 ;
        RECT 518.6600 534.5700 520.2600 750.6700 ;
        RECT 473.6600 534.5700 475.2600 750.6700 ;
        RECT 666.0000 534.5700 669.0000 750.6700 ;
        RECT 461.9000 534.5700 464.9000 750.6700 ;
      LAYER met3 ;
        RECT 666.0000 727.7200 669.0000 728.2000 ;
        RECT 666.0000 733.1600 669.0000 733.6400 ;
        RECT 653.6600 727.7200 655.2600 728.2000 ;
        RECT 653.6600 733.1600 655.2600 733.6400 ;
        RECT 666.0000 738.6000 669.0000 739.0800 ;
        RECT 653.6600 738.6000 655.2600 739.0800 ;
        RECT 666.0000 716.8400 669.0000 717.3200 ;
        RECT 666.0000 722.2800 669.0000 722.7600 ;
        RECT 653.6600 716.8400 655.2600 717.3200 ;
        RECT 653.6600 722.2800 655.2600 722.7600 ;
        RECT 666.0000 700.5200 669.0000 701.0000 ;
        RECT 666.0000 705.9600 669.0000 706.4400 ;
        RECT 653.6600 700.5200 655.2600 701.0000 ;
        RECT 653.6600 705.9600 655.2600 706.4400 ;
        RECT 666.0000 711.4000 669.0000 711.8800 ;
        RECT 653.6600 711.4000 655.2600 711.8800 ;
        RECT 608.6600 727.7200 610.2600 728.2000 ;
        RECT 608.6600 733.1600 610.2600 733.6400 ;
        RECT 608.6600 738.6000 610.2600 739.0800 ;
        RECT 608.6600 716.8400 610.2600 717.3200 ;
        RECT 608.6600 722.2800 610.2600 722.7600 ;
        RECT 608.6600 700.5200 610.2600 701.0000 ;
        RECT 608.6600 705.9600 610.2600 706.4400 ;
        RECT 608.6600 711.4000 610.2600 711.8800 ;
        RECT 666.0000 684.2000 669.0000 684.6800 ;
        RECT 666.0000 689.6400 669.0000 690.1200 ;
        RECT 666.0000 695.0800 669.0000 695.5600 ;
        RECT 653.6600 684.2000 655.2600 684.6800 ;
        RECT 653.6600 689.6400 655.2600 690.1200 ;
        RECT 653.6600 695.0800 655.2600 695.5600 ;
        RECT 666.0000 673.3200 669.0000 673.8000 ;
        RECT 666.0000 678.7600 669.0000 679.2400 ;
        RECT 653.6600 673.3200 655.2600 673.8000 ;
        RECT 653.6600 678.7600 655.2600 679.2400 ;
        RECT 666.0000 657.0000 669.0000 657.4800 ;
        RECT 666.0000 662.4400 669.0000 662.9200 ;
        RECT 666.0000 667.8800 669.0000 668.3600 ;
        RECT 653.6600 657.0000 655.2600 657.4800 ;
        RECT 653.6600 662.4400 655.2600 662.9200 ;
        RECT 653.6600 667.8800 655.2600 668.3600 ;
        RECT 666.0000 646.1200 669.0000 646.6000 ;
        RECT 666.0000 651.5600 669.0000 652.0400 ;
        RECT 653.6600 646.1200 655.2600 646.6000 ;
        RECT 653.6600 651.5600 655.2600 652.0400 ;
        RECT 608.6600 684.2000 610.2600 684.6800 ;
        RECT 608.6600 689.6400 610.2600 690.1200 ;
        RECT 608.6600 695.0800 610.2600 695.5600 ;
        RECT 608.6600 673.3200 610.2600 673.8000 ;
        RECT 608.6600 678.7600 610.2600 679.2400 ;
        RECT 608.6600 657.0000 610.2600 657.4800 ;
        RECT 608.6600 662.4400 610.2600 662.9200 ;
        RECT 608.6600 667.8800 610.2600 668.3600 ;
        RECT 608.6600 646.1200 610.2600 646.6000 ;
        RECT 608.6600 651.5600 610.2600 652.0400 ;
        RECT 563.6600 727.7200 565.2600 728.2000 ;
        RECT 563.6600 733.1600 565.2600 733.6400 ;
        RECT 563.6600 738.6000 565.2600 739.0800 ;
        RECT 518.6600 727.7200 520.2600 728.2000 ;
        RECT 518.6600 733.1600 520.2600 733.6400 ;
        RECT 518.6600 738.6000 520.2600 739.0800 ;
        RECT 563.6600 716.8400 565.2600 717.3200 ;
        RECT 563.6600 722.2800 565.2600 722.7600 ;
        RECT 563.6600 700.5200 565.2600 701.0000 ;
        RECT 563.6600 705.9600 565.2600 706.4400 ;
        RECT 563.6600 711.4000 565.2600 711.8800 ;
        RECT 518.6600 716.8400 520.2600 717.3200 ;
        RECT 518.6600 722.2800 520.2600 722.7600 ;
        RECT 518.6600 700.5200 520.2600 701.0000 ;
        RECT 518.6600 705.9600 520.2600 706.4400 ;
        RECT 518.6600 711.4000 520.2600 711.8800 ;
        RECT 473.6600 727.7200 475.2600 728.2000 ;
        RECT 473.6600 733.1600 475.2600 733.6400 ;
        RECT 461.9000 733.1600 464.9000 733.6400 ;
        RECT 461.9000 727.7200 464.9000 728.2000 ;
        RECT 461.9000 738.6000 464.9000 739.0800 ;
        RECT 473.6600 738.6000 475.2600 739.0800 ;
        RECT 473.6600 716.8400 475.2600 717.3200 ;
        RECT 473.6600 722.2800 475.2600 722.7600 ;
        RECT 461.9000 722.2800 464.9000 722.7600 ;
        RECT 461.9000 716.8400 464.9000 717.3200 ;
        RECT 473.6600 700.5200 475.2600 701.0000 ;
        RECT 473.6600 705.9600 475.2600 706.4400 ;
        RECT 461.9000 705.9600 464.9000 706.4400 ;
        RECT 461.9000 700.5200 464.9000 701.0000 ;
        RECT 461.9000 711.4000 464.9000 711.8800 ;
        RECT 473.6600 711.4000 475.2600 711.8800 ;
        RECT 563.6600 684.2000 565.2600 684.6800 ;
        RECT 563.6600 689.6400 565.2600 690.1200 ;
        RECT 563.6600 695.0800 565.2600 695.5600 ;
        RECT 563.6600 673.3200 565.2600 673.8000 ;
        RECT 563.6600 678.7600 565.2600 679.2400 ;
        RECT 518.6600 684.2000 520.2600 684.6800 ;
        RECT 518.6600 689.6400 520.2600 690.1200 ;
        RECT 518.6600 695.0800 520.2600 695.5600 ;
        RECT 518.6600 673.3200 520.2600 673.8000 ;
        RECT 518.6600 678.7600 520.2600 679.2400 ;
        RECT 563.6600 657.0000 565.2600 657.4800 ;
        RECT 563.6600 662.4400 565.2600 662.9200 ;
        RECT 563.6600 667.8800 565.2600 668.3600 ;
        RECT 563.6600 646.1200 565.2600 646.6000 ;
        RECT 563.6600 651.5600 565.2600 652.0400 ;
        RECT 518.6600 657.0000 520.2600 657.4800 ;
        RECT 518.6600 662.4400 520.2600 662.9200 ;
        RECT 518.6600 667.8800 520.2600 668.3600 ;
        RECT 518.6600 646.1200 520.2600 646.6000 ;
        RECT 518.6600 651.5600 520.2600 652.0400 ;
        RECT 473.6600 684.2000 475.2600 684.6800 ;
        RECT 473.6600 689.6400 475.2600 690.1200 ;
        RECT 473.6600 695.0800 475.2600 695.5600 ;
        RECT 461.9000 684.2000 464.9000 684.6800 ;
        RECT 461.9000 689.6400 464.9000 690.1200 ;
        RECT 461.9000 695.0800 464.9000 695.5600 ;
        RECT 473.6600 673.3200 475.2600 673.8000 ;
        RECT 473.6600 678.7600 475.2600 679.2400 ;
        RECT 461.9000 673.3200 464.9000 673.8000 ;
        RECT 461.9000 678.7600 464.9000 679.2400 ;
        RECT 473.6600 657.0000 475.2600 657.4800 ;
        RECT 473.6600 662.4400 475.2600 662.9200 ;
        RECT 473.6600 667.8800 475.2600 668.3600 ;
        RECT 461.9000 657.0000 464.9000 657.4800 ;
        RECT 461.9000 662.4400 464.9000 662.9200 ;
        RECT 461.9000 667.8800 464.9000 668.3600 ;
        RECT 473.6600 646.1200 475.2600 646.6000 ;
        RECT 473.6600 651.5600 475.2600 652.0400 ;
        RECT 461.9000 646.1200 464.9000 646.6000 ;
        RECT 461.9000 651.5600 464.9000 652.0400 ;
        RECT 666.0000 629.8000 669.0000 630.2800 ;
        RECT 666.0000 635.2400 669.0000 635.7200 ;
        RECT 666.0000 640.6800 669.0000 641.1600 ;
        RECT 653.6600 629.8000 655.2600 630.2800 ;
        RECT 653.6600 635.2400 655.2600 635.7200 ;
        RECT 653.6600 640.6800 655.2600 641.1600 ;
        RECT 666.0000 618.9200 669.0000 619.4000 ;
        RECT 666.0000 624.3600 669.0000 624.8400 ;
        RECT 653.6600 618.9200 655.2600 619.4000 ;
        RECT 653.6600 624.3600 655.2600 624.8400 ;
        RECT 666.0000 602.6000 669.0000 603.0800 ;
        RECT 666.0000 608.0400 669.0000 608.5200 ;
        RECT 666.0000 613.4800 669.0000 613.9600 ;
        RECT 653.6600 602.6000 655.2600 603.0800 ;
        RECT 653.6600 608.0400 655.2600 608.5200 ;
        RECT 653.6600 613.4800 655.2600 613.9600 ;
        RECT 666.0000 591.7200 669.0000 592.2000 ;
        RECT 666.0000 597.1600 669.0000 597.6400 ;
        RECT 653.6600 591.7200 655.2600 592.2000 ;
        RECT 653.6600 597.1600 655.2600 597.6400 ;
        RECT 608.6600 629.8000 610.2600 630.2800 ;
        RECT 608.6600 635.2400 610.2600 635.7200 ;
        RECT 608.6600 640.6800 610.2600 641.1600 ;
        RECT 608.6600 618.9200 610.2600 619.4000 ;
        RECT 608.6600 624.3600 610.2600 624.8400 ;
        RECT 608.6600 602.6000 610.2600 603.0800 ;
        RECT 608.6600 608.0400 610.2600 608.5200 ;
        RECT 608.6600 613.4800 610.2600 613.9600 ;
        RECT 608.6600 591.7200 610.2600 592.2000 ;
        RECT 608.6600 597.1600 610.2600 597.6400 ;
        RECT 666.0000 575.4000 669.0000 575.8800 ;
        RECT 666.0000 580.8400 669.0000 581.3200 ;
        RECT 666.0000 586.2800 669.0000 586.7600 ;
        RECT 653.6600 575.4000 655.2600 575.8800 ;
        RECT 653.6600 580.8400 655.2600 581.3200 ;
        RECT 653.6600 586.2800 655.2600 586.7600 ;
        RECT 666.0000 564.5200 669.0000 565.0000 ;
        RECT 666.0000 569.9600 669.0000 570.4400 ;
        RECT 653.6600 564.5200 655.2600 565.0000 ;
        RECT 653.6600 569.9600 655.2600 570.4400 ;
        RECT 666.0000 548.2000 669.0000 548.6800 ;
        RECT 666.0000 553.6400 669.0000 554.1200 ;
        RECT 666.0000 559.0800 669.0000 559.5600 ;
        RECT 653.6600 548.2000 655.2600 548.6800 ;
        RECT 653.6600 553.6400 655.2600 554.1200 ;
        RECT 653.6600 559.0800 655.2600 559.5600 ;
        RECT 666.0000 542.7600 669.0000 543.2400 ;
        RECT 653.6600 542.7600 655.2600 543.2400 ;
        RECT 608.6600 575.4000 610.2600 575.8800 ;
        RECT 608.6600 580.8400 610.2600 581.3200 ;
        RECT 608.6600 586.2800 610.2600 586.7600 ;
        RECT 608.6600 564.5200 610.2600 565.0000 ;
        RECT 608.6600 569.9600 610.2600 570.4400 ;
        RECT 608.6600 548.2000 610.2600 548.6800 ;
        RECT 608.6600 553.6400 610.2600 554.1200 ;
        RECT 608.6600 559.0800 610.2600 559.5600 ;
        RECT 608.6600 542.7600 610.2600 543.2400 ;
        RECT 563.6600 629.8000 565.2600 630.2800 ;
        RECT 563.6600 635.2400 565.2600 635.7200 ;
        RECT 563.6600 640.6800 565.2600 641.1600 ;
        RECT 563.6600 618.9200 565.2600 619.4000 ;
        RECT 563.6600 624.3600 565.2600 624.8400 ;
        RECT 518.6600 629.8000 520.2600 630.2800 ;
        RECT 518.6600 635.2400 520.2600 635.7200 ;
        RECT 518.6600 640.6800 520.2600 641.1600 ;
        RECT 518.6600 618.9200 520.2600 619.4000 ;
        RECT 518.6600 624.3600 520.2600 624.8400 ;
        RECT 563.6600 602.6000 565.2600 603.0800 ;
        RECT 563.6600 608.0400 565.2600 608.5200 ;
        RECT 563.6600 613.4800 565.2600 613.9600 ;
        RECT 563.6600 591.7200 565.2600 592.2000 ;
        RECT 563.6600 597.1600 565.2600 597.6400 ;
        RECT 518.6600 602.6000 520.2600 603.0800 ;
        RECT 518.6600 608.0400 520.2600 608.5200 ;
        RECT 518.6600 613.4800 520.2600 613.9600 ;
        RECT 518.6600 591.7200 520.2600 592.2000 ;
        RECT 518.6600 597.1600 520.2600 597.6400 ;
        RECT 473.6600 629.8000 475.2600 630.2800 ;
        RECT 473.6600 635.2400 475.2600 635.7200 ;
        RECT 473.6600 640.6800 475.2600 641.1600 ;
        RECT 461.9000 629.8000 464.9000 630.2800 ;
        RECT 461.9000 635.2400 464.9000 635.7200 ;
        RECT 461.9000 640.6800 464.9000 641.1600 ;
        RECT 473.6600 618.9200 475.2600 619.4000 ;
        RECT 473.6600 624.3600 475.2600 624.8400 ;
        RECT 461.9000 618.9200 464.9000 619.4000 ;
        RECT 461.9000 624.3600 464.9000 624.8400 ;
        RECT 473.6600 602.6000 475.2600 603.0800 ;
        RECT 473.6600 608.0400 475.2600 608.5200 ;
        RECT 473.6600 613.4800 475.2600 613.9600 ;
        RECT 461.9000 602.6000 464.9000 603.0800 ;
        RECT 461.9000 608.0400 464.9000 608.5200 ;
        RECT 461.9000 613.4800 464.9000 613.9600 ;
        RECT 473.6600 591.7200 475.2600 592.2000 ;
        RECT 473.6600 597.1600 475.2600 597.6400 ;
        RECT 461.9000 591.7200 464.9000 592.2000 ;
        RECT 461.9000 597.1600 464.9000 597.6400 ;
        RECT 563.6600 575.4000 565.2600 575.8800 ;
        RECT 563.6600 580.8400 565.2600 581.3200 ;
        RECT 563.6600 586.2800 565.2600 586.7600 ;
        RECT 563.6600 564.5200 565.2600 565.0000 ;
        RECT 563.6600 569.9600 565.2600 570.4400 ;
        RECT 518.6600 575.4000 520.2600 575.8800 ;
        RECT 518.6600 580.8400 520.2600 581.3200 ;
        RECT 518.6600 586.2800 520.2600 586.7600 ;
        RECT 518.6600 564.5200 520.2600 565.0000 ;
        RECT 518.6600 569.9600 520.2600 570.4400 ;
        RECT 563.6600 548.2000 565.2600 548.6800 ;
        RECT 563.6600 553.6400 565.2600 554.1200 ;
        RECT 563.6600 559.0800 565.2600 559.5600 ;
        RECT 563.6600 542.7600 565.2600 543.2400 ;
        RECT 518.6600 548.2000 520.2600 548.6800 ;
        RECT 518.6600 553.6400 520.2600 554.1200 ;
        RECT 518.6600 559.0800 520.2600 559.5600 ;
        RECT 518.6600 542.7600 520.2600 543.2400 ;
        RECT 473.6600 575.4000 475.2600 575.8800 ;
        RECT 473.6600 580.8400 475.2600 581.3200 ;
        RECT 473.6600 586.2800 475.2600 586.7600 ;
        RECT 461.9000 575.4000 464.9000 575.8800 ;
        RECT 461.9000 580.8400 464.9000 581.3200 ;
        RECT 461.9000 586.2800 464.9000 586.7600 ;
        RECT 473.6600 564.5200 475.2600 565.0000 ;
        RECT 473.6600 569.9600 475.2600 570.4400 ;
        RECT 461.9000 564.5200 464.9000 565.0000 ;
        RECT 461.9000 569.9600 464.9000 570.4400 ;
        RECT 473.6600 548.2000 475.2600 548.6800 ;
        RECT 473.6600 553.6400 475.2600 554.1200 ;
        RECT 473.6600 559.0800 475.2600 559.5600 ;
        RECT 461.9000 548.2000 464.9000 548.6800 ;
        RECT 461.9000 553.6400 464.9000 554.1200 ;
        RECT 461.9000 559.0800 464.9000 559.5600 ;
        RECT 461.9000 542.7600 464.9000 543.2400 ;
        RECT 473.6600 542.7600 475.2600 543.2400 ;
        RECT 461.9000 747.6700 669.0000 750.6700 ;
        RECT 461.9000 534.5700 669.0000 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 304.9300 655.2600 521.0300 ;
        RECT 608.6600 304.9300 610.2600 521.0300 ;
        RECT 563.6600 304.9300 565.2600 521.0300 ;
        RECT 518.6600 304.9300 520.2600 521.0300 ;
        RECT 473.6600 304.9300 475.2600 521.0300 ;
        RECT 666.0000 304.9300 669.0000 521.0300 ;
        RECT 461.9000 304.9300 464.9000 521.0300 ;
      LAYER met3 ;
        RECT 666.0000 498.0800 669.0000 498.5600 ;
        RECT 666.0000 503.5200 669.0000 504.0000 ;
        RECT 653.6600 498.0800 655.2600 498.5600 ;
        RECT 653.6600 503.5200 655.2600 504.0000 ;
        RECT 666.0000 508.9600 669.0000 509.4400 ;
        RECT 653.6600 508.9600 655.2600 509.4400 ;
        RECT 666.0000 487.2000 669.0000 487.6800 ;
        RECT 666.0000 492.6400 669.0000 493.1200 ;
        RECT 653.6600 487.2000 655.2600 487.6800 ;
        RECT 653.6600 492.6400 655.2600 493.1200 ;
        RECT 666.0000 470.8800 669.0000 471.3600 ;
        RECT 666.0000 476.3200 669.0000 476.8000 ;
        RECT 653.6600 470.8800 655.2600 471.3600 ;
        RECT 653.6600 476.3200 655.2600 476.8000 ;
        RECT 666.0000 481.7600 669.0000 482.2400 ;
        RECT 653.6600 481.7600 655.2600 482.2400 ;
        RECT 608.6600 498.0800 610.2600 498.5600 ;
        RECT 608.6600 503.5200 610.2600 504.0000 ;
        RECT 608.6600 508.9600 610.2600 509.4400 ;
        RECT 608.6600 487.2000 610.2600 487.6800 ;
        RECT 608.6600 492.6400 610.2600 493.1200 ;
        RECT 608.6600 470.8800 610.2600 471.3600 ;
        RECT 608.6600 476.3200 610.2600 476.8000 ;
        RECT 608.6600 481.7600 610.2600 482.2400 ;
        RECT 666.0000 454.5600 669.0000 455.0400 ;
        RECT 666.0000 460.0000 669.0000 460.4800 ;
        RECT 666.0000 465.4400 669.0000 465.9200 ;
        RECT 653.6600 454.5600 655.2600 455.0400 ;
        RECT 653.6600 460.0000 655.2600 460.4800 ;
        RECT 653.6600 465.4400 655.2600 465.9200 ;
        RECT 666.0000 443.6800 669.0000 444.1600 ;
        RECT 666.0000 449.1200 669.0000 449.6000 ;
        RECT 653.6600 443.6800 655.2600 444.1600 ;
        RECT 653.6600 449.1200 655.2600 449.6000 ;
        RECT 666.0000 427.3600 669.0000 427.8400 ;
        RECT 666.0000 432.8000 669.0000 433.2800 ;
        RECT 666.0000 438.2400 669.0000 438.7200 ;
        RECT 653.6600 427.3600 655.2600 427.8400 ;
        RECT 653.6600 432.8000 655.2600 433.2800 ;
        RECT 653.6600 438.2400 655.2600 438.7200 ;
        RECT 666.0000 416.4800 669.0000 416.9600 ;
        RECT 666.0000 421.9200 669.0000 422.4000 ;
        RECT 653.6600 416.4800 655.2600 416.9600 ;
        RECT 653.6600 421.9200 655.2600 422.4000 ;
        RECT 608.6600 454.5600 610.2600 455.0400 ;
        RECT 608.6600 460.0000 610.2600 460.4800 ;
        RECT 608.6600 465.4400 610.2600 465.9200 ;
        RECT 608.6600 443.6800 610.2600 444.1600 ;
        RECT 608.6600 449.1200 610.2600 449.6000 ;
        RECT 608.6600 427.3600 610.2600 427.8400 ;
        RECT 608.6600 432.8000 610.2600 433.2800 ;
        RECT 608.6600 438.2400 610.2600 438.7200 ;
        RECT 608.6600 416.4800 610.2600 416.9600 ;
        RECT 608.6600 421.9200 610.2600 422.4000 ;
        RECT 563.6600 498.0800 565.2600 498.5600 ;
        RECT 563.6600 503.5200 565.2600 504.0000 ;
        RECT 563.6600 508.9600 565.2600 509.4400 ;
        RECT 518.6600 498.0800 520.2600 498.5600 ;
        RECT 518.6600 503.5200 520.2600 504.0000 ;
        RECT 518.6600 508.9600 520.2600 509.4400 ;
        RECT 563.6600 487.2000 565.2600 487.6800 ;
        RECT 563.6600 492.6400 565.2600 493.1200 ;
        RECT 563.6600 470.8800 565.2600 471.3600 ;
        RECT 563.6600 476.3200 565.2600 476.8000 ;
        RECT 563.6600 481.7600 565.2600 482.2400 ;
        RECT 518.6600 487.2000 520.2600 487.6800 ;
        RECT 518.6600 492.6400 520.2600 493.1200 ;
        RECT 518.6600 470.8800 520.2600 471.3600 ;
        RECT 518.6600 476.3200 520.2600 476.8000 ;
        RECT 518.6600 481.7600 520.2600 482.2400 ;
        RECT 473.6600 498.0800 475.2600 498.5600 ;
        RECT 473.6600 503.5200 475.2600 504.0000 ;
        RECT 461.9000 503.5200 464.9000 504.0000 ;
        RECT 461.9000 498.0800 464.9000 498.5600 ;
        RECT 461.9000 508.9600 464.9000 509.4400 ;
        RECT 473.6600 508.9600 475.2600 509.4400 ;
        RECT 473.6600 487.2000 475.2600 487.6800 ;
        RECT 473.6600 492.6400 475.2600 493.1200 ;
        RECT 461.9000 492.6400 464.9000 493.1200 ;
        RECT 461.9000 487.2000 464.9000 487.6800 ;
        RECT 473.6600 470.8800 475.2600 471.3600 ;
        RECT 473.6600 476.3200 475.2600 476.8000 ;
        RECT 461.9000 476.3200 464.9000 476.8000 ;
        RECT 461.9000 470.8800 464.9000 471.3600 ;
        RECT 461.9000 481.7600 464.9000 482.2400 ;
        RECT 473.6600 481.7600 475.2600 482.2400 ;
        RECT 563.6600 454.5600 565.2600 455.0400 ;
        RECT 563.6600 460.0000 565.2600 460.4800 ;
        RECT 563.6600 465.4400 565.2600 465.9200 ;
        RECT 563.6600 443.6800 565.2600 444.1600 ;
        RECT 563.6600 449.1200 565.2600 449.6000 ;
        RECT 518.6600 454.5600 520.2600 455.0400 ;
        RECT 518.6600 460.0000 520.2600 460.4800 ;
        RECT 518.6600 465.4400 520.2600 465.9200 ;
        RECT 518.6600 443.6800 520.2600 444.1600 ;
        RECT 518.6600 449.1200 520.2600 449.6000 ;
        RECT 563.6600 427.3600 565.2600 427.8400 ;
        RECT 563.6600 432.8000 565.2600 433.2800 ;
        RECT 563.6600 438.2400 565.2600 438.7200 ;
        RECT 563.6600 416.4800 565.2600 416.9600 ;
        RECT 563.6600 421.9200 565.2600 422.4000 ;
        RECT 518.6600 427.3600 520.2600 427.8400 ;
        RECT 518.6600 432.8000 520.2600 433.2800 ;
        RECT 518.6600 438.2400 520.2600 438.7200 ;
        RECT 518.6600 416.4800 520.2600 416.9600 ;
        RECT 518.6600 421.9200 520.2600 422.4000 ;
        RECT 473.6600 454.5600 475.2600 455.0400 ;
        RECT 473.6600 460.0000 475.2600 460.4800 ;
        RECT 473.6600 465.4400 475.2600 465.9200 ;
        RECT 461.9000 454.5600 464.9000 455.0400 ;
        RECT 461.9000 460.0000 464.9000 460.4800 ;
        RECT 461.9000 465.4400 464.9000 465.9200 ;
        RECT 473.6600 443.6800 475.2600 444.1600 ;
        RECT 473.6600 449.1200 475.2600 449.6000 ;
        RECT 461.9000 443.6800 464.9000 444.1600 ;
        RECT 461.9000 449.1200 464.9000 449.6000 ;
        RECT 473.6600 427.3600 475.2600 427.8400 ;
        RECT 473.6600 432.8000 475.2600 433.2800 ;
        RECT 473.6600 438.2400 475.2600 438.7200 ;
        RECT 461.9000 427.3600 464.9000 427.8400 ;
        RECT 461.9000 432.8000 464.9000 433.2800 ;
        RECT 461.9000 438.2400 464.9000 438.7200 ;
        RECT 473.6600 416.4800 475.2600 416.9600 ;
        RECT 473.6600 421.9200 475.2600 422.4000 ;
        RECT 461.9000 416.4800 464.9000 416.9600 ;
        RECT 461.9000 421.9200 464.9000 422.4000 ;
        RECT 666.0000 400.1600 669.0000 400.6400 ;
        RECT 666.0000 405.6000 669.0000 406.0800 ;
        RECT 666.0000 411.0400 669.0000 411.5200 ;
        RECT 653.6600 400.1600 655.2600 400.6400 ;
        RECT 653.6600 405.6000 655.2600 406.0800 ;
        RECT 653.6600 411.0400 655.2600 411.5200 ;
        RECT 666.0000 389.2800 669.0000 389.7600 ;
        RECT 666.0000 394.7200 669.0000 395.2000 ;
        RECT 653.6600 389.2800 655.2600 389.7600 ;
        RECT 653.6600 394.7200 655.2600 395.2000 ;
        RECT 666.0000 372.9600 669.0000 373.4400 ;
        RECT 666.0000 378.4000 669.0000 378.8800 ;
        RECT 666.0000 383.8400 669.0000 384.3200 ;
        RECT 653.6600 372.9600 655.2600 373.4400 ;
        RECT 653.6600 378.4000 655.2600 378.8800 ;
        RECT 653.6600 383.8400 655.2600 384.3200 ;
        RECT 666.0000 362.0800 669.0000 362.5600 ;
        RECT 666.0000 367.5200 669.0000 368.0000 ;
        RECT 653.6600 362.0800 655.2600 362.5600 ;
        RECT 653.6600 367.5200 655.2600 368.0000 ;
        RECT 608.6600 400.1600 610.2600 400.6400 ;
        RECT 608.6600 405.6000 610.2600 406.0800 ;
        RECT 608.6600 411.0400 610.2600 411.5200 ;
        RECT 608.6600 389.2800 610.2600 389.7600 ;
        RECT 608.6600 394.7200 610.2600 395.2000 ;
        RECT 608.6600 372.9600 610.2600 373.4400 ;
        RECT 608.6600 378.4000 610.2600 378.8800 ;
        RECT 608.6600 383.8400 610.2600 384.3200 ;
        RECT 608.6600 362.0800 610.2600 362.5600 ;
        RECT 608.6600 367.5200 610.2600 368.0000 ;
        RECT 666.0000 345.7600 669.0000 346.2400 ;
        RECT 666.0000 351.2000 669.0000 351.6800 ;
        RECT 666.0000 356.6400 669.0000 357.1200 ;
        RECT 653.6600 345.7600 655.2600 346.2400 ;
        RECT 653.6600 351.2000 655.2600 351.6800 ;
        RECT 653.6600 356.6400 655.2600 357.1200 ;
        RECT 666.0000 334.8800 669.0000 335.3600 ;
        RECT 666.0000 340.3200 669.0000 340.8000 ;
        RECT 653.6600 334.8800 655.2600 335.3600 ;
        RECT 653.6600 340.3200 655.2600 340.8000 ;
        RECT 666.0000 318.5600 669.0000 319.0400 ;
        RECT 666.0000 324.0000 669.0000 324.4800 ;
        RECT 666.0000 329.4400 669.0000 329.9200 ;
        RECT 653.6600 318.5600 655.2600 319.0400 ;
        RECT 653.6600 324.0000 655.2600 324.4800 ;
        RECT 653.6600 329.4400 655.2600 329.9200 ;
        RECT 666.0000 313.1200 669.0000 313.6000 ;
        RECT 653.6600 313.1200 655.2600 313.6000 ;
        RECT 608.6600 345.7600 610.2600 346.2400 ;
        RECT 608.6600 351.2000 610.2600 351.6800 ;
        RECT 608.6600 356.6400 610.2600 357.1200 ;
        RECT 608.6600 334.8800 610.2600 335.3600 ;
        RECT 608.6600 340.3200 610.2600 340.8000 ;
        RECT 608.6600 318.5600 610.2600 319.0400 ;
        RECT 608.6600 324.0000 610.2600 324.4800 ;
        RECT 608.6600 329.4400 610.2600 329.9200 ;
        RECT 608.6600 313.1200 610.2600 313.6000 ;
        RECT 563.6600 400.1600 565.2600 400.6400 ;
        RECT 563.6600 405.6000 565.2600 406.0800 ;
        RECT 563.6600 411.0400 565.2600 411.5200 ;
        RECT 563.6600 389.2800 565.2600 389.7600 ;
        RECT 563.6600 394.7200 565.2600 395.2000 ;
        RECT 518.6600 400.1600 520.2600 400.6400 ;
        RECT 518.6600 405.6000 520.2600 406.0800 ;
        RECT 518.6600 411.0400 520.2600 411.5200 ;
        RECT 518.6600 389.2800 520.2600 389.7600 ;
        RECT 518.6600 394.7200 520.2600 395.2000 ;
        RECT 563.6600 372.9600 565.2600 373.4400 ;
        RECT 563.6600 378.4000 565.2600 378.8800 ;
        RECT 563.6600 383.8400 565.2600 384.3200 ;
        RECT 563.6600 362.0800 565.2600 362.5600 ;
        RECT 563.6600 367.5200 565.2600 368.0000 ;
        RECT 518.6600 372.9600 520.2600 373.4400 ;
        RECT 518.6600 378.4000 520.2600 378.8800 ;
        RECT 518.6600 383.8400 520.2600 384.3200 ;
        RECT 518.6600 362.0800 520.2600 362.5600 ;
        RECT 518.6600 367.5200 520.2600 368.0000 ;
        RECT 473.6600 400.1600 475.2600 400.6400 ;
        RECT 473.6600 405.6000 475.2600 406.0800 ;
        RECT 473.6600 411.0400 475.2600 411.5200 ;
        RECT 461.9000 400.1600 464.9000 400.6400 ;
        RECT 461.9000 405.6000 464.9000 406.0800 ;
        RECT 461.9000 411.0400 464.9000 411.5200 ;
        RECT 473.6600 389.2800 475.2600 389.7600 ;
        RECT 473.6600 394.7200 475.2600 395.2000 ;
        RECT 461.9000 389.2800 464.9000 389.7600 ;
        RECT 461.9000 394.7200 464.9000 395.2000 ;
        RECT 473.6600 372.9600 475.2600 373.4400 ;
        RECT 473.6600 378.4000 475.2600 378.8800 ;
        RECT 473.6600 383.8400 475.2600 384.3200 ;
        RECT 461.9000 372.9600 464.9000 373.4400 ;
        RECT 461.9000 378.4000 464.9000 378.8800 ;
        RECT 461.9000 383.8400 464.9000 384.3200 ;
        RECT 473.6600 362.0800 475.2600 362.5600 ;
        RECT 473.6600 367.5200 475.2600 368.0000 ;
        RECT 461.9000 362.0800 464.9000 362.5600 ;
        RECT 461.9000 367.5200 464.9000 368.0000 ;
        RECT 563.6600 345.7600 565.2600 346.2400 ;
        RECT 563.6600 351.2000 565.2600 351.6800 ;
        RECT 563.6600 356.6400 565.2600 357.1200 ;
        RECT 563.6600 334.8800 565.2600 335.3600 ;
        RECT 563.6600 340.3200 565.2600 340.8000 ;
        RECT 518.6600 345.7600 520.2600 346.2400 ;
        RECT 518.6600 351.2000 520.2600 351.6800 ;
        RECT 518.6600 356.6400 520.2600 357.1200 ;
        RECT 518.6600 334.8800 520.2600 335.3600 ;
        RECT 518.6600 340.3200 520.2600 340.8000 ;
        RECT 563.6600 318.5600 565.2600 319.0400 ;
        RECT 563.6600 324.0000 565.2600 324.4800 ;
        RECT 563.6600 329.4400 565.2600 329.9200 ;
        RECT 563.6600 313.1200 565.2600 313.6000 ;
        RECT 518.6600 318.5600 520.2600 319.0400 ;
        RECT 518.6600 324.0000 520.2600 324.4800 ;
        RECT 518.6600 329.4400 520.2600 329.9200 ;
        RECT 518.6600 313.1200 520.2600 313.6000 ;
        RECT 473.6600 345.7600 475.2600 346.2400 ;
        RECT 473.6600 351.2000 475.2600 351.6800 ;
        RECT 473.6600 356.6400 475.2600 357.1200 ;
        RECT 461.9000 345.7600 464.9000 346.2400 ;
        RECT 461.9000 351.2000 464.9000 351.6800 ;
        RECT 461.9000 356.6400 464.9000 357.1200 ;
        RECT 473.6600 334.8800 475.2600 335.3600 ;
        RECT 473.6600 340.3200 475.2600 340.8000 ;
        RECT 461.9000 334.8800 464.9000 335.3600 ;
        RECT 461.9000 340.3200 464.9000 340.8000 ;
        RECT 473.6600 318.5600 475.2600 319.0400 ;
        RECT 473.6600 324.0000 475.2600 324.4800 ;
        RECT 473.6600 329.4400 475.2600 329.9200 ;
        RECT 461.9000 318.5600 464.9000 319.0400 ;
        RECT 461.9000 324.0000 464.9000 324.4800 ;
        RECT 461.9000 329.4400 464.9000 329.9200 ;
        RECT 461.9000 313.1200 464.9000 313.6000 ;
        RECT 473.6600 313.1200 475.2600 313.6000 ;
        RECT 461.9000 518.0300 669.0000 521.0300 ;
        RECT 461.9000 304.9300 669.0000 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 75.2900 655.2600 291.3900 ;
        RECT 608.6600 75.2900 610.2600 291.3900 ;
        RECT 563.6600 75.2900 565.2600 291.3900 ;
        RECT 518.6600 75.2900 520.2600 291.3900 ;
        RECT 473.6600 75.2900 475.2600 291.3900 ;
        RECT 666.0000 75.2900 669.0000 291.3900 ;
        RECT 461.9000 75.2900 464.9000 291.3900 ;
      LAYER met3 ;
        RECT 666.0000 268.4400 669.0000 268.9200 ;
        RECT 666.0000 273.8800 669.0000 274.3600 ;
        RECT 653.6600 268.4400 655.2600 268.9200 ;
        RECT 653.6600 273.8800 655.2600 274.3600 ;
        RECT 666.0000 279.3200 669.0000 279.8000 ;
        RECT 653.6600 279.3200 655.2600 279.8000 ;
        RECT 666.0000 257.5600 669.0000 258.0400 ;
        RECT 666.0000 263.0000 669.0000 263.4800 ;
        RECT 653.6600 257.5600 655.2600 258.0400 ;
        RECT 653.6600 263.0000 655.2600 263.4800 ;
        RECT 666.0000 241.2400 669.0000 241.7200 ;
        RECT 666.0000 246.6800 669.0000 247.1600 ;
        RECT 653.6600 241.2400 655.2600 241.7200 ;
        RECT 653.6600 246.6800 655.2600 247.1600 ;
        RECT 666.0000 252.1200 669.0000 252.6000 ;
        RECT 653.6600 252.1200 655.2600 252.6000 ;
        RECT 608.6600 268.4400 610.2600 268.9200 ;
        RECT 608.6600 273.8800 610.2600 274.3600 ;
        RECT 608.6600 279.3200 610.2600 279.8000 ;
        RECT 608.6600 257.5600 610.2600 258.0400 ;
        RECT 608.6600 263.0000 610.2600 263.4800 ;
        RECT 608.6600 241.2400 610.2600 241.7200 ;
        RECT 608.6600 246.6800 610.2600 247.1600 ;
        RECT 608.6600 252.1200 610.2600 252.6000 ;
        RECT 666.0000 224.9200 669.0000 225.4000 ;
        RECT 666.0000 230.3600 669.0000 230.8400 ;
        RECT 666.0000 235.8000 669.0000 236.2800 ;
        RECT 653.6600 224.9200 655.2600 225.4000 ;
        RECT 653.6600 230.3600 655.2600 230.8400 ;
        RECT 653.6600 235.8000 655.2600 236.2800 ;
        RECT 666.0000 214.0400 669.0000 214.5200 ;
        RECT 666.0000 219.4800 669.0000 219.9600 ;
        RECT 653.6600 214.0400 655.2600 214.5200 ;
        RECT 653.6600 219.4800 655.2600 219.9600 ;
        RECT 666.0000 197.7200 669.0000 198.2000 ;
        RECT 666.0000 203.1600 669.0000 203.6400 ;
        RECT 666.0000 208.6000 669.0000 209.0800 ;
        RECT 653.6600 197.7200 655.2600 198.2000 ;
        RECT 653.6600 203.1600 655.2600 203.6400 ;
        RECT 653.6600 208.6000 655.2600 209.0800 ;
        RECT 666.0000 186.8400 669.0000 187.3200 ;
        RECT 666.0000 192.2800 669.0000 192.7600 ;
        RECT 653.6600 186.8400 655.2600 187.3200 ;
        RECT 653.6600 192.2800 655.2600 192.7600 ;
        RECT 608.6600 224.9200 610.2600 225.4000 ;
        RECT 608.6600 230.3600 610.2600 230.8400 ;
        RECT 608.6600 235.8000 610.2600 236.2800 ;
        RECT 608.6600 214.0400 610.2600 214.5200 ;
        RECT 608.6600 219.4800 610.2600 219.9600 ;
        RECT 608.6600 197.7200 610.2600 198.2000 ;
        RECT 608.6600 203.1600 610.2600 203.6400 ;
        RECT 608.6600 208.6000 610.2600 209.0800 ;
        RECT 608.6600 186.8400 610.2600 187.3200 ;
        RECT 608.6600 192.2800 610.2600 192.7600 ;
        RECT 563.6600 268.4400 565.2600 268.9200 ;
        RECT 563.6600 273.8800 565.2600 274.3600 ;
        RECT 563.6600 279.3200 565.2600 279.8000 ;
        RECT 518.6600 268.4400 520.2600 268.9200 ;
        RECT 518.6600 273.8800 520.2600 274.3600 ;
        RECT 518.6600 279.3200 520.2600 279.8000 ;
        RECT 563.6600 257.5600 565.2600 258.0400 ;
        RECT 563.6600 263.0000 565.2600 263.4800 ;
        RECT 563.6600 241.2400 565.2600 241.7200 ;
        RECT 563.6600 246.6800 565.2600 247.1600 ;
        RECT 563.6600 252.1200 565.2600 252.6000 ;
        RECT 518.6600 257.5600 520.2600 258.0400 ;
        RECT 518.6600 263.0000 520.2600 263.4800 ;
        RECT 518.6600 241.2400 520.2600 241.7200 ;
        RECT 518.6600 246.6800 520.2600 247.1600 ;
        RECT 518.6600 252.1200 520.2600 252.6000 ;
        RECT 473.6600 268.4400 475.2600 268.9200 ;
        RECT 473.6600 273.8800 475.2600 274.3600 ;
        RECT 461.9000 273.8800 464.9000 274.3600 ;
        RECT 461.9000 268.4400 464.9000 268.9200 ;
        RECT 461.9000 279.3200 464.9000 279.8000 ;
        RECT 473.6600 279.3200 475.2600 279.8000 ;
        RECT 473.6600 257.5600 475.2600 258.0400 ;
        RECT 473.6600 263.0000 475.2600 263.4800 ;
        RECT 461.9000 263.0000 464.9000 263.4800 ;
        RECT 461.9000 257.5600 464.9000 258.0400 ;
        RECT 473.6600 241.2400 475.2600 241.7200 ;
        RECT 473.6600 246.6800 475.2600 247.1600 ;
        RECT 461.9000 246.6800 464.9000 247.1600 ;
        RECT 461.9000 241.2400 464.9000 241.7200 ;
        RECT 461.9000 252.1200 464.9000 252.6000 ;
        RECT 473.6600 252.1200 475.2600 252.6000 ;
        RECT 563.6600 224.9200 565.2600 225.4000 ;
        RECT 563.6600 230.3600 565.2600 230.8400 ;
        RECT 563.6600 235.8000 565.2600 236.2800 ;
        RECT 563.6600 214.0400 565.2600 214.5200 ;
        RECT 563.6600 219.4800 565.2600 219.9600 ;
        RECT 518.6600 224.9200 520.2600 225.4000 ;
        RECT 518.6600 230.3600 520.2600 230.8400 ;
        RECT 518.6600 235.8000 520.2600 236.2800 ;
        RECT 518.6600 214.0400 520.2600 214.5200 ;
        RECT 518.6600 219.4800 520.2600 219.9600 ;
        RECT 563.6600 197.7200 565.2600 198.2000 ;
        RECT 563.6600 203.1600 565.2600 203.6400 ;
        RECT 563.6600 208.6000 565.2600 209.0800 ;
        RECT 563.6600 186.8400 565.2600 187.3200 ;
        RECT 563.6600 192.2800 565.2600 192.7600 ;
        RECT 518.6600 197.7200 520.2600 198.2000 ;
        RECT 518.6600 203.1600 520.2600 203.6400 ;
        RECT 518.6600 208.6000 520.2600 209.0800 ;
        RECT 518.6600 186.8400 520.2600 187.3200 ;
        RECT 518.6600 192.2800 520.2600 192.7600 ;
        RECT 473.6600 224.9200 475.2600 225.4000 ;
        RECT 473.6600 230.3600 475.2600 230.8400 ;
        RECT 473.6600 235.8000 475.2600 236.2800 ;
        RECT 461.9000 224.9200 464.9000 225.4000 ;
        RECT 461.9000 230.3600 464.9000 230.8400 ;
        RECT 461.9000 235.8000 464.9000 236.2800 ;
        RECT 473.6600 214.0400 475.2600 214.5200 ;
        RECT 473.6600 219.4800 475.2600 219.9600 ;
        RECT 461.9000 214.0400 464.9000 214.5200 ;
        RECT 461.9000 219.4800 464.9000 219.9600 ;
        RECT 473.6600 197.7200 475.2600 198.2000 ;
        RECT 473.6600 203.1600 475.2600 203.6400 ;
        RECT 473.6600 208.6000 475.2600 209.0800 ;
        RECT 461.9000 197.7200 464.9000 198.2000 ;
        RECT 461.9000 203.1600 464.9000 203.6400 ;
        RECT 461.9000 208.6000 464.9000 209.0800 ;
        RECT 473.6600 186.8400 475.2600 187.3200 ;
        RECT 473.6600 192.2800 475.2600 192.7600 ;
        RECT 461.9000 186.8400 464.9000 187.3200 ;
        RECT 461.9000 192.2800 464.9000 192.7600 ;
        RECT 666.0000 170.5200 669.0000 171.0000 ;
        RECT 666.0000 175.9600 669.0000 176.4400 ;
        RECT 666.0000 181.4000 669.0000 181.8800 ;
        RECT 653.6600 170.5200 655.2600 171.0000 ;
        RECT 653.6600 175.9600 655.2600 176.4400 ;
        RECT 653.6600 181.4000 655.2600 181.8800 ;
        RECT 666.0000 159.6400 669.0000 160.1200 ;
        RECT 666.0000 165.0800 669.0000 165.5600 ;
        RECT 653.6600 159.6400 655.2600 160.1200 ;
        RECT 653.6600 165.0800 655.2600 165.5600 ;
        RECT 666.0000 143.3200 669.0000 143.8000 ;
        RECT 666.0000 148.7600 669.0000 149.2400 ;
        RECT 666.0000 154.2000 669.0000 154.6800 ;
        RECT 653.6600 143.3200 655.2600 143.8000 ;
        RECT 653.6600 148.7600 655.2600 149.2400 ;
        RECT 653.6600 154.2000 655.2600 154.6800 ;
        RECT 666.0000 132.4400 669.0000 132.9200 ;
        RECT 666.0000 137.8800 669.0000 138.3600 ;
        RECT 653.6600 132.4400 655.2600 132.9200 ;
        RECT 653.6600 137.8800 655.2600 138.3600 ;
        RECT 608.6600 170.5200 610.2600 171.0000 ;
        RECT 608.6600 175.9600 610.2600 176.4400 ;
        RECT 608.6600 181.4000 610.2600 181.8800 ;
        RECT 608.6600 159.6400 610.2600 160.1200 ;
        RECT 608.6600 165.0800 610.2600 165.5600 ;
        RECT 608.6600 143.3200 610.2600 143.8000 ;
        RECT 608.6600 148.7600 610.2600 149.2400 ;
        RECT 608.6600 154.2000 610.2600 154.6800 ;
        RECT 608.6600 132.4400 610.2600 132.9200 ;
        RECT 608.6600 137.8800 610.2600 138.3600 ;
        RECT 666.0000 116.1200 669.0000 116.6000 ;
        RECT 666.0000 121.5600 669.0000 122.0400 ;
        RECT 666.0000 127.0000 669.0000 127.4800 ;
        RECT 653.6600 116.1200 655.2600 116.6000 ;
        RECT 653.6600 121.5600 655.2600 122.0400 ;
        RECT 653.6600 127.0000 655.2600 127.4800 ;
        RECT 666.0000 105.2400 669.0000 105.7200 ;
        RECT 666.0000 110.6800 669.0000 111.1600 ;
        RECT 653.6600 105.2400 655.2600 105.7200 ;
        RECT 653.6600 110.6800 655.2600 111.1600 ;
        RECT 666.0000 88.9200 669.0000 89.4000 ;
        RECT 666.0000 94.3600 669.0000 94.8400 ;
        RECT 666.0000 99.8000 669.0000 100.2800 ;
        RECT 653.6600 88.9200 655.2600 89.4000 ;
        RECT 653.6600 94.3600 655.2600 94.8400 ;
        RECT 653.6600 99.8000 655.2600 100.2800 ;
        RECT 666.0000 83.4800 669.0000 83.9600 ;
        RECT 653.6600 83.4800 655.2600 83.9600 ;
        RECT 608.6600 116.1200 610.2600 116.6000 ;
        RECT 608.6600 121.5600 610.2600 122.0400 ;
        RECT 608.6600 127.0000 610.2600 127.4800 ;
        RECT 608.6600 105.2400 610.2600 105.7200 ;
        RECT 608.6600 110.6800 610.2600 111.1600 ;
        RECT 608.6600 88.9200 610.2600 89.4000 ;
        RECT 608.6600 94.3600 610.2600 94.8400 ;
        RECT 608.6600 99.8000 610.2600 100.2800 ;
        RECT 608.6600 83.4800 610.2600 83.9600 ;
        RECT 563.6600 170.5200 565.2600 171.0000 ;
        RECT 563.6600 175.9600 565.2600 176.4400 ;
        RECT 563.6600 181.4000 565.2600 181.8800 ;
        RECT 563.6600 159.6400 565.2600 160.1200 ;
        RECT 563.6600 165.0800 565.2600 165.5600 ;
        RECT 518.6600 170.5200 520.2600 171.0000 ;
        RECT 518.6600 175.9600 520.2600 176.4400 ;
        RECT 518.6600 181.4000 520.2600 181.8800 ;
        RECT 518.6600 159.6400 520.2600 160.1200 ;
        RECT 518.6600 165.0800 520.2600 165.5600 ;
        RECT 563.6600 143.3200 565.2600 143.8000 ;
        RECT 563.6600 148.7600 565.2600 149.2400 ;
        RECT 563.6600 154.2000 565.2600 154.6800 ;
        RECT 563.6600 132.4400 565.2600 132.9200 ;
        RECT 563.6600 137.8800 565.2600 138.3600 ;
        RECT 518.6600 143.3200 520.2600 143.8000 ;
        RECT 518.6600 148.7600 520.2600 149.2400 ;
        RECT 518.6600 154.2000 520.2600 154.6800 ;
        RECT 518.6600 132.4400 520.2600 132.9200 ;
        RECT 518.6600 137.8800 520.2600 138.3600 ;
        RECT 473.6600 170.5200 475.2600 171.0000 ;
        RECT 473.6600 175.9600 475.2600 176.4400 ;
        RECT 473.6600 181.4000 475.2600 181.8800 ;
        RECT 461.9000 170.5200 464.9000 171.0000 ;
        RECT 461.9000 175.9600 464.9000 176.4400 ;
        RECT 461.9000 181.4000 464.9000 181.8800 ;
        RECT 473.6600 159.6400 475.2600 160.1200 ;
        RECT 473.6600 165.0800 475.2600 165.5600 ;
        RECT 461.9000 159.6400 464.9000 160.1200 ;
        RECT 461.9000 165.0800 464.9000 165.5600 ;
        RECT 473.6600 143.3200 475.2600 143.8000 ;
        RECT 473.6600 148.7600 475.2600 149.2400 ;
        RECT 473.6600 154.2000 475.2600 154.6800 ;
        RECT 461.9000 143.3200 464.9000 143.8000 ;
        RECT 461.9000 148.7600 464.9000 149.2400 ;
        RECT 461.9000 154.2000 464.9000 154.6800 ;
        RECT 473.6600 132.4400 475.2600 132.9200 ;
        RECT 473.6600 137.8800 475.2600 138.3600 ;
        RECT 461.9000 132.4400 464.9000 132.9200 ;
        RECT 461.9000 137.8800 464.9000 138.3600 ;
        RECT 563.6600 116.1200 565.2600 116.6000 ;
        RECT 563.6600 121.5600 565.2600 122.0400 ;
        RECT 563.6600 127.0000 565.2600 127.4800 ;
        RECT 563.6600 105.2400 565.2600 105.7200 ;
        RECT 563.6600 110.6800 565.2600 111.1600 ;
        RECT 518.6600 116.1200 520.2600 116.6000 ;
        RECT 518.6600 121.5600 520.2600 122.0400 ;
        RECT 518.6600 127.0000 520.2600 127.4800 ;
        RECT 518.6600 105.2400 520.2600 105.7200 ;
        RECT 518.6600 110.6800 520.2600 111.1600 ;
        RECT 563.6600 88.9200 565.2600 89.4000 ;
        RECT 563.6600 94.3600 565.2600 94.8400 ;
        RECT 563.6600 99.8000 565.2600 100.2800 ;
        RECT 563.6600 83.4800 565.2600 83.9600 ;
        RECT 518.6600 88.9200 520.2600 89.4000 ;
        RECT 518.6600 94.3600 520.2600 94.8400 ;
        RECT 518.6600 99.8000 520.2600 100.2800 ;
        RECT 518.6600 83.4800 520.2600 83.9600 ;
        RECT 473.6600 116.1200 475.2600 116.6000 ;
        RECT 473.6600 121.5600 475.2600 122.0400 ;
        RECT 473.6600 127.0000 475.2600 127.4800 ;
        RECT 461.9000 116.1200 464.9000 116.6000 ;
        RECT 461.9000 121.5600 464.9000 122.0400 ;
        RECT 461.9000 127.0000 464.9000 127.4800 ;
        RECT 473.6600 105.2400 475.2600 105.7200 ;
        RECT 473.6600 110.6800 475.2600 111.1600 ;
        RECT 461.9000 105.2400 464.9000 105.7200 ;
        RECT 461.9000 110.6800 464.9000 111.1600 ;
        RECT 473.6600 88.9200 475.2600 89.4000 ;
        RECT 473.6600 94.3600 475.2600 94.8400 ;
        RECT 473.6600 99.8000 475.2600 100.2800 ;
        RECT 461.9000 88.9200 464.9000 89.4000 ;
        RECT 461.9000 94.3600 464.9000 94.8400 ;
        RECT 461.9000 99.8000 464.9000 100.2800 ;
        RECT 461.9000 83.4800 464.9000 83.9600 ;
        RECT 473.6600 83.4800 475.2600 83.9600 ;
        RECT 461.9000 288.3900 669.0000 291.3900 ;
        RECT 461.9000 75.2900 669.0000 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 462.9000 34.6700 464.9000 61.6000 ;
        RECT 666.0000 34.6700 668.0000 61.6000 ;
      LAYER met3 ;
        RECT 666.0000 51.3800 668.0000 51.8600 ;
        RECT 462.9000 51.3800 464.9000 51.8600 ;
        RECT 666.0000 45.9400 668.0000 46.4200 ;
        RECT 666.0000 40.5000 668.0000 40.9800 ;
        RECT 462.9000 45.9400 464.9000 46.4200 ;
        RECT 462.9000 40.5000 464.9000 40.9800 ;
        RECT 462.9000 59.6000 668.0000 61.6000 ;
        RECT 462.9000 34.6700 668.0000 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 2601.3300 655.2600 2817.4300 ;
        RECT 608.6600 2601.3300 610.2600 2817.4300 ;
        RECT 563.6600 2601.3300 565.2600 2817.4300 ;
        RECT 518.6600 2601.3300 520.2600 2817.4300 ;
        RECT 473.6600 2601.3300 475.2600 2817.4300 ;
        RECT 666.0000 2601.3300 669.0000 2817.4300 ;
        RECT 461.9000 2601.3300 464.9000 2817.4300 ;
      LAYER met3 ;
        RECT 666.0000 2794.4800 669.0000 2794.9600 ;
        RECT 666.0000 2799.9200 669.0000 2800.4000 ;
        RECT 653.6600 2794.4800 655.2600 2794.9600 ;
        RECT 653.6600 2799.9200 655.2600 2800.4000 ;
        RECT 666.0000 2805.3600 669.0000 2805.8400 ;
        RECT 653.6600 2805.3600 655.2600 2805.8400 ;
        RECT 666.0000 2783.6000 669.0000 2784.0800 ;
        RECT 666.0000 2789.0400 669.0000 2789.5200 ;
        RECT 653.6600 2783.6000 655.2600 2784.0800 ;
        RECT 653.6600 2789.0400 655.2600 2789.5200 ;
        RECT 666.0000 2767.2800 669.0000 2767.7600 ;
        RECT 666.0000 2772.7200 669.0000 2773.2000 ;
        RECT 653.6600 2767.2800 655.2600 2767.7600 ;
        RECT 653.6600 2772.7200 655.2600 2773.2000 ;
        RECT 666.0000 2778.1600 669.0000 2778.6400 ;
        RECT 653.6600 2778.1600 655.2600 2778.6400 ;
        RECT 608.6600 2794.4800 610.2600 2794.9600 ;
        RECT 608.6600 2799.9200 610.2600 2800.4000 ;
        RECT 608.6600 2805.3600 610.2600 2805.8400 ;
        RECT 608.6600 2783.6000 610.2600 2784.0800 ;
        RECT 608.6600 2789.0400 610.2600 2789.5200 ;
        RECT 608.6600 2767.2800 610.2600 2767.7600 ;
        RECT 608.6600 2772.7200 610.2600 2773.2000 ;
        RECT 608.6600 2778.1600 610.2600 2778.6400 ;
        RECT 666.0000 2750.9600 669.0000 2751.4400 ;
        RECT 666.0000 2756.4000 669.0000 2756.8800 ;
        RECT 666.0000 2761.8400 669.0000 2762.3200 ;
        RECT 653.6600 2750.9600 655.2600 2751.4400 ;
        RECT 653.6600 2756.4000 655.2600 2756.8800 ;
        RECT 653.6600 2761.8400 655.2600 2762.3200 ;
        RECT 666.0000 2740.0800 669.0000 2740.5600 ;
        RECT 666.0000 2745.5200 669.0000 2746.0000 ;
        RECT 653.6600 2740.0800 655.2600 2740.5600 ;
        RECT 653.6600 2745.5200 655.2600 2746.0000 ;
        RECT 666.0000 2723.7600 669.0000 2724.2400 ;
        RECT 666.0000 2729.2000 669.0000 2729.6800 ;
        RECT 666.0000 2734.6400 669.0000 2735.1200 ;
        RECT 653.6600 2723.7600 655.2600 2724.2400 ;
        RECT 653.6600 2729.2000 655.2600 2729.6800 ;
        RECT 653.6600 2734.6400 655.2600 2735.1200 ;
        RECT 666.0000 2712.8800 669.0000 2713.3600 ;
        RECT 666.0000 2718.3200 669.0000 2718.8000 ;
        RECT 653.6600 2712.8800 655.2600 2713.3600 ;
        RECT 653.6600 2718.3200 655.2600 2718.8000 ;
        RECT 608.6600 2750.9600 610.2600 2751.4400 ;
        RECT 608.6600 2756.4000 610.2600 2756.8800 ;
        RECT 608.6600 2761.8400 610.2600 2762.3200 ;
        RECT 608.6600 2740.0800 610.2600 2740.5600 ;
        RECT 608.6600 2745.5200 610.2600 2746.0000 ;
        RECT 608.6600 2723.7600 610.2600 2724.2400 ;
        RECT 608.6600 2729.2000 610.2600 2729.6800 ;
        RECT 608.6600 2734.6400 610.2600 2735.1200 ;
        RECT 608.6600 2712.8800 610.2600 2713.3600 ;
        RECT 608.6600 2718.3200 610.2600 2718.8000 ;
        RECT 563.6600 2794.4800 565.2600 2794.9600 ;
        RECT 563.6600 2799.9200 565.2600 2800.4000 ;
        RECT 563.6600 2805.3600 565.2600 2805.8400 ;
        RECT 518.6600 2794.4800 520.2600 2794.9600 ;
        RECT 518.6600 2799.9200 520.2600 2800.4000 ;
        RECT 518.6600 2805.3600 520.2600 2805.8400 ;
        RECT 563.6600 2783.6000 565.2600 2784.0800 ;
        RECT 563.6600 2789.0400 565.2600 2789.5200 ;
        RECT 563.6600 2767.2800 565.2600 2767.7600 ;
        RECT 563.6600 2772.7200 565.2600 2773.2000 ;
        RECT 563.6600 2778.1600 565.2600 2778.6400 ;
        RECT 518.6600 2783.6000 520.2600 2784.0800 ;
        RECT 518.6600 2789.0400 520.2600 2789.5200 ;
        RECT 518.6600 2767.2800 520.2600 2767.7600 ;
        RECT 518.6600 2772.7200 520.2600 2773.2000 ;
        RECT 518.6600 2778.1600 520.2600 2778.6400 ;
        RECT 473.6600 2794.4800 475.2600 2794.9600 ;
        RECT 473.6600 2799.9200 475.2600 2800.4000 ;
        RECT 461.9000 2799.9200 464.9000 2800.4000 ;
        RECT 461.9000 2794.4800 464.9000 2794.9600 ;
        RECT 461.9000 2805.3600 464.9000 2805.8400 ;
        RECT 473.6600 2805.3600 475.2600 2805.8400 ;
        RECT 473.6600 2783.6000 475.2600 2784.0800 ;
        RECT 473.6600 2789.0400 475.2600 2789.5200 ;
        RECT 461.9000 2789.0400 464.9000 2789.5200 ;
        RECT 461.9000 2783.6000 464.9000 2784.0800 ;
        RECT 473.6600 2767.2800 475.2600 2767.7600 ;
        RECT 473.6600 2772.7200 475.2600 2773.2000 ;
        RECT 461.9000 2772.7200 464.9000 2773.2000 ;
        RECT 461.9000 2767.2800 464.9000 2767.7600 ;
        RECT 461.9000 2778.1600 464.9000 2778.6400 ;
        RECT 473.6600 2778.1600 475.2600 2778.6400 ;
        RECT 563.6600 2750.9600 565.2600 2751.4400 ;
        RECT 563.6600 2756.4000 565.2600 2756.8800 ;
        RECT 563.6600 2761.8400 565.2600 2762.3200 ;
        RECT 563.6600 2740.0800 565.2600 2740.5600 ;
        RECT 563.6600 2745.5200 565.2600 2746.0000 ;
        RECT 518.6600 2750.9600 520.2600 2751.4400 ;
        RECT 518.6600 2756.4000 520.2600 2756.8800 ;
        RECT 518.6600 2761.8400 520.2600 2762.3200 ;
        RECT 518.6600 2740.0800 520.2600 2740.5600 ;
        RECT 518.6600 2745.5200 520.2600 2746.0000 ;
        RECT 563.6600 2723.7600 565.2600 2724.2400 ;
        RECT 563.6600 2729.2000 565.2600 2729.6800 ;
        RECT 563.6600 2734.6400 565.2600 2735.1200 ;
        RECT 563.6600 2712.8800 565.2600 2713.3600 ;
        RECT 563.6600 2718.3200 565.2600 2718.8000 ;
        RECT 518.6600 2723.7600 520.2600 2724.2400 ;
        RECT 518.6600 2729.2000 520.2600 2729.6800 ;
        RECT 518.6600 2734.6400 520.2600 2735.1200 ;
        RECT 518.6600 2712.8800 520.2600 2713.3600 ;
        RECT 518.6600 2718.3200 520.2600 2718.8000 ;
        RECT 473.6600 2750.9600 475.2600 2751.4400 ;
        RECT 473.6600 2756.4000 475.2600 2756.8800 ;
        RECT 473.6600 2761.8400 475.2600 2762.3200 ;
        RECT 461.9000 2750.9600 464.9000 2751.4400 ;
        RECT 461.9000 2756.4000 464.9000 2756.8800 ;
        RECT 461.9000 2761.8400 464.9000 2762.3200 ;
        RECT 473.6600 2740.0800 475.2600 2740.5600 ;
        RECT 473.6600 2745.5200 475.2600 2746.0000 ;
        RECT 461.9000 2740.0800 464.9000 2740.5600 ;
        RECT 461.9000 2745.5200 464.9000 2746.0000 ;
        RECT 473.6600 2723.7600 475.2600 2724.2400 ;
        RECT 473.6600 2729.2000 475.2600 2729.6800 ;
        RECT 473.6600 2734.6400 475.2600 2735.1200 ;
        RECT 461.9000 2723.7600 464.9000 2724.2400 ;
        RECT 461.9000 2729.2000 464.9000 2729.6800 ;
        RECT 461.9000 2734.6400 464.9000 2735.1200 ;
        RECT 473.6600 2712.8800 475.2600 2713.3600 ;
        RECT 473.6600 2718.3200 475.2600 2718.8000 ;
        RECT 461.9000 2712.8800 464.9000 2713.3600 ;
        RECT 461.9000 2718.3200 464.9000 2718.8000 ;
        RECT 666.0000 2696.5600 669.0000 2697.0400 ;
        RECT 666.0000 2702.0000 669.0000 2702.4800 ;
        RECT 666.0000 2707.4400 669.0000 2707.9200 ;
        RECT 653.6600 2696.5600 655.2600 2697.0400 ;
        RECT 653.6600 2702.0000 655.2600 2702.4800 ;
        RECT 653.6600 2707.4400 655.2600 2707.9200 ;
        RECT 666.0000 2685.6800 669.0000 2686.1600 ;
        RECT 666.0000 2691.1200 669.0000 2691.6000 ;
        RECT 653.6600 2685.6800 655.2600 2686.1600 ;
        RECT 653.6600 2691.1200 655.2600 2691.6000 ;
        RECT 666.0000 2669.3600 669.0000 2669.8400 ;
        RECT 666.0000 2674.8000 669.0000 2675.2800 ;
        RECT 666.0000 2680.2400 669.0000 2680.7200 ;
        RECT 653.6600 2669.3600 655.2600 2669.8400 ;
        RECT 653.6600 2674.8000 655.2600 2675.2800 ;
        RECT 653.6600 2680.2400 655.2600 2680.7200 ;
        RECT 666.0000 2658.4800 669.0000 2658.9600 ;
        RECT 666.0000 2663.9200 669.0000 2664.4000 ;
        RECT 653.6600 2658.4800 655.2600 2658.9600 ;
        RECT 653.6600 2663.9200 655.2600 2664.4000 ;
        RECT 608.6600 2696.5600 610.2600 2697.0400 ;
        RECT 608.6600 2702.0000 610.2600 2702.4800 ;
        RECT 608.6600 2707.4400 610.2600 2707.9200 ;
        RECT 608.6600 2685.6800 610.2600 2686.1600 ;
        RECT 608.6600 2691.1200 610.2600 2691.6000 ;
        RECT 608.6600 2669.3600 610.2600 2669.8400 ;
        RECT 608.6600 2674.8000 610.2600 2675.2800 ;
        RECT 608.6600 2680.2400 610.2600 2680.7200 ;
        RECT 608.6600 2658.4800 610.2600 2658.9600 ;
        RECT 608.6600 2663.9200 610.2600 2664.4000 ;
        RECT 666.0000 2642.1600 669.0000 2642.6400 ;
        RECT 666.0000 2647.6000 669.0000 2648.0800 ;
        RECT 666.0000 2653.0400 669.0000 2653.5200 ;
        RECT 653.6600 2642.1600 655.2600 2642.6400 ;
        RECT 653.6600 2647.6000 655.2600 2648.0800 ;
        RECT 653.6600 2653.0400 655.2600 2653.5200 ;
        RECT 666.0000 2631.2800 669.0000 2631.7600 ;
        RECT 666.0000 2636.7200 669.0000 2637.2000 ;
        RECT 653.6600 2631.2800 655.2600 2631.7600 ;
        RECT 653.6600 2636.7200 655.2600 2637.2000 ;
        RECT 666.0000 2614.9600 669.0000 2615.4400 ;
        RECT 666.0000 2620.4000 669.0000 2620.8800 ;
        RECT 666.0000 2625.8400 669.0000 2626.3200 ;
        RECT 653.6600 2614.9600 655.2600 2615.4400 ;
        RECT 653.6600 2620.4000 655.2600 2620.8800 ;
        RECT 653.6600 2625.8400 655.2600 2626.3200 ;
        RECT 666.0000 2609.5200 669.0000 2610.0000 ;
        RECT 653.6600 2609.5200 655.2600 2610.0000 ;
        RECT 608.6600 2642.1600 610.2600 2642.6400 ;
        RECT 608.6600 2647.6000 610.2600 2648.0800 ;
        RECT 608.6600 2653.0400 610.2600 2653.5200 ;
        RECT 608.6600 2631.2800 610.2600 2631.7600 ;
        RECT 608.6600 2636.7200 610.2600 2637.2000 ;
        RECT 608.6600 2614.9600 610.2600 2615.4400 ;
        RECT 608.6600 2620.4000 610.2600 2620.8800 ;
        RECT 608.6600 2625.8400 610.2600 2626.3200 ;
        RECT 608.6600 2609.5200 610.2600 2610.0000 ;
        RECT 563.6600 2696.5600 565.2600 2697.0400 ;
        RECT 563.6600 2702.0000 565.2600 2702.4800 ;
        RECT 563.6600 2707.4400 565.2600 2707.9200 ;
        RECT 563.6600 2685.6800 565.2600 2686.1600 ;
        RECT 563.6600 2691.1200 565.2600 2691.6000 ;
        RECT 518.6600 2696.5600 520.2600 2697.0400 ;
        RECT 518.6600 2702.0000 520.2600 2702.4800 ;
        RECT 518.6600 2707.4400 520.2600 2707.9200 ;
        RECT 518.6600 2685.6800 520.2600 2686.1600 ;
        RECT 518.6600 2691.1200 520.2600 2691.6000 ;
        RECT 563.6600 2669.3600 565.2600 2669.8400 ;
        RECT 563.6600 2674.8000 565.2600 2675.2800 ;
        RECT 563.6600 2680.2400 565.2600 2680.7200 ;
        RECT 563.6600 2658.4800 565.2600 2658.9600 ;
        RECT 563.6600 2663.9200 565.2600 2664.4000 ;
        RECT 518.6600 2669.3600 520.2600 2669.8400 ;
        RECT 518.6600 2674.8000 520.2600 2675.2800 ;
        RECT 518.6600 2680.2400 520.2600 2680.7200 ;
        RECT 518.6600 2658.4800 520.2600 2658.9600 ;
        RECT 518.6600 2663.9200 520.2600 2664.4000 ;
        RECT 473.6600 2696.5600 475.2600 2697.0400 ;
        RECT 473.6600 2702.0000 475.2600 2702.4800 ;
        RECT 473.6600 2707.4400 475.2600 2707.9200 ;
        RECT 461.9000 2696.5600 464.9000 2697.0400 ;
        RECT 461.9000 2702.0000 464.9000 2702.4800 ;
        RECT 461.9000 2707.4400 464.9000 2707.9200 ;
        RECT 473.6600 2685.6800 475.2600 2686.1600 ;
        RECT 473.6600 2691.1200 475.2600 2691.6000 ;
        RECT 461.9000 2685.6800 464.9000 2686.1600 ;
        RECT 461.9000 2691.1200 464.9000 2691.6000 ;
        RECT 473.6600 2669.3600 475.2600 2669.8400 ;
        RECT 473.6600 2674.8000 475.2600 2675.2800 ;
        RECT 473.6600 2680.2400 475.2600 2680.7200 ;
        RECT 461.9000 2669.3600 464.9000 2669.8400 ;
        RECT 461.9000 2674.8000 464.9000 2675.2800 ;
        RECT 461.9000 2680.2400 464.9000 2680.7200 ;
        RECT 473.6600 2658.4800 475.2600 2658.9600 ;
        RECT 473.6600 2663.9200 475.2600 2664.4000 ;
        RECT 461.9000 2658.4800 464.9000 2658.9600 ;
        RECT 461.9000 2663.9200 464.9000 2664.4000 ;
        RECT 563.6600 2642.1600 565.2600 2642.6400 ;
        RECT 563.6600 2647.6000 565.2600 2648.0800 ;
        RECT 563.6600 2653.0400 565.2600 2653.5200 ;
        RECT 563.6600 2631.2800 565.2600 2631.7600 ;
        RECT 563.6600 2636.7200 565.2600 2637.2000 ;
        RECT 518.6600 2642.1600 520.2600 2642.6400 ;
        RECT 518.6600 2647.6000 520.2600 2648.0800 ;
        RECT 518.6600 2653.0400 520.2600 2653.5200 ;
        RECT 518.6600 2631.2800 520.2600 2631.7600 ;
        RECT 518.6600 2636.7200 520.2600 2637.2000 ;
        RECT 563.6600 2614.9600 565.2600 2615.4400 ;
        RECT 563.6600 2620.4000 565.2600 2620.8800 ;
        RECT 563.6600 2625.8400 565.2600 2626.3200 ;
        RECT 563.6600 2609.5200 565.2600 2610.0000 ;
        RECT 518.6600 2614.9600 520.2600 2615.4400 ;
        RECT 518.6600 2620.4000 520.2600 2620.8800 ;
        RECT 518.6600 2625.8400 520.2600 2626.3200 ;
        RECT 518.6600 2609.5200 520.2600 2610.0000 ;
        RECT 473.6600 2642.1600 475.2600 2642.6400 ;
        RECT 473.6600 2647.6000 475.2600 2648.0800 ;
        RECT 473.6600 2653.0400 475.2600 2653.5200 ;
        RECT 461.9000 2642.1600 464.9000 2642.6400 ;
        RECT 461.9000 2647.6000 464.9000 2648.0800 ;
        RECT 461.9000 2653.0400 464.9000 2653.5200 ;
        RECT 473.6600 2631.2800 475.2600 2631.7600 ;
        RECT 473.6600 2636.7200 475.2600 2637.2000 ;
        RECT 461.9000 2631.2800 464.9000 2631.7600 ;
        RECT 461.9000 2636.7200 464.9000 2637.2000 ;
        RECT 473.6600 2614.9600 475.2600 2615.4400 ;
        RECT 473.6600 2620.4000 475.2600 2620.8800 ;
        RECT 473.6600 2625.8400 475.2600 2626.3200 ;
        RECT 461.9000 2614.9600 464.9000 2615.4400 ;
        RECT 461.9000 2620.4000 464.9000 2620.8800 ;
        RECT 461.9000 2625.8400 464.9000 2626.3200 ;
        RECT 461.9000 2609.5200 464.9000 2610.0000 ;
        RECT 473.6600 2609.5200 475.2600 2610.0000 ;
        RECT 461.9000 2814.4300 669.0000 2817.4300 ;
        RECT 461.9000 2601.3300 669.0000 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 2371.6900 655.2600 2587.7900 ;
        RECT 608.6600 2371.6900 610.2600 2587.7900 ;
        RECT 563.6600 2371.6900 565.2600 2587.7900 ;
        RECT 518.6600 2371.6900 520.2600 2587.7900 ;
        RECT 473.6600 2371.6900 475.2600 2587.7900 ;
        RECT 666.0000 2371.6900 669.0000 2587.7900 ;
        RECT 461.9000 2371.6900 464.9000 2587.7900 ;
      LAYER met3 ;
        RECT 666.0000 2564.8400 669.0000 2565.3200 ;
        RECT 666.0000 2570.2800 669.0000 2570.7600 ;
        RECT 653.6600 2564.8400 655.2600 2565.3200 ;
        RECT 653.6600 2570.2800 655.2600 2570.7600 ;
        RECT 666.0000 2575.7200 669.0000 2576.2000 ;
        RECT 653.6600 2575.7200 655.2600 2576.2000 ;
        RECT 666.0000 2553.9600 669.0000 2554.4400 ;
        RECT 666.0000 2559.4000 669.0000 2559.8800 ;
        RECT 653.6600 2553.9600 655.2600 2554.4400 ;
        RECT 653.6600 2559.4000 655.2600 2559.8800 ;
        RECT 666.0000 2537.6400 669.0000 2538.1200 ;
        RECT 666.0000 2543.0800 669.0000 2543.5600 ;
        RECT 653.6600 2537.6400 655.2600 2538.1200 ;
        RECT 653.6600 2543.0800 655.2600 2543.5600 ;
        RECT 666.0000 2548.5200 669.0000 2549.0000 ;
        RECT 653.6600 2548.5200 655.2600 2549.0000 ;
        RECT 608.6600 2564.8400 610.2600 2565.3200 ;
        RECT 608.6600 2570.2800 610.2600 2570.7600 ;
        RECT 608.6600 2575.7200 610.2600 2576.2000 ;
        RECT 608.6600 2553.9600 610.2600 2554.4400 ;
        RECT 608.6600 2559.4000 610.2600 2559.8800 ;
        RECT 608.6600 2537.6400 610.2600 2538.1200 ;
        RECT 608.6600 2543.0800 610.2600 2543.5600 ;
        RECT 608.6600 2548.5200 610.2600 2549.0000 ;
        RECT 666.0000 2521.3200 669.0000 2521.8000 ;
        RECT 666.0000 2526.7600 669.0000 2527.2400 ;
        RECT 666.0000 2532.2000 669.0000 2532.6800 ;
        RECT 653.6600 2521.3200 655.2600 2521.8000 ;
        RECT 653.6600 2526.7600 655.2600 2527.2400 ;
        RECT 653.6600 2532.2000 655.2600 2532.6800 ;
        RECT 666.0000 2510.4400 669.0000 2510.9200 ;
        RECT 666.0000 2515.8800 669.0000 2516.3600 ;
        RECT 653.6600 2510.4400 655.2600 2510.9200 ;
        RECT 653.6600 2515.8800 655.2600 2516.3600 ;
        RECT 666.0000 2494.1200 669.0000 2494.6000 ;
        RECT 666.0000 2499.5600 669.0000 2500.0400 ;
        RECT 666.0000 2505.0000 669.0000 2505.4800 ;
        RECT 653.6600 2494.1200 655.2600 2494.6000 ;
        RECT 653.6600 2499.5600 655.2600 2500.0400 ;
        RECT 653.6600 2505.0000 655.2600 2505.4800 ;
        RECT 666.0000 2483.2400 669.0000 2483.7200 ;
        RECT 666.0000 2488.6800 669.0000 2489.1600 ;
        RECT 653.6600 2483.2400 655.2600 2483.7200 ;
        RECT 653.6600 2488.6800 655.2600 2489.1600 ;
        RECT 608.6600 2521.3200 610.2600 2521.8000 ;
        RECT 608.6600 2526.7600 610.2600 2527.2400 ;
        RECT 608.6600 2532.2000 610.2600 2532.6800 ;
        RECT 608.6600 2510.4400 610.2600 2510.9200 ;
        RECT 608.6600 2515.8800 610.2600 2516.3600 ;
        RECT 608.6600 2494.1200 610.2600 2494.6000 ;
        RECT 608.6600 2499.5600 610.2600 2500.0400 ;
        RECT 608.6600 2505.0000 610.2600 2505.4800 ;
        RECT 608.6600 2483.2400 610.2600 2483.7200 ;
        RECT 608.6600 2488.6800 610.2600 2489.1600 ;
        RECT 563.6600 2564.8400 565.2600 2565.3200 ;
        RECT 563.6600 2570.2800 565.2600 2570.7600 ;
        RECT 563.6600 2575.7200 565.2600 2576.2000 ;
        RECT 518.6600 2564.8400 520.2600 2565.3200 ;
        RECT 518.6600 2570.2800 520.2600 2570.7600 ;
        RECT 518.6600 2575.7200 520.2600 2576.2000 ;
        RECT 563.6600 2553.9600 565.2600 2554.4400 ;
        RECT 563.6600 2559.4000 565.2600 2559.8800 ;
        RECT 563.6600 2537.6400 565.2600 2538.1200 ;
        RECT 563.6600 2543.0800 565.2600 2543.5600 ;
        RECT 563.6600 2548.5200 565.2600 2549.0000 ;
        RECT 518.6600 2553.9600 520.2600 2554.4400 ;
        RECT 518.6600 2559.4000 520.2600 2559.8800 ;
        RECT 518.6600 2537.6400 520.2600 2538.1200 ;
        RECT 518.6600 2543.0800 520.2600 2543.5600 ;
        RECT 518.6600 2548.5200 520.2600 2549.0000 ;
        RECT 473.6600 2564.8400 475.2600 2565.3200 ;
        RECT 473.6600 2570.2800 475.2600 2570.7600 ;
        RECT 461.9000 2570.2800 464.9000 2570.7600 ;
        RECT 461.9000 2564.8400 464.9000 2565.3200 ;
        RECT 461.9000 2575.7200 464.9000 2576.2000 ;
        RECT 473.6600 2575.7200 475.2600 2576.2000 ;
        RECT 473.6600 2553.9600 475.2600 2554.4400 ;
        RECT 473.6600 2559.4000 475.2600 2559.8800 ;
        RECT 461.9000 2559.4000 464.9000 2559.8800 ;
        RECT 461.9000 2553.9600 464.9000 2554.4400 ;
        RECT 473.6600 2537.6400 475.2600 2538.1200 ;
        RECT 473.6600 2543.0800 475.2600 2543.5600 ;
        RECT 461.9000 2543.0800 464.9000 2543.5600 ;
        RECT 461.9000 2537.6400 464.9000 2538.1200 ;
        RECT 461.9000 2548.5200 464.9000 2549.0000 ;
        RECT 473.6600 2548.5200 475.2600 2549.0000 ;
        RECT 563.6600 2521.3200 565.2600 2521.8000 ;
        RECT 563.6600 2526.7600 565.2600 2527.2400 ;
        RECT 563.6600 2532.2000 565.2600 2532.6800 ;
        RECT 563.6600 2510.4400 565.2600 2510.9200 ;
        RECT 563.6600 2515.8800 565.2600 2516.3600 ;
        RECT 518.6600 2521.3200 520.2600 2521.8000 ;
        RECT 518.6600 2526.7600 520.2600 2527.2400 ;
        RECT 518.6600 2532.2000 520.2600 2532.6800 ;
        RECT 518.6600 2510.4400 520.2600 2510.9200 ;
        RECT 518.6600 2515.8800 520.2600 2516.3600 ;
        RECT 563.6600 2494.1200 565.2600 2494.6000 ;
        RECT 563.6600 2499.5600 565.2600 2500.0400 ;
        RECT 563.6600 2505.0000 565.2600 2505.4800 ;
        RECT 563.6600 2483.2400 565.2600 2483.7200 ;
        RECT 563.6600 2488.6800 565.2600 2489.1600 ;
        RECT 518.6600 2494.1200 520.2600 2494.6000 ;
        RECT 518.6600 2499.5600 520.2600 2500.0400 ;
        RECT 518.6600 2505.0000 520.2600 2505.4800 ;
        RECT 518.6600 2483.2400 520.2600 2483.7200 ;
        RECT 518.6600 2488.6800 520.2600 2489.1600 ;
        RECT 473.6600 2521.3200 475.2600 2521.8000 ;
        RECT 473.6600 2526.7600 475.2600 2527.2400 ;
        RECT 473.6600 2532.2000 475.2600 2532.6800 ;
        RECT 461.9000 2521.3200 464.9000 2521.8000 ;
        RECT 461.9000 2526.7600 464.9000 2527.2400 ;
        RECT 461.9000 2532.2000 464.9000 2532.6800 ;
        RECT 473.6600 2510.4400 475.2600 2510.9200 ;
        RECT 473.6600 2515.8800 475.2600 2516.3600 ;
        RECT 461.9000 2510.4400 464.9000 2510.9200 ;
        RECT 461.9000 2515.8800 464.9000 2516.3600 ;
        RECT 473.6600 2494.1200 475.2600 2494.6000 ;
        RECT 473.6600 2499.5600 475.2600 2500.0400 ;
        RECT 473.6600 2505.0000 475.2600 2505.4800 ;
        RECT 461.9000 2494.1200 464.9000 2494.6000 ;
        RECT 461.9000 2499.5600 464.9000 2500.0400 ;
        RECT 461.9000 2505.0000 464.9000 2505.4800 ;
        RECT 473.6600 2483.2400 475.2600 2483.7200 ;
        RECT 473.6600 2488.6800 475.2600 2489.1600 ;
        RECT 461.9000 2483.2400 464.9000 2483.7200 ;
        RECT 461.9000 2488.6800 464.9000 2489.1600 ;
        RECT 666.0000 2466.9200 669.0000 2467.4000 ;
        RECT 666.0000 2472.3600 669.0000 2472.8400 ;
        RECT 666.0000 2477.8000 669.0000 2478.2800 ;
        RECT 653.6600 2466.9200 655.2600 2467.4000 ;
        RECT 653.6600 2472.3600 655.2600 2472.8400 ;
        RECT 653.6600 2477.8000 655.2600 2478.2800 ;
        RECT 666.0000 2456.0400 669.0000 2456.5200 ;
        RECT 666.0000 2461.4800 669.0000 2461.9600 ;
        RECT 653.6600 2456.0400 655.2600 2456.5200 ;
        RECT 653.6600 2461.4800 655.2600 2461.9600 ;
        RECT 666.0000 2439.7200 669.0000 2440.2000 ;
        RECT 666.0000 2445.1600 669.0000 2445.6400 ;
        RECT 666.0000 2450.6000 669.0000 2451.0800 ;
        RECT 653.6600 2439.7200 655.2600 2440.2000 ;
        RECT 653.6600 2445.1600 655.2600 2445.6400 ;
        RECT 653.6600 2450.6000 655.2600 2451.0800 ;
        RECT 666.0000 2428.8400 669.0000 2429.3200 ;
        RECT 666.0000 2434.2800 669.0000 2434.7600 ;
        RECT 653.6600 2428.8400 655.2600 2429.3200 ;
        RECT 653.6600 2434.2800 655.2600 2434.7600 ;
        RECT 608.6600 2466.9200 610.2600 2467.4000 ;
        RECT 608.6600 2472.3600 610.2600 2472.8400 ;
        RECT 608.6600 2477.8000 610.2600 2478.2800 ;
        RECT 608.6600 2456.0400 610.2600 2456.5200 ;
        RECT 608.6600 2461.4800 610.2600 2461.9600 ;
        RECT 608.6600 2439.7200 610.2600 2440.2000 ;
        RECT 608.6600 2445.1600 610.2600 2445.6400 ;
        RECT 608.6600 2450.6000 610.2600 2451.0800 ;
        RECT 608.6600 2428.8400 610.2600 2429.3200 ;
        RECT 608.6600 2434.2800 610.2600 2434.7600 ;
        RECT 666.0000 2412.5200 669.0000 2413.0000 ;
        RECT 666.0000 2417.9600 669.0000 2418.4400 ;
        RECT 666.0000 2423.4000 669.0000 2423.8800 ;
        RECT 653.6600 2412.5200 655.2600 2413.0000 ;
        RECT 653.6600 2417.9600 655.2600 2418.4400 ;
        RECT 653.6600 2423.4000 655.2600 2423.8800 ;
        RECT 666.0000 2401.6400 669.0000 2402.1200 ;
        RECT 666.0000 2407.0800 669.0000 2407.5600 ;
        RECT 653.6600 2401.6400 655.2600 2402.1200 ;
        RECT 653.6600 2407.0800 655.2600 2407.5600 ;
        RECT 666.0000 2385.3200 669.0000 2385.8000 ;
        RECT 666.0000 2390.7600 669.0000 2391.2400 ;
        RECT 666.0000 2396.2000 669.0000 2396.6800 ;
        RECT 653.6600 2385.3200 655.2600 2385.8000 ;
        RECT 653.6600 2390.7600 655.2600 2391.2400 ;
        RECT 653.6600 2396.2000 655.2600 2396.6800 ;
        RECT 666.0000 2379.8800 669.0000 2380.3600 ;
        RECT 653.6600 2379.8800 655.2600 2380.3600 ;
        RECT 608.6600 2412.5200 610.2600 2413.0000 ;
        RECT 608.6600 2417.9600 610.2600 2418.4400 ;
        RECT 608.6600 2423.4000 610.2600 2423.8800 ;
        RECT 608.6600 2401.6400 610.2600 2402.1200 ;
        RECT 608.6600 2407.0800 610.2600 2407.5600 ;
        RECT 608.6600 2385.3200 610.2600 2385.8000 ;
        RECT 608.6600 2390.7600 610.2600 2391.2400 ;
        RECT 608.6600 2396.2000 610.2600 2396.6800 ;
        RECT 608.6600 2379.8800 610.2600 2380.3600 ;
        RECT 563.6600 2466.9200 565.2600 2467.4000 ;
        RECT 563.6600 2472.3600 565.2600 2472.8400 ;
        RECT 563.6600 2477.8000 565.2600 2478.2800 ;
        RECT 563.6600 2456.0400 565.2600 2456.5200 ;
        RECT 563.6600 2461.4800 565.2600 2461.9600 ;
        RECT 518.6600 2466.9200 520.2600 2467.4000 ;
        RECT 518.6600 2472.3600 520.2600 2472.8400 ;
        RECT 518.6600 2477.8000 520.2600 2478.2800 ;
        RECT 518.6600 2456.0400 520.2600 2456.5200 ;
        RECT 518.6600 2461.4800 520.2600 2461.9600 ;
        RECT 563.6600 2439.7200 565.2600 2440.2000 ;
        RECT 563.6600 2445.1600 565.2600 2445.6400 ;
        RECT 563.6600 2450.6000 565.2600 2451.0800 ;
        RECT 563.6600 2428.8400 565.2600 2429.3200 ;
        RECT 563.6600 2434.2800 565.2600 2434.7600 ;
        RECT 518.6600 2439.7200 520.2600 2440.2000 ;
        RECT 518.6600 2445.1600 520.2600 2445.6400 ;
        RECT 518.6600 2450.6000 520.2600 2451.0800 ;
        RECT 518.6600 2428.8400 520.2600 2429.3200 ;
        RECT 518.6600 2434.2800 520.2600 2434.7600 ;
        RECT 473.6600 2466.9200 475.2600 2467.4000 ;
        RECT 473.6600 2472.3600 475.2600 2472.8400 ;
        RECT 473.6600 2477.8000 475.2600 2478.2800 ;
        RECT 461.9000 2466.9200 464.9000 2467.4000 ;
        RECT 461.9000 2472.3600 464.9000 2472.8400 ;
        RECT 461.9000 2477.8000 464.9000 2478.2800 ;
        RECT 473.6600 2456.0400 475.2600 2456.5200 ;
        RECT 473.6600 2461.4800 475.2600 2461.9600 ;
        RECT 461.9000 2456.0400 464.9000 2456.5200 ;
        RECT 461.9000 2461.4800 464.9000 2461.9600 ;
        RECT 473.6600 2439.7200 475.2600 2440.2000 ;
        RECT 473.6600 2445.1600 475.2600 2445.6400 ;
        RECT 473.6600 2450.6000 475.2600 2451.0800 ;
        RECT 461.9000 2439.7200 464.9000 2440.2000 ;
        RECT 461.9000 2445.1600 464.9000 2445.6400 ;
        RECT 461.9000 2450.6000 464.9000 2451.0800 ;
        RECT 473.6600 2428.8400 475.2600 2429.3200 ;
        RECT 473.6600 2434.2800 475.2600 2434.7600 ;
        RECT 461.9000 2428.8400 464.9000 2429.3200 ;
        RECT 461.9000 2434.2800 464.9000 2434.7600 ;
        RECT 563.6600 2412.5200 565.2600 2413.0000 ;
        RECT 563.6600 2417.9600 565.2600 2418.4400 ;
        RECT 563.6600 2423.4000 565.2600 2423.8800 ;
        RECT 563.6600 2401.6400 565.2600 2402.1200 ;
        RECT 563.6600 2407.0800 565.2600 2407.5600 ;
        RECT 518.6600 2412.5200 520.2600 2413.0000 ;
        RECT 518.6600 2417.9600 520.2600 2418.4400 ;
        RECT 518.6600 2423.4000 520.2600 2423.8800 ;
        RECT 518.6600 2401.6400 520.2600 2402.1200 ;
        RECT 518.6600 2407.0800 520.2600 2407.5600 ;
        RECT 563.6600 2385.3200 565.2600 2385.8000 ;
        RECT 563.6600 2390.7600 565.2600 2391.2400 ;
        RECT 563.6600 2396.2000 565.2600 2396.6800 ;
        RECT 563.6600 2379.8800 565.2600 2380.3600 ;
        RECT 518.6600 2385.3200 520.2600 2385.8000 ;
        RECT 518.6600 2390.7600 520.2600 2391.2400 ;
        RECT 518.6600 2396.2000 520.2600 2396.6800 ;
        RECT 518.6600 2379.8800 520.2600 2380.3600 ;
        RECT 473.6600 2412.5200 475.2600 2413.0000 ;
        RECT 473.6600 2417.9600 475.2600 2418.4400 ;
        RECT 473.6600 2423.4000 475.2600 2423.8800 ;
        RECT 461.9000 2412.5200 464.9000 2413.0000 ;
        RECT 461.9000 2417.9600 464.9000 2418.4400 ;
        RECT 461.9000 2423.4000 464.9000 2423.8800 ;
        RECT 473.6600 2401.6400 475.2600 2402.1200 ;
        RECT 473.6600 2407.0800 475.2600 2407.5600 ;
        RECT 461.9000 2401.6400 464.9000 2402.1200 ;
        RECT 461.9000 2407.0800 464.9000 2407.5600 ;
        RECT 473.6600 2385.3200 475.2600 2385.8000 ;
        RECT 473.6600 2390.7600 475.2600 2391.2400 ;
        RECT 473.6600 2396.2000 475.2600 2396.6800 ;
        RECT 461.9000 2385.3200 464.9000 2385.8000 ;
        RECT 461.9000 2390.7600 464.9000 2391.2400 ;
        RECT 461.9000 2396.2000 464.9000 2396.6800 ;
        RECT 461.9000 2379.8800 464.9000 2380.3600 ;
        RECT 473.6600 2379.8800 475.2600 2380.3600 ;
        RECT 461.9000 2584.7900 669.0000 2587.7900 ;
        RECT 461.9000 2371.6900 669.0000 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 2142.0500 655.2600 2358.1500 ;
        RECT 608.6600 2142.0500 610.2600 2358.1500 ;
        RECT 563.6600 2142.0500 565.2600 2358.1500 ;
        RECT 518.6600 2142.0500 520.2600 2358.1500 ;
        RECT 473.6600 2142.0500 475.2600 2358.1500 ;
        RECT 666.0000 2142.0500 669.0000 2358.1500 ;
        RECT 461.9000 2142.0500 464.9000 2358.1500 ;
      LAYER met3 ;
        RECT 666.0000 2335.2000 669.0000 2335.6800 ;
        RECT 666.0000 2340.6400 669.0000 2341.1200 ;
        RECT 653.6600 2335.2000 655.2600 2335.6800 ;
        RECT 653.6600 2340.6400 655.2600 2341.1200 ;
        RECT 666.0000 2346.0800 669.0000 2346.5600 ;
        RECT 653.6600 2346.0800 655.2600 2346.5600 ;
        RECT 666.0000 2324.3200 669.0000 2324.8000 ;
        RECT 666.0000 2329.7600 669.0000 2330.2400 ;
        RECT 653.6600 2324.3200 655.2600 2324.8000 ;
        RECT 653.6600 2329.7600 655.2600 2330.2400 ;
        RECT 666.0000 2308.0000 669.0000 2308.4800 ;
        RECT 666.0000 2313.4400 669.0000 2313.9200 ;
        RECT 653.6600 2308.0000 655.2600 2308.4800 ;
        RECT 653.6600 2313.4400 655.2600 2313.9200 ;
        RECT 666.0000 2318.8800 669.0000 2319.3600 ;
        RECT 653.6600 2318.8800 655.2600 2319.3600 ;
        RECT 608.6600 2335.2000 610.2600 2335.6800 ;
        RECT 608.6600 2340.6400 610.2600 2341.1200 ;
        RECT 608.6600 2346.0800 610.2600 2346.5600 ;
        RECT 608.6600 2324.3200 610.2600 2324.8000 ;
        RECT 608.6600 2329.7600 610.2600 2330.2400 ;
        RECT 608.6600 2308.0000 610.2600 2308.4800 ;
        RECT 608.6600 2313.4400 610.2600 2313.9200 ;
        RECT 608.6600 2318.8800 610.2600 2319.3600 ;
        RECT 666.0000 2291.6800 669.0000 2292.1600 ;
        RECT 666.0000 2297.1200 669.0000 2297.6000 ;
        RECT 666.0000 2302.5600 669.0000 2303.0400 ;
        RECT 653.6600 2291.6800 655.2600 2292.1600 ;
        RECT 653.6600 2297.1200 655.2600 2297.6000 ;
        RECT 653.6600 2302.5600 655.2600 2303.0400 ;
        RECT 666.0000 2280.8000 669.0000 2281.2800 ;
        RECT 666.0000 2286.2400 669.0000 2286.7200 ;
        RECT 653.6600 2280.8000 655.2600 2281.2800 ;
        RECT 653.6600 2286.2400 655.2600 2286.7200 ;
        RECT 666.0000 2264.4800 669.0000 2264.9600 ;
        RECT 666.0000 2269.9200 669.0000 2270.4000 ;
        RECT 666.0000 2275.3600 669.0000 2275.8400 ;
        RECT 653.6600 2264.4800 655.2600 2264.9600 ;
        RECT 653.6600 2269.9200 655.2600 2270.4000 ;
        RECT 653.6600 2275.3600 655.2600 2275.8400 ;
        RECT 666.0000 2253.6000 669.0000 2254.0800 ;
        RECT 666.0000 2259.0400 669.0000 2259.5200 ;
        RECT 653.6600 2253.6000 655.2600 2254.0800 ;
        RECT 653.6600 2259.0400 655.2600 2259.5200 ;
        RECT 608.6600 2291.6800 610.2600 2292.1600 ;
        RECT 608.6600 2297.1200 610.2600 2297.6000 ;
        RECT 608.6600 2302.5600 610.2600 2303.0400 ;
        RECT 608.6600 2280.8000 610.2600 2281.2800 ;
        RECT 608.6600 2286.2400 610.2600 2286.7200 ;
        RECT 608.6600 2264.4800 610.2600 2264.9600 ;
        RECT 608.6600 2269.9200 610.2600 2270.4000 ;
        RECT 608.6600 2275.3600 610.2600 2275.8400 ;
        RECT 608.6600 2253.6000 610.2600 2254.0800 ;
        RECT 608.6600 2259.0400 610.2600 2259.5200 ;
        RECT 563.6600 2335.2000 565.2600 2335.6800 ;
        RECT 563.6600 2340.6400 565.2600 2341.1200 ;
        RECT 563.6600 2346.0800 565.2600 2346.5600 ;
        RECT 518.6600 2335.2000 520.2600 2335.6800 ;
        RECT 518.6600 2340.6400 520.2600 2341.1200 ;
        RECT 518.6600 2346.0800 520.2600 2346.5600 ;
        RECT 563.6600 2324.3200 565.2600 2324.8000 ;
        RECT 563.6600 2329.7600 565.2600 2330.2400 ;
        RECT 563.6600 2308.0000 565.2600 2308.4800 ;
        RECT 563.6600 2313.4400 565.2600 2313.9200 ;
        RECT 563.6600 2318.8800 565.2600 2319.3600 ;
        RECT 518.6600 2324.3200 520.2600 2324.8000 ;
        RECT 518.6600 2329.7600 520.2600 2330.2400 ;
        RECT 518.6600 2308.0000 520.2600 2308.4800 ;
        RECT 518.6600 2313.4400 520.2600 2313.9200 ;
        RECT 518.6600 2318.8800 520.2600 2319.3600 ;
        RECT 473.6600 2335.2000 475.2600 2335.6800 ;
        RECT 473.6600 2340.6400 475.2600 2341.1200 ;
        RECT 461.9000 2340.6400 464.9000 2341.1200 ;
        RECT 461.9000 2335.2000 464.9000 2335.6800 ;
        RECT 461.9000 2346.0800 464.9000 2346.5600 ;
        RECT 473.6600 2346.0800 475.2600 2346.5600 ;
        RECT 473.6600 2324.3200 475.2600 2324.8000 ;
        RECT 473.6600 2329.7600 475.2600 2330.2400 ;
        RECT 461.9000 2329.7600 464.9000 2330.2400 ;
        RECT 461.9000 2324.3200 464.9000 2324.8000 ;
        RECT 473.6600 2308.0000 475.2600 2308.4800 ;
        RECT 473.6600 2313.4400 475.2600 2313.9200 ;
        RECT 461.9000 2313.4400 464.9000 2313.9200 ;
        RECT 461.9000 2308.0000 464.9000 2308.4800 ;
        RECT 461.9000 2318.8800 464.9000 2319.3600 ;
        RECT 473.6600 2318.8800 475.2600 2319.3600 ;
        RECT 563.6600 2291.6800 565.2600 2292.1600 ;
        RECT 563.6600 2297.1200 565.2600 2297.6000 ;
        RECT 563.6600 2302.5600 565.2600 2303.0400 ;
        RECT 563.6600 2280.8000 565.2600 2281.2800 ;
        RECT 563.6600 2286.2400 565.2600 2286.7200 ;
        RECT 518.6600 2291.6800 520.2600 2292.1600 ;
        RECT 518.6600 2297.1200 520.2600 2297.6000 ;
        RECT 518.6600 2302.5600 520.2600 2303.0400 ;
        RECT 518.6600 2280.8000 520.2600 2281.2800 ;
        RECT 518.6600 2286.2400 520.2600 2286.7200 ;
        RECT 563.6600 2264.4800 565.2600 2264.9600 ;
        RECT 563.6600 2269.9200 565.2600 2270.4000 ;
        RECT 563.6600 2275.3600 565.2600 2275.8400 ;
        RECT 563.6600 2253.6000 565.2600 2254.0800 ;
        RECT 563.6600 2259.0400 565.2600 2259.5200 ;
        RECT 518.6600 2264.4800 520.2600 2264.9600 ;
        RECT 518.6600 2269.9200 520.2600 2270.4000 ;
        RECT 518.6600 2275.3600 520.2600 2275.8400 ;
        RECT 518.6600 2253.6000 520.2600 2254.0800 ;
        RECT 518.6600 2259.0400 520.2600 2259.5200 ;
        RECT 473.6600 2291.6800 475.2600 2292.1600 ;
        RECT 473.6600 2297.1200 475.2600 2297.6000 ;
        RECT 473.6600 2302.5600 475.2600 2303.0400 ;
        RECT 461.9000 2291.6800 464.9000 2292.1600 ;
        RECT 461.9000 2297.1200 464.9000 2297.6000 ;
        RECT 461.9000 2302.5600 464.9000 2303.0400 ;
        RECT 473.6600 2280.8000 475.2600 2281.2800 ;
        RECT 473.6600 2286.2400 475.2600 2286.7200 ;
        RECT 461.9000 2280.8000 464.9000 2281.2800 ;
        RECT 461.9000 2286.2400 464.9000 2286.7200 ;
        RECT 473.6600 2264.4800 475.2600 2264.9600 ;
        RECT 473.6600 2269.9200 475.2600 2270.4000 ;
        RECT 473.6600 2275.3600 475.2600 2275.8400 ;
        RECT 461.9000 2264.4800 464.9000 2264.9600 ;
        RECT 461.9000 2269.9200 464.9000 2270.4000 ;
        RECT 461.9000 2275.3600 464.9000 2275.8400 ;
        RECT 473.6600 2253.6000 475.2600 2254.0800 ;
        RECT 473.6600 2259.0400 475.2600 2259.5200 ;
        RECT 461.9000 2253.6000 464.9000 2254.0800 ;
        RECT 461.9000 2259.0400 464.9000 2259.5200 ;
        RECT 666.0000 2237.2800 669.0000 2237.7600 ;
        RECT 666.0000 2242.7200 669.0000 2243.2000 ;
        RECT 666.0000 2248.1600 669.0000 2248.6400 ;
        RECT 653.6600 2237.2800 655.2600 2237.7600 ;
        RECT 653.6600 2242.7200 655.2600 2243.2000 ;
        RECT 653.6600 2248.1600 655.2600 2248.6400 ;
        RECT 666.0000 2226.4000 669.0000 2226.8800 ;
        RECT 666.0000 2231.8400 669.0000 2232.3200 ;
        RECT 653.6600 2226.4000 655.2600 2226.8800 ;
        RECT 653.6600 2231.8400 655.2600 2232.3200 ;
        RECT 666.0000 2210.0800 669.0000 2210.5600 ;
        RECT 666.0000 2215.5200 669.0000 2216.0000 ;
        RECT 666.0000 2220.9600 669.0000 2221.4400 ;
        RECT 653.6600 2210.0800 655.2600 2210.5600 ;
        RECT 653.6600 2215.5200 655.2600 2216.0000 ;
        RECT 653.6600 2220.9600 655.2600 2221.4400 ;
        RECT 666.0000 2199.2000 669.0000 2199.6800 ;
        RECT 666.0000 2204.6400 669.0000 2205.1200 ;
        RECT 653.6600 2199.2000 655.2600 2199.6800 ;
        RECT 653.6600 2204.6400 655.2600 2205.1200 ;
        RECT 608.6600 2237.2800 610.2600 2237.7600 ;
        RECT 608.6600 2242.7200 610.2600 2243.2000 ;
        RECT 608.6600 2248.1600 610.2600 2248.6400 ;
        RECT 608.6600 2226.4000 610.2600 2226.8800 ;
        RECT 608.6600 2231.8400 610.2600 2232.3200 ;
        RECT 608.6600 2210.0800 610.2600 2210.5600 ;
        RECT 608.6600 2215.5200 610.2600 2216.0000 ;
        RECT 608.6600 2220.9600 610.2600 2221.4400 ;
        RECT 608.6600 2199.2000 610.2600 2199.6800 ;
        RECT 608.6600 2204.6400 610.2600 2205.1200 ;
        RECT 666.0000 2182.8800 669.0000 2183.3600 ;
        RECT 666.0000 2188.3200 669.0000 2188.8000 ;
        RECT 666.0000 2193.7600 669.0000 2194.2400 ;
        RECT 653.6600 2182.8800 655.2600 2183.3600 ;
        RECT 653.6600 2188.3200 655.2600 2188.8000 ;
        RECT 653.6600 2193.7600 655.2600 2194.2400 ;
        RECT 666.0000 2172.0000 669.0000 2172.4800 ;
        RECT 666.0000 2177.4400 669.0000 2177.9200 ;
        RECT 653.6600 2172.0000 655.2600 2172.4800 ;
        RECT 653.6600 2177.4400 655.2600 2177.9200 ;
        RECT 666.0000 2155.6800 669.0000 2156.1600 ;
        RECT 666.0000 2161.1200 669.0000 2161.6000 ;
        RECT 666.0000 2166.5600 669.0000 2167.0400 ;
        RECT 653.6600 2155.6800 655.2600 2156.1600 ;
        RECT 653.6600 2161.1200 655.2600 2161.6000 ;
        RECT 653.6600 2166.5600 655.2600 2167.0400 ;
        RECT 666.0000 2150.2400 669.0000 2150.7200 ;
        RECT 653.6600 2150.2400 655.2600 2150.7200 ;
        RECT 608.6600 2182.8800 610.2600 2183.3600 ;
        RECT 608.6600 2188.3200 610.2600 2188.8000 ;
        RECT 608.6600 2193.7600 610.2600 2194.2400 ;
        RECT 608.6600 2172.0000 610.2600 2172.4800 ;
        RECT 608.6600 2177.4400 610.2600 2177.9200 ;
        RECT 608.6600 2155.6800 610.2600 2156.1600 ;
        RECT 608.6600 2161.1200 610.2600 2161.6000 ;
        RECT 608.6600 2166.5600 610.2600 2167.0400 ;
        RECT 608.6600 2150.2400 610.2600 2150.7200 ;
        RECT 563.6600 2237.2800 565.2600 2237.7600 ;
        RECT 563.6600 2242.7200 565.2600 2243.2000 ;
        RECT 563.6600 2248.1600 565.2600 2248.6400 ;
        RECT 563.6600 2226.4000 565.2600 2226.8800 ;
        RECT 563.6600 2231.8400 565.2600 2232.3200 ;
        RECT 518.6600 2237.2800 520.2600 2237.7600 ;
        RECT 518.6600 2242.7200 520.2600 2243.2000 ;
        RECT 518.6600 2248.1600 520.2600 2248.6400 ;
        RECT 518.6600 2226.4000 520.2600 2226.8800 ;
        RECT 518.6600 2231.8400 520.2600 2232.3200 ;
        RECT 563.6600 2210.0800 565.2600 2210.5600 ;
        RECT 563.6600 2215.5200 565.2600 2216.0000 ;
        RECT 563.6600 2220.9600 565.2600 2221.4400 ;
        RECT 563.6600 2199.2000 565.2600 2199.6800 ;
        RECT 563.6600 2204.6400 565.2600 2205.1200 ;
        RECT 518.6600 2210.0800 520.2600 2210.5600 ;
        RECT 518.6600 2215.5200 520.2600 2216.0000 ;
        RECT 518.6600 2220.9600 520.2600 2221.4400 ;
        RECT 518.6600 2199.2000 520.2600 2199.6800 ;
        RECT 518.6600 2204.6400 520.2600 2205.1200 ;
        RECT 473.6600 2237.2800 475.2600 2237.7600 ;
        RECT 473.6600 2242.7200 475.2600 2243.2000 ;
        RECT 473.6600 2248.1600 475.2600 2248.6400 ;
        RECT 461.9000 2237.2800 464.9000 2237.7600 ;
        RECT 461.9000 2242.7200 464.9000 2243.2000 ;
        RECT 461.9000 2248.1600 464.9000 2248.6400 ;
        RECT 473.6600 2226.4000 475.2600 2226.8800 ;
        RECT 473.6600 2231.8400 475.2600 2232.3200 ;
        RECT 461.9000 2226.4000 464.9000 2226.8800 ;
        RECT 461.9000 2231.8400 464.9000 2232.3200 ;
        RECT 473.6600 2210.0800 475.2600 2210.5600 ;
        RECT 473.6600 2215.5200 475.2600 2216.0000 ;
        RECT 473.6600 2220.9600 475.2600 2221.4400 ;
        RECT 461.9000 2210.0800 464.9000 2210.5600 ;
        RECT 461.9000 2215.5200 464.9000 2216.0000 ;
        RECT 461.9000 2220.9600 464.9000 2221.4400 ;
        RECT 473.6600 2199.2000 475.2600 2199.6800 ;
        RECT 473.6600 2204.6400 475.2600 2205.1200 ;
        RECT 461.9000 2199.2000 464.9000 2199.6800 ;
        RECT 461.9000 2204.6400 464.9000 2205.1200 ;
        RECT 563.6600 2182.8800 565.2600 2183.3600 ;
        RECT 563.6600 2188.3200 565.2600 2188.8000 ;
        RECT 563.6600 2193.7600 565.2600 2194.2400 ;
        RECT 563.6600 2172.0000 565.2600 2172.4800 ;
        RECT 563.6600 2177.4400 565.2600 2177.9200 ;
        RECT 518.6600 2182.8800 520.2600 2183.3600 ;
        RECT 518.6600 2188.3200 520.2600 2188.8000 ;
        RECT 518.6600 2193.7600 520.2600 2194.2400 ;
        RECT 518.6600 2172.0000 520.2600 2172.4800 ;
        RECT 518.6600 2177.4400 520.2600 2177.9200 ;
        RECT 563.6600 2155.6800 565.2600 2156.1600 ;
        RECT 563.6600 2161.1200 565.2600 2161.6000 ;
        RECT 563.6600 2166.5600 565.2600 2167.0400 ;
        RECT 563.6600 2150.2400 565.2600 2150.7200 ;
        RECT 518.6600 2155.6800 520.2600 2156.1600 ;
        RECT 518.6600 2161.1200 520.2600 2161.6000 ;
        RECT 518.6600 2166.5600 520.2600 2167.0400 ;
        RECT 518.6600 2150.2400 520.2600 2150.7200 ;
        RECT 473.6600 2182.8800 475.2600 2183.3600 ;
        RECT 473.6600 2188.3200 475.2600 2188.8000 ;
        RECT 473.6600 2193.7600 475.2600 2194.2400 ;
        RECT 461.9000 2182.8800 464.9000 2183.3600 ;
        RECT 461.9000 2188.3200 464.9000 2188.8000 ;
        RECT 461.9000 2193.7600 464.9000 2194.2400 ;
        RECT 473.6600 2172.0000 475.2600 2172.4800 ;
        RECT 473.6600 2177.4400 475.2600 2177.9200 ;
        RECT 461.9000 2172.0000 464.9000 2172.4800 ;
        RECT 461.9000 2177.4400 464.9000 2177.9200 ;
        RECT 473.6600 2155.6800 475.2600 2156.1600 ;
        RECT 473.6600 2161.1200 475.2600 2161.6000 ;
        RECT 473.6600 2166.5600 475.2600 2167.0400 ;
        RECT 461.9000 2155.6800 464.9000 2156.1600 ;
        RECT 461.9000 2161.1200 464.9000 2161.6000 ;
        RECT 461.9000 2166.5600 464.9000 2167.0400 ;
        RECT 461.9000 2150.2400 464.9000 2150.7200 ;
        RECT 473.6600 2150.2400 475.2600 2150.7200 ;
        RECT 461.9000 2355.1500 669.0000 2358.1500 ;
        RECT 461.9000 2142.0500 669.0000 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 1912.4100 655.2600 2128.5100 ;
        RECT 608.6600 1912.4100 610.2600 2128.5100 ;
        RECT 563.6600 1912.4100 565.2600 2128.5100 ;
        RECT 518.6600 1912.4100 520.2600 2128.5100 ;
        RECT 473.6600 1912.4100 475.2600 2128.5100 ;
        RECT 666.0000 1912.4100 669.0000 2128.5100 ;
        RECT 461.9000 1912.4100 464.9000 2128.5100 ;
      LAYER met3 ;
        RECT 666.0000 2105.5600 669.0000 2106.0400 ;
        RECT 666.0000 2111.0000 669.0000 2111.4800 ;
        RECT 653.6600 2105.5600 655.2600 2106.0400 ;
        RECT 653.6600 2111.0000 655.2600 2111.4800 ;
        RECT 666.0000 2116.4400 669.0000 2116.9200 ;
        RECT 653.6600 2116.4400 655.2600 2116.9200 ;
        RECT 666.0000 2094.6800 669.0000 2095.1600 ;
        RECT 666.0000 2100.1200 669.0000 2100.6000 ;
        RECT 653.6600 2094.6800 655.2600 2095.1600 ;
        RECT 653.6600 2100.1200 655.2600 2100.6000 ;
        RECT 666.0000 2078.3600 669.0000 2078.8400 ;
        RECT 666.0000 2083.8000 669.0000 2084.2800 ;
        RECT 653.6600 2078.3600 655.2600 2078.8400 ;
        RECT 653.6600 2083.8000 655.2600 2084.2800 ;
        RECT 666.0000 2089.2400 669.0000 2089.7200 ;
        RECT 653.6600 2089.2400 655.2600 2089.7200 ;
        RECT 608.6600 2105.5600 610.2600 2106.0400 ;
        RECT 608.6600 2111.0000 610.2600 2111.4800 ;
        RECT 608.6600 2116.4400 610.2600 2116.9200 ;
        RECT 608.6600 2094.6800 610.2600 2095.1600 ;
        RECT 608.6600 2100.1200 610.2600 2100.6000 ;
        RECT 608.6600 2078.3600 610.2600 2078.8400 ;
        RECT 608.6600 2083.8000 610.2600 2084.2800 ;
        RECT 608.6600 2089.2400 610.2600 2089.7200 ;
        RECT 666.0000 2062.0400 669.0000 2062.5200 ;
        RECT 666.0000 2067.4800 669.0000 2067.9600 ;
        RECT 666.0000 2072.9200 669.0000 2073.4000 ;
        RECT 653.6600 2062.0400 655.2600 2062.5200 ;
        RECT 653.6600 2067.4800 655.2600 2067.9600 ;
        RECT 653.6600 2072.9200 655.2600 2073.4000 ;
        RECT 666.0000 2051.1600 669.0000 2051.6400 ;
        RECT 666.0000 2056.6000 669.0000 2057.0800 ;
        RECT 653.6600 2051.1600 655.2600 2051.6400 ;
        RECT 653.6600 2056.6000 655.2600 2057.0800 ;
        RECT 666.0000 2034.8400 669.0000 2035.3200 ;
        RECT 666.0000 2040.2800 669.0000 2040.7600 ;
        RECT 666.0000 2045.7200 669.0000 2046.2000 ;
        RECT 653.6600 2034.8400 655.2600 2035.3200 ;
        RECT 653.6600 2040.2800 655.2600 2040.7600 ;
        RECT 653.6600 2045.7200 655.2600 2046.2000 ;
        RECT 666.0000 2023.9600 669.0000 2024.4400 ;
        RECT 666.0000 2029.4000 669.0000 2029.8800 ;
        RECT 653.6600 2023.9600 655.2600 2024.4400 ;
        RECT 653.6600 2029.4000 655.2600 2029.8800 ;
        RECT 608.6600 2062.0400 610.2600 2062.5200 ;
        RECT 608.6600 2067.4800 610.2600 2067.9600 ;
        RECT 608.6600 2072.9200 610.2600 2073.4000 ;
        RECT 608.6600 2051.1600 610.2600 2051.6400 ;
        RECT 608.6600 2056.6000 610.2600 2057.0800 ;
        RECT 608.6600 2034.8400 610.2600 2035.3200 ;
        RECT 608.6600 2040.2800 610.2600 2040.7600 ;
        RECT 608.6600 2045.7200 610.2600 2046.2000 ;
        RECT 608.6600 2023.9600 610.2600 2024.4400 ;
        RECT 608.6600 2029.4000 610.2600 2029.8800 ;
        RECT 563.6600 2105.5600 565.2600 2106.0400 ;
        RECT 563.6600 2111.0000 565.2600 2111.4800 ;
        RECT 563.6600 2116.4400 565.2600 2116.9200 ;
        RECT 518.6600 2105.5600 520.2600 2106.0400 ;
        RECT 518.6600 2111.0000 520.2600 2111.4800 ;
        RECT 518.6600 2116.4400 520.2600 2116.9200 ;
        RECT 563.6600 2094.6800 565.2600 2095.1600 ;
        RECT 563.6600 2100.1200 565.2600 2100.6000 ;
        RECT 563.6600 2078.3600 565.2600 2078.8400 ;
        RECT 563.6600 2083.8000 565.2600 2084.2800 ;
        RECT 563.6600 2089.2400 565.2600 2089.7200 ;
        RECT 518.6600 2094.6800 520.2600 2095.1600 ;
        RECT 518.6600 2100.1200 520.2600 2100.6000 ;
        RECT 518.6600 2078.3600 520.2600 2078.8400 ;
        RECT 518.6600 2083.8000 520.2600 2084.2800 ;
        RECT 518.6600 2089.2400 520.2600 2089.7200 ;
        RECT 473.6600 2105.5600 475.2600 2106.0400 ;
        RECT 473.6600 2111.0000 475.2600 2111.4800 ;
        RECT 461.9000 2111.0000 464.9000 2111.4800 ;
        RECT 461.9000 2105.5600 464.9000 2106.0400 ;
        RECT 461.9000 2116.4400 464.9000 2116.9200 ;
        RECT 473.6600 2116.4400 475.2600 2116.9200 ;
        RECT 473.6600 2094.6800 475.2600 2095.1600 ;
        RECT 473.6600 2100.1200 475.2600 2100.6000 ;
        RECT 461.9000 2100.1200 464.9000 2100.6000 ;
        RECT 461.9000 2094.6800 464.9000 2095.1600 ;
        RECT 473.6600 2078.3600 475.2600 2078.8400 ;
        RECT 473.6600 2083.8000 475.2600 2084.2800 ;
        RECT 461.9000 2083.8000 464.9000 2084.2800 ;
        RECT 461.9000 2078.3600 464.9000 2078.8400 ;
        RECT 461.9000 2089.2400 464.9000 2089.7200 ;
        RECT 473.6600 2089.2400 475.2600 2089.7200 ;
        RECT 563.6600 2062.0400 565.2600 2062.5200 ;
        RECT 563.6600 2067.4800 565.2600 2067.9600 ;
        RECT 563.6600 2072.9200 565.2600 2073.4000 ;
        RECT 563.6600 2051.1600 565.2600 2051.6400 ;
        RECT 563.6600 2056.6000 565.2600 2057.0800 ;
        RECT 518.6600 2062.0400 520.2600 2062.5200 ;
        RECT 518.6600 2067.4800 520.2600 2067.9600 ;
        RECT 518.6600 2072.9200 520.2600 2073.4000 ;
        RECT 518.6600 2051.1600 520.2600 2051.6400 ;
        RECT 518.6600 2056.6000 520.2600 2057.0800 ;
        RECT 563.6600 2034.8400 565.2600 2035.3200 ;
        RECT 563.6600 2040.2800 565.2600 2040.7600 ;
        RECT 563.6600 2045.7200 565.2600 2046.2000 ;
        RECT 563.6600 2023.9600 565.2600 2024.4400 ;
        RECT 563.6600 2029.4000 565.2600 2029.8800 ;
        RECT 518.6600 2034.8400 520.2600 2035.3200 ;
        RECT 518.6600 2040.2800 520.2600 2040.7600 ;
        RECT 518.6600 2045.7200 520.2600 2046.2000 ;
        RECT 518.6600 2023.9600 520.2600 2024.4400 ;
        RECT 518.6600 2029.4000 520.2600 2029.8800 ;
        RECT 473.6600 2062.0400 475.2600 2062.5200 ;
        RECT 473.6600 2067.4800 475.2600 2067.9600 ;
        RECT 473.6600 2072.9200 475.2600 2073.4000 ;
        RECT 461.9000 2062.0400 464.9000 2062.5200 ;
        RECT 461.9000 2067.4800 464.9000 2067.9600 ;
        RECT 461.9000 2072.9200 464.9000 2073.4000 ;
        RECT 473.6600 2051.1600 475.2600 2051.6400 ;
        RECT 473.6600 2056.6000 475.2600 2057.0800 ;
        RECT 461.9000 2051.1600 464.9000 2051.6400 ;
        RECT 461.9000 2056.6000 464.9000 2057.0800 ;
        RECT 473.6600 2034.8400 475.2600 2035.3200 ;
        RECT 473.6600 2040.2800 475.2600 2040.7600 ;
        RECT 473.6600 2045.7200 475.2600 2046.2000 ;
        RECT 461.9000 2034.8400 464.9000 2035.3200 ;
        RECT 461.9000 2040.2800 464.9000 2040.7600 ;
        RECT 461.9000 2045.7200 464.9000 2046.2000 ;
        RECT 473.6600 2023.9600 475.2600 2024.4400 ;
        RECT 473.6600 2029.4000 475.2600 2029.8800 ;
        RECT 461.9000 2023.9600 464.9000 2024.4400 ;
        RECT 461.9000 2029.4000 464.9000 2029.8800 ;
        RECT 666.0000 2007.6400 669.0000 2008.1200 ;
        RECT 666.0000 2013.0800 669.0000 2013.5600 ;
        RECT 666.0000 2018.5200 669.0000 2019.0000 ;
        RECT 653.6600 2007.6400 655.2600 2008.1200 ;
        RECT 653.6600 2013.0800 655.2600 2013.5600 ;
        RECT 653.6600 2018.5200 655.2600 2019.0000 ;
        RECT 666.0000 1996.7600 669.0000 1997.2400 ;
        RECT 666.0000 2002.2000 669.0000 2002.6800 ;
        RECT 653.6600 1996.7600 655.2600 1997.2400 ;
        RECT 653.6600 2002.2000 655.2600 2002.6800 ;
        RECT 666.0000 1980.4400 669.0000 1980.9200 ;
        RECT 666.0000 1985.8800 669.0000 1986.3600 ;
        RECT 666.0000 1991.3200 669.0000 1991.8000 ;
        RECT 653.6600 1980.4400 655.2600 1980.9200 ;
        RECT 653.6600 1985.8800 655.2600 1986.3600 ;
        RECT 653.6600 1991.3200 655.2600 1991.8000 ;
        RECT 666.0000 1969.5600 669.0000 1970.0400 ;
        RECT 666.0000 1975.0000 669.0000 1975.4800 ;
        RECT 653.6600 1969.5600 655.2600 1970.0400 ;
        RECT 653.6600 1975.0000 655.2600 1975.4800 ;
        RECT 608.6600 2007.6400 610.2600 2008.1200 ;
        RECT 608.6600 2013.0800 610.2600 2013.5600 ;
        RECT 608.6600 2018.5200 610.2600 2019.0000 ;
        RECT 608.6600 1996.7600 610.2600 1997.2400 ;
        RECT 608.6600 2002.2000 610.2600 2002.6800 ;
        RECT 608.6600 1980.4400 610.2600 1980.9200 ;
        RECT 608.6600 1985.8800 610.2600 1986.3600 ;
        RECT 608.6600 1991.3200 610.2600 1991.8000 ;
        RECT 608.6600 1969.5600 610.2600 1970.0400 ;
        RECT 608.6600 1975.0000 610.2600 1975.4800 ;
        RECT 666.0000 1953.2400 669.0000 1953.7200 ;
        RECT 666.0000 1958.6800 669.0000 1959.1600 ;
        RECT 666.0000 1964.1200 669.0000 1964.6000 ;
        RECT 653.6600 1953.2400 655.2600 1953.7200 ;
        RECT 653.6600 1958.6800 655.2600 1959.1600 ;
        RECT 653.6600 1964.1200 655.2600 1964.6000 ;
        RECT 666.0000 1942.3600 669.0000 1942.8400 ;
        RECT 666.0000 1947.8000 669.0000 1948.2800 ;
        RECT 653.6600 1942.3600 655.2600 1942.8400 ;
        RECT 653.6600 1947.8000 655.2600 1948.2800 ;
        RECT 666.0000 1926.0400 669.0000 1926.5200 ;
        RECT 666.0000 1931.4800 669.0000 1931.9600 ;
        RECT 666.0000 1936.9200 669.0000 1937.4000 ;
        RECT 653.6600 1926.0400 655.2600 1926.5200 ;
        RECT 653.6600 1931.4800 655.2600 1931.9600 ;
        RECT 653.6600 1936.9200 655.2600 1937.4000 ;
        RECT 666.0000 1920.6000 669.0000 1921.0800 ;
        RECT 653.6600 1920.6000 655.2600 1921.0800 ;
        RECT 608.6600 1953.2400 610.2600 1953.7200 ;
        RECT 608.6600 1958.6800 610.2600 1959.1600 ;
        RECT 608.6600 1964.1200 610.2600 1964.6000 ;
        RECT 608.6600 1942.3600 610.2600 1942.8400 ;
        RECT 608.6600 1947.8000 610.2600 1948.2800 ;
        RECT 608.6600 1926.0400 610.2600 1926.5200 ;
        RECT 608.6600 1931.4800 610.2600 1931.9600 ;
        RECT 608.6600 1936.9200 610.2600 1937.4000 ;
        RECT 608.6600 1920.6000 610.2600 1921.0800 ;
        RECT 563.6600 2007.6400 565.2600 2008.1200 ;
        RECT 563.6600 2013.0800 565.2600 2013.5600 ;
        RECT 563.6600 2018.5200 565.2600 2019.0000 ;
        RECT 563.6600 1996.7600 565.2600 1997.2400 ;
        RECT 563.6600 2002.2000 565.2600 2002.6800 ;
        RECT 518.6600 2007.6400 520.2600 2008.1200 ;
        RECT 518.6600 2013.0800 520.2600 2013.5600 ;
        RECT 518.6600 2018.5200 520.2600 2019.0000 ;
        RECT 518.6600 1996.7600 520.2600 1997.2400 ;
        RECT 518.6600 2002.2000 520.2600 2002.6800 ;
        RECT 563.6600 1980.4400 565.2600 1980.9200 ;
        RECT 563.6600 1985.8800 565.2600 1986.3600 ;
        RECT 563.6600 1991.3200 565.2600 1991.8000 ;
        RECT 563.6600 1969.5600 565.2600 1970.0400 ;
        RECT 563.6600 1975.0000 565.2600 1975.4800 ;
        RECT 518.6600 1980.4400 520.2600 1980.9200 ;
        RECT 518.6600 1985.8800 520.2600 1986.3600 ;
        RECT 518.6600 1991.3200 520.2600 1991.8000 ;
        RECT 518.6600 1969.5600 520.2600 1970.0400 ;
        RECT 518.6600 1975.0000 520.2600 1975.4800 ;
        RECT 473.6600 2007.6400 475.2600 2008.1200 ;
        RECT 473.6600 2013.0800 475.2600 2013.5600 ;
        RECT 473.6600 2018.5200 475.2600 2019.0000 ;
        RECT 461.9000 2007.6400 464.9000 2008.1200 ;
        RECT 461.9000 2013.0800 464.9000 2013.5600 ;
        RECT 461.9000 2018.5200 464.9000 2019.0000 ;
        RECT 473.6600 1996.7600 475.2600 1997.2400 ;
        RECT 473.6600 2002.2000 475.2600 2002.6800 ;
        RECT 461.9000 1996.7600 464.9000 1997.2400 ;
        RECT 461.9000 2002.2000 464.9000 2002.6800 ;
        RECT 473.6600 1980.4400 475.2600 1980.9200 ;
        RECT 473.6600 1985.8800 475.2600 1986.3600 ;
        RECT 473.6600 1991.3200 475.2600 1991.8000 ;
        RECT 461.9000 1980.4400 464.9000 1980.9200 ;
        RECT 461.9000 1985.8800 464.9000 1986.3600 ;
        RECT 461.9000 1991.3200 464.9000 1991.8000 ;
        RECT 473.6600 1969.5600 475.2600 1970.0400 ;
        RECT 473.6600 1975.0000 475.2600 1975.4800 ;
        RECT 461.9000 1969.5600 464.9000 1970.0400 ;
        RECT 461.9000 1975.0000 464.9000 1975.4800 ;
        RECT 563.6600 1953.2400 565.2600 1953.7200 ;
        RECT 563.6600 1958.6800 565.2600 1959.1600 ;
        RECT 563.6600 1964.1200 565.2600 1964.6000 ;
        RECT 563.6600 1942.3600 565.2600 1942.8400 ;
        RECT 563.6600 1947.8000 565.2600 1948.2800 ;
        RECT 518.6600 1953.2400 520.2600 1953.7200 ;
        RECT 518.6600 1958.6800 520.2600 1959.1600 ;
        RECT 518.6600 1964.1200 520.2600 1964.6000 ;
        RECT 518.6600 1942.3600 520.2600 1942.8400 ;
        RECT 518.6600 1947.8000 520.2600 1948.2800 ;
        RECT 563.6600 1926.0400 565.2600 1926.5200 ;
        RECT 563.6600 1931.4800 565.2600 1931.9600 ;
        RECT 563.6600 1936.9200 565.2600 1937.4000 ;
        RECT 563.6600 1920.6000 565.2600 1921.0800 ;
        RECT 518.6600 1926.0400 520.2600 1926.5200 ;
        RECT 518.6600 1931.4800 520.2600 1931.9600 ;
        RECT 518.6600 1936.9200 520.2600 1937.4000 ;
        RECT 518.6600 1920.6000 520.2600 1921.0800 ;
        RECT 473.6600 1953.2400 475.2600 1953.7200 ;
        RECT 473.6600 1958.6800 475.2600 1959.1600 ;
        RECT 473.6600 1964.1200 475.2600 1964.6000 ;
        RECT 461.9000 1953.2400 464.9000 1953.7200 ;
        RECT 461.9000 1958.6800 464.9000 1959.1600 ;
        RECT 461.9000 1964.1200 464.9000 1964.6000 ;
        RECT 473.6600 1942.3600 475.2600 1942.8400 ;
        RECT 473.6600 1947.8000 475.2600 1948.2800 ;
        RECT 461.9000 1942.3600 464.9000 1942.8400 ;
        RECT 461.9000 1947.8000 464.9000 1948.2800 ;
        RECT 473.6600 1926.0400 475.2600 1926.5200 ;
        RECT 473.6600 1931.4800 475.2600 1931.9600 ;
        RECT 473.6600 1936.9200 475.2600 1937.4000 ;
        RECT 461.9000 1926.0400 464.9000 1926.5200 ;
        RECT 461.9000 1931.4800 464.9000 1931.9600 ;
        RECT 461.9000 1936.9200 464.9000 1937.4000 ;
        RECT 461.9000 1920.6000 464.9000 1921.0800 ;
        RECT 473.6600 1920.6000 475.2600 1921.0800 ;
        RECT 461.9000 2125.5100 669.0000 2128.5100 ;
        RECT 461.9000 1912.4100 669.0000 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 1682.7700 655.2600 1898.8700 ;
        RECT 608.6600 1682.7700 610.2600 1898.8700 ;
        RECT 563.6600 1682.7700 565.2600 1898.8700 ;
        RECT 518.6600 1682.7700 520.2600 1898.8700 ;
        RECT 473.6600 1682.7700 475.2600 1898.8700 ;
        RECT 666.0000 1682.7700 669.0000 1898.8700 ;
        RECT 461.9000 1682.7700 464.9000 1898.8700 ;
      LAYER met3 ;
        RECT 666.0000 1875.9200 669.0000 1876.4000 ;
        RECT 666.0000 1881.3600 669.0000 1881.8400 ;
        RECT 653.6600 1875.9200 655.2600 1876.4000 ;
        RECT 653.6600 1881.3600 655.2600 1881.8400 ;
        RECT 666.0000 1886.8000 669.0000 1887.2800 ;
        RECT 653.6600 1886.8000 655.2600 1887.2800 ;
        RECT 666.0000 1865.0400 669.0000 1865.5200 ;
        RECT 666.0000 1870.4800 669.0000 1870.9600 ;
        RECT 653.6600 1865.0400 655.2600 1865.5200 ;
        RECT 653.6600 1870.4800 655.2600 1870.9600 ;
        RECT 666.0000 1848.7200 669.0000 1849.2000 ;
        RECT 666.0000 1854.1600 669.0000 1854.6400 ;
        RECT 653.6600 1848.7200 655.2600 1849.2000 ;
        RECT 653.6600 1854.1600 655.2600 1854.6400 ;
        RECT 666.0000 1859.6000 669.0000 1860.0800 ;
        RECT 653.6600 1859.6000 655.2600 1860.0800 ;
        RECT 608.6600 1875.9200 610.2600 1876.4000 ;
        RECT 608.6600 1881.3600 610.2600 1881.8400 ;
        RECT 608.6600 1886.8000 610.2600 1887.2800 ;
        RECT 608.6600 1865.0400 610.2600 1865.5200 ;
        RECT 608.6600 1870.4800 610.2600 1870.9600 ;
        RECT 608.6600 1848.7200 610.2600 1849.2000 ;
        RECT 608.6600 1854.1600 610.2600 1854.6400 ;
        RECT 608.6600 1859.6000 610.2600 1860.0800 ;
        RECT 666.0000 1832.4000 669.0000 1832.8800 ;
        RECT 666.0000 1837.8400 669.0000 1838.3200 ;
        RECT 666.0000 1843.2800 669.0000 1843.7600 ;
        RECT 653.6600 1832.4000 655.2600 1832.8800 ;
        RECT 653.6600 1837.8400 655.2600 1838.3200 ;
        RECT 653.6600 1843.2800 655.2600 1843.7600 ;
        RECT 666.0000 1821.5200 669.0000 1822.0000 ;
        RECT 666.0000 1826.9600 669.0000 1827.4400 ;
        RECT 653.6600 1821.5200 655.2600 1822.0000 ;
        RECT 653.6600 1826.9600 655.2600 1827.4400 ;
        RECT 666.0000 1805.2000 669.0000 1805.6800 ;
        RECT 666.0000 1810.6400 669.0000 1811.1200 ;
        RECT 666.0000 1816.0800 669.0000 1816.5600 ;
        RECT 653.6600 1805.2000 655.2600 1805.6800 ;
        RECT 653.6600 1810.6400 655.2600 1811.1200 ;
        RECT 653.6600 1816.0800 655.2600 1816.5600 ;
        RECT 666.0000 1794.3200 669.0000 1794.8000 ;
        RECT 666.0000 1799.7600 669.0000 1800.2400 ;
        RECT 653.6600 1794.3200 655.2600 1794.8000 ;
        RECT 653.6600 1799.7600 655.2600 1800.2400 ;
        RECT 608.6600 1832.4000 610.2600 1832.8800 ;
        RECT 608.6600 1837.8400 610.2600 1838.3200 ;
        RECT 608.6600 1843.2800 610.2600 1843.7600 ;
        RECT 608.6600 1821.5200 610.2600 1822.0000 ;
        RECT 608.6600 1826.9600 610.2600 1827.4400 ;
        RECT 608.6600 1805.2000 610.2600 1805.6800 ;
        RECT 608.6600 1810.6400 610.2600 1811.1200 ;
        RECT 608.6600 1816.0800 610.2600 1816.5600 ;
        RECT 608.6600 1794.3200 610.2600 1794.8000 ;
        RECT 608.6600 1799.7600 610.2600 1800.2400 ;
        RECT 563.6600 1875.9200 565.2600 1876.4000 ;
        RECT 563.6600 1881.3600 565.2600 1881.8400 ;
        RECT 563.6600 1886.8000 565.2600 1887.2800 ;
        RECT 518.6600 1875.9200 520.2600 1876.4000 ;
        RECT 518.6600 1881.3600 520.2600 1881.8400 ;
        RECT 518.6600 1886.8000 520.2600 1887.2800 ;
        RECT 563.6600 1865.0400 565.2600 1865.5200 ;
        RECT 563.6600 1870.4800 565.2600 1870.9600 ;
        RECT 563.6600 1848.7200 565.2600 1849.2000 ;
        RECT 563.6600 1854.1600 565.2600 1854.6400 ;
        RECT 563.6600 1859.6000 565.2600 1860.0800 ;
        RECT 518.6600 1865.0400 520.2600 1865.5200 ;
        RECT 518.6600 1870.4800 520.2600 1870.9600 ;
        RECT 518.6600 1848.7200 520.2600 1849.2000 ;
        RECT 518.6600 1854.1600 520.2600 1854.6400 ;
        RECT 518.6600 1859.6000 520.2600 1860.0800 ;
        RECT 473.6600 1875.9200 475.2600 1876.4000 ;
        RECT 473.6600 1881.3600 475.2600 1881.8400 ;
        RECT 461.9000 1881.3600 464.9000 1881.8400 ;
        RECT 461.9000 1875.9200 464.9000 1876.4000 ;
        RECT 461.9000 1886.8000 464.9000 1887.2800 ;
        RECT 473.6600 1886.8000 475.2600 1887.2800 ;
        RECT 473.6600 1865.0400 475.2600 1865.5200 ;
        RECT 473.6600 1870.4800 475.2600 1870.9600 ;
        RECT 461.9000 1870.4800 464.9000 1870.9600 ;
        RECT 461.9000 1865.0400 464.9000 1865.5200 ;
        RECT 473.6600 1848.7200 475.2600 1849.2000 ;
        RECT 473.6600 1854.1600 475.2600 1854.6400 ;
        RECT 461.9000 1854.1600 464.9000 1854.6400 ;
        RECT 461.9000 1848.7200 464.9000 1849.2000 ;
        RECT 461.9000 1859.6000 464.9000 1860.0800 ;
        RECT 473.6600 1859.6000 475.2600 1860.0800 ;
        RECT 563.6600 1832.4000 565.2600 1832.8800 ;
        RECT 563.6600 1837.8400 565.2600 1838.3200 ;
        RECT 563.6600 1843.2800 565.2600 1843.7600 ;
        RECT 563.6600 1821.5200 565.2600 1822.0000 ;
        RECT 563.6600 1826.9600 565.2600 1827.4400 ;
        RECT 518.6600 1832.4000 520.2600 1832.8800 ;
        RECT 518.6600 1837.8400 520.2600 1838.3200 ;
        RECT 518.6600 1843.2800 520.2600 1843.7600 ;
        RECT 518.6600 1821.5200 520.2600 1822.0000 ;
        RECT 518.6600 1826.9600 520.2600 1827.4400 ;
        RECT 563.6600 1805.2000 565.2600 1805.6800 ;
        RECT 563.6600 1810.6400 565.2600 1811.1200 ;
        RECT 563.6600 1816.0800 565.2600 1816.5600 ;
        RECT 563.6600 1794.3200 565.2600 1794.8000 ;
        RECT 563.6600 1799.7600 565.2600 1800.2400 ;
        RECT 518.6600 1805.2000 520.2600 1805.6800 ;
        RECT 518.6600 1810.6400 520.2600 1811.1200 ;
        RECT 518.6600 1816.0800 520.2600 1816.5600 ;
        RECT 518.6600 1794.3200 520.2600 1794.8000 ;
        RECT 518.6600 1799.7600 520.2600 1800.2400 ;
        RECT 473.6600 1832.4000 475.2600 1832.8800 ;
        RECT 473.6600 1837.8400 475.2600 1838.3200 ;
        RECT 473.6600 1843.2800 475.2600 1843.7600 ;
        RECT 461.9000 1832.4000 464.9000 1832.8800 ;
        RECT 461.9000 1837.8400 464.9000 1838.3200 ;
        RECT 461.9000 1843.2800 464.9000 1843.7600 ;
        RECT 473.6600 1821.5200 475.2600 1822.0000 ;
        RECT 473.6600 1826.9600 475.2600 1827.4400 ;
        RECT 461.9000 1821.5200 464.9000 1822.0000 ;
        RECT 461.9000 1826.9600 464.9000 1827.4400 ;
        RECT 473.6600 1805.2000 475.2600 1805.6800 ;
        RECT 473.6600 1810.6400 475.2600 1811.1200 ;
        RECT 473.6600 1816.0800 475.2600 1816.5600 ;
        RECT 461.9000 1805.2000 464.9000 1805.6800 ;
        RECT 461.9000 1810.6400 464.9000 1811.1200 ;
        RECT 461.9000 1816.0800 464.9000 1816.5600 ;
        RECT 473.6600 1794.3200 475.2600 1794.8000 ;
        RECT 473.6600 1799.7600 475.2600 1800.2400 ;
        RECT 461.9000 1794.3200 464.9000 1794.8000 ;
        RECT 461.9000 1799.7600 464.9000 1800.2400 ;
        RECT 666.0000 1778.0000 669.0000 1778.4800 ;
        RECT 666.0000 1783.4400 669.0000 1783.9200 ;
        RECT 666.0000 1788.8800 669.0000 1789.3600 ;
        RECT 653.6600 1778.0000 655.2600 1778.4800 ;
        RECT 653.6600 1783.4400 655.2600 1783.9200 ;
        RECT 653.6600 1788.8800 655.2600 1789.3600 ;
        RECT 666.0000 1767.1200 669.0000 1767.6000 ;
        RECT 666.0000 1772.5600 669.0000 1773.0400 ;
        RECT 653.6600 1767.1200 655.2600 1767.6000 ;
        RECT 653.6600 1772.5600 655.2600 1773.0400 ;
        RECT 666.0000 1750.8000 669.0000 1751.2800 ;
        RECT 666.0000 1756.2400 669.0000 1756.7200 ;
        RECT 666.0000 1761.6800 669.0000 1762.1600 ;
        RECT 653.6600 1750.8000 655.2600 1751.2800 ;
        RECT 653.6600 1756.2400 655.2600 1756.7200 ;
        RECT 653.6600 1761.6800 655.2600 1762.1600 ;
        RECT 666.0000 1739.9200 669.0000 1740.4000 ;
        RECT 666.0000 1745.3600 669.0000 1745.8400 ;
        RECT 653.6600 1739.9200 655.2600 1740.4000 ;
        RECT 653.6600 1745.3600 655.2600 1745.8400 ;
        RECT 608.6600 1778.0000 610.2600 1778.4800 ;
        RECT 608.6600 1783.4400 610.2600 1783.9200 ;
        RECT 608.6600 1788.8800 610.2600 1789.3600 ;
        RECT 608.6600 1767.1200 610.2600 1767.6000 ;
        RECT 608.6600 1772.5600 610.2600 1773.0400 ;
        RECT 608.6600 1750.8000 610.2600 1751.2800 ;
        RECT 608.6600 1756.2400 610.2600 1756.7200 ;
        RECT 608.6600 1761.6800 610.2600 1762.1600 ;
        RECT 608.6600 1739.9200 610.2600 1740.4000 ;
        RECT 608.6600 1745.3600 610.2600 1745.8400 ;
        RECT 666.0000 1723.6000 669.0000 1724.0800 ;
        RECT 666.0000 1729.0400 669.0000 1729.5200 ;
        RECT 666.0000 1734.4800 669.0000 1734.9600 ;
        RECT 653.6600 1723.6000 655.2600 1724.0800 ;
        RECT 653.6600 1729.0400 655.2600 1729.5200 ;
        RECT 653.6600 1734.4800 655.2600 1734.9600 ;
        RECT 666.0000 1712.7200 669.0000 1713.2000 ;
        RECT 666.0000 1718.1600 669.0000 1718.6400 ;
        RECT 653.6600 1712.7200 655.2600 1713.2000 ;
        RECT 653.6600 1718.1600 655.2600 1718.6400 ;
        RECT 666.0000 1696.4000 669.0000 1696.8800 ;
        RECT 666.0000 1701.8400 669.0000 1702.3200 ;
        RECT 666.0000 1707.2800 669.0000 1707.7600 ;
        RECT 653.6600 1696.4000 655.2600 1696.8800 ;
        RECT 653.6600 1701.8400 655.2600 1702.3200 ;
        RECT 653.6600 1707.2800 655.2600 1707.7600 ;
        RECT 666.0000 1690.9600 669.0000 1691.4400 ;
        RECT 653.6600 1690.9600 655.2600 1691.4400 ;
        RECT 608.6600 1723.6000 610.2600 1724.0800 ;
        RECT 608.6600 1729.0400 610.2600 1729.5200 ;
        RECT 608.6600 1734.4800 610.2600 1734.9600 ;
        RECT 608.6600 1712.7200 610.2600 1713.2000 ;
        RECT 608.6600 1718.1600 610.2600 1718.6400 ;
        RECT 608.6600 1696.4000 610.2600 1696.8800 ;
        RECT 608.6600 1701.8400 610.2600 1702.3200 ;
        RECT 608.6600 1707.2800 610.2600 1707.7600 ;
        RECT 608.6600 1690.9600 610.2600 1691.4400 ;
        RECT 563.6600 1778.0000 565.2600 1778.4800 ;
        RECT 563.6600 1783.4400 565.2600 1783.9200 ;
        RECT 563.6600 1788.8800 565.2600 1789.3600 ;
        RECT 563.6600 1767.1200 565.2600 1767.6000 ;
        RECT 563.6600 1772.5600 565.2600 1773.0400 ;
        RECT 518.6600 1778.0000 520.2600 1778.4800 ;
        RECT 518.6600 1783.4400 520.2600 1783.9200 ;
        RECT 518.6600 1788.8800 520.2600 1789.3600 ;
        RECT 518.6600 1767.1200 520.2600 1767.6000 ;
        RECT 518.6600 1772.5600 520.2600 1773.0400 ;
        RECT 563.6600 1750.8000 565.2600 1751.2800 ;
        RECT 563.6600 1756.2400 565.2600 1756.7200 ;
        RECT 563.6600 1761.6800 565.2600 1762.1600 ;
        RECT 563.6600 1739.9200 565.2600 1740.4000 ;
        RECT 563.6600 1745.3600 565.2600 1745.8400 ;
        RECT 518.6600 1750.8000 520.2600 1751.2800 ;
        RECT 518.6600 1756.2400 520.2600 1756.7200 ;
        RECT 518.6600 1761.6800 520.2600 1762.1600 ;
        RECT 518.6600 1739.9200 520.2600 1740.4000 ;
        RECT 518.6600 1745.3600 520.2600 1745.8400 ;
        RECT 473.6600 1778.0000 475.2600 1778.4800 ;
        RECT 473.6600 1783.4400 475.2600 1783.9200 ;
        RECT 473.6600 1788.8800 475.2600 1789.3600 ;
        RECT 461.9000 1778.0000 464.9000 1778.4800 ;
        RECT 461.9000 1783.4400 464.9000 1783.9200 ;
        RECT 461.9000 1788.8800 464.9000 1789.3600 ;
        RECT 473.6600 1767.1200 475.2600 1767.6000 ;
        RECT 473.6600 1772.5600 475.2600 1773.0400 ;
        RECT 461.9000 1767.1200 464.9000 1767.6000 ;
        RECT 461.9000 1772.5600 464.9000 1773.0400 ;
        RECT 473.6600 1750.8000 475.2600 1751.2800 ;
        RECT 473.6600 1756.2400 475.2600 1756.7200 ;
        RECT 473.6600 1761.6800 475.2600 1762.1600 ;
        RECT 461.9000 1750.8000 464.9000 1751.2800 ;
        RECT 461.9000 1756.2400 464.9000 1756.7200 ;
        RECT 461.9000 1761.6800 464.9000 1762.1600 ;
        RECT 473.6600 1739.9200 475.2600 1740.4000 ;
        RECT 473.6600 1745.3600 475.2600 1745.8400 ;
        RECT 461.9000 1739.9200 464.9000 1740.4000 ;
        RECT 461.9000 1745.3600 464.9000 1745.8400 ;
        RECT 563.6600 1723.6000 565.2600 1724.0800 ;
        RECT 563.6600 1729.0400 565.2600 1729.5200 ;
        RECT 563.6600 1734.4800 565.2600 1734.9600 ;
        RECT 563.6600 1712.7200 565.2600 1713.2000 ;
        RECT 563.6600 1718.1600 565.2600 1718.6400 ;
        RECT 518.6600 1723.6000 520.2600 1724.0800 ;
        RECT 518.6600 1729.0400 520.2600 1729.5200 ;
        RECT 518.6600 1734.4800 520.2600 1734.9600 ;
        RECT 518.6600 1712.7200 520.2600 1713.2000 ;
        RECT 518.6600 1718.1600 520.2600 1718.6400 ;
        RECT 563.6600 1696.4000 565.2600 1696.8800 ;
        RECT 563.6600 1701.8400 565.2600 1702.3200 ;
        RECT 563.6600 1707.2800 565.2600 1707.7600 ;
        RECT 563.6600 1690.9600 565.2600 1691.4400 ;
        RECT 518.6600 1696.4000 520.2600 1696.8800 ;
        RECT 518.6600 1701.8400 520.2600 1702.3200 ;
        RECT 518.6600 1707.2800 520.2600 1707.7600 ;
        RECT 518.6600 1690.9600 520.2600 1691.4400 ;
        RECT 473.6600 1723.6000 475.2600 1724.0800 ;
        RECT 473.6600 1729.0400 475.2600 1729.5200 ;
        RECT 473.6600 1734.4800 475.2600 1734.9600 ;
        RECT 461.9000 1723.6000 464.9000 1724.0800 ;
        RECT 461.9000 1729.0400 464.9000 1729.5200 ;
        RECT 461.9000 1734.4800 464.9000 1734.9600 ;
        RECT 473.6600 1712.7200 475.2600 1713.2000 ;
        RECT 473.6600 1718.1600 475.2600 1718.6400 ;
        RECT 461.9000 1712.7200 464.9000 1713.2000 ;
        RECT 461.9000 1718.1600 464.9000 1718.6400 ;
        RECT 473.6600 1696.4000 475.2600 1696.8800 ;
        RECT 473.6600 1701.8400 475.2600 1702.3200 ;
        RECT 473.6600 1707.2800 475.2600 1707.7600 ;
        RECT 461.9000 1696.4000 464.9000 1696.8800 ;
        RECT 461.9000 1701.8400 464.9000 1702.3200 ;
        RECT 461.9000 1707.2800 464.9000 1707.7600 ;
        RECT 461.9000 1690.9600 464.9000 1691.4400 ;
        RECT 473.6600 1690.9600 475.2600 1691.4400 ;
        RECT 461.9000 1895.8700 669.0000 1898.8700 ;
        RECT 461.9000 1682.7700 669.0000 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 1453.1300 655.2600 1669.2300 ;
        RECT 608.6600 1453.1300 610.2600 1669.2300 ;
        RECT 563.6600 1453.1300 565.2600 1669.2300 ;
        RECT 518.6600 1453.1300 520.2600 1669.2300 ;
        RECT 473.6600 1453.1300 475.2600 1669.2300 ;
        RECT 666.0000 1453.1300 669.0000 1669.2300 ;
        RECT 461.9000 1453.1300 464.9000 1669.2300 ;
      LAYER met3 ;
        RECT 666.0000 1646.2800 669.0000 1646.7600 ;
        RECT 666.0000 1651.7200 669.0000 1652.2000 ;
        RECT 653.6600 1646.2800 655.2600 1646.7600 ;
        RECT 653.6600 1651.7200 655.2600 1652.2000 ;
        RECT 666.0000 1657.1600 669.0000 1657.6400 ;
        RECT 653.6600 1657.1600 655.2600 1657.6400 ;
        RECT 666.0000 1635.4000 669.0000 1635.8800 ;
        RECT 666.0000 1640.8400 669.0000 1641.3200 ;
        RECT 653.6600 1635.4000 655.2600 1635.8800 ;
        RECT 653.6600 1640.8400 655.2600 1641.3200 ;
        RECT 666.0000 1619.0800 669.0000 1619.5600 ;
        RECT 666.0000 1624.5200 669.0000 1625.0000 ;
        RECT 653.6600 1619.0800 655.2600 1619.5600 ;
        RECT 653.6600 1624.5200 655.2600 1625.0000 ;
        RECT 666.0000 1629.9600 669.0000 1630.4400 ;
        RECT 653.6600 1629.9600 655.2600 1630.4400 ;
        RECT 608.6600 1646.2800 610.2600 1646.7600 ;
        RECT 608.6600 1651.7200 610.2600 1652.2000 ;
        RECT 608.6600 1657.1600 610.2600 1657.6400 ;
        RECT 608.6600 1635.4000 610.2600 1635.8800 ;
        RECT 608.6600 1640.8400 610.2600 1641.3200 ;
        RECT 608.6600 1619.0800 610.2600 1619.5600 ;
        RECT 608.6600 1624.5200 610.2600 1625.0000 ;
        RECT 608.6600 1629.9600 610.2600 1630.4400 ;
        RECT 666.0000 1602.7600 669.0000 1603.2400 ;
        RECT 666.0000 1608.2000 669.0000 1608.6800 ;
        RECT 666.0000 1613.6400 669.0000 1614.1200 ;
        RECT 653.6600 1602.7600 655.2600 1603.2400 ;
        RECT 653.6600 1608.2000 655.2600 1608.6800 ;
        RECT 653.6600 1613.6400 655.2600 1614.1200 ;
        RECT 666.0000 1591.8800 669.0000 1592.3600 ;
        RECT 666.0000 1597.3200 669.0000 1597.8000 ;
        RECT 653.6600 1591.8800 655.2600 1592.3600 ;
        RECT 653.6600 1597.3200 655.2600 1597.8000 ;
        RECT 666.0000 1575.5600 669.0000 1576.0400 ;
        RECT 666.0000 1581.0000 669.0000 1581.4800 ;
        RECT 666.0000 1586.4400 669.0000 1586.9200 ;
        RECT 653.6600 1575.5600 655.2600 1576.0400 ;
        RECT 653.6600 1581.0000 655.2600 1581.4800 ;
        RECT 653.6600 1586.4400 655.2600 1586.9200 ;
        RECT 666.0000 1564.6800 669.0000 1565.1600 ;
        RECT 666.0000 1570.1200 669.0000 1570.6000 ;
        RECT 653.6600 1564.6800 655.2600 1565.1600 ;
        RECT 653.6600 1570.1200 655.2600 1570.6000 ;
        RECT 608.6600 1602.7600 610.2600 1603.2400 ;
        RECT 608.6600 1608.2000 610.2600 1608.6800 ;
        RECT 608.6600 1613.6400 610.2600 1614.1200 ;
        RECT 608.6600 1591.8800 610.2600 1592.3600 ;
        RECT 608.6600 1597.3200 610.2600 1597.8000 ;
        RECT 608.6600 1575.5600 610.2600 1576.0400 ;
        RECT 608.6600 1581.0000 610.2600 1581.4800 ;
        RECT 608.6600 1586.4400 610.2600 1586.9200 ;
        RECT 608.6600 1564.6800 610.2600 1565.1600 ;
        RECT 608.6600 1570.1200 610.2600 1570.6000 ;
        RECT 563.6600 1646.2800 565.2600 1646.7600 ;
        RECT 563.6600 1651.7200 565.2600 1652.2000 ;
        RECT 563.6600 1657.1600 565.2600 1657.6400 ;
        RECT 518.6600 1646.2800 520.2600 1646.7600 ;
        RECT 518.6600 1651.7200 520.2600 1652.2000 ;
        RECT 518.6600 1657.1600 520.2600 1657.6400 ;
        RECT 563.6600 1635.4000 565.2600 1635.8800 ;
        RECT 563.6600 1640.8400 565.2600 1641.3200 ;
        RECT 563.6600 1619.0800 565.2600 1619.5600 ;
        RECT 563.6600 1624.5200 565.2600 1625.0000 ;
        RECT 563.6600 1629.9600 565.2600 1630.4400 ;
        RECT 518.6600 1635.4000 520.2600 1635.8800 ;
        RECT 518.6600 1640.8400 520.2600 1641.3200 ;
        RECT 518.6600 1619.0800 520.2600 1619.5600 ;
        RECT 518.6600 1624.5200 520.2600 1625.0000 ;
        RECT 518.6600 1629.9600 520.2600 1630.4400 ;
        RECT 473.6600 1646.2800 475.2600 1646.7600 ;
        RECT 473.6600 1651.7200 475.2600 1652.2000 ;
        RECT 461.9000 1651.7200 464.9000 1652.2000 ;
        RECT 461.9000 1646.2800 464.9000 1646.7600 ;
        RECT 461.9000 1657.1600 464.9000 1657.6400 ;
        RECT 473.6600 1657.1600 475.2600 1657.6400 ;
        RECT 473.6600 1635.4000 475.2600 1635.8800 ;
        RECT 473.6600 1640.8400 475.2600 1641.3200 ;
        RECT 461.9000 1640.8400 464.9000 1641.3200 ;
        RECT 461.9000 1635.4000 464.9000 1635.8800 ;
        RECT 473.6600 1619.0800 475.2600 1619.5600 ;
        RECT 473.6600 1624.5200 475.2600 1625.0000 ;
        RECT 461.9000 1624.5200 464.9000 1625.0000 ;
        RECT 461.9000 1619.0800 464.9000 1619.5600 ;
        RECT 461.9000 1629.9600 464.9000 1630.4400 ;
        RECT 473.6600 1629.9600 475.2600 1630.4400 ;
        RECT 563.6600 1602.7600 565.2600 1603.2400 ;
        RECT 563.6600 1608.2000 565.2600 1608.6800 ;
        RECT 563.6600 1613.6400 565.2600 1614.1200 ;
        RECT 563.6600 1591.8800 565.2600 1592.3600 ;
        RECT 563.6600 1597.3200 565.2600 1597.8000 ;
        RECT 518.6600 1602.7600 520.2600 1603.2400 ;
        RECT 518.6600 1608.2000 520.2600 1608.6800 ;
        RECT 518.6600 1613.6400 520.2600 1614.1200 ;
        RECT 518.6600 1591.8800 520.2600 1592.3600 ;
        RECT 518.6600 1597.3200 520.2600 1597.8000 ;
        RECT 563.6600 1575.5600 565.2600 1576.0400 ;
        RECT 563.6600 1581.0000 565.2600 1581.4800 ;
        RECT 563.6600 1586.4400 565.2600 1586.9200 ;
        RECT 563.6600 1564.6800 565.2600 1565.1600 ;
        RECT 563.6600 1570.1200 565.2600 1570.6000 ;
        RECT 518.6600 1575.5600 520.2600 1576.0400 ;
        RECT 518.6600 1581.0000 520.2600 1581.4800 ;
        RECT 518.6600 1586.4400 520.2600 1586.9200 ;
        RECT 518.6600 1564.6800 520.2600 1565.1600 ;
        RECT 518.6600 1570.1200 520.2600 1570.6000 ;
        RECT 473.6600 1602.7600 475.2600 1603.2400 ;
        RECT 473.6600 1608.2000 475.2600 1608.6800 ;
        RECT 473.6600 1613.6400 475.2600 1614.1200 ;
        RECT 461.9000 1602.7600 464.9000 1603.2400 ;
        RECT 461.9000 1608.2000 464.9000 1608.6800 ;
        RECT 461.9000 1613.6400 464.9000 1614.1200 ;
        RECT 473.6600 1591.8800 475.2600 1592.3600 ;
        RECT 473.6600 1597.3200 475.2600 1597.8000 ;
        RECT 461.9000 1591.8800 464.9000 1592.3600 ;
        RECT 461.9000 1597.3200 464.9000 1597.8000 ;
        RECT 473.6600 1575.5600 475.2600 1576.0400 ;
        RECT 473.6600 1581.0000 475.2600 1581.4800 ;
        RECT 473.6600 1586.4400 475.2600 1586.9200 ;
        RECT 461.9000 1575.5600 464.9000 1576.0400 ;
        RECT 461.9000 1581.0000 464.9000 1581.4800 ;
        RECT 461.9000 1586.4400 464.9000 1586.9200 ;
        RECT 473.6600 1564.6800 475.2600 1565.1600 ;
        RECT 473.6600 1570.1200 475.2600 1570.6000 ;
        RECT 461.9000 1564.6800 464.9000 1565.1600 ;
        RECT 461.9000 1570.1200 464.9000 1570.6000 ;
        RECT 666.0000 1548.3600 669.0000 1548.8400 ;
        RECT 666.0000 1553.8000 669.0000 1554.2800 ;
        RECT 666.0000 1559.2400 669.0000 1559.7200 ;
        RECT 653.6600 1548.3600 655.2600 1548.8400 ;
        RECT 653.6600 1553.8000 655.2600 1554.2800 ;
        RECT 653.6600 1559.2400 655.2600 1559.7200 ;
        RECT 666.0000 1537.4800 669.0000 1537.9600 ;
        RECT 666.0000 1542.9200 669.0000 1543.4000 ;
        RECT 653.6600 1537.4800 655.2600 1537.9600 ;
        RECT 653.6600 1542.9200 655.2600 1543.4000 ;
        RECT 666.0000 1521.1600 669.0000 1521.6400 ;
        RECT 666.0000 1526.6000 669.0000 1527.0800 ;
        RECT 666.0000 1532.0400 669.0000 1532.5200 ;
        RECT 653.6600 1521.1600 655.2600 1521.6400 ;
        RECT 653.6600 1526.6000 655.2600 1527.0800 ;
        RECT 653.6600 1532.0400 655.2600 1532.5200 ;
        RECT 666.0000 1510.2800 669.0000 1510.7600 ;
        RECT 666.0000 1515.7200 669.0000 1516.2000 ;
        RECT 653.6600 1510.2800 655.2600 1510.7600 ;
        RECT 653.6600 1515.7200 655.2600 1516.2000 ;
        RECT 608.6600 1548.3600 610.2600 1548.8400 ;
        RECT 608.6600 1553.8000 610.2600 1554.2800 ;
        RECT 608.6600 1559.2400 610.2600 1559.7200 ;
        RECT 608.6600 1537.4800 610.2600 1537.9600 ;
        RECT 608.6600 1542.9200 610.2600 1543.4000 ;
        RECT 608.6600 1521.1600 610.2600 1521.6400 ;
        RECT 608.6600 1526.6000 610.2600 1527.0800 ;
        RECT 608.6600 1532.0400 610.2600 1532.5200 ;
        RECT 608.6600 1510.2800 610.2600 1510.7600 ;
        RECT 608.6600 1515.7200 610.2600 1516.2000 ;
        RECT 666.0000 1493.9600 669.0000 1494.4400 ;
        RECT 666.0000 1499.4000 669.0000 1499.8800 ;
        RECT 666.0000 1504.8400 669.0000 1505.3200 ;
        RECT 653.6600 1493.9600 655.2600 1494.4400 ;
        RECT 653.6600 1499.4000 655.2600 1499.8800 ;
        RECT 653.6600 1504.8400 655.2600 1505.3200 ;
        RECT 666.0000 1483.0800 669.0000 1483.5600 ;
        RECT 666.0000 1488.5200 669.0000 1489.0000 ;
        RECT 653.6600 1483.0800 655.2600 1483.5600 ;
        RECT 653.6600 1488.5200 655.2600 1489.0000 ;
        RECT 666.0000 1466.7600 669.0000 1467.2400 ;
        RECT 666.0000 1472.2000 669.0000 1472.6800 ;
        RECT 666.0000 1477.6400 669.0000 1478.1200 ;
        RECT 653.6600 1466.7600 655.2600 1467.2400 ;
        RECT 653.6600 1472.2000 655.2600 1472.6800 ;
        RECT 653.6600 1477.6400 655.2600 1478.1200 ;
        RECT 666.0000 1461.3200 669.0000 1461.8000 ;
        RECT 653.6600 1461.3200 655.2600 1461.8000 ;
        RECT 608.6600 1493.9600 610.2600 1494.4400 ;
        RECT 608.6600 1499.4000 610.2600 1499.8800 ;
        RECT 608.6600 1504.8400 610.2600 1505.3200 ;
        RECT 608.6600 1483.0800 610.2600 1483.5600 ;
        RECT 608.6600 1488.5200 610.2600 1489.0000 ;
        RECT 608.6600 1466.7600 610.2600 1467.2400 ;
        RECT 608.6600 1472.2000 610.2600 1472.6800 ;
        RECT 608.6600 1477.6400 610.2600 1478.1200 ;
        RECT 608.6600 1461.3200 610.2600 1461.8000 ;
        RECT 563.6600 1548.3600 565.2600 1548.8400 ;
        RECT 563.6600 1553.8000 565.2600 1554.2800 ;
        RECT 563.6600 1559.2400 565.2600 1559.7200 ;
        RECT 563.6600 1537.4800 565.2600 1537.9600 ;
        RECT 563.6600 1542.9200 565.2600 1543.4000 ;
        RECT 518.6600 1548.3600 520.2600 1548.8400 ;
        RECT 518.6600 1553.8000 520.2600 1554.2800 ;
        RECT 518.6600 1559.2400 520.2600 1559.7200 ;
        RECT 518.6600 1537.4800 520.2600 1537.9600 ;
        RECT 518.6600 1542.9200 520.2600 1543.4000 ;
        RECT 563.6600 1521.1600 565.2600 1521.6400 ;
        RECT 563.6600 1526.6000 565.2600 1527.0800 ;
        RECT 563.6600 1532.0400 565.2600 1532.5200 ;
        RECT 563.6600 1510.2800 565.2600 1510.7600 ;
        RECT 563.6600 1515.7200 565.2600 1516.2000 ;
        RECT 518.6600 1521.1600 520.2600 1521.6400 ;
        RECT 518.6600 1526.6000 520.2600 1527.0800 ;
        RECT 518.6600 1532.0400 520.2600 1532.5200 ;
        RECT 518.6600 1510.2800 520.2600 1510.7600 ;
        RECT 518.6600 1515.7200 520.2600 1516.2000 ;
        RECT 473.6600 1548.3600 475.2600 1548.8400 ;
        RECT 473.6600 1553.8000 475.2600 1554.2800 ;
        RECT 473.6600 1559.2400 475.2600 1559.7200 ;
        RECT 461.9000 1548.3600 464.9000 1548.8400 ;
        RECT 461.9000 1553.8000 464.9000 1554.2800 ;
        RECT 461.9000 1559.2400 464.9000 1559.7200 ;
        RECT 473.6600 1537.4800 475.2600 1537.9600 ;
        RECT 473.6600 1542.9200 475.2600 1543.4000 ;
        RECT 461.9000 1537.4800 464.9000 1537.9600 ;
        RECT 461.9000 1542.9200 464.9000 1543.4000 ;
        RECT 473.6600 1521.1600 475.2600 1521.6400 ;
        RECT 473.6600 1526.6000 475.2600 1527.0800 ;
        RECT 473.6600 1532.0400 475.2600 1532.5200 ;
        RECT 461.9000 1521.1600 464.9000 1521.6400 ;
        RECT 461.9000 1526.6000 464.9000 1527.0800 ;
        RECT 461.9000 1532.0400 464.9000 1532.5200 ;
        RECT 473.6600 1510.2800 475.2600 1510.7600 ;
        RECT 473.6600 1515.7200 475.2600 1516.2000 ;
        RECT 461.9000 1510.2800 464.9000 1510.7600 ;
        RECT 461.9000 1515.7200 464.9000 1516.2000 ;
        RECT 563.6600 1493.9600 565.2600 1494.4400 ;
        RECT 563.6600 1499.4000 565.2600 1499.8800 ;
        RECT 563.6600 1504.8400 565.2600 1505.3200 ;
        RECT 563.6600 1483.0800 565.2600 1483.5600 ;
        RECT 563.6600 1488.5200 565.2600 1489.0000 ;
        RECT 518.6600 1493.9600 520.2600 1494.4400 ;
        RECT 518.6600 1499.4000 520.2600 1499.8800 ;
        RECT 518.6600 1504.8400 520.2600 1505.3200 ;
        RECT 518.6600 1483.0800 520.2600 1483.5600 ;
        RECT 518.6600 1488.5200 520.2600 1489.0000 ;
        RECT 563.6600 1466.7600 565.2600 1467.2400 ;
        RECT 563.6600 1472.2000 565.2600 1472.6800 ;
        RECT 563.6600 1477.6400 565.2600 1478.1200 ;
        RECT 563.6600 1461.3200 565.2600 1461.8000 ;
        RECT 518.6600 1466.7600 520.2600 1467.2400 ;
        RECT 518.6600 1472.2000 520.2600 1472.6800 ;
        RECT 518.6600 1477.6400 520.2600 1478.1200 ;
        RECT 518.6600 1461.3200 520.2600 1461.8000 ;
        RECT 473.6600 1493.9600 475.2600 1494.4400 ;
        RECT 473.6600 1499.4000 475.2600 1499.8800 ;
        RECT 473.6600 1504.8400 475.2600 1505.3200 ;
        RECT 461.9000 1493.9600 464.9000 1494.4400 ;
        RECT 461.9000 1499.4000 464.9000 1499.8800 ;
        RECT 461.9000 1504.8400 464.9000 1505.3200 ;
        RECT 473.6600 1483.0800 475.2600 1483.5600 ;
        RECT 473.6600 1488.5200 475.2600 1489.0000 ;
        RECT 461.9000 1483.0800 464.9000 1483.5600 ;
        RECT 461.9000 1488.5200 464.9000 1489.0000 ;
        RECT 473.6600 1466.7600 475.2600 1467.2400 ;
        RECT 473.6600 1472.2000 475.2600 1472.6800 ;
        RECT 473.6600 1477.6400 475.2600 1478.1200 ;
        RECT 461.9000 1466.7600 464.9000 1467.2400 ;
        RECT 461.9000 1472.2000 464.9000 1472.6800 ;
        RECT 461.9000 1477.6400 464.9000 1478.1200 ;
        RECT 461.9000 1461.3200 464.9000 1461.8000 ;
        RECT 473.6600 1461.3200 475.2600 1461.8000 ;
        RECT 461.9000 1666.2300 669.0000 1669.2300 ;
        RECT 461.9000 1453.1300 669.0000 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 1223.4900 655.2600 1439.5900 ;
        RECT 608.6600 1223.4900 610.2600 1439.5900 ;
        RECT 563.6600 1223.4900 565.2600 1439.5900 ;
        RECT 518.6600 1223.4900 520.2600 1439.5900 ;
        RECT 473.6600 1223.4900 475.2600 1439.5900 ;
        RECT 666.0000 1223.4900 669.0000 1439.5900 ;
        RECT 461.9000 1223.4900 464.9000 1439.5900 ;
      LAYER met3 ;
        RECT 666.0000 1416.6400 669.0000 1417.1200 ;
        RECT 666.0000 1422.0800 669.0000 1422.5600 ;
        RECT 653.6600 1416.6400 655.2600 1417.1200 ;
        RECT 653.6600 1422.0800 655.2600 1422.5600 ;
        RECT 666.0000 1427.5200 669.0000 1428.0000 ;
        RECT 653.6600 1427.5200 655.2600 1428.0000 ;
        RECT 666.0000 1405.7600 669.0000 1406.2400 ;
        RECT 666.0000 1411.2000 669.0000 1411.6800 ;
        RECT 653.6600 1405.7600 655.2600 1406.2400 ;
        RECT 653.6600 1411.2000 655.2600 1411.6800 ;
        RECT 666.0000 1389.4400 669.0000 1389.9200 ;
        RECT 666.0000 1394.8800 669.0000 1395.3600 ;
        RECT 653.6600 1389.4400 655.2600 1389.9200 ;
        RECT 653.6600 1394.8800 655.2600 1395.3600 ;
        RECT 666.0000 1400.3200 669.0000 1400.8000 ;
        RECT 653.6600 1400.3200 655.2600 1400.8000 ;
        RECT 608.6600 1416.6400 610.2600 1417.1200 ;
        RECT 608.6600 1422.0800 610.2600 1422.5600 ;
        RECT 608.6600 1427.5200 610.2600 1428.0000 ;
        RECT 608.6600 1405.7600 610.2600 1406.2400 ;
        RECT 608.6600 1411.2000 610.2600 1411.6800 ;
        RECT 608.6600 1389.4400 610.2600 1389.9200 ;
        RECT 608.6600 1394.8800 610.2600 1395.3600 ;
        RECT 608.6600 1400.3200 610.2600 1400.8000 ;
        RECT 666.0000 1373.1200 669.0000 1373.6000 ;
        RECT 666.0000 1378.5600 669.0000 1379.0400 ;
        RECT 666.0000 1384.0000 669.0000 1384.4800 ;
        RECT 653.6600 1373.1200 655.2600 1373.6000 ;
        RECT 653.6600 1378.5600 655.2600 1379.0400 ;
        RECT 653.6600 1384.0000 655.2600 1384.4800 ;
        RECT 666.0000 1362.2400 669.0000 1362.7200 ;
        RECT 666.0000 1367.6800 669.0000 1368.1600 ;
        RECT 653.6600 1362.2400 655.2600 1362.7200 ;
        RECT 653.6600 1367.6800 655.2600 1368.1600 ;
        RECT 666.0000 1345.9200 669.0000 1346.4000 ;
        RECT 666.0000 1351.3600 669.0000 1351.8400 ;
        RECT 666.0000 1356.8000 669.0000 1357.2800 ;
        RECT 653.6600 1345.9200 655.2600 1346.4000 ;
        RECT 653.6600 1351.3600 655.2600 1351.8400 ;
        RECT 653.6600 1356.8000 655.2600 1357.2800 ;
        RECT 666.0000 1335.0400 669.0000 1335.5200 ;
        RECT 666.0000 1340.4800 669.0000 1340.9600 ;
        RECT 653.6600 1335.0400 655.2600 1335.5200 ;
        RECT 653.6600 1340.4800 655.2600 1340.9600 ;
        RECT 608.6600 1373.1200 610.2600 1373.6000 ;
        RECT 608.6600 1378.5600 610.2600 1379.0400 ;
        RECT 608.6600 1384.0000 610.2600 1384.4800 ;
        RECT 608.6600 1362.2400 610.2600 1362.7200 ;
        RECT 608.6600 1367.6800 610.2600 1368.1600 ;
        RECT 608.6600 1345.9200 610.2600 1346.4000 ;
        RECT 608.6600 1351.3600 610.2600 1351.8400 ;
        RECT 608.6600 1356.8000 610.2600 1357.2800 ;
        RECT 608.6600 1335.0400 610.2600 1335.5200 ;
        RECT 608.6600 1340.4800 610.2600 1340.9600 ;
        RECT 563.6600 1416.6400 565.2600 1417.1200 ;
        RECT 563.6600 1422.0800 565.2600 1422.5600 ;
        RECT 563.6600 1427.5200 565.2600 1428.0000 ;
        RECT 518.6600 1416.6400 520.2600 1417.1200 ;
        RECT 518.6600 1422.0800 520.2600 1422.5600 ;
        RECT 518.6600 1427.5200 520.2600 1428.0000 ;
        RECT 563.6600 1405.7600 565.2600 1406.2400 ;
        RECT 563.6600 1411.2000 565.2600 1411.6800 ;
        RECT 563.6600 1389.4400 565.2600 1389.9200 ;
        RECT 563.6600 1394.8800 565.2600 1395.3600 ;
        RECT 563.6600 1400.3200 565.2600 1400.8000 ;
        RECT 518.6600 1405.7600 520.2600 1406.2400 ;
        RECT 518.6600 1411.2000 520.2600 1411.6800 ;
        RECT 518.6600 1389.4400 520.2600 1389.9200 ;
        RECT 518.6600 1394.8800 520.2600 1395.3600 ;
        RECT 518.6600 1400.3200 520.2600 1400.8000 ;
        RECT 473.6600 1416.6400 475.2600 1417.1200 ;
        RECT 473.6600 1422.0800 475.2600 1422.5600 ;
        RECT 461.9000 1422.0800 464.9000 1422.5600 ;
        RECT 461.9000 1416.6400 464.9000 1417.1200 ;
        RECT 461.9000 1427.5200 464.9000 1428.0000 ;
        RECT 473.6600 1427.5200 475.2600 1428.0000 ;
        RECT 473.6600 1405.7600 475.2600 1406.2400 ;
        RECT 473.6600 1411.2000 475.2600 1411.6800 ;
        RECT 461.9000 1411.2000 464.9000 1411.6800 ;
        RECT 461.9000 1405.7600 464.9000 1406.2400 ;
        RECT 473.6600 1389.4400 475.2600 1389.9200 ;
        RECT 473.6600 1394.8800 475.2600 1395.3600 ;
        RECT 461.9000 1394.8800 464.9000 1395.3600 ;
        RECT 461.9000 1389.4400 464.9000 1389.9200 ;
        RECT 461.9000 1400.3200 464.9000 1400.8000 ;
        RECT 473.6600 1400.3200 475.2600 1400.8000 ;
        RECT 563.6600 1373.1200 565.2600 1373.6000 ;
        RECT 563.6600 1378.5600 565.2600 1379.0400 ;
        RECT 563.6600 1384.0000 565.2600 1384.4800 ;
        RECT 563.6600 1362.2400 565.2600 1362.7200 ;
        RECT 563.6600 1367.6800 565.2600 1368.1600 ;
        RECT 518.6600 1373.1200 520.2600 1373.6000 ;
        RECT 518.6600 1378.5600 520.2600 1379.0400 ;
        RECT 518.6600 1384.0000 520.2600 1384.4800 ;
        RECT 518.6600 1362.2400 520.2600 1362.7200 ;
        RECT 518.6600 1367.6800 520.2600 1368.1600 ;
        RECT 563.6600 1345.9200 565.2600 1346.4000 ;
        RECT 563.6600 1351.3600 565.2600 1351.8400 ;
        RECT 563.6600 1356.8000 565.2600 1357.2800 ;
        RECT 563.6600 1335.0400 565.2600 1335.5200 ;
        RECT 563.6600 1340.4800 565.2600 1340.9600 ;
        RECT 518.6600 1345.9200 520.2600 1346.4000 ;
        RECT 518.6600 1351.3600 520.2600 1351.8400 ;
        RECT 518.6600 1356.8000 520.2600 1357.2800 ;
        RECT 518.6600 1335.0400 520.2600 1335.5200 ;
        RECT 518.6600 1340.4800 520.2600 1340.9600 ;
        RECT 473.6600 1373.1200 475.2600 1373.6000 ;
        RECT 473.6600 1378.5600 475.2600 1379.0400 ;
        RECT 473.6600 1384.0000 475.2600 1384.4800 ;
        RECT 461.9000 1373.1200 464.9000 1373.6000 ;
        RECT 461.9000 1378.5600 464.9000 1379.0400 ;
        RECT 461.9000 1384.0000 464.9000 1384.4800 ;
        RECT 473.6600 1362.2400 475.2600 1362.7200 ;
        RECT 473.6600 1367.6800 475.2600 1368.1600 ;
        RECT 461.9000 1362.2400 464.9000 1362.7200 ;
        RECT 461.9000 1367.6800 464.9000 1368.1600 ;
        RECT 473.6600 1345.9200 475.2600 1346.4000 ;
        RECT 473.6600 1351.3600 475.2600 1351.8400 ;
        RECT 473.6600 1356.8000 475.2600 1357.2800 ;
        RECT 461.9000 1345.9200 464.9000 1346.4000 ;
        RECT 461.9000 1351.3600 464.9000 1351.8400 ;
        RECT 461.9000 1356.8000 464.9000 1357.2800 ;
        RECT 473.6600 1335.0400 475.2600 1335.5200 ;
        RECT 473.6600 1340.4800 475.2600 1340.9600 ;
        RECT 461.9000 1335.0400 464.9000 1335.5200 ;
        RECT 461.9000 1340.4800 464.9000 1340.9600 ;
        RECT 666.0000 1318.7200 669.0000 1319.2000 ;
        RECT 666.0000 1324.1600 669.0000 1324.6400 ;
        RECT 666.0000 1329.6000 669.0000 1330.0800 ;
        RECT 653.6600 1318.7200 655.2600 1319.2000 ;
        RECT 653.6600 1324.1600 655.2600 1324.6400 ;
        RECT 653.6600 1329.6000 655.2600 1330.0800 ;
        RECT 666.0000 1307.8400 669.0000 1308.3200 ;
        RECT 666.0000 1313.2800 669.0000 1313.7600 ;
        RECT 653.6600 1307.8400 655.2600 1308.3200 ;
        RECT 653.6600 1313.2800 655.2600 1313.7600 ;
        RECT 666.0000 1291.5200 669.0000 1292.0000 ;
        RECT 666.0000 1296.9600 669.0000 1297.4400 ;
        RECT 666.0000 1302.4000 669.0000 1302.8800 ;
        RECT 653.6600 1291.5200 655.2600 1292.0000 ;
        RECT 653.6600 1296.9600 655.2600 1297.4400 ;
        RECT 653.6600 1302.4000 655.2600 1302.8800 ;
        RECT 666.0000 1280.6400 669.0000 1281.1200 ;
        RECT 666.0000 1286.0800 669.0000 1286.5600 ;
        RECT 653.6600 1280.6400 655.2600 1281.1200 ;
        RECT 653.6600 1286.0800 655.2600 1286.5600 ;
        RECT 608.6600 1318.7200 610.2600 1319.2000 ;
        RECT 608.6600 1324.1600 610.2600 1324.6400 ;
        RECT 608.6600 1329.6000 610.2600 1330.0800 ;
        RECT 608.6600 1307.8400 610.2600 1308.3200 ;
        RECT 608.6600 1313.2800 610.2600 1313.7600 ;
        RECT 608.6600 1291.5200 610.2600 1292.0000 ;
        RECT 608.6600 1296.9600 610.2600 1297.4400 ;
        RECT 608.6600 1302.4000 610.2600 1302.8800 ;
        RECT 608.6600 1280.6400 610.2600 1281.1200 ;
        RECT 608.6600 1286.0800 610.2600 1286.5600 ;
        RECT 666.0000 1264.3200 669.0000 1264.8000 ;
        RECT 666.0000 1269.7600 669.0000 1270.2400 ;
        RECT 666.0000 1275.2000 669.0000 1275.6800 ;
        RECT 653.6600 1264.3200 655.2600 1264.8000 ;
        RECT 653.6600 1269.7600 655.2600 1270.2400 ;
        RECT 653.6600 1275.2000 655.2600 1275.6800 ;
        RECT 666.0000 1253.4400 669.0000 1253.9200 ;
        RECT 666.0000 1258.8800 669.0000 1259.3600 ;
        RECT 653.6600 1253.4400 655.2600 1253.9200 ;
        RECT 653.6600 1258.8800 655.2600 1259.3600 ;
        RECT 666.0000 1237.1200 669.0000 1237.6000 ;
        RECT 666.0000 1242.5600 669.0000 1243.0400 ;
        RECT 666.0000 1248.0000 669.0000 1248.4800 ;
        RECT 653.6600 1237.1200 655.2600 1237.6000 ;
        RECT 653.6600 1242.5600 655.2600 1243.0400 ;
        RECT 653.6600 1248.0000 655.2600 1248.4800 ;
        RECT 666.0000 1231.6800 669.0000 1232.1600 ;
        RECT 653.6600 1231.6800 655.2600 1232.1600 ;
        RECT 608.6600 1264.3200 610.2600 1264.8000 ;
        RECT 608.6600 1269.7600 610.2600 1270.2400 ;
        RECT 608.6600 1275.2000 610.2600 1275.6800 ;
        RECT 608.6600 1253.4400 610.2600 1253.9200 ;
        RECT 608.6600 1258.8800 610.2600 1259.3600 ;
        RECT 608.6600 1237.1200 610.2600 1237.6000 ;
        RECT 608.6600 1242.5600 610.2600 1243.0400 ;
        RECT 608.6600 1248.0000 610.2600 1248.4800 ;
        RECT 608.6600 1231.6800 610.2600 1232.1600 ;
        RECT 563.6600 1318.7200 565.2600 1319.2000 ;
        RECT 563.6600 1324.1600 565.2600 1324.6400 ;
        RECT 563.6600 1329.6000 565.2600 1330.0800 ;
        RECT 563.6600 1307.8400 565.2600 1308.3200 ;
        RECT 563.6600 1313.2800 565.2600 1313.7600 ;
        RECT 518.6600 1318.7200 520.2600 1319.2000 ;
        RECT 518.6600 1324.1600 520.2600 1324.6400 ;
        RECT 518.6600 1329.6000 520.2600 1330.0800 ;
        RECT 518.6600 1307.8400 520.2600 1308.3200 ;
        RECT 518.6600 1313.2800 520.2600 1313.7600 ;
        RECT 563.6600 1291.5200 565.2600 1292.0000 ;
        RECT 563.6600 1296.9600 565.2600 1297.4400 ;
        RECT 563.6600 1302.4000 565.2600 1302.8800 ;
        RECT 563.6600 1280.6400 565.2600 1281.1200 ;
        RECT 563.6600 1286.0800 565.2600 1286.5600 ;
        RECT 518.6600 1291.5200 520.2600 1292.0000 ;
        RECT 518.6600 1296.9600 520.2600 1297.4400 ;
        RECT 518.6600 1302.4000 520.2600 1302.8800 ;
        RECT 518.6600 1280.6400 520.2600 1281.1200 ;
        RECT 518.6600 1286.0800 520.2600 1286.5600 ;
        RECT 473.6600 1318.7200 475.2600 1319.2000 ;
        RECT 473.6600 1324.1600 475.2600 1324.6400 ;
        RECT 473.6600 1329.6000 475.2600 1330.0800 ;
        RECT 461.9000 1318.7200 464.9000 1319.2000 ;
        RECT 461.9000 1324.1600 464.9000 1324.6400 ;
        RECT 461.9000 1329.6000 464.9000 1330.0800 ;
        RECT 473.6600 1307.8400 475.2600 1308.3200 ;
        RECT 473.6600 1313.2800 475.2600 1313.7600 ;
        RECT 461.9000 1307.8400 464.9000 1308.3200 ;
        RECT 461.9000 1313.2800 464.9000 1313.7600 ;
        RECT 473.6600 1291.5200 475.2600 1292.0000 ;
        RECT 473.6600 1296.9600 475.2600 1297.4400 ;
        RECT 473.6600 1302.4000 475.2600 1302.8800 ;
        RECT 461.9000 1291.5200 464.9000 1292.0000 ;
        RECT 461.9000 1296.9600 464.9000 1297.4400 ;
        RECT 461.9000 1302.4000 464.9000 1302.8800 ;
        RECT 473.6600 1280.6400 475.2600 1281.1200 ;
        RECT 473.6600 1286.0800 475.2600 1286.5600 ;
        RECT 461.9000 1280.6400 464.9000 1281.1200 ;
        RECT 461.9000 1286.0800 464.9000 1286.5600 ;
        RECT 563.6600 1264.3200 565.2600 1264.8000 ;
        RECT 563.6600 1269.7600 565.2600 1270.2400 ;
        RECT 563.6600 1275.2000 565.2600 1275.6800 ;
        RECT 563.6600 1253.4400 565.2600 1253.9200 ;
        RECT 563.6600 1258.8800 565.2600 1259.3600 ;
        RECT 518.6600 1264.3200 520.2600 1264.8000 ;
        RECT 518.6600 1269.7600 520.2600 1270.2400 ;
        RECT 518.6600 1275.2000 520.2600 1275.6800 ;
        RECT 518.6600 1253.4400 520.2600 1253.9200 ;
        RECT 518.6600 1258.8800 520.2600 1259.3600 ;
        RECT 563.6600 1237.1200 565.2600 1237.6000 ;
        RECT 563.6600 1242.5600 565.2600 1243.0400 ;
        RECT 563.6600 1248.0000 565.2600 1248.4800 ;
        RECT 563.6600 1231.6800 565.2600 1232.1600 ;
        RECT 518.6600 1237.1200 520.2600 1237.6000 ;
        RECT 518.6600 1242.5600 520.2600 1243.0400 ;
        RECT 518.6600 1248.0000 520.2600 1248.4800 ;
        RECT 518.6600 1231.6800 520.2600 1232.1600 ;
        RECT 473.6600 1264.3200 475.2600 1264.8000 ;
        RECT 473.6600 1269.7600 475.2600 1270.2400 ;
        RECT 473.6600 1275.2000 475.2600 1275.6800 ;
        RECT 461.9000 1264.3200 464.9000 1264.8000 ;
        RECT 461.9000 1269.7600 464.9000 1270.2400 ;
        RECT 461.9000 1275.2000 464.9000 1275.6800 ;
        RECT 473.6600 1253.4400 475.2600 1253.9200 ;
        RECT 473.6600 1258.8800 475.2600 1259.3600 ;
        RECT 461.9000 1253.4400 464.9000 1253.9200 ;
        RECT 461.9000 1258.8800 464.9000 1259.3600 ;
        RECT 473.6600 1237.1200 475.2600 1237.6000 ;
        RECT 473.6600 1242.5600 475.2600 1243.0400 ;
        RECT 473.6600 1248.0000 475.2600 1248.4800 ;
        RECT 461.9000 1237.1200 464.9000 1237.6000 ;
        RECT 461.9000 1242.5600 464.9000 1243.0400 ;
        RECT 461.9000 1248.0000 464.9000 1248.4800 ;
        RECT 461.9000 1231.6800 464.9000 1232.1600 ;
        RECT 473.6600 1231.6800 475.2600 1232.1600 ;
        RECT 461.9000 1436.5900 669.0000 1439.5900 ;
        RECT 461.9000 1223.4900 669.0000 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 993.8500 655.2600 1209.9500 ;
        RECT 608.6600 993.8500 610.2600 1209.9500 ;
        RECT 563.6600 993.8500 565.2600 1209.9500 ;
        RECT 518.6600 993.8500 520.2600 1209.9500 ;
        RECT 473.6600 993.8500 475.2600 1209.9500 ;
        RECT 666.0000 993.8500 669.0000 1209.9500 ;
        RECT 461.9000 993.8500 464.9000 1209.9500 ;
      LAYER met3 ;
        RECT 666.0000 1187.0000 669.0000 1187.4800 ;
        RECT 666.0000 1192.4400 669.0000 1192.9200 ;
        RECT 653.6600 1187.0000 655.2600 1187.4800 ;
        RECT 653.6600 1192.4400 655.2600 1192.9200 ;
        RECT 666.0000 1197.8800 669.0000 1198.3600 ;
        RECT 653.6600 1197.8800 655.2600 1198.3600 ;
        RECT 666.0000 1176.1200 669.0000 1176.6000 ;
        RECT 666.0000 1181.5600 669.0000 1182.0400 ;
        RECT 653.6600 1176.1200 655.2600 1176.6000 ;
        RECT 653.6600 1181.5600 655.2600 1182.0400 ;
        RECT 666.0000 1159.8000 669.0000 1160.2800 ;
        RECT 666.0000 1165.2400 669.0000 1165.7200 ;
        RECT 653.6600 1159.8000 655.2600 1160.2800 ;
        RECT 653.6600 1165.2400 655.2600 1165.7200 ;
        RECT 666.0000 1170.6800 669.0000 1171.1600 ;
        RECT 653.6600 1170.6800 655.2600 1171.1600 ;
        RECT 608.6600 1187.0000 610.2600 1187.4800 ;
        RECT 608.6600 1192.4400 610.2600 1192.9200 ;
        RECT 608.6600 1197.8800 610.2600 1198.3600 ;
        RECT 608.6600 1176.1200 610.2600 1176.6000 ;
        RECT 608.6600 1181.5600 610.2600 1182.0400 ;
        RECT 608.6600 1159.8000 610.2600 1160.2800 ;
        RECT 608.6600 1165.2400 610.2600 1165.7200 ;
        RECT 608.6600 1170.6800 610.2600 1171.1600 ;
        RECT 666.0000 1143.4800 669.0000 1143.9600 ;
        RECT 666.0000 1148.9200 669.0000 1149.4000 ;
        RECT 666.0000 1154.3600 669.0000 1154.8400 ;
        RECT 653.6600 1143.4800 655.2600 1143.9600 ;
        RECT 653.6600 1148.9200 655.2600 1149.4000 ;
        RECT 653.6600 1154.3600 655.2600 1154.8400 ;
        RECT 666.0000 1132.6000 669.0000 1133.0800 ;
        RECT 666.0000 1138.0400 669.0000 1138.5200 ;
        RECT 653.6600 1132.6000 655.2600 1133.0800 ;
        RECT 653.6600 1138.0400 655.2600 1138.5200 ;
        RECT 666.0000 1116.2800 669.0000 1116.7600 ;
        RECT 666.0000 1121.7200 669.0000 1122.2000 ;
        RECT 666.0000 1127.1600 669.0000 1127.6400 ;
        RECT 653.6600 1116.2800 655.2600 1116.7600 ;
        RECT 653.6600 1121.7200 655.2600 1122.2000 ;
        RECT 653.6600 1127.1600 655.2600 1127.6400 ;
        RECT 666.0000 1105.4000 669.0000 1105.8800 ;
        RECT 666.0000 1110.8400 669.0000 1111.3200 ;
        RECT 653.6600 1105.4000 655.2600 1105.8800 ;
        RECT 653.6600 1110.8400 655.2600 1111.3200 ;
        RECT 608.6600 1143.4800 610.2600 1143.9600 ;
        RECT 608.6600 1148.9200 610.2600 1149.4000 ;
        RECT 608.6600 1154.3600 610.2600 1154.8400 ;
        RECT 608.6600 1132.6000 610.2600 1133.0800 ;
        RECT 608.6600 1138.0400 610.2600 1138.5200 ;
        RECT 608.6600 1116.2800 610.2600 1116.7600 ;
        RECT 608.6600 1121.7200 610.2600 1122.2000 ;
        RECT 608.6600 1127.1600 610.2600 1127.6400 ;
        RECT 608.6600 1105.4000 610.2600 1105.8800 ;
        RECT 608.6600 1110.8400 610.2600 1111.3200 ;
        RECT 563.6600 1187.0000 565.2600 1187.4800 ;
        RECT 563.6600 1192.4400 565.2600 1192.9200 ;
        RECT 563.6600 1197.8800 565.2600 1198.3600 ;
        RECT 518.6600 1187.0000 520.2600 1187.4800 ;
        RECT 518.6600 1192.4400 520.2600 1192.9200 ;
        RECT 518.6600 1197.8800 520.2600 1198.3600 ;
        RECT 563.6600 1176.1200 565.2600 1176.6000 ;
        RECT 563.6600 1181.5600 565.2600 1182.0400 ;
        RECT 563.6600 1159.8000 565.2600 1160.2800 ;
        RECT 563.6600 1165.2400 565.2600 1165.7200 ;
        RECT 563.6600 1170.6800 565.2600 1171.1600 ;
        RECT 518.6600 1176.1200 520.2600 1176.6000 ;
        RECT 518.6600 1181.5600 520.2600 1182.0400 ;
        RECT 518.6600 1159.8000 520.2600 1160.2800 ;
        RECT 518.6600 1165.2400 520.2600 1165.7200 ;
        RECT 518.6600 1170.6800 520.2600 1171.1600 ;
        RECT 473.6600 1187.0000 475.2600 1187.4800 ;
        RECT 473.6600 1192.4400 475.2600 1192.9200 ;
        RECT 461.9000 1192.4400 464.9000 1192.9200 ;
        RECT 461.9000 1187.0000 464.9000 1187.4800 ;
        RECT 461.9000 1197.8800 464.9000 1198.3600 ;
        RECT 473.6600 1197.8800 475.2600 1198.3600 ;
        RECT 473.6600 1176.1200 475.2600 1176.6000 ;
        RECT 473.6600 1181.5600 475.2600 1182.0400 ;
        RECT 461.9000 1181.5600 464.9000 1182.0400 ;
        RECT 461.9000 1176.1200 464.9000 1176.6000 ;
        RECT 473.6600 1159.8000 475.2600 1160.2800 ;
        RECT 473.6600 1165.2400 475.2600 1165.7200 ;
        RECT 461.9000 1165.2400 464.9000 1165.7200 ;
        RECT 461.9000 1159.8000 464.9000 1160.2800 ;
        RECT 461.9000 1170.6800 464.9000 1171.1600 ;
        RECT 473.6600 1170.6800 475.2600 1171.1600 ;
        RECT 563.6600 1143.4800 565.2600 1143.9600 ;
        RECT 563.6600 1148.9200 565.2600 1149.4000 ;
        RECT 563.6600 1154.3600 565.2600 1154.8400 ;
        RECT 563.6600 1132.6000 565.2600 1133.0800 ;
        RECT 563.6600 1138.0400 565.2600 1138.5200 ;
        RECT 518.6600 1143.4800 520.2600 1143.9600 ;
        RECT 518.6600 1148.9200 520.2600 1149.4000 ;
        RECT 518.6600 1154.3600 520.2600 1154.8400 ;
        RECT 518.6600 1132.6000 520.2600 1133.0800 ;
        RECT 518.6600 1138.0400 520.2600 1138.5200 ;
        RECT 563.6600 1116.2800 565.2600 1116.7600 ;
        RECT 563.6600 1121.7200 565.2600 1122.2000 ;
        RECT 563.6600 1127.1600 565.2600 1127.6400 ;
        RECT 563.6600 1105.4000 565.2600 1105.8800 ;
        RECT 563.6600 1110.8400 565.2600 1111.3200 ;
        RECT 518.6600 1116.2800 520.2600 1116.7600 ;
        RECT 518.6600 1121.7200 520.2600 1122.2000 ;
        RECT 518.6600 1127.1600 520.2600 1127.6400 ;
        RECT 518.6600 1105.4000 520.2600 1105.8800 ;
        RECT 518.6600 1110.8400 520.2600 1111.3200 ;
        RECT 473.6600 1143.4800 475.2600 1143.9600 ;
        RECT 473.6600 1148.9200 475.2600 1149.4000 ;
        RECT 473.6600 1154.3600 475.2600 1154.8400 ;
        RECT 461.9000 1143.4800 464.9000 1143.9600 ;
        RECT 461.9000 1148.9200 464.9000 1149.4000 ;
        RECT 461.9000 1154.3600 464.9000 1154.8400 ;
        RECT 473.6600 1132.6000 475.2600 1133.0800 ;
        RECT 473.6600 1138.0400 475.2600 1138.5200 ;
        RECT 461.9000 1132.6000 464.9000 1133.0800 ;
        RECT 461.9000 1138.0400 464.9000 1138.5200 ;
        RECT 473.6600 1116.2800 475.2600 1116.7600 ;
        RECT 473.6600 1121.7200 475.2600 1122.2000 ;
        RECT 473.6600 1127.1600 475.2600 1127.6400 ;
        RECT 461.9000 1116.2800 464.9000 1116.7600 ;
        RECT 461.9000 1121.7200 464.9000 1122.2000 ;
        RECT 461.9000 1127.1600 464.9000 1127.6400 ;
        RECT 473.6600 1105.4000 475.2600 1105.8800 ;
        RECT 473.6600 1110.8400 475.2600 1111.3200 ;
        RECT 461.9000 1105.4000 464.9000 1105.8800 ;
        RECT 461.9000 1110.8400 464.9000 1111.3200 ;
        RECT 666.0000 1089.0800 669.0000 1089.5600 ;
        RECT 666.0000 1094.5200 669.0000 1095.0000 ;
        RECT 666.0000 1099.9600 669.0000 1100.4400 ;
        RECT 653.6600 1089.0800 655.2600 1089.5600 ;
        RECT 653.6600 1094.5200 655.2600 1095.0000 ;
        RECT 653.6600 1099.9600 655.2600 1100.4400 ;
        RECT 666.0000 1078.2000 669.0000 1078.6800 ;
        RECT 666.0000 1083.6400 669.0000 1084.1200 ;
        RECT 653.6600 1078.2000 655.2600 1078.6800 ;
        RECT 653.6600 1083.6400 655.2600 1084.1200 ;
        RECT 666.0000 1061.8800 669.0000 1062.3600 ;
        RECT 666.0000 1067.3200 669.0000 1067.8000 ;
        RECT 666.0000 1072.7600 669.0000 1073.2400 ;
        RECT 653.6600 1061.8800 655.2600 1062.3600 ;
        RECT 653.6600 1067.3200 655.2600 1067.8000 ;
        RECT 653.6600 1072.7600 655.2600 1073.2400 ;
        RECT 666.0000 1051.0000 669.0000 1051.4800 ;
        RECT 666.0000 1056.4400 669.0000 1056.9200 ;
        RECT 653.6600 1051.0000 655.2600 1051.4800 ;
        RECT 653.6600 1056.4400 655.2600 1056.9200 ;
        RECT 608.6600 1089.0800 610.2600 1089.5600 ;
        RECT 608.6600 1094.5200 610.2600 1095.0000 ;
        RECT 608.6600 1099.9600 610.2600 1100.4400 ;
        RECT 608.6600 1078.2000 610.2600 1078.6800 ;
        RECT 608.6600 1083.6400 610.2600 1084.1200 ;
        RECT 608.6600 1061.8800 610.2600 1062.3600 ;
        RECT 608.6600 1067.3200 610.2600 1067.8000 ;
        RECT 608.6600 1072.7600 610.2600 1073.2400 ;
        RECT 608.6600 1051.0000 610.2600 1051.4800 ;
        RECT 608.6600 1056.4400 610.2600 1056.9200 ;
        RECT 666.0000 1034.6800 669.0000 1035.1600 ;
        RECT 666.0000 1040.1200 669.0000 1040.6000 ;
        RECT 666.0000 1045.5600 669.0000 1046.0400 ;
        RECT 653.6600 1034.6800 655.2600 1035.1600 ;
        RECT 653.6600 1040.1200 655.2600 1040.6000 ;
        RECT 653.6600 1045.5600 655.2600 1046.0400 ;
        RECT 666.0000 1023.8000 669.0000 1024.2800 ;
        RECT 666.0000 1029.2400 669.0000 1029.7200 ;
        RECT 653.6600 1023.8000 655.2600 1024.2800 ;
        RECT 653.6600 1029.2400 655.2600 1029.7200 ;
        RECT 666.0000 1007.4800 669.0000 1007.9600 ;
        RECT 666.0000 1012.9200 669.0000 1013.4000 ;
        RECT 666.0000 1018.3600 669.0000 1018.8400 ;
        RECT 653.6600 1007.4800 655.2600 1007.9600 ;
        RECT 653.6600 1012.9200 655.2600 1013.4000 ;
        RECT 653.6600 1018.3600 655.2600 1018.8400 ;
        RECT 666.0000 1002.0400 669.0000 1002.5200 ;
        RECT 653.6600 1002.0400 655.2600 1002.5200 ;
        RECT 608.6600 1034.6800 610.2600 1035.1600 ;
        RECT 608.6600 1040.1200 610.2600 1040.6000 ;
        RECT 608.6600 1045.5600 610.2600 1046.0400 ;
        RECT 608.6600 1023.8000 610.2600 1024.2800 ;
        RECT 608.6600 1029.2400 610.2600 1029.7200 ;
        RECT 608.6600 1007.4800 610.2600 1007.9600 ;
        RECT 608.6600 1012.9200 610.2600 1013.4000 ;
        RECT 608.6600 1018.3600 610.2600 1018.8400 ;
        RECT 608.6600 1002.0400 610.2600 1002.5200 ;
        RECT 563.6600 1089.0800 565.2600 1089.5600 ;
        RECT 563.6600 1094.5200 565.2600 1095.0000 ;
        RECT 563.6600 1099.9600 565.2600 1100.4400 ;
        RECT 563.6600 1078.2000 565.2600 1078.6800 ;
        RECT 563.6600 1083.6400 565.2600 1084.1200 ;
        RECT 518.6600 1089.0800 520.2600 1089.5600 ;
        RECT 518.6600 1094.5200 520.2600 1095.0000 ;
        RECT 518.6600 1099.9600 520.2600 1100.4400 ;
        RECT 518.6600 1078.2000 520.2600 1078.6800 ;
        RECT 518.6600 1083.6400 520.2600 1084.1200 ;
        RECT 563.6600 1061.8800 565.2600 1062.3600 ;
        RECT 563.6600 1067.3200 565.2600 1067.8000 ;
        RECT 563.6600 1072.7600 565.2600 1073.2400 ;
        RECT 563.6600 1051.0000 565.2600 1051.4800 ;
        RECT 563.6600 1056.4400 565.2600 1056.9200 ;
        RECT 518.6600 1061.8800 520.2600 1062.3600 ;
        RECT 518.6600 1067.3200 520.2600 1067.8000 ;
        RECT 518.6600 1072.7600 520.2600 1073.2400 ;
        RECT 518.6600 1051.0000 520.2600 1051.4800 ;
        RECT 518.6600 1056.4400 520.2600 1056.9200 ;
        RECT 473.6600 1089.0800 475.2600 1089.5600 ;
        RECT 473.6600 1094.5200 475.2600 1095.0000 ;
        RECT 473.6600 1099.9600 475.2600 1100.4400 ;
        RECT 461.9000 1089.0800 464.9000 1089.5600 ;
        RECT 461.9000 1094.5200 464.9000 1095.0000 ;
        RECT 461.9000 1099.9600 464.9000 1100.4400 ;
        RECT 473.6600 1078.2000 475.2600 1078.6800 ;
        RECT 473.6600 1083.6400 475.2600 1084.1200 ;
        RECT 461.9000 1078.2000 464.9000 1078.6800 ;
        RECT 461.9000 1083.6400 464.9000 1084.1200 ;
        RECT 473.6600 1061.8800 475.2600 1062.3600 ;
        RECT 473.6600 1067.3200 475.2600 1067.8000 ;
        RECT 473.6600 1072.7600 475.2600 1073.2400 ;
        RECT 461.9000 1061.8800 464.9000 1062.3600 ;
        RECT 461.9000 1067.3200 464.9000 1067.8000 ;
        RECT 461.9000 1072.7600 464.9000 1073.2400 ;
        RECT 473.6600 1051.0000 475.2600 1051.4800 ;
        RECT 473.6600 1056.4400 475.2600 1056.9200 ;
        RECT 461.9000 1051.0000 464.9000 1051.4800 ;
        RECT 461.9000 1056.4400 464.9000 1056.9200 ;
        RECT 563.6600 1034.6800 565.2600 1035.1600 ;
        RECT 563.6600 1040.1200 565.2600 1040.6000 ;
        RECT 563.6600 1045.5600 565.2600 1046.0400 ;
        RECT 563.6600 1023.8000 565.2600 1024.2800 ;
        RECT 563.6600 1029.2400 565.2600 1029.7200 ;
        RECT 518.6600 1034.6800 520.2600 1035.1600 ;
        RECT 518.6600 1040.1200 520.2600 1040.6000 ;
        RECT 518.6600 1045.5600 520.2600 1046.0400 ;
        RECT 518.6600 1023.8000 520.2600 1024.2800 ;
        RECT 518.6600 1029.2400 520.2600 1029.7200 ;
        RECT 563.6600 1007.4800 565.2600 1007.9600 ;
        RECT 563.6600 1012.9200 565.2600 1013.4000 ;
        RECT 563.6600 1018.3600 565.2600 1018.8400 ;
        RECT 563.6600 1002.0400 565.2600 1002.5200 ;
        RECT 518.6600 1007.4800 520.2600 1007.9600 ;
        RECT 518.6600 1012.9200 520.2600 1013.4000 ;
        RECT 518.6600 1018.3600 520.2600 1018.8400 ;
        RECT 518.6600 1002.0400 520.2600 1002.5200 ;
        RECT 473.6600 1034.6800 475.2600 1035.1600 ;
        RECT 473.6600 1040.1200 475.2600 1040.6000 ;
        RECT 473.6600 1045.5600 475.2600 1046.0400 ;
        RECT 461.9000 1034.6800 464.9000 1035.1600 ;
        RECT 461.9000 1040.1200 464.9000 1040.6000 ;
        RECT 461.9000 1045.5600 464.9000 1046.0400 ;
        RECT 473.6600 1023.8000 475.2600 1024.2800 ;
        RECT 473.6600 1029.2400 475.2600 1029.7200 ;
        RECT 461.9000 1023.8000 464.9000 1024.2800 ;
        RECT 461.9000 1029.2400 464.9000 1029.7200 ;
        RECT 473.6600 1007.4800 475.2600 1007.9600 ;
        RECT 473.6600 1012.9200 475.2600 1013.4000 ;
        RECT 473.6600 1018.3600 475.2600 1018.8400 ;
        RECT 461.9000 1007.4800 464.9000 1007.9600 ;
        RECT 461.9000 1012.9200 464.9000 1013.4000 ;
        RECT 461.9000 1018.3600 464.9000 1018.8400 ;
        RECT 461.9000 1002.0400 464.9000 1002.5200 ;
        RECT 473.6600 1002.0400 475.2600 1002.5200 ;
        RECT 461.9000 1206.9500 669.0000 1209.9500 ;
        RECT 461.9000 993.8500 669.0000 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 653.6600 764.2100 655.2600 980.3100 ;
        RECT 608.6600 764.2100 610.2600 980.3100 ;
        RECT 563.6600 764.2100 565.2600 980.3100 ;
        RECT 518.6600 764.2100 520.2600 980.3100 ;
        RECT 473.6600 764.2100 475.2600 980.3100 ;
        RECT 666.0000 764.2100 669.0000 980.3100 ;
        RECT 461.9000 764.2100 464.9000 980.3100 ;
      LAYER met3 ;
        RECT 666.0000 957.3600 669.0000 957.8400 ;
        RECT 666.0000 962.8000 669.0000 963.2800 ;
        RECT 653.6600 957.3600 655.2600 957.8400 ;
        RECT 653.6600 962.8000 655.2600 963.2800 ;
        RECT 666.0000 968.2400 669.0000 968.7200 ;
        RECT 653.6600 968.2400 655.2600 968.7200 ;
        RECT 666.0000 946.4800 669.0000 946.9600 ;
        RECT 666.0000 951.9200 669.0000 952.4000 ;
        RECT 653.6600 946.4800 655.2600 946.9600 ;
        RECT 653.6600 951.9200 655.2600 952.4000 ;
        RECT 666.0000 930.1600 669.0000 930.6400 ;
        RECT 666.0000 935.6000 669.0000 936.0800 ;
        RECT 653.6600 930.1600 655.2600 930.6400 ;
        RECT 653.6600 935.6000 655.2600 936.0800 ;
        RECT 666.0000 941.0400 669.0000 941.5200 ;
        RECT 653.6600 941.0400 655.2600 941.5200 ;
        RECT 608.6600 957.3600 610.2600 957.8400 ;
        RECT 608.6600 962.8000 610.2600 963.2800 ;
        RECT 608.6600 968.2400 610.2600 968.7200 ;
        RECT 608.6600 946.4800 610.2600 946.9600 ;
        RECT 608.6600 951.9200 610.2600 952.4000 ;
        RECT 608.6600 930.1600 610.2600 930.6400 ;
        RECT 608.6600 935.6000 610.2600 936.0800 ;
        RECT 608.6600 941.0400 610.2600 941.5200 ;
        RECT 666.0000 913.8400 669.0000 914.3200 ;
        RECT 666.0000 919.2800 669.0000 919.7600 ;
        RECT 666.0000 924.7200 669.0000 925.2000 ;
        RECT 653.6600 913.8400 655.2600 914.3200 ;
        RECT 653.6600 919.2800 655.2600 919.7600 ;
        RECT 653.6600 924.7200 655.2600 925.2000 ;
        RECT 666.0000 902.9600 669.0000 903.4400 ;
        RECT 666.0000 908.4000 669.0000 908.8800 ;
        RECT 653.6600 902.9600 655.2600 903.4400 ;
        RECT 653.6600 908.4000 655.2600 908.8800 ;
        RECT 666.0000 886.6400 669.0000 887.1200 ;
        RECT 666.0000 892.0800 669.0000 892.5600 ;
        RECT 666.0000 897.5200 669.0000 898.0000 ;
        RECT 653.6600 886.6400 655.2600 887.1200 ;
        RECT 653.6600 892.0800 655.2600 892.5600 ;
        RECT 653.6600 897.5200 655.2600 898.0000 ;
        RECT 666.0000 875.7600 669.0000 876.2400 ;
        RECT 666.0000 881.2000 669.0000 881.6800 ;
        RECT 653.6600 875.7600 655.2600 876.2400 ;
        RECT 653.6600 881.2000 655.2600 881.6800 ;
        RECT 608.6600 913.8400 610.2600 914.3200 ;
        RECT 608.6600 919.2800 610.2600 919.7600 ;
        RECT 608.6600 924.7200 610.2600 925.2000 ;
        RECT 608.6600 902.9600 610.2600 903.4400 ;
        RECT 608.6600 908.4000 610.2600 908.8800 ;
        RECT 608.6600 886.6400 610.2600 887.1200 ;
        RECT 608.6600 892.0800 610.2600 892.5600 ;
        RECT 608.6600 897.5200 610.2600 898.0000 ;
        RECT 608.6600 875.7600 610.2600 876.2400 ;
        RECT 608.6600 881.2000 610.2600 881.6800 ;
        RECT 563.6600 957.3600 565.2600 957.8400 ;
        RECT 563.6600 962.8000 565.2600 963.2800 ;
        RECT 563.6600 968.2400 565.2600 968.7200 ;
        RECT 518.6600 957.3600 520.2600 957.8400 ;
        RECT 518.6600 962.8000 520.2600 963.2800 ;
        RECT 518.6600 968.2400 520.2600 968.7200 ;
        RECT 563.6600 946.4800 565.2600 946.9600 ;
        RECT 563.6600 951.9200 565.2600 952.4000 ;
        RECT 563.6600 930.1600 565.2600 930.6400 ;
        RECT 563.6600 935.6000 565.2600 936.0800 ;
        RECT 563.6600 941.0400 565.2600 941.5200 ;
        RECT 518.6600 946.4800 520.2600 946.9600 ;
        RECT 518.6600 951.9200 520.2600 952.4000 ;
        RECT 518.6600 930.1600 520.2600 930.6400 ;
        RECT 518.6600 935.6000 520.2600 936.0800 ;
        RECT 518.6600 941.0400 520.2600 941.5200 ;
        RECT 473.6600 957.3600 475.2600 957.8400 ;
        RECT 473.6600 962.8000 475.2600 963.2800 ;
        RECT 461.9000 962.8000 464.9000 963.2800 ;
        RECT 461.9000 957.3600 464.9000 957.8400 ;
        RECT 461.9000 968.2400 464.9000 968.7200 ;
        RECT 473.6600 968.2400 475.2600 968.7200 ;
        RECT 473.6600 946.4800 475.2600 946.9600 ;
        RECT 473.6600 951.9200 475.2600 952.4000 ;
        RECT 461.9000 951.9200 464.9000 952.4000 ;
        RECT 461.9000 946.4800 464.9000 946.9600 ;
        RECT 473.6600 930.1600 475.2600 930.6400 ;
        RECT 473.6600 935.6000 475.2600 936.0800 ;
        RECT 461.9000 935.6000 464.9000 936.0800 ;
        RECT 461.9000 930.1600 464.9000 930.6400 ;
        RECT 461.9000 941.0400 464.9000 941.5200 ;
        RECT 473.6600 941.0400 475.2600 941.5200 ;
        RECT 563.6600 913.8400 565.2600 914.3200 ;
        RECT 563.6600 919.2800 565.2600 919.7600 ;
        RECT 563.6600 924.7200 565.2600 925.2000 ;
        RECT 563.6600 902.9600 565.2600 903.4400 ;
        RECT 563.6600 908.4000 565.2600 908.8800 ;
        RECT 518.6600 913.8400 520.2600 914.3200 ;
        RECT 518.6600 919.2800 520.2600 919.7600 ;
        RECT 518.6600 924.7200 520.2600 925.2000 ;
        RECT 518.6600 902.9600 520.2600 903.4400 ;
        RECT 518.6600 908.4000 520.2600 908.8800 ;
        RECT 563.6600 886.6400 565.2600 887.1200 ;
        RECT 563.6600 892.0800 565.2600 892.5600 ;
        RECT 563.6600 897.5200 565.2600 898.0000 ;
        RECT 563.6600 875.7600 565.2600 876.2400 ;
        RECT 563.6600 881.2000 565.2600 881.6800 ;
        RECT 518.6600 886.6400 520.2600 887.1200 ;
        RECT 518.6600 892.0800 520.2600 892.5600 ;
        RECT 518.6600 897.5200 520.2600 898.0000 ;
        RECT 518.6600 875.7600 520.2600 876.2400 ;
        RECT 518.6600 881.2000 520.2600 881.6800 ;
        RECT 473.6600 913.8400 475.2600 914.3200 ;
        RECT 473.6600 919.2800 475.2600 919.7600 ;
        RECT 473.6600 924.7200 475.2600 925.2000 ;
        RECT 461.9000 913.8400 464.9000 914.3200 ;
        RECT 461.9000 919.2800 464.9000 919.7600 ;
        RECT 461.9000 924.7200 464.9000 925.2000 ;
        RECT 473.6600 902.9600 475.2600 903.4400 ;
        RECT 473.6600 908.4000 475.2600 908.8800 ;
        RECT 461.9000 902.9600 464.9000 903.4400 ;
        RECT 461.9000 908.4000 464.9000 908.8800 ;
        RECT 473.6600 886.6400 475.2600 887.1200 ;
        RECT 473.6600 892.0800 475.2600 892.5600 ;
        RECT 473.6600 897.5200 475.2600 898.0000 ;
        RECT 461.9000 886.6400 464.9000 887.1200 ;
        RECT 461.9000 892.0800 464.9000 892.5600 ;
        RECT 461.9000 897.5200 464.9000 898.0000 ;
        RECT 473.6600 875.7600 475.2600 876.2400 ;
        RECT 473.6600 881.2000 475.2600 881.6800 ;
        RECT 461.9000 875.7600 464.9000 876.2400 ;
        RECT 461.9000 881.2000 464.9000 881.6800 ;
        RECT 666.0000 859.4400 669.0000 859.9200 ;
        RECT 666.0000 864.8800 669.0000 865.3600 ;
        RECT 666.0000 870.3200 669.0000 870.8000 ;
        RECT 653.6600 859.4400 655.2600 859.9200 ;
        RECT 653.6600 864.8800 655.2600 865.3600 ;
        RECT 653.6600 870.3200 655.2600 870.8000 ;
        RECT 666.0000 848.5600 669.0000 849.0400 ;
        RECT 666.0000 854.0000 669.0000 854.4800 ;
        RECT 653.6600 848.5600 655.2600 849.0400 ;
        RECT 653.6600 854.0000 655.2600 854.4800 ;
        RECT 666.0000 832.2400 669.0000 832.7200 ;
        RECT 666.0000 837.6800 669.0000 838.1600 ;
        RECT 666.0000 843.1200 669.0000 843.6000 ;
        RECT 653.6600 832.2400 655.2600 832.7200 ;
        RECT 653.6600 837.6800 655.2600 838.1600 ;
        RECT 653.6600 843.1200 655.2600 843.6000 ;
        RECT 666.0000 821.3600 669.0000 821.8400 ;
        RECT 666.0000 826.8000 669.0000 827.2800 ;
        RECT 653.6600 821.3600 655.2600 821.8400 ;
        RECT 653.6600 826.8000 655.2600 827.2800 ;
        RECT 608.6600 859.4400 610.2600 859.9200 ;
        RECT 608.6600 864.8800 610.2600 865.3600 ;
        RECT 608.6600 870.3200 610.2600 870.8000 ;
        RECT 608.6600 848.5600 610.2600 849.0400 ;
        RECT 608.6600 854.0000 610.2600 854.4800 ;
        RECT 608.6600 832.2400 610.2600 832.7200 ;
        RECT 608.6600 837.6800 610.2600 838.1600 ;
        RECT 608.6600 843.1200 610.2600 843.6000 ;
        RECT 608.6600 821.3600 610.2600 821.8400 ;
        RECT 608.6600 826.8000 610.2600 827.2800 ;
        RECT 666.0000 805.0400 669.0000 805.5200 ;
        RECT 666.0000 810.4800 669.0000 810.9600 ;
        RECT 666.0000 815.9200 669.0000 816.4000 ;
        RECT 653.6600 805.0400 655.2600 805.5200 ;
        RECT 653.6600 810.4800 655.2600 810.9600 ;
        RECT 653.6600 815.9200 655.2600 816.4000 ;
        RECT 666.0000 794.1600 669.0000 794.6400 ;
        RECT 666.0000 799.6000 669.0000 800.0800 ;
        RECT 653.6600 794.1600 655.2600 794.6400 ;
        RECT 653.6600 799.6000 655.2600 800.0800 ;
        RECT 666.0000 777.8400 669.0000 778.3200 ;
        RECT 666.0000 783.2800 669.0000 783.7600 ;
        RECT 666.0000 788.7200 669.0000 789.2000 ;
        RECT 653.6600 777.8400 655.2600 778.3200 ;
        RECT 653.6600 783.2800 655.2600 783.7600 ;
        RECT 653.6600 788.7200 655.2600 789.2000 ;
        RECT 666.0000 772.4000 669.0000 772.8800 ;
        RECT 653.6600 772.4000 655.2600 772.8800 ;
        RECT 608.6600 805.0400 610.2600 805.5200 ;
        RECT 608.6600 810.4800 610.2600 810.9600 ;
        RECT 608.6600 815.9200 610.2600 816.4000 ;
        RECT 608.6600 794.1600 610.2600 794.6400 ;
        RECT 608.6600 799.6000 610.2600 800.0800 ;
        RECT 608.6600 777.8400 610.2600 778.3200 ;
        RECT 608.6600 783.2800 610.2600 783.7600 ;
        RECT 608.6600 788.7200 610.2600 789.2000 ;
        RECT 608.6600 772.4000 610.2600 772.8800 ;
        RECT 563.6600 859.4400 565.2600 859.9200 ;
        RECT 563.6600 864.8800 565.2600 865.3600 ;
        RECT 563.6600 870.3200 565.2600 870.8000 ;
        RECT 563.6600 848.5600 565.2600 849.0400 ;
        RECT 563.6600 854.0000 565.2600 854.4800 ;
        RECT 518.6600 859.4400 520.2600 859.9200 ;
        RECT 518.6600 864.8800 520.2600 865.3600 ;
        RECT 518.6600 870.3200 520.2600 870.8000 ;
        RECT 518.6600 848.5600 520.2600 849.0400 ;
        RECT 518.6600 854.0000 520.2600 854.4800 ;
        RECT 563.6600 832.2400 565.2600 832.7200 ;
        RECT 563.6600 837.6800 565.2600 838.1600 ;
        RECT 563.6600 843.1200 565.2600 843.6000 ;
        RECT 563.6600 821.3600 565.2600 821.8400 ;
        RECT 563.6600 826.8000 565.2600 827.2800 ;
        RECT 518.6600 832.2400 520.2600 832.7200 ;
        RECT 518.6600 837.6800 520.2600 838.1600 ;
        RECT 518.6600 843.1200 520.2600 843.6000 ;
        RECT 518.6600 821.3600 520.2600 821.8400 ;
        RECT 518.6600 826.8000 520.2600 827.2800 ;
        RECT 473.6600 859.4400 475.2600 859.9200 ;
        RECT 473.6600 864.8800 475.2600 865.3600 ;
        RECT 473.6600 870.3200 475.2600 870.8000 ;
        RECT 461.9000 859.4400 464.9000 859.9200 ;
        RECT 461.9000 864.8800 464.9000 865.3600 ;
        RECT 461.9000 870.3200 464.9000 870.8000 ;
        RECT 473.6600 848.5600 475.2600 849.0400 ;
        RECT 473.6600 854.0000 475.2600 854.4800 ;
        RECT 461.9000 848.5600 464.9000 849.0400 ;
        RECT 461.9000 854.0000 464.9000 854.4800 ;
        RECT 473.6600 832.2400 475.2600 832.7200 ;
        RECT 473.6600 837.6800 475.2600 838.1600 ;
        RECT 473.6600 843.1200 475.2600 843.6000 ;
        RECT 461.9000 832.2400 464.9000 832.7200 ;
        RECT 461.9000 837.6800 464.9000 838.1600 ;
        RECT 461.9000 843.1200 464.9000 843.6000 ;
        RECT 473.6600 821.3600 475.2600 821.8400 ;
        RECT 473.6600 826.8000 475.2600 827.2800 ;
        RECT 461.9000 821.3600 464.9000 821.8400 ;
        RECT 461.9000 826.8000 464.9000 827.2800 ;
        RECT 563.6600 805.0400 565.2600 805.5200 ;
        RECT 563.6600 810.4800 565.2600 810.9600 ;
        RECT 563.6600 815.9200 565.2600 816.4000 ;
        RECT 563.6600 794.1600 565.2600 794.6400 ;
        RECT 563.6600 799.6000 565.2600 800.0800 ;
        RECT 518.6600 805.0400 520.2600 805.5200 ;
        RECT 518.6600 810.4800 520.2600 810.9600 ;
        RECT 518.6600 815.9200 520.2600 816.4000 ;
        RECT 518.6600 794.1600 520.2600 794.6400 ;
        RECT 518.6600 799.6000 520.2600 800.0800 ;
        RECT 563.6600 777.8400 565.2600 778.3200 ;
        RECT 563.6600 783.2800 565.2600 783.7600 ;
        RECT 563.6600 788.7200 565.2600 789.2000 ;
        RECT 563.6600 772.4000 565.2600 772.8800 ;
        RECT 518.6600 777.8400 520.2600 778.3200 ;
        RECT 518.6600 783.2800 520.2600 783.7600 ;
        RECT 518.6600 788.7200 520.2600 789.2000 ;
        RECT 518.6600 772.4000 520.2600 772.8800 ;
        RECT 473.6600 805.0400 475.2600 805.5200 ;
        RECT 473.6600 810.4800 475.2600 810.9600 ;
        RECT 473.6600 815.9200 475.2600 816.4000 ;
        RECT 461.9000 805.0400 464.9000 805.5200 ;
        RECT 461.9000 810.4800 464.9000 810.9600 ;
        RECT 461.9000 815.9200 464.9000 816.4000 ;
        RECT 473.6600 794.1600 475.2600 794.6400 ;
        RECT 473.6600 799.6000 475.2600 800.0800 ;
        RECT 461.9000 794.1600 464.9000 794.6400 ;
        RECT 461.9000 799.6000 464.9000 800.0800 ;
        RECT 473.6600 777.8400 475.2600 778.3200 ;
        RECT 473.6600 783.2800 475.2600 783.7600 ;
        RECT 473.6600 788.7200 475.2600 789.2000 ;
        RECT 461.9000 777.8400 464.9000 778.3200 ;
        RECT 461.9000 783.2800 464.9000 783.7600 ;
        RECT 461.9000 788.7200 464.9000 789.2000 ;
        RECT 461.9000 772.4000 464.9000 772.8800 ;
        RECT 473.6600 772.4000 475.2600 772.8800 ;
        RECT 461.9000 977.3100 669.0000 980.3100 ;
        RECT 461.9000 764.2100 669.0000 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 683.1200 2830.6100 685.1200 2857.5400 ;
        RECT 886.2200 2830.6100 888.2200 2857.5400 ;
      LAYER met3 ;
        RECT 886.2200 2847.3200 888.2200 2847.8000 ;
        RECT 683.1200 2847.3200 685.1200 2847.8000 ;
        RECT 886.2200 2841.8800 888.2200 2842.3600 ;
        RECT 886.2200 2836.4400 888.2200 2836.9200 ;
        RECT 683.1200 2841.8800 685.1200 2842.3600 ;
        RECT 683.1200 2836.4400 685.1200 2836.9200 ;
        RECT 683.1200 2855.5400 888.2200 2857.5400 ;
        RECT 683.1200 2830.6100 888.2200 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 534.5700 875.4800 750.6700 ;
        RECT 828.8800 534.5700 830.4800 750.6700 ;
        RECT 783.8800 534.5700 785.4800 750.6700 ;
        RECT 738.8800 534.5700 740.4800 750.6700 ;
        RECT 693.8800 534.5700 695.4800 750.6700 ;
        RECT 886.2200 534.5700 889.2200 750.6700 ;
        RECT 682.1200 534.5700 685.1200 750.6700 ;
      LAYER met3 ;
        RECT 886.2200 727.7200 889.2200 728.2000 ;
        RECT 886.2200 733.1600 889.2200 733.6400 ;
        RECT 873.8800 727.7200 875.4800 728.2000 ;
        RECT 873.8800 733.1600 875.4800 733.6400 ;
        RECT 886.2200 738.6000 889.2200 739.0800 ;
        RECT 873.8800 738.6000 875.4800 739.0800 ;
        RECT 886.2200 716.8400 889.2200 717.3200 ;
        RECT 886.2200 722.2800 889.2200 722.7600 ;
        RECT 873.8800 716.8400 875.4800 717.3200 ;
        RECT 873.8800 722.2800 875.4800 722.7600 ;
        RECT 886.2200 700.5200 889.2200 701.0000 ;
        RECT 886.2200 705.9600 889.2200 706.4400 ;
        RECT 873.8800 700.5200 875.4800 701.0000 ;
        RECT 873.8800 705.9600 875.4800 706.4400 ;
        RECT 886.2200 711.4000 889.2200 711.8800 ;
        RECT 873.8800 711.4000 875.4800 711.8800 ;
        RECT 828.8800 727.7200 830.4800 728.2000 ;
        RECT 828.8800 733.1600 830.4800 733.6400 ;
        RECT 828.8800 738.6000 830.4800 739.0800 ;
        RECT 828.8800 716.8400 830.4800 717.3200 ;
        RECT 828.8800 722.2800 830.4800 722.7600 ;
        RECT 828.8800 700.5200 830.4800 701.0000 ;
        RECT 828.8800 705.9600 830.4800 706.4400 ;
        RECT 828.8800 711.4000 830.4800 711.8800 ;
        RECT 886.2200 684.2000 889.2200 684.6800 ;
        RECT 886.2200 689.6400 889.2200 690.1200 ;
        RECT 886.2200 695.0800 889.2200 695.5600 ;
        RECT 873.8800 684.2000 875.4800 684.6800 ;
        RECT 873.8800 689.6400 875.4800 690.1200 ;
        RECT 873.8800 695.0800 875.4800 695.5600 ;
        RECT 886.2200 673.3200 889.2200 673.8000 ;
        RECT 886.2200 678.7600 889.2200 679.2400 ;
        RECT 873.8800 673.3200 875.4800 673.8000 ;
        RECT 873.8800 678.7600 875.4800 679.2400 ;
        RECT 886.2200 657.0000 889.2200 657.4800 ;
        RECT 886.2200 662.4400 889.2200 662.9200 ;
        RECT 886.2200 667.8800 889.2200 668.3600 ;
        RECT 873.8800 657.0000 875.4800 657.4800 ;
        RECT 873.8800 662.4400 875.4800 662.9200 ;
        RECT 873.8800 667.8800 875.4800 668.3600 ;
        RECT 886.2200 646.1200 889.2200 646.6000 ;
        RECT 886.2200 651.5600 889.2200 652.0400 ;
        RECT 873.8800 646.1200 875.4800 646.6000 ;
        RECT 873.8800 651.5600 875.4800 652.0400 ;
        RECT 828.8800 684.2000 830.4800 684.6800 ;
        RECT 828.8800 689.6400 830.4800 690.1200 ;
        RECT 828.8800 695.0800 830.4800 695.5600 ;
        RECT 828.8800 673.3200 830.4800 673.8000 ;
        RECT 828.8800 678.7600 830.4800 679.2400 ;
        RECT 828.8800 657.0000 830.4800 657.4800 ;
        RECT 828.8800 662.4400 830.4800 662.9200 ;
        RECT 828.8800 667.8800 830.4800 668.3600 ;
        RECT 828.8800 646.1200 830.4800 646.6000 ;
        RECT 828.8800 651.5600 830.4800 652.0400 ;
        RECT 783.8800 727.7200 785.4800 728.2000 ;
        RECT 783.8800 733.1600 785.4800 733.6400 ;
        RECT 783.8800 738.6000 785.4800 739.0800 ;
        RECT 738.8800 727.7200 740.4800 728.2000 ;
        RECT 738.8800 733.1600 740.4800 733.6400 ;
        RECT 738.8800 738.6000 740.4800 739.0800 ;
        RECT 783.8800 716.8400 785.4800 717.3200 ;
        RECT 783.8800 722.2800 785.4800 722.7600 ;
        RECT 783.8800 700.5200 785.4800 701.0000 ;
        RECT 783.8800 705.9600 785.4800 706.4400 ;
        RECT 783.8800 711.4000 785.4800 711.8800 ;
        RECT 738.8800 716.8400 740.4800 717.3200 ;
        RECT 738.8800 722.2800 740.4800 722.7600 ;
        RECT 738.8800 700.5200 740.4800 701.0000 ;
        RECT 738.8800 705.9600 740.4800 706.4400 ;
        RECT 738.8800 711.4000 740.4800 711.8800 ;
        RECT 693.8800 727.7200 695.4800 728.2000 ;
        RECT 693.8800 733.1600 695.4800 733.6400 ;
        RECT 682.1200 733.1600 685.1200 733.6400 ;
        RECT 682.1200 727.7200 685.1200 728.2000 ;
        RECT 682.1200 738.6000 685.1200 739.0800 ;
        RECT 693.8800 738.6000 695.4800 739.0800 ;
        RECT 693.8800 716.8400 695.4800 717.3200 ;
        RECT 693.8800 722.2800 695.4800 722.7600 ;
        RECT 682.1200 722.2800 685.1200 722.7600 ;
        RECT 682.1200 716.8400 685.1200 717.3200 ;
        RECT 693.8800 700.5200 695.4800 701.0000 ;
        RECT 693.8800 705.9600 695.4800 706.4400 ;
        RECT 682.1200 705.9600 685.1200 706.4400 ;
        RECT 682.1200 700.5200 685.1200 701.0000 ;
        RECT 682.1200 711.4000 685.1200 711.8800 ;
        RECT 693.8800 711.4000 695.4800 711.8800 ;
        RECT 783.8800 684.2000 785.4800 684.6800 ;
        RECT 783.8800 689.6400 785.4800 690.1200 ;
        RECT 783.8800 695.0800 785.4800 695.5600 ;
        RECT 783.8800 673.3200 785.4800 673.8000 ;
        RECT 783.8800 678.7600 785.4800 679.2400 ;
        RECT 738.8800 684.2000 740.4800 684.6800 ;
        RECT 738.8800 689.6400 740.4800 690.1200 ;
        RECT 738.8800 695.0800 740.4800 695.5600 ;
        RECT 738.8800 673.3200 740.4800 673.8000 ;
        RECT 738.8800 678.7600 740.4800 679.2400 ;
        RECT 783.8800 657.0000 785.4800 657.4800 ;
        RECT 783.8800 662.4400 785.4800 662.9200 ;
        RECT 783.8800 667.8800 785.4800 668.3600 ;
        RECT 783.8800 646.1200 785.4800 646.6000 ;
        RECT 783.8800 651.5600 785.4800 652.0400 ;
        RECT 738.8800 657.0000 740.4800 657.4800 ;
        RECT 738.8800 662.4400 740.4800 662.9200 ;
        RECT 738.8800 667.8800 740.4800 668.3600 ;
        RECT 738.8800 646.1200 740.4800 646.6000 ;
        RECT 738.8800 651.5600 740.4800 652.0400 ;
        RECT 693.8800 684.2000 695.4800 684.6800 ;
        RECT 693.8800 689.6400 695.4800 690.1200 ;
        RECT 693.8800 695.0800 695.4800 695.5600 ;
        RECT 682.1200 684.2000 685.1200 684.6800 ;
        RECT 682.1200 689.6400 685.1200 690.1200 ;
        RECT 682.1200 695.0800 685.1200 695.5600 ;
        RECT 693.8800 673.3200 695.4800 673.8000 ;
        RECT 693.8800 678.7600 695.4800 679.2400 ;
        RECT 682.1200 673.3200 685.1200 673.8000 ;
        RECT 682.1200 678.7600 685.1200 679.2400 ;
        RECT 693.8800 657.0000 695.4800 657.4800 ;
        RECT 693.8800 662.4400 695.4800 662.9200 ;
        RECT 693.8800 667.8800 695.4800 668.3600 ;
        RECT 682.1200 657.0000 685.1200 657.4800 ;
        RECT 682.1200 662.4400 685.1200 662.9200 ;
        RECT 682.1200 667.8800 685.1200 668.3600 ;
        RECT 693.8800 646.1200 695.4800 646.6000 ;
        RECT 693.8800 651.5600 695.4800 652.0400 ;
        RECT 682.1200 646.1200 685.1200 646.6000 ;
        RECT 682.1200 651.5600 685.1200 652.0400 ;
        RECT 886.2200 629.8000 889.2200 630.2800 ;
        RECT 886.2200 635.2400 889.2200 635.7200 ;
        RECT 886.2200 640.6800 889.2200 641.1600 ;
        RECT 873.8800 629.8000 875.4800 630.2800 ;
        RECT 873.8800 635.2400 875.4800 635.7200 ;
        RECT 873.8800 640.6800 875.4800 641.1600 ;
        RECT 886.2200 618.9200 889.2200 619.4000 ;
        RECT 886.2200 624.3600 889.2200 624.8400 ;
        RECT 873.8800 618.9200 875.4800 619.4000 ;
        RECT 873.8800 624.3600 875.4800 624.8400 ;
        RECT 886.2200 602.6000 889.2200 603.0800 ;
        RECT 886.2200 608.0400 889.2200 608.5200 ;
        RECT 886.2200 613.4800 889.2200 613.9600 ;
        RECT 873.8800 602.6000 875.4800 603.0800 ;
        RECT 873.8800 608.0400 875.4800 608.5200 ;
        RECT 873.8800 613.4800 875.4800 613.9600 ;
        RECT 886.2200 591.7200 889.2200 592.2000 ;
        RECT 886.2200 597.1600 889.2200 597.6400 ;
        RECT 873.8800 591.7200 875.4800 592.2000 ;
        RECT 873.8800 597.1600 875.4800 597.6400 ;
        RECT 828.8800 629.8000 830.4800 630.2800 ;
        RECT 828.8800 635.2400 830.4800 635.7200 ;
        RECT 828.8800 640.6800 830.4800 641.1600 ;
        RECT 828.8800 618.9200 830.4800 619.4000 ;
        RECT 828.8800 624.3600 830.4800 624.8400 ;
        RECT 828.8800 602.6000 830.4800 603.0800 ;
        RECT 828.8800 608.0400 830.4800 608.5200 ;
        RECT 828.8800 613.4800 830.4800 613.9600 ;
        RECT 828.8800 591.7200 830.4800 592.2000 ;
        RECT 828.8800 597.1600 830.4800 597.6400 ;
        RECT 886.2200 575.4000 889.2200 575.8800 ;
        RECT 886.2200 580.8400 889.2200 581.3200 ;
        RECT 886.2200 586.2800 889.2200 586.7600 ;
        RECT 873.8800 575.4000 875.4800 575.8800 ;
        RECT 873.8800 580.8400 875.4800 581.3200 ;
        RECT 873.8800 586.2800 875.4800 586.7600 ;
        RECT 886.2200 564.5200 889.2200 565.0000 ;
        RECT 886.2200 569.9600 889.2200 570.4400 ;
        RECT 873.8800 564.5200 875.4800 565.0000 ;
        RECT 873.8800 569.9600 875.4800 570.4400 ;
        RECT 886.2200 548.2000 889.2200 548.6800 ;
        RECT 886.2200 553.6400 889.2200 554.1200 ;
        RECT 886.2200 559.0800 889.2200 559.5600 ;
        RECT 873.8800 548.2000 875.4800 548.6800 ;
        RECT 873.8800 553.6400 875.4800 554.1200 ;
        RECT 873.8800 559.0800 875.4800 559.5600 ;
        RECT 886.2200 542.7600 889.2200 543.2400 ;
        RECT 873.8800 542.7600 875.4800 543.2400 ;
        RECT 828.8800 575.4000 830.4800 575.8800 ;
        RECT 828.8800 580.8400 830.4800 581.3200 ;
        RECT 828.8800 586.2800 830.4800 586.7600 ;
        RECT 828.8800 564.5200 830.4800 565.0000 ;
        RECT 828.8800 569.9600 830.4800 570.4400 ;
        RECT 828.8800 548.2000 830.4800 548.6800 ;
        RECT 828.8800 553.6400 830.4800 554.1200 ;
        RECT 828.8800 559.0800 830.4800 559.5600 ;
        RECT 828.8800 542.7600 830.4800 543.2400 ;
        RECT 783.8800 629.8000 785.4800 630.2800 ;
        RECT 783.8800 635.2400 785.4800 635.7200 ;
        RECT 783.8800 640.6800 785.4800 641.1600 ;
        RECT 783.8800 618.9200 785.4800 619.4000 ;
        RECT 783.8800 624.3600 785.4800 624.8400 ;
        RECT 738.8800 629.8000 740.4800 630.2800 ;
        RECT 738.8800 635.2400 740.4800 635.7200 ;
        RECT 738.8800 640.6800 740.4800 641.1600 ;
        RECT 738.8800 618.9200 740.4800 619.4000 ;
        RECT 738.8800 624.3600 740.4800 624.8400 ;
        RECT 783.8800 602.6000 785.4800 603.0800 ;
        RECT 783.8800 608.0400 785.4800 608.5200 ;
        RECT 783.8800 613.4800 785.4800 613.9600 ;
        RECT 783.8800 591.7200 785.4800 592.2000 ;
        RECT 783.8800 597.1600 785.4800 597.6400 ;
        RECT 738.8800 602.6000 740.4800 603.0800 ;
        RECT 738.8800 608.0400 740.4800 608.5200 ;
        RECT 738.8800 613.4800 740.4800 613.9600 ;
        RECT 738.8800 591.7200 740.4800 592.2000 ;
        RECT 738.8800 597.1600 740.4800 597.6400 ;
        RECT 693.8800 629.8000 695.4800 630.2800 ;
        RECT 693.8800 635.2400 695.4800 635.7200 ;
        RECT 693.8800 640.6800 695.4800 641.1600 ;
        RECT 682.1200 629.8000 685.1200 630.2800 ;
        RECT 682.1200 635.2400 685.1200 635.7200 ;
        RECT 682.1200 640.6800 685.1200 641.1600 ;
        RECT 693.8800 618.9200 695.4800 619.4000 ;
        RECT 693.8800 624.3600 695.4800 624.8400 ;
        RECT 682.1200 618.9200 685.1200 619.4000 ;
        RECT 682.1200 624.3600 685.1200 624.8400 ;
        RECT 693.8800 602.6000 695.4800 603.0800 ;
        RECT 693.8800 608.0400 695.4800 608.5200 ;
        RECT 693.8800 613.4800 695.4800 613.9600 ;
        RECT 682.1200 602.6000 685.1200 603.0800 ;
        RECT 682.1200 608.0400 685.1200 608.5200 ;
        RECT 682.1200 613.4800 685.1200 613.9600 ;
        RECT 693.8800 591.7200 695.4800 592.2000 ;
        RECT 693.8800 597.1600 695.4800 597.6400 ;
        RECT 682.1200 591.7200 685.1200 592.2000 ;
        RECT 682.1200 597.1600 685.1200 597.6400 ;
        RECT 783.8800 575.4000 785.4800 575.8800 ;
        RECT 783.8800 580.8400 785.4800 581.3200 ;
        RECT 783.8800 586.2800 785.4800 586.7600 ;
        RECT 783.8800 564.5200 785.4800 565.0000 ;
        RECT 783.8800 569.9600 785.4800 570.4400 ;
        RECT 738.8800 575.4000 740.4800 575.8800 ;
        RECT 738.8800 580.8400 740.4800 581.3200 ;
        RECT 738.8800 586.2800 740.4800 586.7600 ;
        RECT 738.8800 564.5200 740.4800 565.0000 ;
        RECT 738.8800 569.9600 740.4800 570.4400 ;
        RECT 783.8800 548.2000 785.4800 548.6800 ;
        RECT 783.8800 553.6400 785.4800 554.1200 ;
        RECT 783.8800 559.0800 785.4800 559.5600 ;
        RECT 783.8800 542.7600 785.4800 543.2400 ;
        RECT 738.8800 548.2000 740.4800 548.6800 ;
        RECT 738.8800 553.6400 740.4800 554.1200 ;
        RECT 738.8800 559.0800 740.4800 559.5600 ;
        RECT 738.8800 542.7600 740.4800 543.2400 ;
        RECT 693.8800 575.4000 695.4800 575.8800 ;
        RECT 693.8800 580.8400 695.4800 581.3200 ;
        RECT 693.8800 586.2800 695.4800 586.7600 ;
        RECT 682.1200 575.4000 685.1200 575.8800 ;
        RECT 682.1200 580.8400 685.1200 581.3200 ;
        RECT 682.1200 586.2800 685.1200 586.7600 ;
        RECT 693.8800 564.5200 695.4800 565.0000 ;
        RECT 693.8800 569.9600 695.4800 570.4400 ;
        RECT 682.1200 564.5200 685.1200 565.0000 ;
        RECT 682.1200 569.9600 685.1200 570.4400 ;
        RECT 693.8800 548.2000 695.4800 548.6800 ;
        RECT 693.8800 553.6400 695.4800 554.1200 ;
        RECT 693.8800 559.0800 695.4800 559.5600 ;
        RECT 682.1200 548.2000 685.1200 548.6800 ;
        RECT 682.1200 553.6400 685.1200 554.1200 ;
        RECT 682.1200 559.0800 685.1200 559.5600 ;
        RECT 682.1200 542.7600 685.1200 543.2400 ;
        RECT 693.8800 542.7600 695.4800 543.2400 ;
        RECT 682.1200 747.6700 889.2200 750.6700 ;
        RECT 682.1200 534.5700 889.2200 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 304.9300 875.4800 521.0300 ;
        RECT 828.8800 304.9300 830.4800 521.0300 ;
        RECT 783.8800 304.9300 785.4800 521.0300 ;
        RECT 738.8800 304.9300 740.4800 521.0300 ;
        RECT 693.8800 304.9300 695.4800 521.0300 ;
        RECT 886.2200 304.9300 889.2200 521.0300 ;
        RECT 682.1200 304.9300 685.1200 521.0300 ;
      LAYER met3 ;
        RECT 886.2200 498.0800 889.2200 498.5600 ;
        RECT 886.2200 503.5200 889.2200 504.0000 ;
        RECT 873.8800 498.0800 875.4800 498.5600 ;
        RECT 873.8800 503.5200 875.4800 504.0000 ;
        RECT 886.2200 508.9600 889.2200 509.4400 ;
        RECT 873.8800 508.9600 875.4800 509.4400 ;
        RECT 886.2200 487.2000 889.2200 487.6800 ;
        RECT 886.2200 492.6400 889.2200 493.1200 ;
        RECT 873.8800 487.2000 875.4800 487.6800 ;
        RECT 873.8800 492.6400 875.4800 493.1200 ;
        RECT 886.2200 470.8800 889.2200 471.3600 ;
        RECT 886.2200 476.3200 889.2200 476.8000 ;
        RECT 873.8800 470.8800 875.4800 471.3600 ;
        RECT 873.8800 476.3200 875.4800 476.8000 ;
        RECT 886.2200 481.7600 889.2200 482.2400 ;
        RECT 873.8800 481.7600 875.4800 482.2400 ;
        RECT 828.8800 498.0800 830.4800 498.5600 ;
        RECT 828.8800 503.5200 830.4800 504.0000 ;
        RECT 828.8800 508.9600 830.4800 509.4400 ;
        RECT 828.8800 487.2000 830.4800 487.6800 ;
        RECT 828.8800 492.6400 830.4800 493.1200 ;
        RECT 828.8800 470.8800 830.4800 471.3600 ;
        RECT 828.8800 476.3200 830.4800 476.8000 ;
        RECT 828.8800 481.7600 830.4800 482.2400 ;
        RECT 886.2200 454.5600 889.2200 455.0400 ;
        RECT 886.2200 460.0000 889.2200 460.4800 ;
        RECT 886.2200 465.4400 889.2200 465.9200 ;
        RECT 873.8800 454.5600 875.4800 455.0400 ;
        RECT 873.8800 460.0000 875.4800 460.4800 ;
        RECT 873.8800 465.4400 875.4800 465.9200 ;
        RECT 886.2200 443.6800 889.2200 444.1600 ;
        RECT 886.2200 449.1200 889.2200 449.6000 ;
        RECT 873.8800 443.6800 875.4800 444.1600 ;
        RECT 873.8800 449.1200 875.4800 449.6000 ;
        RECT 886.2200 427.3600 889.2200 427.8400 ;
        RECT 886.2200 432.8000 889.2200 433.2800 ;
        RECT 886.2200 438.2400 889.2200 438.7200 ;
        RECT 873.8800 427.3600 875.4800 427.8400 ;
        RECT 873.8800 432.8000 875.4800 433.2800 ;
        RECT 873.8800 438.2400 875.4800 438.7200 ;
        RECT 886.2200 416.4800 889.2200 416.9600 ;
        RECT 886.2200 421.9200 889.2200 422.4000 ;
        RECT 873.8800 416.4800 875.4800 416.9600 ;
        RECT 873.8800 421.9200 875.4800 422.4000 ;
        RECT 828.8800 454.5600 830.4800 455.0400 ;
        RECT 828.8800 460.0000 830.4800 460.4800 ;
        RECT 828.8800 465.4400 830.4800 465.9200 ;
        RECT 828.8800 443.6800 830.4800 444.1600 ;
        RECT 828.8800 449.1200 830.4800 449.6000 ;
        RECT 828.8800 427.3600 830.4800 427.8400 ;
        RECT 828.8800 432.8000 830.4800 433.2800 ;
        RECT 828.8800 438.2400 830.4800 438.7200 ;
        RECT 828.8800 416.4800 830.4800 416.9600 ;
        RECT 828.8800 421.9200 830.4800 422.4000 ;
        RECT 783.8800 498.0800 785.4800 498.5600 ;
        RECT 783.8800 503.5200 785.4800 504.0000 ;
        RECT 783.8800 508.9600 785.4800 509.4400 ;
        RECT 738.8800 498.0800 740.4800 498.5600 ;
        RECT 738.8800 503.5200 740.4800 504.0000 ;
        RECT 738.8800 508.9600 740.4800 509.4400 ;
        RECT 783.8800 487.2000 785.4800 487.6800 ;
        RECT 783.8800 492.6400 785.4800 493.1200 ;
        RECT 783.8800 470.8800 785.4800 471.3600 ;
        RECT 783.8800 476.3200 785.4800 476.8000 ;
        RECT 783.8800 481.7600 785.4800 482.2400 ;
        RECT 738.8800 487.2000 740.4800 487.6800 ;
        RECT 738.8800 492.6400 740.4800 493.1200 ;
        RECT 738.8800 470.8800 740.4800 471.3600 ;
        RECT 738.8800 476.3200 740.4800 476.8000 ;
        RECT 738.8800 481.7600 740.4800 482.2400 ;
        RECT 693.8800 498.0800 695.4800 498.5600 ;
        RECT 693.8800 503.5200 695.4800 504.0000 ;
        RECT 682.1200 503.5200 685.1200 504.0000 ;
        RECT 682.1200 498.0800 685.1200 498.5600 ;
        RECT 682.1200 508.9600 685.1200 509.4400 ;
        RECT 693.8800 508.9600 695.4800 509.4400 ;
        RECT 693.8800 487.2000 695.4800 487.6800 ;
        RECT 693.8800 492.6400 695.4800 493.1200 ;
        RECT 682.1200 492.6400 685.1200 493.1200 ;
        RECT 682.1200 487.2000 685.1200 487.6800 ;
        RECT 693.8800 470.8800 695.4800 471.3600 ;
        RECT 693.8800 476.3200 695.4800 476.8000 ;
        RECT 682.1200 476.3200 685.1200 476.8000 ;
        RECT 682.1200 470.8800 685.1200 471.3600 ;
        RECT 682.1200 481.7600 685.1200 482.2400 ;
        RECT 693.8800 481.7600 695.4800 482.2400 ;
        RECT 783.8800 454.5600 785.4800 455.0400 ;
        RECT 783.8800 460.0000 785.4800 460.4800 ;
        RECT 783.8800 465.4400 785.4800 465.9200 ;
        RECT 783.8800 443.6800 785.4800 444.1600 ;
        RECT 783.8800 449.1200 785.4800 449.6000 ;
        RECT 738.8800 454.5600 740.4800 455.0400 ;
        RECT 738.8800 460.0000 740.4800 460.4800 ;
        RECT 738.8800 465.4400 740.4800 465.9200 ;
        RECT 738.8800 443.6800 740.4800 444.1600 ;
        RECT 738.8800 449.1200 740.4800 449.6000 ;
        RECT 783.8800 427.3600 785.4800 427.8400 ;
        RECT 783.8800 432.8000 785.4800 433.2800 ;
        RECT 783.8800 438.2400 785.4800 438.7200 ;
        RECT 783.8800 416.4800 785.4800 416.9600 ;
        RECT 783.8800 421.9200 785.4800 422.4000 ;
        RECT 738.8800 427.3600 740.4800 427.8400 ;
        RECT 738.8800 432.8000 740.4800 433.2800 ;
        RECT 738.8800 438.2400 740.4800 438.7200 ;
        RECT 738.8800 416.4800 740.4800 416.9600 ;
        RECT 738.8800 421.9200 740.4800 422.4000 ;
        RECT 693.8800 454.5600 695.4800 455.0400 ;
        RECT 693.8800 460.0000 695.4800 460.4800 ;
        RECT 693.8800 465.4400 695.4800 465.9200 ;
        RECT 682.1200 454.5600 685.1200 455.0400 ;
        RECT 682.1200 460.0000 685.1200 460.4800 ;
        RECT 682.1200 465.4400 685.1200 465.9200 ;
        RECT 693.8800 443.6800 695.4800 444.1600 ;
        RECT 693.8800 449.1200 695.4800 449.6000 ;
        RECT 682.1200 443.6800 685.1200 444.1600 ;
        RECT 682.1200 449.1200 685.1200 449.6000 ;
        RECT 693.8800 427.3600 695.4800 427.8400 ;
        RECT 693.8800 432.8000 695.4800 433.2800 ;
        RECT 693.8800 438.2400 695.4800 438.7200 ;
        RECT 682.1200 427.3600 685.1200 427.8400 ;
        RECT 682.1200 432.8000 685.1200 433.2800 ;
        RECT 682.1200 438.2400 685.1200 438.7200 ;
        RECT 693.8800 416.4800 695.4800 416.9600 ;
        RECT 693.8800 421.9200 695.4800 422.4000 ;
        RECT 682.1200 416.4800 685.1200 416.9600 ;
        RECT 682.1200 421.9200 685.1200 422.4000 ;
        RECT 886.2200 400.1600 889.2200 400.6400 ;
        RECT 886.2200 405.6000 889.2200 406.0800 ;
        RECT 886.2200 411.0400 889.2200 411.5200 ;
        RECT 873.8800 400.1600 875.4800 400.6400 ;
        RECT 873.8800 405.6000 875.4800 406.0800 ;
        RECT 873.8800 411.0400 875.4800 411.5200 ;
        RECT 886.2200 389.2800 889.2200 389.7600 ;
        RECT 886.2200 394.7200 889.2200 395.2000 ;
        RECT 873.8800 389.2800 875.4800 389.7600 ;
        RECT 873.8800 394.7200 875.4800 395.2000 ;
        RECT 886.2200 372.9600 889.2200 373.4400 ;
        RECT 886.2200 378.4000 889.2200 378.8800 ;
        RECT 886.2200 383.8400 889.2200 384.3200 ;
        RECT 873.8800 372.9600 875.4800 373.4400 ;
        RECT 873.8800 378.4000 875.4800 378.8800 ;
        RECT 873.8800 383.8400 875.4800 384.3200 ;
        RECT 886.2200 362.0800 889.2200 362.5600 ;
        RECT 886.2200 367.5200 889.2200 368.0000 ;
        RECT 873.8800 362.0800 875.4800 362.5600 ;
        RECT 873.8800 367.5200 875.4800 368.0000 ;
        RECT 828.8800 400.1600 830.4800 400.6400 ;
        RECT 828.8800 405.6000 830.4800 406.0800 ;
        RECT 828.8800 411.0400 830.4800 411.5200 ;
        RECT 828.8800 389.2800 830.4800 389.7600 ;
        RECT 828.8800 394.7200 830.4800 395.2000 ;
        RECT 828.8800 372.9600 830.4800 373.4400 ;
        RECT 828.8800 378.4000 830.4800 378.8800 ;
        RECT 828.8800 383.8400 830.4800 384.3200 ;
        RECT 828.8800 362.0800 830.4800 362.5600 ;
        RECT 828.8800 367.5200 830.4800 368.0000 ;
        RECT 886.2200 345.7600 889.2200 346.2400 ;
        RECT 886.2200 351.2000 889.2200 351.6800 ;
        RECT 886.2200 356.6400 889.2200 357.1200 ;
        RECT 873.8800 345.7600 875.4800 346.2400 ;
        RECT 873.8800 351.2000 875.4800 351.6800 ;
        RECT 873.8800 356.6400 875.4800 357.1200 ;
        RECT 886.2200 334.8800 889.2200 335.3600 ;
        RECT 886.2200 340.3200 889.2200 340.8000 ;
        RECT 873.8800 334.8800 875.4800 335.3600 ;
        RECT 873.8800 340.3200 875.4800 340.8000 ;
        RECT 886.2200 318.5600 889.2200 319.0400 ;
        RECT 886.2200 324.0000 889.2200 324.4800 ;
        RECT 886.2200 329.4400 889.2200 329.9200 ;
        RECT 873.8800 318.5600 875.4800 319.0400 ;
        RECT 873.8800 324.0000 875.4800 324.4800 ;
        RECT 873.8800 329.4400 875.4800 329.9200 ;
        RECT 886.2200 313.1200 889.2200 313.6000 ;
        RECT 873.8800 313.1200 875.4800 313.6000 ;
        RECT 828.8800 345.7600 830.4800 346.2400 ;
        RECT 828.8800 351.2000 830.4800 351.6800 ;
        RECT 828.8800 356.6400 830.4800 357.1200 ;
        RECT 828.8800 334.8800 830.4800 335.3600 ;
        RECT 828.8800 340.3200 830.4800 340.8000 ;
        RECT 828.8800 318.5600 830.4800 319.0400 ;
        RECT 828.8800 324.0000 830.4800 324.4800 ;
        RECT 828.8800 329.4400 830.4800 329.9200 ;
        RECT 828.8800 313.1200 830.4800 313.6000 ;
        RECT 783.8800 400.1600 785.4800 400.6400 ;
        RECT 783.8800 405.6000 785.4800 406.0800 ;
        RECT 783.8800 411.0400 785.4800 411.5200 ;
        RECT 783.8800 389.2800 785.4800 389.7600 ;
        RECT 783.8800 394.7200 785.4800 395.2000 ;
        RECT 738.8800 400.1600 740.4800 400.6400 ;
        RECT 738.8800 405.6000 740.4800 406.0800 ;
        RECT 738.8800 411.0400 740.4800 411.5200 ;
        RECT 738.8800 389.2800 740.4800 389.7600 ;
        RECT 738.8800 394.7200 740.4800 395.2000 ;
        RECT 783.8800 372.9600 785.4800 373.4400 ;
        RECT 783.8800 378.4000 785.4800 378.8800 ;
        RECT 783.8800 383.8400 785.4800 384.3200 ;
        RECT 783.8800 362.0800 785.4800 362.5600 ;
        RECT 783.8800 367.5200 785.4800 368.0000 ;
        RECT 738.8800 372.9600 740.4800 373.4400 ;
        RECT 738.8800 378.4000 740.4800 378.8800 ;
        RECT 738.8800 383.8400 740.4800 384.3200 ;
        RECT 738.8800 362.0800 740.4800 362.5600 ;
        RECT 738.8800 367.5200 740.4800 368.0000 ;
        RECT 693.8800 400.1600 695.4800 400.6400 ;
        RECT 693.8800 405.6000 695.4800 406.0800 ;
        RECT 693.8800 411.0400 695.4800 411.5200 ;
        RECT 682.1200 400.1600 685.1200 400.6400 ;
        RECT 682.1200 405.6000 685.1200 406.0800 ;
        RECT 682.1200 411.0400 685.1200 411.5200 ;
        RECT 693.8800 389.2800 695.4800 389.7600 ;
        RECT 693.8800 394.7200 695.4800 395.2000 ;
        RECT 682.1200 389.2800 685.1200 389.7600 ;
        RECT 682.1200 394.7200 685.1200 395.2000 ;
        RECT 693.8800 372.9600 695.4800 373.4400 ;
        RECT 693.8800 378.4000 695.4800 378.8800 ;
        RECT 693.8800 383.8400 695.4800 384.3200 ;
        RECT 682.1200 372.9600 685.1200 373.4400 ;
        RECT 682.1200 378.4000 685.1200 378.8800 ;
        RECT 682.1200 383.8400 685.1200 384.3200 ;
        RECT 693.8800 362.0800 695.4800 362.5600 ;
        RECT 693.8800 367.5200 695.4800 368.0000 ;
        RECT 682.1200 362.0800 685.1200 362.5600 ;
        RECT 682.1200 367.5200 685.1200 368.0000 ;
        RECT 783.8800 345.7600 785.4800 346.2400 ;
        RECT 783.8800 351.2000 785.4800 351.6800 ;
        RECT 783.8800 356.6400 785.4800 357.1200 ;
        RECT 783.8800 334.8800 785.4800 335.3600 ;
        RECT 783.8800 340.3200 785.4800 340.8000 ;
        RECT 738.8800 345.7600 740.4800 346.2400 ;
        RECT 738.8800 351.2000 740.4800 351.6800 ;
        RECT 738.8800 356.6400 740.4800 357.1200 ;
        RECT 738.8800 334.8800 740.4800 335.3600 ;
        RECT 738.8800 340.3200 740.4800 340.8000 ;
        RECT 783.8800 318.5600 785.4800 319.0400 ;
        RECT 783.8800 324.0000 785.4800 324.4800 ;
        RECT 783.8800 329.4400 785.4800 329.9200 ;
        RECT 783.8800 313.1200 785.4800 313.6000 ;
        RECT 738.8800 318.5600 740.4800 319.0400 ;
        RECT 738.8800 324.0000 740.4800 324.4800 ;
        RECT 738.8800 329.4400 740.4800 329.9200 ;
        RECT 738.8800 313.1200 740.4800 313.6000 ;
        RECT 693.8800 345.7600 695.4800 346.2400 ;
        RECT 693.8800 351.2000 695.4800 351.6800 ;
        RECT 693.8800 356.6400 695.4800 357.1200 ;
        RECT 682.1200 345.7600 685.1200 346.2400 ;
        RECT 682.1200 351.2000 685.1200 351.6800 ;
        RECT 682.1200 356.6400 685.1200 357.1200 ;
        RECT 693.8800 334.8800 695.4800 335.3600 ;
        RECT 693.8800 340.3200 695.4800 340.8000 ;
        RECT 682.1200 334.8800 685.1200 335.3600 ;
        RECT 682.1200 340.3200 685.1200 340.8000 ;
        RECT 693.8800 318.5600 695.4800 319.0400 ;
        RECT 693.8800 324.0000 695.4800 324.4800 ;
        RECT 693.8800 329.4400 695.4800 329.9200 ;
        RECT 682.1200 318.5600 685.1200 319.0400 ;
        RECT 682.1200 324.0000 685.1200 324.4800 ;
        RECT 682.1200 329.4400 685.1200 329.9200 ;
        RECT 682.1200 313.1200 685.1200 313.6000 ;
        RECT 693.8800 313.1200 695.4800 313.6000 ;
        RECT 682.1200 518.0300 889.2200 521.0300 ;
        RECT 682.1200 304.9300 889.2200 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 75.2900 875.4800 291.3900 ;
        RECT 828.8800 75.2900 830.4800 291.3900 ;
        RECT 783.8800 75.2900 785.4800 291.3900 ;
        RECT 738.8800 75.2900 740.4800 291.3900 ;
        RECT 693.8800 75.2900 695.4800 291.3900 ;
        RECT 886.2200 75.2900 889.2200 291.3900 ;
        RECT 682.1200 75.2900 685.1200 291.3900 ;
      LAYER met3 ;
        RECT 886.2200 268.4400 889.2200 268.9200 ;
        RECT 886.2200 273.8800 889.2200 274.3600 ;
        RECT 873.8800 268.4400 875.4800 268.9200 ;
        RECT 873.8800 273.8800 875.4800 274.3600 ;
        RECT 886.2200 279.3200 889.2200 279.8000 ;
        RECT 873.8800 279.3200 875.4800 279.8000 ;
        RECT 886.2200 257.5600 889.2200 258.0400 ;
        RECT 886.2200 263.0000 889.2200 263.4800 ;
        RECT 873.8800 257.5600 875.4800 258.0400 ;
        RECT 873.8800 263.0000 875.4800 263.4800 ;
        RECT 886.2200 241.2400 889.2200 241.7200 ;
        RECT 886.2200 246.6800 889.2200 247.1600 ;
        RECT 873.8800 241.2400 875.4800 241.7200 ;
        RECT 873.8800 246.6800 875.4800 247.1600 ;
        RECT 886.2200 252.1200 889.2200 252.6000 ;
        RECT 873.8800 252.1200 875.4800 252.6000 ;
        RECT 828.8800 268.4400 830.4800 268.9200 ;
        RECT 828.8800 273.8800 830.4800 274.3600 ;
        RECT 828.8800 279.3200 830.4800 279.8000 ;
        RECT 828.8800 257.5600 830.4800 258.0400 ;
        RECT 828.8800 263.0000 830.4800 263.4800 ;
        RECT 828.8800 241.2400 830.4800 241.7200 ;
        RECT 828.8800 246.6800 830.4800 247.1600 ;
        RECT 828.8800 252.1200 830.4800 252.6000 ;
        RECT 886.2200 224.9200 889.2200 225.4000 ;
        RECT 886.2200 230.3600 889.2200 230.8400 ;
        RECT 886.2200 235.8000 889.2200 236.2800 ;
        RECT 873.8800 224.9200 875.4800 225.4000 ;
        RECT 873.8800 230.3600 875.4800 230.8400 ;
        RECT 873.8800 235.8000 875.4800 236.2800 ;
        RECT 886.2200 214.0400 889.2200 214.5200 ;
        RECT 886.2200 219.4800 889.2200 219.9600 ;
        RECT 873.8800 214.0400 875.4800 214.5200 ;
        RECT 873.8800 219.4800 875.4800 219.9600 ;
        RECT 886.2200 197.7200 889.2200 198.2000 ;
        RECT 886.2200 203.1600 889.2200 203.6400 ;
        RECT 886.2200 208.6000 889.2200 209.0800 ;
        RECT 873.8800 197.7200 875.4800 198.2000 ;
        RECT 873.8800 203.1600 875.4800 203.6400 ;
        RECT 873.8800 208.6000 875.4800 209.0800 ;
        RECT 886.2200 186.8400 889.2200 187.3200 ;
        RECT 886.2200 192.2800 889.2200 192.7600 ;
        RECT 873.8800 186.8400 875.4800 187.3200 ;
        RECT 873.8800 192.2800 875.4800 192.7600 ;
        RECT 828.8800 224.9200 830.4800 225.4000 ;
        RECT 828.8800 230.3600 830.4800 230.8400 ;
        RECT 828.8800 235.8000 830.4800 236.2800 ;
        RECT 828.8800 214.0400 830.4800 214.5200 ;
        RECT 828.8800 219.4800 830.4800 219.9600 ;
        RECT 828.8800 197.7200 830.4800 198.2000 ;
        RECT 828.8800 203.1600 830.4800 203.6400 ;
        RECT 828.8800 208.6000 830.4800 209.0800 ;
        RECT 828.8800 186.8400 830.4800 187.3200 ;
        RECT 828.8800 192.2800 830.4800 192.7600 ;
        RECT 783.8800 268.4400 785.4800 268.9200 ;
        RECT 783.8800 273.8800 785.4800 274.3600 ;
        RECT 783.8800 279.3200 785.4800 279.8000 ;
        RECT 738.8800 268.4400 740.4800 268.9200 ;
        RECT 738.8800 273.8800 740.4800 274.3600 ;
        RECT 738.8800 279.3200 740.4800 279.8000 ;
        RECT 783.8800 257.5600 785.4800 258.0400 ;
        RECT 783.8800 263.0000 785.4800 263.4800 ;
        RECT 783.8800 241.2400 785.4800 241.7200 ;
        RECT 783.8800 246.6800 785.4800 247.1600 ;
        RECT 783.8800 252.1200 785.4800 252.6000 ;
        RECT 738.8800 257.5600 740.4800 258.0400 ;
        RECT 738.8800 263.0000 740.4800 263.4800 ;
        RECT 738.8800 241.2400 740.4800 241.7200 ;
        RECT 738.8800 246.6800 740.4800 247.1600 ;
        RECT 738.8800 252.1200 740.4800 252.6000 ;
        RECT 693.8800 268.4400 695.4800 268.9200 ;
        RECT 693.8800 273.8800 695.4800 274.3600 ;
        RECT 682.1200 273.8800 685.1200 274.3600 ;
        RECT 682.1200 268.4400 685.1200 268.9200 ;
        RECT 682.1200 279.3200 685.1200 279.8000 ;
        RECT 693.8800 279.3200 695.4800 279.8000 ;
        RECT 693.8800 257.5600 695.4800 258.0400 ;
        RECT 693.8800 263.0000 695.4800 263.4800 ;
        RECT 682.1200 263.0000 685.1200 263.4800 ;
        RECT 682.1200 257.5600 685.1200 258.0400 ;
        RECT 693.8800 241.2400 695.4800 241.7200 ;
        RECT 693.8800 246.6800 695.4800 247.1600 ;
        RECT 682.1200 246.6800 685.1200 247.1600 ;
        RECT 682.1200 241.2400 685.1200 241.7200 ;
        RECT 682.1200 252.1200 685.1200 252.6000 ;
        RECT 693.8800 252.1200 695.4800 252.6000 ;
        RECT 783.8800 224.9200 785.4800 225.4000 ;
        RECT 783.8800 230.3600 785.4800 230.8400 ;
        RECT 783.8800 235.8000 785.4800 236.2800 ;
        RECT 783.8800 214.0400 785.4800 214.5200 ;
        RECT 783.8800 219.4800 785.4800 219.9600 ;
        RECT 738.8800 224.9200 740.4800 225.4000 ;
        RECT 738.8800 230.3600 740.4800 230.8400 ;
        RECT 738.8800 235.8000 740.4800 236.2800 ;
        RECT 738.8800 214.0400 740.4800 214.5200 ;
        RECT 738.8800 219.4800 740.4800 219.9600 ;
        RECT 783.8800 197.7200 785.4800 198.2000 ;
        RECT 783.8800 203.1600 785.4800 203.6400 ;
        RECT 783.8800 208.6000 785.4800 209.0800 ;
        RECT 783.8800 186.8400 785.4800 187.3200 ;
        RECT 783.8800 192.2800 785.4800 192.7600 ;
        RECT 738.8800 197.7200 740.4800 198.2000 ;
        RECT 738.8800 203.1600 740.4800 203.6400 ;
        RECT 738.8800 208.6000 740.4800 209.0800 ;
        RECT 738.8800 186.8400 740.4800 187.3200 ;
        RECT 738.8800 192.2800 740.4800 192.7600 ;
        RECT 693.8800 224.9200 695.4800 225.4000 ;
        RECT 693.8800 230.3600 695.4800 230.8400 ;
        RECT 693.8800 235.8000 695.4800 236.2800 ;
        RECT 682.1200 224.9200 685.1200 225.4000 ;
        RECT 682.1200 230.3600 685.1200 230.8400 ;
        RECT 682.1200 235.8000 685.1200 236.2800 ;
        RECT 693.8800 214.0400 695.4800 214.5200 ;
        RECT 693.8800 219.4800 695.4800 219.9600 ;
        RECT 682.1200 214.0400 685.1200 214.5200 ;
        RECT 682.1200 219.4800 685.1200 219.9600 ;
        RECT 693.8800 197.7200 695.4800 198.2000 ;
        RECT 693.8800 203.1600 695.4800 203.6400 ;
        RECT 693.8800 208.6000 695.4800 209.0800 ;
        RECT 682.1200 197.7200 685.1200 198.2000 ;
        RECT 682.1200 203.1600 685.1200 203.6400 ;
        RECT 682.1200 208.6000 685.1200 209.0800 ;
        RECT 693.8800 186.8400 695.4800 187.3200 ;
        RECT 693.8800 192.2800 695.4800 192.7600 ;
        RECT 682.1200 186.8400 685.1200 187.3200 ;
        RECT 682.1200 192.2800 685.1200 192.7600 ;
        RECT 886.2200 170.5200 889.2200 171.0000 ;
        RECT 886.2200 175.9600 889.2200 176.4400 ;
        RECT 886.2200 181.4000 889.2200 181.8800 ;
        RECT 873.8800 170.5200 875.4800 171.0000 ;
        RECT 873.8800 175.9600 875.4800 176.4400 ;
        RECT 873.8800 181.4000 875.4800 181.8800 ;
        RECT 886.2200 159.6400 889.2200 160.1200 ;
        RECT 886.2200 165.0800 889.2200 165.5600 ;
        RECT 873.8800 159.6400 875.4800 160.1200 ;
        RECT 873.8800 165.0800 875.4800 165.5600 ;
        RECT 886.2200 143.3200 889.2200 143.8000 ;
        RECT 886.2200 148.7600 889.2200 149.2400 ;
        RECT 886.2200 154.2000 889.2200 154.6800 ;
        RECT 873.8800 143.3200 875.4800 143.8000 ;
        RECT 873.8800 148.7600 875.4800 149.2400 ;
        RECT 873.8800 154.2000 875.4800 154.6800 ;
        RECT 886.2200 132.4400 889.2200 132.9200 ;
        RECT 886.2200 137.8800 889.2200 138.3600 ;
        RECT 873.8800 132.4400 875.4800 132.9200 ;
        RECT 873.8800 137.8800 875.4800 138.3600 ;
        RECT 828.8800 170.5200 830.4800 171.0000 ;
        RECT 828.8800 175.9600 830.4800 176.4400 ;
        RECT 828.8800 181.4000 830.4800 181.8800 ;
        RECT 828.8800 159.6400 830.4800 160.1200 ;
        RECT 828.8800 165.0800 830.4800 165.5600 ;
        RECT 828.8800 143.3200 830.4800 143.8000 ;
        RECT 828.8800 148.7600 830.4800 149.2400 ;
        RECT 828.8800 154.2000 830.4800 154.6800 ;
        RECT 828.8800 132.4400 830.4800 132.9200 ;
        RECT 828.8800 137.8800 830.4800 138.3600 ;
        RECT 886.2200 116.1200 889.2200 116.6000 ;
        RECT 886.2200 121.5600 889.2200 122.0400 ;
        RECT 886.2200 127.0000 889.2200 127.4800 ;
        RECT 873.8800 116.1200 875.4800 116.6000 ;
        RECT 873.8800 121.5600 875.4800 122.0400 ;
        RECT 873.8800 127.0000 875.4800 127.4800 ;
        RECT 886.2200 105.2400 889.2200 105.7200 ;
        RECT 886.2200 110.6800 889.2200 111.1600 ;
        RECT 873.8800 105.2400 875.4800 105.7200 ;
        RECT 873.8800 110.6800 875.4800 111.1600 ;
        RECT 886.2200 88.9200 889.2200 89.4000 ;
        RECT 886.2200 94.3600 889.2200 94.8400 ;
        RECT 886.2200 99.8000 889.2200 100.2800 ;
        RECT 873.8800 88.9200 875.4800 89.4000 ;
        RECT 873.8800 94.3600 875.4800 94.8400 ;
        RECT 873.8800 99.8000 875.4800 100.2800 ;
        RECT 886.2200 83.4800 889.2200 83.9600 ;
        RECT 873.8800 83.4800 875.4800 83.9600 ;
        RECT 828.8800 116.1200 830.4800 116.6000 ;
        RECT 828.8800 121.5600 830.4800 122.0400 ;
        RECT 828.8800 127.0000 830.4800 127.4800 ;
        RECT 828.8800 105.2400 830.4800 105.7200 ;
        RECT 828.8800 110.6800 830.4800 111.1600 ;
        RECT 828.8800 88.9200 830.4800 89.4000 ;
        RECT 828.8800 94.3600 830.4800 94.8400 ;
        RECT 828.8800 99.8000 830.4800 100.2800 ;
        RECT 828.8800 83.4800 830.4800 83.9600 ;
        RECT 783.8800 170.5200 785.4800 171.0000 ;
        RECT 783.8800 175.9600 785.4800 176.4400 ;
        RECT 783.8800 181.4000 785.4800 181.8800 ;
        RECT 783.8800 159.6400 785.4800 160.1200 ;
        RECT 783.8800 165.0800 785.4800 165.5600 ;
        RECT 738.8800 170.5200 740.4800 171.0000 ;
        RECT 738.8800 175.9600 740.4800 176.4400 ;
        RECT 738.8800 181.4000 740.4800 181.8800 ;
        RECT 738.8800 159.6400 740.4800 160.1200 ;
        RECT 738.8800 165.0800 740.4800 165.5600 ;
        RECT 783.8800 143.3200 785.4800 143.8000 ;
        RECT 783.8800 148.7600 785.4800 149.2400 ;
        RECT 783.8800 154.2000 785.4800 154.6800 ;
        RECT 783.8800 132.4400 785.4800 132.9200 ;
        RECT 783.8800 137.8800 785.4800 138.3600 ;
        RECT 738.8800 143.3200 740.4800 143.8000 ;
        RECT 738.8800 148.7600 740.4800 149.2400 ;
        RECT 738.8800 154.2000 740.4800 154.6800 ;
        RECT 738.8800 132.4400 740.4800 132.9200 ;
        RECT 738.8800 137.8800 740.4800 138.3600 ;
        RECT 693.8800 170.5200 695.4800 171.0000 ;
        RECT 693.8800 175.9600 695.4800 176.4400 ;
        RECT 693.8800 181.4000 695.4800 181.8800 ;
        RECT 682.1200 170.5200 685.1200 171.0000 ;
        RECT 682.1200 175.9600 685.1200 176.4400 ;
        RECT 682.1200 181.4000 685.1200 181.8800 ;
        RECT 693.8800 159.6400 695.4800 160.1200 ;
        RECT 693.8800 165.0800 695.4800 165.5600 ;
        RECT 682.1200 159.6400 685.1200 160.1200 ;
        RECT 682.1200 165.0800 685.1200 165.5600 ;
        RECT 693.8800 143.3200 695.4800 143.8000 ;
        RECT 693.8800 148.7600 695.4800 149.2400 ;
        RECT 693.8800 154.2000 695.4800 154.6800 ;
        RECT 682.1200 143.3200 685.1200 143.8000 ;
        RECT 682.1200 148.7600 685.1200 149.2400 ;
        RECT 682.1200 154.2000 685.1200 154.6800 ;
        RECT 693.8800 132.4400 695.4800 132.9200 ;
        RECT 693.8800 137.8800 695.4800 138.3600 ;
        RECT 682.1200 132.4400 685.1200 132.9200 ;
        RECT 682.1200 137.8800 685.1200 138.3600 ;
        RECT 783.8800 116.1200 785.4800 116.6000 ;
        RECT 783.8800 121.5600 785.4800 122.0400 ;
        RECT 783.8800 127.0000 785.4800 127.4800 ;
        RECT 783.8800 105.2400 785.4800 105.7200 ;
        RECT 783.8800 110.6800 785.4800 111.1600 ;
        RECT 738.8800 116.1200 740.4800 116.6000 ;
        RECT 738.8800 121.5600 740.4800 122.0400 ;
        RECT 738.8800 127.0000 740.4800 127.4800 ;
        RECT 738.8800 105.2400 740.4800 105.7200 ;
        RECT 738.8800 110.6800 740.4800 111.1600 ;
        RECT 783.8800 88.9200 785.4800 89.4000 ;
        RECT 783.8800 94.3600 785.4800 94.8400 ;
        RECT 783.8800 99.8000 785.4800 100.2800 ;
        RECT 783.8800 83.4800 785.4800 83.9600 ;
        RECT 738.8800 88.9200 740.4800 89.4000 ;
        RECT 738.8800 94.3600 740.4800 94.8400 ;
        RECT 738.8800 99.8000 740.4800 100.2800 ;
        RECT 738.8800 83.4800 740.4800 83.9600 ;
        RECT 693.8800 116.1200 695.4800 116.6000 ;
        RECT 693.8800 121.5600 695.4800 122.0400 ;
        RECT 693.8800 127.0000 695.4800 127.4800 ;
        RECT 682.1200 116.1200 685.1200 116.6000 ;
        RECT 682.1200 121.5600 685.1200 122.0400 ;
        RECT 682.1200 127.0000 685.1200 127.4800 ;
        RECT 693.8800 105.2400 695.4800 105.7200 ;
        RECT 693.8800 110.6800 695.4800 111.1600 ;
        RECT 682.1200 105.2400 685.1200 105.7200 ;
        RECT 682.1200 110.6800 685.1200 111.1600 ;
        RECT 693.8800 88.9200 695.4800 89.4000 ;
        RECT 693.8800 94.3600 695.4800 94.8400 ;
        RECT 693.8800 99.8000 695.4800 100.2800 ;
        RECT 682.1200 88.9200 685.1200 89.4000 ;
        RECT 682.1200 94.3600 685.1200 94.8400 ;
        RECT 682.1200 99.8000 685.1200 100.2800 ;
        RECT 682.1200 83.4800 685.1200 83.9600 ;
        RECT 693.8800 83.4800 695.4800 83.9600 ;
        RECT 682.1200 288.3900 889.2200 291.3900 ;
        RECT 682.1200 75.2900 889.2200 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 683.1200 34.6700 685.1200 61.6000 ;
        RECT 886.2200 34.6700 888.2200 61.6000 ;
      LAYER met3 ;
        RECT 886.2200 51.3800 888.2200 51.8600 ;
        RECT 683.1200 51.3800 685.1200 51.8600 ;
        RECT 886.2200 45.9400 888.2200 46.4200 ;
        RECT 886.2200 40.5000 888.2200 40.9800 ;
        RECT 683.1200 45.9400 685.1200 46.4200 ;
        RECT 683.1200 40.5000 685.1200 40.9800 ;
        RECT 683.1200 59.6000 888.2200 61.6000 ;
        RECT 683.1200 34.6700 888.2200 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 2601.3300 875.4800 2817.4300 ;
        RECT 828.8800 2601.3300 830.4800 2817.4300 ;
        RECT 783.8800 2601.3300 785.4800 2817.4300 ;
        RECT 738.8800 2601.3300 740.4800 2817.4300 ;
        RECT 693.8800 2601.3300 695.4800 2817.4300 ;
        RECT 886.2200 2601.3300 889.2200 2817.4300 ;
        RECT 682.1200 2601.3300 685.1200 2817.4300 ;
      LAYER met3 ;
        RECT 886.2200 2794.4800 889.2200 2794.9600 ;
        RECT 886.2200 2799.9200 889.2200 2800.4000 ;
        RECT 873.8800 2794.4800 875.4800 2794.9600 ;
        RECT 873.8800 2799.9200 875.4800 2800.4000 ;
        RECT 886.2200 2805.3600 889.2200 2805.8400 ;
        RECT 873.8800 2805.3600 875.4800 2805.8400 ;
        RECT 886.2200 2783.6000 889.2200 2784.0800 ;
        RECT 886.2200 2789.0400 889.2200 2789.5200 ;
        RECT 873.8800 2783.6000 875.4800 2784.0800 ;
        RECT 873.8800 2789.0400 875.4800 2789.5200 ;
        RECT 886.2200 2767.2800 889.2200 2767.7600 ;
        RECT 886.2200 2772.7200 889.2200 2773.2000 ;
        RECT 873.8800 2767.2800 875.4800 2767.7600 ;
        RECT 873.8800 2772.7200 875.4800 2773.2000 ;
        RECT 886.2200 2778.1600 889.2200 2778.6400 ;
        RECT 873.8800 2778.1600 875.4800 2778.6400 ;
        RECT 828.8800 2794.4800 830.4800 2794.9600 ;
        RECT 828.8800 2799.9200 830.4800 2800.4000 ;
        RECT 828.8800 2805.3600 830.4800 2805.8400 ;
        RECT 828.8800 2783.6000 830.4800 2784.0800 ;
        RECT 828.8800 2789.0400 830.4800 2789.5200 ;
        RECT 828.8800 2767.2800 830.4800 2767.7600 ;
        RECT 828.8800 2772.7200 830.4800 2773.2000 ;
        RECT 828.8800 2778.1600 830.4800 2778.6400 ;
        RECT 886.2200 2750.9600 889.2200 2751.4400 ;
        RECT 886.2200 2756.4000 889.2200 2756.8800 ;
        RECT 886.2200 2761.8400 889.2200 2762.3200 ;
        RECT 873.8800 2750.9600 875.4800 2751.4400 ;
        RECT 873.8800 2756.4000 875.4800 2756.8800 ;
        RECT 873.8800 2761.8400 875.4800 2762.3200 ;
        RECT 886.2200 2740.0800 889.2200 2740.5600 ;
        RECT 886.2200 2745.5200 889.2200 2746.0000 ;
        RECT 873.8800 2740.0800 875.4800 2740.5600 ;
        RECT 873.8800 2745.5200 875.4800 2746.0000 ;
        RECT 886.2200 2723.7600 889.2200 2724.2400 ;
        RECT 886.2200 2729.2000 889.2200 2729.6800 ;
        RECT 886.2200 2734.6400 889.2200 2735.1200 ;
        RECT 873.8800 2723.7600 875.4800 2724.2400 ;
        RECT 873.8800 2729.2000 875.4800 2729.6800 ;
        RECT 873.8800 2734.6400 875.4800 2735.1200 ;
        RECT 886.2200 2712.8800 889.2200 2713.3600 ;
        RECT 886.2200 2718.3200 889.2200 2718.8000 ;
        RECT 873.8800 2712.8800 875.4800 2713.3600 ;
        RECT 873.8800 2718.3200 875.4800 2718.8000 ;
        RECT 828.8800 2750.9600 830.4800 2751.4400 ;
        RECT 828.8800 2756.4000 830.4800 2756.8800 ;
        RECT 828.8800 2761.8400 830.4800 2762.3200 ;
        RECT 828.8800 2740.0800 830.4800 2740.5600 ;
        RECT 828.8800 2745.5200 830.4800 2746.0000 ;
        RECT 828.8800 2723.7600 830.4800 2724.2400 ;
        RECT 828.8800 2729.2000 830.4800 2729.6800 ;
        RECT 828.8800 2734.6400 830.4800 2735.1200 ;
        RECT 828.8800 2712.8800 830.4800 2713.3600 ;
        RECT 828.8800 2718.3200 830.4800 2718.8000 ;
        RECT 783.8800 2794.4800 785.4800 2794.9600 ;
        RECT 783.8800 2799.9200 785.4800 2800.4000 ;
        RECT 783.8800 2805.3600 785.4800 2805.8400 ;
        RECT 738.8800 2794.4800 740.4800 2794.9600 ;
        RECT 738.8800 2799.9200 740.4800 2800.4000 ;
        RECT 738.8800 2805.3600 740.4800 2805.8400 ;
        RECT 783.8800 2783.6000 785.4800 2784.0800 ;
        RECT 783.8800 2789.0400 785.4800 2789.5200 ;
        RECT 783.8800 2767.2800 785.4800 2767.7600 ;
        RECT 783.8800 2772.7200 785.4800 2773.2000 ;
        RECT 783.8800 2778.1600 785.4800 2778.6400 ;
        RECT 738.8800 2783.6000 740.4800 2784.0800 ;
        RECT 738.8800 2789.0400 740.4800 2789.5200 ;
        RECT 738.8800 2767.2800 740.4800 2767.7600 ;
        RECT 738.8800 2772.7200 740.4800 2773.2000 ;
        RECT 738.8800 2778.1600 740.4800 2778.6400 ;
        RECT 693.8800 2794.4800 695.4800 2794.9600 ;
        RECT 693.8800 2799.9200 695.4800 2800.4000 ;
        RECT 682.1200 2799.9200 685.1200 2800.4000 ;
        RECT 682.1200 2794.4800 685.1200 2794.9600 ;
        RECT 682.1200 2805.3600 685.1200 2805.8400 ;
        RECT 693.8800 2805.3600 695.4800 2805.8400 ;
        RECT 693.8800 2783.6000 695.4800 2784.0800 ;
        RECT 693.8800 2789.0400 695.4800 2789.5200 ;
        RECT 682.1200 2789.0400 685.1200 2789.5200 ;
        RECT 682.1200 2783.6000 685.1200 2784.0800 ;
        RECT 693.8800 2767.2800 695.4800 2767.7600 ;
        RECT 693.8800 2772.7200 695.4800 2773.2000 ;
        RECT 682.1200 2772.7200 685.1200 2773.2000 ;
        RECT 682.1200 2767.2800 685.1200 2767.7600 ;
        RECT 682.1200 2778.1600 685.1200 2778.6400 ;
        RECT 693.8800 2778.1600 695.4800 2778.6400 ;
        RECT 783.8800 2750.9600 785.4800 2751.4400 ;
        RECT 783.8800 2756.4000 785.4800 2756.8800 ;
        RECT 783.8800 2761.8400 785.4800 2762.3200 ;
        RECT 783.8800 2740.0800 785.4800 2740.5600 ;
        RECT 783.8800 2745.5200 785.4800 2746.0000 ;
        RECT 738.8800 2750.9600 740.4800 2751.4400 ;
        RECT 738.8800 2756.4000 740.4800 2756.8800 ;
        RECT 738.8800 2761.8400 740.4800 2762.3200 ;
        RECT 738.8800 2740.0800 740.4800 2740.5600 ;
        RECT 738.8800 2745.5200 740.4800 2746.0000 ;
        RECT 783.8800 2723.7600 785.4800 2724.2400 ;
        RECT 783.8800 2729.2000 785.4800 2729.6800 ;
        RECT 783.8800 2734.6400 785.4800 2735.1200 ;
        RECT 783.8800 2712.8800 785.4800 2713.3600 ;
        RECT 783.8800 2718.3200 785.4800 2718.8000 ;
        RECT 738.8800 2723.7600 740.4800 2724.2400 ;
        RECT 738.8800 2729.2000 740.4800 2729.6800 ;
        RECT 738.8800 2734.6400 740.4800 2735.1200 ;
        RECT 738.8800 2712.8800 740.4800 2713.3600 ;
        RECT 738.8800 2718.3200 740.4800 2718.8000 ;
        RECT 693.8800 2750.9600 695.4800 2751.4400 ;
        RECT 693.8800 2756.4000 695.4800 2756.8800 ;
        RECT 693.8800 2761.8400 695.4800 2762.3200 ;
        RECT 682.1200 2750.9600 685.1200 2751.4400 ;
        RECT 682.1200 2756.4000 685.1200 2756.8800 ;
        RECT 682.1200 2761.8400 685.1200 2762.3200 ;
        RECT 693.8800 2740.0800 695.4800 2740.5600 ;
        RECT 693.8800 2745.5200 695.4800 2746.0000 ;
        RECT 682.1200 2740.0800 685.1200 2740.5600 ;
        RECT 682.1200 2745.5200 685.1200 2746.0000 ;
        RECT 693.8800 2723.7600 695.4800 2724.2400 ;
        RECT 693.8800 2729.2000 695.4800 2729.6800 ;
        RECT 693.8800 2734.6400 695.4800 2735.1200 ;
        RECT 682.1200 2723.7600 685.1200 2724.2400 ;
        RECT 682.1200 2729.2000 685.1200 2729.6800 ;
        RECT 682.1200 2734.6400 685.1200 2735.1200 ;
        RECT 693.8800 2712.8800 695.4800 2713.3600 ;
        RECT 693.8800 2718.3200 695.4800 2718.8000 ;
        RECT 682.1200 2712.8800 685.1200 2713.3600 ;
        RECT 682.1200 2718.3200 685.1200 2718.8000 ;
        RECT 886.2200 2696.5600 889.2200 2697.0400 ;
        RECT 886.2200 2702.0000 889.2200 2702.4800 ;
        RECT 886.2200 2707.4400 889.2200 2707.9200 ;
        RECT 873.8800 2696.5600 875.4800 2697.0400 ;
        RECT 873.8800 2702.0000 875.4800 2702.4800 ;
        RECT 873.8800 2707.4400 875.4800 2707.9200 ;
        RECT 886.2200 2685.6800 889.2200 2686.1600 ;
        RECT 886.2200 2691.1200 889.2200 2691.6000 ;
        RECT 873.8800 2685.6800 875.4800 2686.1600 ;
        RECT 873.8800 2691.1200 875.4800 2691.6000 ;
        RECT 886.2200 2669.3600 889.2200 2669.8400 ;
        RECT 886.2200 2674.8000 889.2200 2675.2800 ;
        RECT 886.2200 2680.2400 889.2200 2680.7200 ;
        RECT 873.8800 2669.3600 875.4800 2669.8400 ;
        RECT 873.8800 2674.8000 875.4800 2675.2800 ;
        RECT 873.8800 2680.2400 875.4800 2680.7200 ;
        RECT 886.2200 2658.4800 889.2200 2658.9600 ;
        RECT 886.2200 2663.9200 889.2200 2664.4000 ;
        RECT 873.8800 2658.4800 875.4800 2658.9600 ;
        RECT 873.8800 2663.9200 875.4800 2664.4000 ;
        RECT 828.8800 2696.5600 830.4800 2697.0400 ;
        RECT 828.8800 2702.0000 830.4800 2702.4800 ;
        RECT 828.8800 2707.4400 830.4800 2707.9200 ;
        RECT 828.8800 2685.6800 830.4800 2686.1600 ;
        RECT 828.8800 2691.1200 830.4800 2691.6000 ;
        RECT 828.8800 2669.3600 830.4800 2669.8400 ;
        RECT 828.8800 2674.8000 830.4800 2675.2800 ;
        RECT 828.8800 2680.2400 830.4800 2680.7200 ;
        RECT 828.8800 2658.4800 830.4800 2658.9600 ;
        RECT 828.8800 2663.9200 830.4800 2664.4000 ;
        RECT 886.2200 2642.1600 889.2200 2642.6400 ;
        RECT 886.2200 2647.6000 889.2200 2648.0800 ;
        RECT 886.2200 2653.0400 889.2200 2653.5200 ;
        RECT 873.8800 2642.1600 875.4800 2642.6400 ;
        RECT 873.8800 2647.6000 875.4800 2648.0800 ;
        RECT 873.8800 2653.0400 875.4800 2653.5200 ;
        RECT 886.2200 2631.2800 889.2200 2631.7600 ;
        RECT 886.2200 2636.7200 889.2200 2637.2000 ;
        RECT 873.8800 2631.2800 875.4800 2631.7600 ;
        RECT 873.8800 2636.7200 875.4800 2637.2000 ;
        RECT 886.2200 2614.9600 889.2200 2615.4400 ;
        RECT 886.2200 2620.4000 889.2200 2620.8800 ;
        RECT 886.2200 2625.8400 889.2200 2626.3200 ;
        RECT 873.8800 2614.9600 875.4800 2615.4400 ;
        RECT 873.8800 2620.4000 875.4800 2620.8800 ;
        RECT 873.8800 2625.8400 875.4800 2626.3200 ;
        RECT 886.2200 2609.5200 889.2200 2610.0000 ;
        RECT 873.8800 2609.5200 875.4800 2610.0000 ;
        RECT 828.8800 2642.1600 830.4800 2642.6400 ;
        RECT 828.8800 2647.6000 830.4800 2648.0800 ;
        RECT 828.8800 2653.0400 830.4800 2653.5200 ;
        RECT 828.8800 2631.2800 830.4800 2631.7600 ;
        RECT 828.8800 2636.7200 830.4800 2637.2000 ;
        RECT 828.8800 2614.9600 830.4800 2615.4400 ;
        RECT 828.8800 2620.4000 830.4800 2620.8800 ;
        RECT 828.8800 2625.8400 830.4800 2626.3200 ;
        RECT 828.8800 2609.5200 830.4800 2610.0000 ;
        RECT 783.8800 2696.5600 785.4800 2697.0400 ;
        RECT 783.8800 2702.0000 785.4800 2702.4800 ;
        RECT 783.8800 2707.4400 785.4800 2707.9200 ;
        RECT 783.8800 2685.6800 785.4800 2686.1600 ;
        RECT 783.8800 2691.1200 785.4800 2691.6000 ;
        RECT 738.8800 2696.5600 740.4800 2697.0400 ;
        RECT 738.8800 2702.0000 740.4800 2702.4800 ;
        RECT 738.8800 2707.4400 740.4800 2707.9200 ;
        RECT 738.8800 2685.6800 740.4800 2686.1600 ;
        RECT 738.8800 2691.1200 740.4800 2691.6000 ;
        RECT 783.8800 2669.3600 785.4800 2669.8400 ;
        RECT 783.8800 2674.8000 785.4800 2675.2800 ;
        RECT 783.8800 2680.2400 785.4800 2680.7200 ;
        RECT 783.8800 2658.4800 785.4800 2658.9600 ;
        RECT 783.8800 2663.9200 785.4800 2664.4000 ;
        RECT 738.8800 2669.3600 740.4800 2669.8400 ;
        RECT 738.8800 2674.8000 740.4800 2675.2800 ;
        RECT 738.8800 2680.2400 740.4800 2680.7200 ;
        RECT 738.8800 2658.4800 740.4800 2658.9600 ;
        RECT 738.8800 2663.9200 740.4800 2664.4000 ;
        RECT 693.8800 2696.5600 695.4800 2697.0400 ;
        RECT 693.8800 2702.0000 695.4800 2702.4800 ;
        RECT 693.8800 2707.4400 695.4800 2707.9200 ;
        RECT 682.1200 2696.5600 685.1200 2697.0400 ;
        RECT 682.1200 2702.0000 685.1200 2702.4800 ;
        RECT 682.1200 2707.4400 685.1200 2707.9200 ;
        RECT 693.8800 2685.6800 695.4800 2686.1600 ;
        RECT 693.8800 2691.1200 695.4800 2691.6000 ;
        RECT 682.1200 2685.6800 685.1200 2686.1600 ;
        RECT 682.1200 2691.1200 685.1200 2691.6000 ;
        RECT 693.8800 2669.3600 695.4800 2669.8400 ;
        RECT 693.8800 2674.8000 695.4800 2675.2800 ;
        RECT 693.8800 2680.2400 695.4800 2680.7200 ;
        RECT 682.1200 2669.3600 685.1200 2669.8400 ;
        RECT 682.1200 2674.8000 685.1200 2675.2800 ;
        RECT 682.1200 2680.2400 685.1200 2680.7200 ;
        RECT 693.8800 2658.4800 695.4800 2658.9600 ;
        RECT 693.8800 2663.9200 695.4800 2664.4000 ;
        RECT 682.1200 2658.4800 685.1200 2658.9600 ;
        RECT 682.1200 2663.9200 685.1200 2664.4000 ;
        RECT 783.8800 2642.1600 785.4800 2642.6400 ;
        RECT 783.8800 2647.6000 785.4800 2648.0800 ;
        RECT 783.8800 2653.0400 785.4800 2653.5200 ;
        RECT 783.8800 2631.2800 785.4800 2631.7600 ;
        RECT 783.8800 2636.7200 785.4800 2637.2000 ;
        RECT 738.8800 2642.1600 740.4800 2642.6400 ;
        RECT 738.8800 2647.6000 740.4800 2648.0800 ;
        RECT 738.8800 2653.0400 740.4800 2653.5200 ;
        RECT 738.8800 2631.2800 740.4800 2631.7600 ;
        RECT 738.8800 2636.7200 740.4800 2637.2000 ;
        RECT 783.8800 2614.9600 785.4800 2615.4400 ;
        RECT 783.8800 2620.4000 785.4800 2620.8800 ;
        RECT 783.8800 2625.8400 785.4800 2626.3200 ;
        RECT 783.8800 2609.5200 785.4800 2610.0000 ;
        RECT 738.8800 2614.9600 740.4800 2615.4400 ;
        RECT 738.8800 2620.4000 740.4800 2620.8800 ;
        RECT 738.8800 2625.8400 740.4800 2626.3200 ;
        RECT 738.8800 2609.5200 740.4800 2610.0000 ;
        RECT 693.8800 2642.1600 695.4800 2642.6400 ;
        RECT 693.8800 2647.6000 695.4800 2648.0800 ;
        RECT 693.8800 2653.0400 695.4800 2653.5200 ;
        RECT 682.1200 2642.1600 685.1200 2642.6400 ;
        RECT 682.1200 2647.6000 685.1200 2648.0800 ;
        RECT 682.1200 2653.0400 685.1200 2653.5200 ;
        RECT 693.8800 2631.2800 695.4800 2631.7600 ;
        RECT 693.8800 2636.7200 695.4800 2637.2000 ;
        RECT 682.1200 2631.2800 685.1200 2631.7600 ;
        RECT 682.1200 2636.7200 685.1200 2637.2000 ;
        RECT 693.8800 2614.9600 695.4800 2615.4400 ;
        RECT 693.8800 2620.4000 695.4800 2620.8800 ;
        RECT 693.8800 2625.8400 695.4800 2626.3200 ;
        RECT 682.1200 2614.9600 685.1200 2615.4400 ;
        RECT 682.1200 2620.4000 685.1200 2620.8800 ;
        RECT 682.1200 2625.8400 685.1200 2626.3200 ;
        RECT 682.1200 2609.5200 685.1200 2610.0000 ;
        RECT 693.8800 2609.5200 695.4800 2610.0000 ;
        RECT 682.1200 2814.4300 889.2200 2817.4300 ;
        RECT 682.1200 2601.3300 889.2200 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 2371.6900 875.4800 2587.7900 ;
        RECT 828.8800 2371.6900 830.4800 2587.7900 ;
        RECT 783.8800 2371.6900 785.4800 2587.7900 ;
        RECT 738.8800 2371.6900 740.4800 2587.7900 ;
        RECT 693.8800 2371.6900 695.4800 2587.7900 ;
        RECT 886.2200 2371.6900 889.2200 2587.7900 ;
        RECT 682.1200 2371.6900 685.1200 2587.7900 ;
      LAYER met3 ;
        RECT 886.2200 2564.8400 889.2200 2565.3200 ;
        RECT 886.2200 2570.2800 889.2200 2570.7600 ;
        RECT 873.8800 2564.8400 875.4800 2565.3200 ;
        RECT 873.8800 2570.2800 875.4800 2570.7600 ;
        RECT 886.2200 2575.7200 889.2200 2576.2000 ;
        RECT 873.8800 2575.7200 875.4800 2576.2000 ;
        RECT 886.2200 2553.9600 889.2200 2554.4400 ;
        RECT 886.2200 2559.4000 889.2200 2559.8800 ;
        RECT 873.8800 2553.9600 875.4800 2554.4400 ;
        RECT 873.8800 2559.4000 875.4800 2559.8800 ;
        RECT 886.2200 2537.6400 889.2200 2538.1200 ;
        RECT 886.2200 2543.0800 889.2200 2543.5600 ;
        RECT 873.8800 2537.6400 875.4800 2538.1200 ;
        RECT 873.8800 2543.0800 875.4800 2543.5600 ;
        RECT 886.2200 2548.5200 889.2200 2549.0000 ;
        RECT 873.8800 2548.5200 875.4800 2549.0000 ;
        RECT 828.8800 2564.8400 830.4800 2565.3200 ;
        RECT 828.8800 2570.2800 830.4800 2570.7600 ;
        RECT 828.8800 2575.7200 830.4800 2576.2000 ;
        RECT 828.8800 2553.9600 830.4800 2554.4400 ;
        RECT 828.8800 2559.4000 830.4800 2559.8800 ;
        RECT 828.8800 2537.6400 830.4800 2538.1200 ;
        RECT 828.8800 2543.0800 830.4800 2543.5600 ;
        RECT 828.8800 2548.5200 830.4800 2549.0000 ;
        RECT 886.2200 2521.3200 889.2200 2521.8000 ;
        RECT 886.2200 2526.7600 889.2200 2527.2400 ;
        RECT 886.2200 2532.2000 889.2200 2532.6800 ;
        RECT 873.8800 2521.3200 875.4800 2521.8000 ;
        RECT 873.8800 2526.7600 875.4800 2527.2400 ;
        RECT 873.8800 2532.2000 875.4800 2532.6800 ;
        RECT 886.2200 2510.4400 889.2200 2510.9200 ;
        RECT 886.2200 2515.8800 889.2200 2516.3600 ;
        RECT 873.8800 2510.4400 875.4800 2510.9200 ;
        RECT 873.8800 2515.8800 875.4800 2516.3600 ;
        RECT 886.2200 2494.1200 889.2200 2494.6000 ;
        RECT 886.2200 2499.5600 889.2200 2500.0400 ;
        RECT 886.2200 2505.0000 889.2200 2505.4800 ;
        RECT 873.8800 2494.1200 875.4800 2494.6000 ;
        RECT 873.8800 2499.5600 875.4800 2500.0400 ;
        RECT 873.8800 2505.0000 875.4800 2505.4800 ;
        RECT 886.2200 2483.2400 889.2200 2483.7200 ;
        RECT 886.2200 2488.6800 889.2200 2489.1600 ;
        RECT 873.8800 2483.2400 875.4800 2483.7200 ;
        RECT 873.8800 2488.6800 875.4800 2489.1600 ;
        RECT 828.8800 2521.3200 830.4800 2521.8000 ;
        RECT 828.8800 2526.7600 830.4800 2527.2400 ;
        RECT 828.8800 2532.2000 830.4800 2532.6800 ;
        RECT 828.8800 2510.4400 830.4800 2510.9200 ;
        RECT 828.8800 2515.8800 830.4800 2516.3600 ;
        RECT 828.8800 2494.1200 830.4800 2494.6000 ;
        RECT 828.8800 2499.5600 830.4800 2500.0400 ;
        RECT 828.8800 2505.0000 830.4800 2505.4800 ;
        RECT 828.8800 2483.2400 830.4800 2483.7200 ;
        RECT 828.8800 2488.6800 830.4800 2489.1600 ;
        RECT 783.8800 2564.8400 785.4800 2565.3200 ;
        RECT 783.8800 2570.2800 785.4800 2570.7600 ;
        RECT 783.8800 2575.7200 785.4800 2576.2000 ;
        RECT 738.8800 2564.8400 740.4800 2565.3200 ;
        RECT 738.8800 2570.2800 740.4800 2570.7600 ;
        RECT 738.8800 2575.7200 740.4800 2576.2000 ;
        RECT 783.8800 2553.9600 785.4800 2554.4400 ;
        RECT 783.8800 2559.4000 785.4800 2559.8800 ;
        RECT 783.8800 2537.6400 785.4800 2538.1200 ;
        RECT 783.8800 2543.0800 785.4800 2543.5600 ;
        RECT 783.8800 2548.5200 785.4800 2549.0000 ;
        RECT 738.8800 2553.9600 740.4800 2554.4400 ;
        RECT 738.8800 2559.4000 740.4800 2559.8800 ;
        RECT 738.8800 2537.6400 740.4800 2538.1200 ;
        RECT 738.8800 2543.0800 740.4800 2543.5600 ;
        RECT 738.8800 2548.5200 740.4800 2549.0000 ;
        RECT 693.8800 2564.8400 695.4800 2565.3200 ;
        RECT 693.8800 2570.2800 695.4800 2570.7600 ;
        RECT 682.1200 2570.2800 685.1200 2570.7600 ;
        RECT 682.1200 2564.8400 685.1200 2565.3200 ;
        RECT 682.1200 2575.7200 685.1200 2576.2000 ;
        RECT 693.8800 2575.7200 695.4800 2576.2000 ;
        RECT 693.8800 2553.9600 695.4800 2554.4400 ;
        RECT 693.8800 2559.4000 695.4800 2559.8800 ;
        RECT 682.1200 2559.4000 685.1200 2559.8800 ;
        RECT 682.1200 2553.9600 685.1200 2554.4400 ;
        RECT 693.8800 2537.6400 695.4800 2538.1200 ;
        RECT 693.8800 2543.0800 695.4800 2543.5600 ;
        RECT 682.1200 2543.0800 685.1200 2543.5600 ;
        RECT 682.1200 2537.6400 685.1200 2538.1200 ;
        RECT 682.1200 2548.5200 685.1200 2549.0000 ;
        RECT 693.8800 2548.5200 695.4800 2549.0000 ;
        RECT 783.8800 2521.3200 785.4800 2521.8000 ;
        RECT 783.8800 2526.7600 785.4800 2527.2400 ;
        RECT 783.8800 2532.2000 785.4800 2532.6800 ;
        RECT 783.8800 2510.4400 785.4800 2510.9200 ;
        RECT 783.8800 2515.8800 785.4800 2516.3600 ;
        RECT 738.8800 2521.3200 740.4800 2521.8000 ;
        RECT 738.8800 2526.7600 740.4800 2527.2400 ;
        RECT 738.8800 2532.2000 740.4800 2532.6800 ;
        RECT 738.8800 2510.4400 740.4800 2510.9200 ;
        RECT 738.8800 2515.8800 740.4800 2516.3600 ;
        RECT 783.8800 2494.1200 785.4800 2494.6000 ;
        RECT 783.8800 2499.5600 785.4800 2500.0400 ;
        RECT 783.8800 2505.0000 785.4800 2505.4800 ;
        RECT 783.8800 2483.2400 785.4800 2483.7200 ;
        RECT 783.8800 2488.6800 785.4800 2489.1600 ;
        RECT 738.8800 2494.1200 740.4800 2494.6000 ;
        RECT 738.8800 2499.5600 740.4800 2500.0400 ;
        RECT 738.8800 2505.0000 740.4800 2505.4800 ;
        RECT 738.8800 2483.2400 740.4800 2483.7200 ;
        RECT 738.8800 2488.6800 740.4800 2489.1600 ;
        RECT 693.8800 2521.3200 695.4800 2521.8000 ;
        RECT 693.8800 2526.7600 695.4800 2527.2400 ;
        RECT 693.8800 2532.2000 695.4800 2532.6800 ;
        RECT 682.1200 2521.3200 685.1200 2521.8000 ;
        RECT 682.1200 2526.7600 685.1200 2527.2400 ;
        RECT 682.1200 2532.2000 685.1200 2532.6800 ;
        RECT 693.8800 2510.4400 695.4800 2510.9200 ;
        RECT 693.8800 2515.8800 695.4800 2516.3600 ;
        RECT 682.1200 2510.4400 685.1200 2510.9200 ;
        RECT 682.1200 2515.8800 685.1200 2516.3600 ;
        RECT 693.8800 2494.1200 695.4800 2494.6000 ;
        RECT 693.8800 2499.5600 695.4800 2500.0400 ;
        RECT 693.8800 2505.0000 695.4800 2505.4800 ;
        RECT 682.1200 2494.1200 685.1200 2494.6000 ;
        RECT 682.1200 2499.5600 685.1200 2500.0400 ;
        RECT 682.1200 2505.0000 685.1200 2505.4800 ;
        RECT 693.8800 2483.2400 695.4800 2483.7200 ;
        RECT 693.8800 2488.6800 695.4800 2489.1600 ;
        RECT 682.1200 2483.2400 685.1200 2483.7200 ;
        RECT 682.1200 2488.6800 685.1200 2489.1600 ;
        RECT 886.2200 2466.9200 889.2200 2467.4000 ;
        RECT 886.2200 2472.3600 889.2200 2472.8400 ;
        RECT 886.2200 2477.8000 889.2200 2478.2800 ;
        RECT 873.8800 2466.9200 875.4800 2467.4000 ;
        RECT 873.8800 2472.3600 875.4800 2472.8400 ;
        RECT 873.8800 2477.8000 875.4800 2478.2800 ;
        RECT 886.2200 2456.0400 889.2200 2456.5200 ;
        RECT 886.2200 2461.4800 889.2200 2461.9600 ;
        RECT 873.8800 2456.0400 875.4800 2456.5200 ;
        RECT 873.8800 2461.4800 875.4800 2461.9600 ;
        RECT 886.2200 2439.7200 889.2200 2440.2000 ;
        RECT 886.2200 2445.1600 889.2200 2445.6400 ;
        RECT 886.2200 2450.6000 889.2200 2451.0800 ;
        RECT 873.8800 2439.7200 875.4800 2440.2000 ;
        RECT 873.8800 2445.1600 875.4800 2445.6400 ;
        RECT 873.8800 2450.6000 875.4800 2451.0800 ;
        RECT 886.2200 2428.8400 889.2200 2429.3200 ;
        RECT 886.2200 2434.2800 889.2200 2434.7600 ;
        RECT 873.8800 2428.8400 875.4800 2429.3200 ;
        RECT 873.8800 2434.2800 875.4800 2434.7600 ;
        RECT 828.8800 2466.9200 830.4800 2467.4000 ;
        RECT 828.8800 2472.3600 830.4800 2472.8400 ;
        RECT 828.8800 2477.8000 830.4800 2478.2800 ;
        RECT 828.8800 2456.0400 830.4800 2456.5200 ;
        RECT 828.8800 2461.4800 830.4800 2461.9600 ;
        RECT 828.8800 2439.7200 830.4800 2440.2000 ;
        RECT 828.8800 2445.1600 830.4800 2445.6400 ;
        RECT 828.8800 2450.6000 830.4800 2451.0800 ;
        RECT 828.8800 2428.8400 830.4800 2429.3200 ;
        RECT 828.8800 2434.2800 830.4800 2434.7600 ;
        RECT 886.2200 2412.5200 889.2200 2413.0000 ;
        RECT 886.2200 2417.9600 889.2200 2418.4400 ;
        RECT 886.2200 2423.4000 889.2200 2423.8800 ;
        RECT 873.8800 2412.5200 875.4800 2413.0000 ;
        RECT 873.8800 2417.9600 875.4800 2418.4400 ;
        RECT 873.8800 2423.4000 875.4800 2423.8800 ;
        RECT 886.2200 2401.6400 889.2200 2402.1200 ;
        RECT 886.2200 2407.0800 889.2200 2407.5600 ;
        RECT 873.8800 2401.6400 875.4800 2402.1200 ;
        RECT 873.8800 2407.0800 875.4800 2407.5600 ;
        RECT 886.2200 2385.3200 889.2200 2385.8000 ;
        RECT 886.2200 2390.7600 889.2200 2391.2400 ;
        RECT 886.2200 2396.2000 889.2200 2396.6800 ;
        RECT 873.8800 2385.3200 875.4800 2385.8000 ;
        RECT 873.8800 2390.7600 875.4800 2391.2400 ;
        RECT 873.8800 2396.2000 875.4800 2396.6800 ;
        RECT 886.2200 2379.8800 889.2200 2380.3600 ;
        RECT 873.8800 2379.8800 875.4800 2380.3600 ;
        RECT 828.8800 2412.5200 830.4800 2413.0000 ;
        RECT 828.8800 2417.9600 830.4800 2418.4400 ;
        RECT 828.8800 2423.4000 830.4800 2423.8800 ;
        RECT 828.8800 2401.6400 830.4800 2402.1200 ;
        RECT 828.8800 2407.0800 830.4800 2407.5600 ;
        RECT 828.8800 2385.3200 830.4800 2385.8000 ;
        RECT 828.8800 2390.7600 830.4800 2391.2400 ;
        RECT 828.8800 2396.2000 830.4800 2396.6800 ;
        RECT 828.8800 2379.8800 830.4800 2380.3600 ;
        RECT 783.8800 2466.9200 785.4800 2467.4000 ;
        RECT 783.8800 2472.3600 785.4800 2472.8400 ;
        RECT 783.8800 2477.8000 785.4800 2478.2800 ;
        RECT 783.8800 2456.0400 785.4800 2456.5200 ;
        RECT 783.8800 2461.4800 785.4800 2461.9600 ;
        RECT 738.8800 2466.9200 740.4800 2467.4000 ;
        RECT 738.8800 2472.3600 740.4800 2472.8400 ;
        RECT 738.8800 2477.8000 740.4800 2478.2800 ;
        RECT 738.8800 2456.0400 740.4800 2456.5200 ;
        RECT 738.8800 2461.4800 740.4800 2461.9600 ;
        RECT 783.8800 2439.7200 785.4800 2440.2000 ;
        RECT 783.8800 2445.1600 785.4800 2445.6400 ;
        RECT 783.8800 2450.6000 785.4800 2451.0800 ;
        RECT 783.8800 2428.8400 785.4800 2429.3200 ;
        RECT 783.8800 2434.2800 785.4800 2434.7600 ;
        RECT 738.8800 2439.7200 740.4800 2440.2000 ;
        RECT 738.8800 2445.1600 740.4800 2445.6400 ;
        RECT 738.8800 2450.6000 740.4800 2451.0800 ;
        RECT 738.8800 2428.8400 740.4800 2429.3200 ;
        RECT 738.8800 2434.2800 740.4800 2434.7600 ;
        RECT 693.8800 2466.9200 695.4800 2467.4000 ;
        RECT 693.8800 2472.3600 695.4800 2472.8400 ;
        RECT 693.8800 2477.8000 695.4800 2478.2800 ;
        RECT 682.1200 2466.9200 685.1200 2467.4000 ;
        RECT 682.1200 2472.3600 685.1200 2472.8400 ;
        RECT 682.1200 2477.8000 685.1200 2478.2800 ;
        RECT 693.8800 2456.0400 695.4800 2456.5200 ;
        RECT 693.8800 2461.4800 695.4800 2461.9600 ;
        RECT 682.1200 2456.0400 685.1200 2456.5200 ;
        RECT 682.1200 2461.4800 685.1200 2461.9600 ;
        RECT 693.8800 2439.7200 695.4800 2440.2000 ;
        RECT 693.8800 2445.1600 695.4800 2445.6400 ;
        RECT 693.8800 2450.6000 695.4800 2451.0800 ;
        RECT 682.1200 2439.7200 685.1200 2440.2000 ;
        RECT 682.1200 2445.1600 685.1200 2445.6400 ;
        RECT 682.1200 2450.6000 685.1200 2451.0800 ;
        RECT 693.8800 2428.8400 695.4800 2429.3200 ;
        RECT 693.8800 2434.2800 695.4800 2434.7600 ;
        RECT 682.1200 2428.8400 685.1200 2429.3200 ;
        RECT 682.1200 2434.2800 685.1200 2434.7600 ;
        RECT 783.8800 2412.5200 785.4800 2413.0000 ;
        RECT 783.8800 2417.9600 785.4800 2418.4400 ;
        RECT 783.8800 2423.4000 785.4800 2423.8800 ;
        RECT 783.8800 2401.6400 785.4800 2402.1200 ;
        RECT 783.8800 2407.0800 785.4800 2407.5600 ;
        RECT 738.8800 2412.5200 740.4800 2413.0000 ;
        RECT 738.8800 2417.9600 740.4800 2418.4400 ;
        RECT 738.8800 2423.4000 740.4800 2423.8800 ;
        RECT 738.8800 2401.6400 740.4800 2402.1200 ;
        RECT 738.8800 2407.0800 740.4800 2407.5600 ;
        RECT 783.8800 2385.3200 785.4800 2385.8000 ;
        RECT 783.8800 2390.7600 785.4800 2391.2400 ;
        RECT 783.8800 2396.2000 785.4800 2396.6800 ;
        RECT 783.8800 2379.8800 785.4800 2380.3600 ;
        RECT 738.8800 2385.3200 740.4800 2385.8000 ;
        RECT 738.8800 2390.7600 740.4800 2391.2400 ;
        RECT 738.8800 2396.2000 740.4800 2396.6800 ;
        RECT 738.8800 2379.8800 740.4800 2380.3600 ;
        RECT 693.8800 2412.5200 695.4800 2413.0000 ;
        RECT 693.8800 2417.9600 695.4800 2418.4400 ;
        RECT 693.8800 2423.4000 695.4800 2423.8800 ;
        RECT 682.1200 2412.5200 685.1200 2413.0000 ;
        RECT 682.1200 2417.9600 685.1200 2418.4400 ;
        RECT 682.1200 2423.4000 685.1200 2423.8800 ;
        RECT 693.8800 2401.6400 695.4800 2402.1200 ;
        RECT 693.8800 2407.0800 695.4800 2407.5600 ;
        RECT 682.1200 2401.6400 685.1200 2402.1200 ;
        RECT 682.1200 2407.0800 685.1200 2407.5600 ;
        RECT 693.8800 2385.3200 695.4800 2385.8000 ;
        RECT 693.8800 2390.7600 695.4800 2391.2400 ;
        RECT 693.8800 2396.2000 695.4800 2396.6800 ;
        RECT 682.1200 2385.3200 685.1200 2385.8000 ;
        RECT 682.1200 2390.7600 685.1200 2391.2400 ;
        RECT 682.1200 2396.2000 685.1200 2396.6800 ;
        RECT 682.1200 2379.8800 685.1200 2380.3600 ;
        RECT 693.8800 2379.8800 695.4800 2380.3600 ;
        RECT 682.1200 2584.7900 889.2200 2587.7900 ;
        RECT 682.1200 2371.6900 889.2200 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 2142.0500 875.4800 2358.1500 ;
        RECT 828.8800 2142.0500 830.4800 2358.1500 ;
        RECT 783.8800 2142.0500 785.4800 2358.1500 ;
        RECT 738.8800 2142.0500 740.4800 2358.1500 ;
        RECT 693.8800 2142.0500 695.4800 2358.1500 ;
        RECT 886.2200 2142.0500 889.2200 2358.1500 ;
        RECT 682.1200 2142.0500 685.1200 2358.1500 ;
      LAYER met3 ;
        RECT 886.2200 2335.2000 889.2200 2335.6800 ;
        RECT 886.2200 2340.6400 889.2200 2341.1200 ;
        RECT 873.8800 2335.2000 875.4800 2335.6800 ;
        RECT 873.8800 2340.6400 875.4800 2341.1200 ;
        RECT 886.2200 2346.0800 889.2200 2346.5600 ;
        RECT 873.8800 2346.0800 875.4800 2346.5600 ;
        RECT 886.2200 2324.3200 889.2200 2324.8000 ;
        RECT 886.2200 2329.7600 889.2200 2330.2400 ;
        RECT 873.8800 2324.3200 875.4800 2324.8000 ;
        RECT 873.8800 2329.7600 875.4800 2330.2400 ;
        RECT 886.2200 2308.0000 889.2200 2308.4800 ;
        RECT 886.2200 2313.4400 889.2200 2313.9200 ;
        RECT 873.8800 2308.0000 875.4800 2308.4800 ;
        RECT 873.8800 2313.4400 875.4800 2313.9200 ;
        RECT 886.2200 2318.8800 889.2200 2319.3600 ;
        RECT 873.8800 2318.8800 875.4800 2319.3600 ;
        RECT 828.8800 2335.2000 830.4800 2335.6800 ;
        RECT 828.8800 2340.6400 830.4800 2341.1200 ;
        RECT 828.8800 2346.0800 830.4800 2346.5600 ;
        RECT 828.8800 2324.3200 830.4800 2324.8000 ;
        RECT 828.8800 2329.7600 830.4800 2330.2400 ;
        RECT 828.8800 2308.0000 830.4800 2308.4800 ;
        RECT 828.8800 2313.4400 830.4800 2313.9200 ;
        RECT 828.8800 2318.8800 830.4800 2319.3600 ;
        RECT 886.2200 2291.6800 889.2200 2292.1600 ;
        RECT 886.2200 2297.1200 889.2200 2297.6000 ;
        RECT 886.2200 2302.5600 889.2200 2303.0400 ;
        RECT 873.8800 2291.6800 875.4800 2292.1600 ;
        RECT 873.8800 2297.1200 875.4800 2297.6000 ;
        RECT 873.8800 2302.5600 875.4800 2303.0400 ;
        RECT 886.2200 2280.8000 889.2200 2281.2800 ;
        RECT 886.2200 2286.2400 889.2200 2286.7200 ;
        RECT 873.8800 2280.8000 875.4800 2281.2800 ;
        RECT 873.8800 2286.2400 875.4800 2286.7200 ;
        RECT 886.2200 2264.4800 889.2200 2264.9600 ;
        RECT 886.2200 2269.9200 889.2200 2270.4000 ;
        RECT 886.2200 2275.3600 889.2200 2275.8400 ;
        RECT 873.8800 2264.4800 875.4800 2264.9600 ;
        RECT 873.8800 2269.9200 875.4800 2270.4000 ;
        RECT 873.8800 2275.3600 875.4800 2275.8400 ;
        RECT 886.2200 2253.6000 889.2200 2254.0800 ;
        RECT 886.2200 2259.0400 889.2200 2259.5200 ;
        RECT 873.8800 2253.6000 875.4800 2254.0800 ;
        RECT 873.8800 2259.0400 875.4800 2259.5200 ;
        RECT 828.8800 2291.6800 830.4800 2292.1600 ;
        RECT 828.8800 2297.1200 830.4800 2297.6000 ;
        RECT 828.8800 2302.5600 830.4800 2303.0400 ;
        RECT 828.8800 2280.8000 830.4800 2281.2800 ;
        RECT 828.8800 2286.2400 830.4800 2286.7200 ;
        RECT 828.8800 2264.4800 830.4800 2264.9600 ;
        RECT 828.8800 2269.9200 830.4800 2270.4000 ;
        RECT 828.8800 2275.3600 830.4800 2275.8400 ;
        RECT 828.8800 2253.6000 830.4800 2254.0800 ;
        RECT 828.8800 2259.0400 830.4800 2259.5200 ;
        RECT 783.8800 2335.2000 785.4800 2335.6800 ;
        RECT 783.8800 2340.6400 785.4800 2341.1200 ;
        RECT 783.8800 2346.0800 785.4800 2346.5600 ;
        RECT 738.8800 2335.2000 740.4800 2335.6800 ;
        RECT 738.8800 2340.6400 740.4800 2341.1200 ;
        RECT 738.8800 2346.0800 740.4800 2346.5600 ;
        RECT 783.8800 2324.3200 785.4800 2324.8000 ;
        RECT 783.8800 2329.7600 785.4800 2330.2400 ;
        RECT 783.8800 2308.0000 785.4800 2308.4800 ;
        RECT 783.8800 2313.4400 785.4800 2313.9200 ;
        RECT 783.8800 2318.8800 785.4800 2319.3600 ;
        RECT 738.8800 2324.3200 740.4800 2324.8000 ;
        RECT 738.8800 2329.7600 740.4800 2330.2400 ;
        RECT 738.8800 2308.0000 740.4800 2308.4800 ;
        RECT 738.8800 2313.4400 740.4800 2313.9200 ;
        RECT 738.8800 2318.8800 740.4800 2319.3600 ;
        RECT 693.8800 2335.2000 695.4800 2335.6800 ;
        RECT 693.8800 2340.6400 695.4800 2341.1200 ;
        RECT 682.1200 2340.6400 685.1200 2341.1200 ;
        RECT 682.1200 2335.2000 685.1200 2335.6800 ;
        RECT 682.1200 2346.0800 685.1200 2346.5600 ;
        RECT 693.8800 2346.0800 695.4800 2346.5600 ;
        RECT 693.8800 2324.3200 695.4800 2324.8000 ;
        RECT 693.8800 2329.7600 695.4800 2330.2400 ;
        RECT 682.1200 2329.7600 685.1200 2330.2400 ;
        RECT 682.1200 2324.3200 685.1200 2324.8000 ;
        RECT 693.8800 2308.0000 695.4800 2308.4800 ;
        RECT 693.8800 2313.4400 695.4800 2313.9200 ;
        RECT 682.1200 2313.4400 685.1200 2313.9200 ;
        RECT 682.1200 2308.0000 685.1200 2308.4800 ;
        RECT 682.1200 2318.8800 685.1200 2319.3600 ;
        RECT 693.8800 2318.8800 695.4800 2319.3600 ;
        RECT 783.8800 2291.6800 785.4800 2292.1600 ;
        RECT 783.8800 2297.1200 785.4800 2297.6000 ;
        RECT 783.8800 2302.5600 785.4800 2303.0400 ;
        RECT 783.8800 2280.8000 785.4800 2281.2800 ;
        RECT 783.8800 2286.2400 785.4800 2286.7200 ;
        RECT 738.8800 2291.6800 740.4800 2292.1600 ;
        RECT 738.8800 2297.1200 740.4800 2297.6000 ;
        RECT 738.8800 2302.5600 740.4800 2303.0400 ;
        RECT 738.8800 2280.8000 740.4800 2281.2800 ;
        RECT 738.8800 2286.2400 740.4800 2286.7200 ;
        RECT 783.8800 2264.4800 785.4800 2264.9600 ;
        RECT 783.8800 2269.9200 785.4800 2270.4000 ;
        RECT 783.8800 2275.3600 785.4800 2275.8400 ;
        RECT 783.8800 2253.6000 785.4800 2254.0800 ;
        RECT 783.8800 2259.0400 785.4800 2259.5200 ;
        RECT 738.8800 2264.4800 740.4800 2264.9600 ;
        RECT 738.8800 2269.9200 740.4800 2270.4000 ;
        RECT 738.8800 2275.3600 740.4800 2275.8400 ;
        RECT 738.8800 2253.6000 740.4800 2254.0800 ;
        RECT 738.8800 2259.0400 740.4800 2259.5200 ;
        RECT 693.8800 2291.6800 695.4800 2292.1600 ;
        RECT 693.8800 2297.1200 695.4800 2297.6000 ;
        RECT 693.8800 2302.5600 695.4800 2303.0400 ;
        RECT 682.1200 2291.6800 685.1200 2292.1600 ;
        RECT 682.1200 2297.1200 685.1200 2297.6000 ;
        RECT 682.1200 2302.5600 685.1200 2303.0400 ;
        RECT 693.8800 2280.8000 695.4800 2281.2800 ;
        RECT 693.8800 2286.2400 695.4800 2286.7200 ;
        RECT 682.1200 2280.8000 685.1200 2281.2800 ;
        RECT 682.1200 2286.2400 685.1200 2286.7200 ;
        RECT 693.8800 2264.4800 695.4800 2264.9600 ;
        RECT 693.8800 2269.9200 695.4800 2270.4000 ;
        RECT 693.8800 2275.3600 695.4800 2275.8400 ;
        RECT 682.1200 2264.4800 685.1200 2264.9600 ;
        RECT 682.1200 2269.9200 685.1200 2270.4000 ;
        RECT 682.1200 2275.3600 685.1200 2275.8400 ;
        RECT 693.8800 2253.6000 695.4800 2254.0800 ;
        RECT 693.8800 2259.0400 695.4800 2259.5200 ;
        RECT 682.1200 2253.6000 685.1200 2254.0800 ;
        RECT 682.1200 2259.0400 685.1200 2259.5200 ;
        RECT 886.2200 2237.2800 889.2200 2237.7600 ;
        RECT 886.2200 2242.7200 889.2200 2243.2000 ;
        RECT 886.2200 2248.1600 889.2200 2248.6400 ;
        RECT 873.8800 2237.2800 875.4800 2237.7600 ;
        RECT 873.8800 2242.7200 875.4800 2243.2000 ;
        RECT 873.8800 2248.1600 875.4800 2248.6400 ;
        RECT 886.2200 2226.4000 889.2200 2226.8800 ;
        RECT 886.2200 2231.8400 889.2200 2232.3200 ;
        RECT 873.8800 2226.4000 875.4800 2226.8800 ;
        RECT 873.8800 2231.8400 875.4800 2232.3200 ;
        RECT 886.2200 2210.0800 889.2200 2210.5600 ;
        RECT 886.2200 2215.5200 889.2200 2216.0000 ;
        RECT 886.2200 2220.9600 889.2200 2221.4400 ;
        RECT 873.8800 2210.0800 875.4800 2210.5600 ;
        RECT 873.8800 2215.5200 875.4800 2216.0000 ;
        RECT 873.8800 2220.9600 875.4800 2221.4400 ;
        RECT 886.2200 2199.2000 889.2200 2199.6800 ;
        RECT 886.2200 2204.6400 889.2200 2205.1200 ;
        RECT 873.8800 2199.2000 875.4800 2199.6800 ;
        RECT 873.8800 2204.6400 875.4800 2205.1200 ;
        RECT 828.8800 2237.2800 830.4800 2237.7600 ;
        RECT 828.8800 2242.7200 830.4800 2243.2000 ;
        RECT 828.8800 2248.1600 830.4800 2248.6400 ;
        RECT 828.8800 2226.4000 830.4800 2226.8800 ;
        RECT 828.8800 2231.8400 830.4800 2232.3200 ;
        RECT 828.8800 2210.0800 830.4800 2210.5600 ;
        RECT 828.8800 2215.5200 830.4800 2216.0000 ;
        RECT 828.8800 2220.9600 830.4800 2221.4400 ;
        RECT 828.8800 2199.2000 830.4800 2199.6800 ;
        RECT 828.8800 2204.6400 830.4800 2205.1200 ;
        RECT 886.2200 2182.8800 889.2200 2183.3600 ;
        RECT 886.2200 2188.3200 889.2200 2188.8000 ;
        RECT 886.2200 2193.7600 889.2200 2194.2400 ;
        RECT 873.8800 2182.8800 875.4800 2183.3600 ;
        RECT 873.8800 2188.3200 875.4800 2188.8000 ;
        RECT 873.8800 2193.7600 875.4800 2194.2400 ;
        RECT 886.2200 2172.0000 889.2200 2172.4800 ;
        RECT 886.2200 2177.4400 889.2200 2177.9200 ;
        RECT 873.8800 2172.0000 875.4800 2172.4800 ;
        RECT 873.8800 2177.4400 875.4800 2177.9200 ;
        RECT 886.2200 2155.6800 889.2200 2156.1600 ;
        RECT 886.2200 2161.1200 889.2200 2161.6000 ;
        RECT 886.2200 2166.5600 889.2200 2167.0400 ;
        RECT 873.8800 2155.6800 875.4800 2156.1600 ;
        RECT 873.8800 2161.1200 875.4800 2161.6000 ;
        RECT 873.8800 2166.5600 875.4800 2167.0400 ;
        RECT 886.2200 2150.2400 889.2200 2150.7200 ;
        RECT 873.8800 2150.2400 875.4800 2150.7200 ;
        RECT 828.8800 2182.8800 830.4800 2183.3600 ;
        RECT 828.8800 2188.3200 830.4800 2188.8000 ;
        RECT 828.8800 2193.7600 830.4800 2194.2400 ;
        RECT 828.8800 2172.0000 830.4800 2172.4800 ;
        RECT 828.8800 2177.4400 830.4800 2177.9200 ;
        RECT 828.8800 2155.6800 830.4800 2156.1600 ;
        RECT 828.8800 2161.1200 830.4800 2161.6000 ;
        RECT 828.8800 2166.5600 830.4800 2167.0400 ;
        RECT 828.8800 2150.2400 830.4800 2150.7200 ;
        RECT 783.8800 2237.2800 785.4800 2237.7600 ;
        RECT 783.8800 2242.7200 785.4800 2243.2000 ;
        RECT 783.8800 2248.1600 785.4800 2248.6400 ;
        RECT 783.8800 2226.4000 785.4800 2226.8800 ;
        RECT 783.8800 2231.8400 785.4800 2232.3200 ;
        RECT 738.8800 2237.2800 740.4800 2237.7600 ;
        RECT 738.8800 2242.7200 740.4800 2243.2000 ;
        RECT 738.8800 2248.1600 740.4800 2248.6400 ;
        RECT 738.8800 2226.4000 740.4800 2226.8800 ;
        RECT 738.8800 2231.8400 740.4800 2232.3200 ;
        RECT 783.8800 2210.0800 785.4800 2210.5600 ;
        RECT 783.8800 2215.5200 785.4800 2216.0000 ;
        RECT 783.8800 2220.9600 785.4800 2221.4400 ;
        RECT 783.8800 2199.2000 785.4800 2199.6800 ;
        RECT 783.8800 2204.6400 785.4800 2205.1200 ;
        RECT 738.8800 2210.0800 740.4800 2210.5600 ;
        RECT 738.8800 2215.5200 740.4800 2216.0000 ;
        RECT 738.8800 2220.9600 740.4800 2221.4400 ;
        RECT 738.8800 2199.2000 740.4800 2199.6800 ;
        RECT 738.8800 2204.6400 740.4800 2205.1200 ;
        RECT 693.8800 2237.2800 695.4800 2237.7600 ;
        RECT 693.8800 2242.7200 695.4800 2243.2000 ;
        RECT 693.8800 2248.1600 695.4800 2248.6400 ;
        RECT 682.1200 2237.2800 685.1200 2237.7600 ;
        RECT 682.1200 2242.7200 685.1200 2243.2000 ;
        RECT 682.1200 2248.1600 685.1200 2248.6400 ;
        RECT 693.8800 2226.4000 695.4800 2226.8800 ;
        RECT 693.8800 2231.8400 695.4800 2232.3200 ;
        RECT 682.1200 2226.4000 685.1200 2226.8800 ;
        RECT 682.1200 2231.8400 685.1200 2232.3200 ;
        RECT 693.8800 2210.0800 695.4800 2210.5600 ;
        RECT 693.8800 2215.5200 695.4800 2216.0000 ;
        RECT 693.8800 2220.9600 695.4800 2221.4400 ;
        RECT 682.1200 2210.0800 685.1200 2210.5600 ;
        RECT 682.1200 2215.5200 685.1200 2216.0000 ;
        RECT 682.1200 2220.9600 685.1200 2221.4400 ;
        RECT 693.8800 2199.2000 695.4800 2199.6800 ;
        RECT 693.8800 2204.6400 695.4800 2205.1200 ;
        RECT 682.1200 2199.2000 685.1200 2199.6800 ;
        RECT 682.1200 2204.6400 685.1200 2205.1200 ;
        RECT 783.8800 2182.8800 785.4800 2183.3600 ;
        RECT 783.8800 2188.3200 785.4800 2188.8000 ;
        RECT 783.8800 2193.7600 785.4800 2194.2400 ;
        RECT 783.8800 2172.0000 785.4800 2172.4800 ;
        RECT 783.8800 2177.4400 785.4800 2177.9200 ;
        RECT 738.8800 2182.8800 740.4800 2183.3600 ;
        RECT 738.8800 2188.3200 740.4800 2188.8000 ;
        RECT 738.8800 2193.7600 740.4800 2194.2400 ;
        RECT 738.8800 2172.0000 740.4800 2172.4800 ;
        RECT 738.8800 2177.4400 740.4800 2177.9200 ;
        RECT 783.8800 2155.6800 785.4800 2156.1600 ;
        RECT 783.8800 2161.1200 785.4800 2161.6000 ;
        RECT 783.8800 2166.5600 785.4800 2167.0400 ;
        RECT 783.8800 2150.2400 785.4800 2150.7200 ;
        RECT 738.8800 2155.6800 740.4800 2156.1600 ;
        RECT 738.8800 2161.1200 740.4800 2161.6000 ;
        RECT 738.8800 2166.5600 740.4800 2167.0400 ;
        RECT 738.8800 2150.2400 740.4800 2150.7200 ;
        RECT 693.8800 2182.8800 695.4800 2183.3600 ;
        RECT 693.8800 2188.3200 695.4800 2188.8000 ;
        RECT 693.8800 2193.7600 695.4800 2194.2400 ;
        RECT 682.1200 2182.8800 685.1200 2183.3600 ;
        RECT 682.1200 2188.3200 685.1200 2188.8000 ;
        RECT 682.1200 2193.7600 685.1200 2194.2400 ;
        RECT 693.8800 2172.0000 695.4800 2172.4800 ;
        RECT 693.8800 2177.4400 695.4800 2177.9200 ;
        RECT 682.1200 2172.0000 685.1200 2172.4800 ;
        RECT 682.1200 2177.4400 685.1200 2177.9200 ;
        RECT 693.8800 2155.6800 695.4800 2156.1600 ;
        RECT 693.8800 2161.1200 695.4800 2161.6000 ;
        RECT 693.8800 2166.5600 695.4800 2167.0400 ;
        RECT 682.1200 2155.6800 685.1200 2156.1600 ;
        RECT 682.1200 2161.1200 685.1200 2161.6000 ;
        RECT 682.1200 2166.5600 685.1200 2167.0400 ;
        RECT 682.1200 2150.2400 685.1200 2150.7200 ;
        RECT 693.8800 2150.2400 695.4800 2150.7200 ;
        RECT 682.1200 2355.1500 889.2200 2358.1500 ;
        RECT 682.1200 2142.0500 889.2200 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 1912.4100 875.4800 2128.5100 ;
        RECT 828.8800 1912.4100 830.4800 2128.5100 ;
        RECT 783.8800 1912.4100 785.4800 2128.5100 ;
        RECT 738.8800 1912.4100 740.4800 2128.5100 ;
        RECT 693.8800 1912.4100 695.4800 2128.5100 ;
        RECT 886.2200 1912.4100 889.2200 2128.5100 ;
        RECT 682.1200 1912.4100 685.1200 2128.5100 ;
      LAYER met3 ;
        RECT 886.2200 2105.5600 889.2200 2106.0400 ;
        RECT 886.2200 2111.0000 889.2200 2111.4800 ;
        RECT 873.8800 2105.5600 875.4800 2106.0400 ;
        RECT 873.8800 2111.0000 875.4800 2111.4800 ;
        RECT 886.2200 2116.4400 889.2200 2116.9200 ;
        RECT 873.8800 2116.4400 875.4800 2116.9200 ;
        RECT 886.2200 2094.6800 889.2200 2095.1600 ;
        RECT 886.2200 2100.1200 889.2200 2100.6000 ;
        RECT 873.8800 2094.6800 875.4800 2095.1600 ;
        RECT 873.8800 2100.1200 875.4800 2100.6000 ;
        RECT 886.2200 2078.3600 889.2200 2078.8400 ;
        RECT 886.2200 2083.8000 889.2200 2084.2800 ;
        RECT 873.8800 2078.3600 875.4800 2078.8400 ;
        RECT 873.8800 2083.8000 875.4800 2084.2800 ;
        RECT 886.2200 2089.2400 889.2200 2089.7200 ;
        RECT 873.8800 2089.2400 875.4800 2089.7200 ;
        RECT 828.8800 2105.5600 830.4800 2106.0400 ;
        RECT 828.8800 2111.0000 830.4800 2111.4800 ;
        RECT 828.8800 2116.4400 830.4800 2116.9200 ;
        RECT 828.8800 2094.6800 830.4800 2095.1600 ;
        RECT 828.8800 2100.1200 830.4800 2100.6000 ;
        RECT 828.8800 2078.3600 830.4800 2078.8400 ;
        RECT 828.8800 2083.8000 830.4800 2084.2800 ;
        RECT 828.8800 2089.2400 830.4800 2089.7200 ;
        RECT 886.2200 2062.0400 889.2200 2062.5200 ;
        RECT 886.2200 2067.4800 889.2200 2067.9600 ;
        RECT 886.2200 2072.9200 889.2200 2073.4000 ;
        RECT 873.8800 2062.0400 875.4800 2062.5200 ;
        RECT 873.8800 2067.4800 875.4800 2067.9600 ;
        RECT 873.8800 2072.9200 875.4800 2073.4000 ;
        RECT 886.2200 2051.1600 889.2200 2051.6400 ;
        RECT 886.2200 2056.6000 889.2200 2057.0800 ;
        RECT 873.8800 2051.1600 875.4800 2051.6400 ;
        RECT 873.8800 2056.6000 875.4800 2057.0800 ;
        RECT 886.2200 2034.8400 889.2200 2035.3200 ;
        RECT 886.2200 2040.2800 889.2200 2040.7600 ;
        RECT 886.2200 2045.7200 889.2200 2046.2000 ;
        RECT 873.8800 2034.8400 875.4800 2035.3200 ;
        RECT 873.8800 2040.2800 875.4800 2040.7600 ;
        RECT 873.8800 2045.7200 875.4800 2046.2000 ;
        RECT 886.2200 2023.9600 889.2200 2024.4400 ;
        RECT 886.2200 2029.4000 889.2200 2029.8800 ;
        RECT 873.8800 2023.9600 875.4800 2024.4400 ;
        RECT 873.8800 2029.4000 875.4800 2029.8800 ;
        RECT 828.8800 2062.0400 830.4800 2062.5200 ;
        RECT 828.8800 2067.4800 830.4800 2067.9600 ;
        RECT 828.8800 2072.9200 830.4800 2073.4000 ;
        RECT 828.8800 2051.1600 830.4800 2051.6400 ;
        RECT 828.8800 2056.6000 830.4800 2057.0800 ;
        RECT 828.8800 2034.8400 830.4800 2035.3200 ;
        RECT 828.8800 2040.2800 830.4800 2040.7600 ;
        RECT 828.8800 2045.7200 830.4800 2046.2000 ;
        RECT 828.8800 2023.9600 830.4800 2024.4400 ;
        RECT 828.8800 2029.4000 830.4800 2029.8800 ;
        RECT 783.8800 2105.5600 785.4800 2106.0400 ;
        RECT 783.8800 2111.0000 785.4800 2111.4800 ;
        RECT 783.8800 2116.4400 785.4800 2116.9200 ;
        RECT 738.8800 2105.5600 740.4800 2106.0400 ;
        RECT 738.8800 2111.0000 740.4800 2111.4800 ;
        RECT 738.8800 2116.4400 740.4800 2116.9200 ;
        RECT 783.8800 2094.6800 785.4800 2095.1600 ;
        RECT 783.8800 2100.1200 785.4800 2100.6000 ;
        RECT 783.8800 2078.3600 785.4800 2078.8400 ;
        RECT 783.8800 2083.8000 785.4800 2084.2800 ;
        RECT 783.8800 2089.2400 785.4800 2089.7200 ;
        RECT 738.8800 2094.6800 740.4800 2095.1600 ;
        RECT 738.8800 2100.1200 740.4800 2100.6000 ;
        RECT 738.8800 2078.3600 740.4800 2078.8400 ;
        RECT 738.8800 2083.8000 740.4800 2084.2800 ;
        RECT 738.8800 2089.2400 740.4800 2089.7200 ;
        RECT 693.8800 2105.5600 695.4800 2106.0400 ;
        RECT 693.8800 2111.0000 695.4800 2111.4800 ;
        RECT 682.1200 2111.0000 685.1200 2111.4800 ;
        RECT 682.1200 2105.5600 685.1200 2106.0400 ;
        RECT 682.1200 2116.4400 685.1200 2116.9200 ;
        RECT 693.8800 2116.4400 695.4800 2116.9200 ;
        RECT 693.8800 2094.6800 695.4800 2095.1600 ;
        RECT 693.8800 2100.1200 695.4800 2100.6000 ;
        RECT 682.1200 2100.1200 685.1200 2100.6000 ;
        RECT 682.1200 2094.6800 685.1200 2095.1600 ;
        RECT 693.8800 2078.3600 695.4800 2078.8400 ;
        RECT 693.8800 2083.8000 695.4800 2084.2800 ;
        RECT 682.1200 2083.8000 685.1200 2084.2800 ;
        RECT 682.1200 2078.3600 685.1200 2078.8400 ;
        RECT 682.1200 2089.2400 685.1200 2089.7200 ;
        RECT 693.8800 2089.2400 695.4800 2089.7200 ;
        RECT 783.8800 2062.0400 785.4800 2062.5200 ;
        RECT 783.8800 2067.4800 785.4800 2067.9600 ;
        RECT 783.8800 2072.9200 785.4800 2073.4000 ;
        RECT 783.8800 2051.1600 785.4800 2051.6400 ;
        RECT 783.8800 2056.6000 785.4800 2057.0800 ;
        RECT 738.8800 2062.0400 740.4800 2062.5200 ;
        RECT 738.8800 2067.4800 740.4800 2067.9600 ;
        RECT 738.8800 2072.9200 740.4800 2073.4000 ;
        RECT 738.8800 2051.1600 740.4800 2051.6400 ;
        RECT 738.8800 2056.6000 740.4800 2057.0800 ;
        RECT 783.8800 2034.8400 785.4800 2035.3200 ;
        RECT 783.8800 2040.2800 785.4800 2040.7600 ;
        RECT 783.8800 2045.7200 785.4800 2046.2000 ;
        RECT 783.8800 2023.9600 785.4800 2024.4400 ;
        RECT 783.8800 2029.4000 785.4800 2029.8800 ;
        RECT 738.8800 2034.8400 740.4800 2035.3200 ;
        RECT 738.8800 2040.2800 740.4800 2040.7600 ;
        RECT 738.8800 2045.7200 740.4800 2046.2000 ;
        RECT 738.8800 2023.9600 740.4800 2024.4400 ;
        RECT 738.8800 2029.4000 740.4800 2029.8800 ;
        RECT 693.8800 2062.0400 695.4800 2062.5200 ;
        RECT 693.8800 2067.4800 695.4800 2067.9600 ;
        RECT 693.8800 2072.9200 695.4800 2073.4000 ;
        RECT 682.1200 2062.0400 685.1200 2062.5200 ;
        RECT 682.1200 2067.4800 685.1200 2067.9600 ;
        RECT 682.1200 2072.9200 685.1200 2073.4000 ;
        RECT 693.8800 2051.1600 695.4800 2051.6400 ;
        RECT 693.8800 2056.6000 695.4800 2057.0800 ;
        RECT 682.1200 2051.1600 685.1200 2051.6400 ;
        RECT 682.1200 2056.6000 685.1200 2057.0800 ;
        RECT 693.8800 2034.8400 695.4800 2035.3200 ;
        RECT 693.8800 2040.2800 695.4800 2040.7600 ;
        RECT 693.8800 2045.7200 695.4800 2046.2000 ;
        RECT 682.1200 2034.8400 685.1200 2035.3200 ;
        RECT 682.1200 2040.2800 685.1200 2040.7600 ;
        RECT 682.1200 2045.7200 685.1200 2046.2000 ;
        RECT 693.8800 2023.9600 695.4800 2024.4400 ;
        RECT 693.8800 2029.4000 695.4800 2029.8800 ;
        RECT 682.1200 2023.9600 685.1200 2024.4400 ;
        RECT 682.1200 2029.4000 685.1200 2029.8800 ;
        RECT 886.2200 2007.6400 889.2200 2008.1200 ;
        RECT 886.2200 2013.0800 889.2200 2013.5600 ;
        RECT 886.2200 2018.5200 889.2200 2019.0000 ;
        RECT 873.8800 2007.6400 875.4800 2008.1200 ;
        RECT 873.8800 2013.0800 875.4800 2013.5600 ;
        RECT 873.8800 2018.5200 875.4800 2019.0000 ;
        RECT 886.2200 1996.7600 889.2200 1997.2400 ;
        RECT 886.2200 2002.2000 889.2200 2002.6800 ;
        RECT 873.8800 1996.7600 875.4800 1997.2400 ;
        RECT 873.8800 2002.2000 875.4800 2002.6800 ;
        RECT 886.2200 1980.4400 889.2200 1980.9200 ;
        RECT 886.2200 1985.8800 889.2200 1986.3600 ;
        RECT 886.2200 1991.3200 889.2200 1991.8000 ;
        RECT 873.8800 1980.4400 875.4800 1980.9200 ;
        RECT 873.8800 1985.8800 875.4800 1986.3600 ;
        RECT 873.8800 1991.3200 875.4800 1991.8000 ;
        RECT 886.2200 1969.5600 889.2200 1970.0400 ;
        RECT 886.2200 1975.0000 889.2200 1975.4800 ;
        RECT 873.8800 1969.5600 875.4800 1970.0400 ;
        RECT 873.8800 1975.0000 875.4800 1975.4800 ;
        RECT 828.8800 2007.6400 830.4800 2008.1200 ;
        RECT 828.8800 2013.0800 830.4800 2013.5600 ;
        RECT 828.8800 2018.5200 830.4800 2019.0000 ;
        RECT 828.8800 1996.7600 830.4800 1997.2400 ;
        RECT 828.8800 2002.2000 830.4800 2002.6800 ;
        RECT 828.8800 1980.4400 830.4800 1980.9200 ;
        RECT 828.8800 1985.8800 830.4800 1986.3600 ;
        RECT 828.8800 1991.3200 830.4800 1991.8000 ;
        RECT 828.8800 1969.5600 830.4800 1970.0400 ;
        RECT 828.8800 1975.0000 830.4800 1975.4800 ;
        RECT 886.2200 1953.2400 889.2200 1953.7200 ;
        RECT 886.2200 1958.6800 889.2200 1959.1600 ;
        RECT 886.2200 1964.1200 889.2200 1964.6000 ;
        RECT 873.8800 1953.2400 875.4800 1953.7200 ;
        RECT 873.8800 1958.6800 875.4800 1959.1600 ;
        RECT 873.8800 1964.1200 875.4800 1964.6000 ;
        RECT 886.2200 1942.3600 889.2200 1942.8400 ;
        RECT 886.2200 1947.8000 889.2200 1948.2800 ;
        RECT 873.8800 1942.3600 875.4800 1942.8400 ;
        RECT 873.8800 1947.8000 875.4800 1948.2800 ;
        RECT 886.2200 1926.0400 889.2200 1926.5200 ;
        RECT 886.2200 1931.4800 889.2200 1931.9600 ;
        RECT 886.2200 1936.9200 889.2200 1937.4000 ;
        RECT 873.8800 1926.0400 875.4800 1926.5200 ;
        RECT 873.8800 1931.4800 875.4800 1931.9600 ;
        RECT 873.8800 1936.9200 875.4800 1937.4000 ;
        RECT 886.2200 1920.6000 889.2200 1921.0800 ;
        RECT 873.8800 1920.6000 875.4800 1921.0800 ;
        RECT 828.8800 1953.2400 830.4800 1953.7200 ;
        RECT 828.8800 1958.6800 830.4800 1959.1600 ;
        RECT 828.8800 1964.1200 830.4800 1964.6000 ;
        RECT 828.8800 1942.3600 830.4800 1942.8400 ;
        RECT 828.8800 1947.8000 830.4800 1948.2800 ;
        RECT 828.8800 1926.0400 830.4800 1926.5200 ;
        RECT 828.8800 1931.4800 830.4800 1931.9600 ;
        RECT 828.8800 1936.9200 830.4800 1937.4000 ;
        RECT 828.8800 1920.6000 830.4800 1921.0800 ;
        RECT 783.8800 2007.6400 785.4800 2008.1200 ;
        RECT 783.8800 2013.0800 785.4800 2013.5600 ;
        RECT 783.8800 2018.5200 785.4800 2019.0000 ;
        RECT 783.8800 1996.7600 785.4800 1997.2400 ;
        RECT 783.8800 2002.2000 785.4800 2002.6800 ;
        RECT 738.8800 2007.6400 740.4800 2008.1200 ;
        RECT 738.8800 2013.0800 740.4800 2013.5600 ;
        RECT 738.8800 2018.5200 740.4800 2019.0000 ;
        RECT 738.8800 1996.7600 740.4800 1997.2400 ;
        RECT 738.8800 2002.2000 740.4800 2002.6800 ;
        RECT 783.8800 1980.4400 785.4800 1980.9200 ;
        RECT 783.8800 1985.8800 785.4800 1986.3600 ;
        RECT 783.8800 1991.3200 785.4800 1991.8000 ;
        RECT 783.8800 1969.5600 785.4800 1970.0400 ;
        RECT 783.8800 1975.0000 785.4800 1975.4800 ;
        RECT 738.8800 1980.4400 740.4800 1980.9200 ;
        RECT 738.8800 1985.8800 740.4800 1986.3600 ;
        RECT 738.8800 1991.3200 740.4800 1991.8000 ;
        RECT 738.8800 1969.5600 740.4800 1970.0400 ;
        RECT 738.8800 1975.0000 740.4800 1975.4800 ;
        RECT 693.8800 2007.6400 695.4800 2008.1200 ;
        RECT 693.8800 2013.0800 695.4800 2013.5600 ;
        RECT 693.8800 2018.5200 695.4800 2019.0000 ;
        RECT 682.1200 2007.6400 685.1200 2008.1200 ;
        RECT 682.1200 2013.0800 685.1200 2013.5600 ;
        RECT 682.1200 2018.5200 685.1200 2019.0000 ;
        RECT 693.8800 1996.7600 695.4800 1997.2400 ;
        RECT 693.8800 2002.2000 695.4800 2002.6800 ;
        RECT 682.1200 1996.7600 685.1200 1997.2400 ;
        RECT 682.1200 2002.2000 685.1200 2002.6800 ;
        RECT 693.8800 1980.4400 695.4800 1980.9200 ;
        RECT 693.8800 1985.8800 695.4800 1986.3600 ;
        RECT 693.8800 1991.3200 695.4800 1991.8000 ;
        RECT 682.1200 1980.4400 685.1200 1980.9200 ;
        RECT 682.1200 1985.8800 685.1200 1986.3600 ;
        RECT 682.1200 1991.3200 685.1200 1991.8000 ;
        RECT 693.8800 1969.5600 695.4800 1970.0400 ;
        RECT 693.8800 1975.0000 695.4800 1975.4800 ;
        RECT 682.1200 1969.5600 685.1200 1970.0400 ;
        RECT 682.1200 1975.0000 685.1200 1975.4800 ;
        RECT 783.8800 1953.2400 785.4800 1953.7200 ;
        RECT 783.8800 1958.6800 785.4800 1959.1600 ;
        RECT 783.8800 1964.1200 785.4800 1964.6000 ;
        RECT 783.8800 1942.3600 785.4800 1942.8400 ;
        RECT 783.8800 1947.8000 785.4800 1948.2800 ;
        RECT 738.8800 1953.2400 740.4800 1953.7200 ;
        RECT 738.8800 1958.6800 740.4800 1959.1600 ;
        RECT 738.8800 1964.1200 740.4800 1964.6000 ;
        RECT 738.8800 1942.3600 740.4800 1942.8400 ;
        RECT 738.8800 1947.8000 740.4800 1948.2800 ;
        RECT 783.8800 1926.0400 785.4800 1926.5200 ;
        RECT 783.8800 1931.4800 785.4800 1931.9600 ;
        RECT 783.8800 1936.9200 785.4800 1937.4000 ;
        RECT 783.8800 1920.6000 785.4800 1921.0800 ;
        RECT 738.8800 1926.0400 740.4800 1926.5200 ;
        RECT 738.8800 1931.4800 740.4800 1931.9600 ;
        RECT 738.8800 1936.9200 740.4800 1937.4000 ;
        RECT 738.8800 1920.6000 740.4800 1921.0800 ;
        RECT 693.8800 1953.2400 695.4800 1953.7200 ;
        RECT 693.8800 1958.6800 695.4800 1959.1600 ;
        RECT 693.8800 1964.1200 695.4800 1964.6000 ;
        RECT 682.1200 1953.2400 685.1200 1953.7200 ;
        RECT 682.1200 1958.6800 685.1200 1959.1600 ;
        RECT 682.1200 1964.1200 685.1200 1964.6000 ;
        RECT 693.8800 1942.3600 695.4800 1942.8400 ;
        RECT 693.8800 1947.8000 695.4800 1948.2800 ;
        RECT 682.1200 1942.3600 685.1200 1942.8400 ;
        RECT 682.1200 1947.8000 685.1200 1948.2800 ;
        RECT 693.8800 1926.0400 695.4800 1926.5200 ;
        RECT 693.8800 1931.4800 695.4800 1931.9600 ;
        RECT 693.8800 1936.9200 695.4800 1937.4000 ;
        RECT 682.1200 1926.0400 685.1200 1926.5200 ;
        RECT 682.1200 1931.4800 685.1200 1931.9600 ;
        RECT 682.1200 1936.9200 685.1200 1937.4000 ;
        RECT 682.1200 1920.6000 685.1200 1921.0800 ;
        RECT 693.8800 1920.6000 695.4800 1921.0800 ;
        RECT 682.1200 2125.5100 889.2200 2128.5100 ;
        RECT 682.1200 1912.4100 889.2200 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 1682.7700 875.4800 1898.8700 ;
        RECT 828.8800 1682.7700 830.4800 1898.8700 ;
        RECT 783.8800 1682.7700 785.4800 1898.8700 ;
        RECT 738.8800 1682.7700 740.4800 1898.8700 ;
        RECT 693.8800 1682.7700 695.4800 1898.8700 ;
        RECT 886.2200 1682.7700 889.2200 1898.8700 ;
        RECT 682.1200 1682.7700 685.1200 1898.8700 ;
      LAYER met3 ;
        RECT 886.2200 1875.9200 889.2200 1876.4000 ;
        RECT 886.2200 1881.3600 889.2200 1881.8400 ;
        RECT 873.8800 1875.9200 875.4800 1876.4000 ;
        RECT 873.8800 1881.3600 875.4800 1881.8400 ;
        RECT 886.2200 1886.8000 889.2200 1887.2800 ;
        RECT 873.8800 1886.8000 875.4800 1887.2800 ;
        RECT 886.2200 1865.0400 889.2200 1865.5200 ;
        RECT 886.2200 1870.4800 889.2200 1870.9600 ;
        RECT 873.8800 1865.0400 875.4800 1865.5200 ;
        RECT 873.8800 1870.4800 875.4800 1870.9600 ;
        RECT 886.2200 1848.7200 889.2200 1849.2000 ;
        RECT 886.2200 1854.1600 889.2200 1854.6400 ;
        RECT 873.8800 1848.7200 875.4800 1849.2000 ;
        RECT 873.8800 1854.1600 875.4800 1854.6400 ;
        RECT 886.2200 1859.6000 889.2200 1860.0800 ;
        RECT 873.8800 1859.6000 875.4800 1860.0800 ;
        RECT 828.8800 1875.9200 830.4800 1876.4000 ;
        RECT 828.8800 1881.3600 830.4800 1881.8400 ;
        RECT 828.8800 1886.8000 830.4800 1887.2800 ;
        RECT 828.8800 1865.0400 830.4800 1865.5200 ;
        RECT 828.8800 1870.4800 830.4800 1870.9600 ;
        RECT 828.8800 1848.7200 830.4800 1849.2000 ;
        RECT 828.8800 1854.1600 830.4800 1854.6400 ;
        RECT 828.8800 1859.6000 830.4800 1860.0800 ;
        RECT 886.2200 1832.4000 889.2200 1832.8800 ;
        RECT 886.2200 1837.8400 889.2200 1838.3200 ;
        RECT 886.2200 1843.2800 889.2200 1843.7600 ;
        RECT 873.8800 1832.4000 875.4800 1832.8800 ;
        RECT 873.8800 1837.8400 875.4800 1838.3200 ;
        RECT 873.8800 1843.2800 875.4800 1843.7600 ;
        RECT 886.2200 1821.5200 889.2200 1822.0000 ;
        RECT 886.2200 1826.9600 889.2200 1827.4400 ;
        RECT 873.8800 1821.5200 875.4800 1822.0000 ;
        RECT 873.8800 1826.9600 875.4800 1827.4400 ;
        RECT 886.2200 1805.2000 889.2200 1805.6800 ;
        RECT 886.2200 1810.6400 889.2200 1811.1200 ;
        RECT 886.2200 1816.0800 889.2200 1816.5600 ;
        RECT 873.8800 1805.2000 875.4800 1805.6800 ;
        RECT 873.8800 1810.6400 875.4800 1811.1200 ;
        RECT 873.8800 1816.0800 875.4800 1816.5600 ;
        RECT 886.2200 1794.3200 889.2200 1794.8000 ;
        RECT 886.2200 1799.7600 889.2200 1800.2400 ;
        RECT 873.8800 1794.3200 875.4800 1794.8000 ;
        RECT 873.8800 1799.7600 875.4800 1800.2400 ;
        RECT 828.8800 1832.4000 830.4800 1832.8800 ;
        RECT 828.8800 1837.8400 830.4800 1838.3200 ;
        RECT 828.8800 1843.2800 830.4800 1843.7600 ;
        RECT 828.8800 1821.5200 830.4800 1822.0000 ;
        RECT 828.8800 1826.9600 830.4800 1827.4400 ;
        RECT 828.8800 1805.2000 830.4800 1805.6800 ;
        RECT 828.8800 1810.6400 830.4800 1811.1200 ;
        RECT 828.8800 1816.0800 830.4800 1816.5600 ;
        RECT 828.8800 1794.3200 830.4800 1794.8000 ;
        RECT 828.8800 1799.7600 830.4800 1800.2400 ;
        RECT 783.8800 1875.9200 785.4800 1876.4000 ;
        RECT 783.8800 1881.3600 785.4800 1881.8400 ;
        RECT 783.8800 1886.8000 785.4800 1887.2800 ;
        RECT 738.8800 1875.9200 740.4800 1876.4000 ;
        RECT 738.8800 1881.3600 740.4800 1881.8400 ;
        RECT 738.8800 1886.8000 740.4800 1887.2800 ;
        RECT 783.8800 1865.0400 785.4800 1865.5200 ;
        RECT 783.8800 1870.4800 785.4800 1870.9600 ;
        RECT 783.8800 1848.7200 785.4800 1849.2000 ;
        RECT 783.8800 1854.1600 785.4800 1854.6400 ;
        RECT 783.8800 1859.6000 785.4800 1860.0800 ;
        RECT 738.8800 1865.0400 740.4800 1865.5200 ;
        RECT 738.8800 1870.4800 740.4800 1870.9600 ;
        RECT 738.8800 1848.7200 740.4800 1849.2000 ;
        RECT 738.8800 1854.1600 740.4800 1854.6400 ;
        RECT 738.8800 1859.6000 740.4800 1860.0800 ;
        RECT 693.8800 1875.9200 695.4800 1876.4000 ;
        RECT 693.8800 1881.3600 695.4800 1881.8400 ;
        RECT 682.1200 1881.3600 685.1200 1881.8400 ;
        RECT 682.1200 1875.9200 685.1200 1876.4000 ;
        RECT 682.1200 1886.8000 685.1200 1887.2800 ;
        RECT 693.8800 1886.8000 695.4800 1887.2800 ;
        RECT 693.8800 1865.0400 695.4800 1865.5200 ;
        RECT 693.8800 1870.4800 695.4800 1870.9600 ;
        RECT 682.1200 1870.4800 685.1200 1870.9600 ;
        RECT 682.1200 1865.0400 685.1200 1865.5200 ;
        RECT 693.8800 1848.7200 695.4800 1849.2000 ;
        RECT 693.8800 1854.1600 695.4800 1854.6400 ;
        RECT 682.1200 1854.1600 685.1200 1854.6400 ;
        RECT 682.1200 1848.7200 685.1200 1849.2000 ;
        RECT 682.1200 1859.6000 685.1200 1860.0800 ;
        RECT 693.8800 1859.6000 695.4800 1860.0800 ;
        RECT 783.8800 1832.4000 785.4800 1832.8800 ;
        RECT 783.8800 1837.8400 785.4800 1838.3200 ;
        RECT 783.8800 1843.2800 785.4800 1843.7600 ;
        RECT 783.8800 1821.5200 785.4800 1822.0000 ;
        RECT 783.8800 1826.9600 785.4800 1827.4400 ;
        RECT 738.8800 1832.4000 740.4800 1832.8800 ;
        RECT 738.8800 1837.8400 740.4800 1838.3200 ;
        RECT 738.8800 1843.2800 740.4800 1843.7600 ;
        RECT 738.8800 1821.5200 740.4800 1822.0000 ;
        RECT 738.8800 1826.9600 740.4800 1827.4400 ;
        RECT 783.8800 1805.2000 785.4800 1805.6800 ;
        RECT 783.8800 1810.6400 785.4800 1811.1200 ;
        RECT 783.8800 1816.0800 785.4800 1816.5600 ;
        RECT 783.8800 1794.3200 785.4800 1794.8000 ;
        RECT 783.8800 1799.7600 785.4800 1800.2400 ;
        RECT 738.8800 1805.2000 740.4800 1805.6800 ;
        RECT 738.8800 1810.6400 740.4800 1811.1200 ;
        RECT 738.8800 1816.0800 740.4800 1816.5600 ;
        RECT 738.8800 1794.3200 740.4800 1794.8000 ;
        RECT 738.8800 1799.7600 740.4800 1800.2400 ;
        RECT 693.8800 1832.4000 695.4800 1832.8800 ;
        RECT 693.8800 1837.8400 695.4800 1838.3200 ;
        RECT 693.8800 1843.2800 695.4800 1843.7600 ;
        RECT 682.1200 1832.4000 685.1200 1832.8800 ;
        RECT 682.1200 1837.8400 685.1200 1838.3200 ;
        RECT 682.1200 1843.2800 685.1200 1843.7600 ;
        RECT 693.8800 1821.5200 695.4800 1822.0000 ;
        RECT 693.8800 1826.9600 695.4800 1827.4400 ;
        RECT 682.1200 1821.5200 685.1200 1822.0000 ;
        RECT 682.1200 1826.9600 685.1200 1827.4400 ;
        RECT 693.8800 1805.2000 695.4800 1805.6800 ;
        RECT 693.8800 1810.6400 695.4800 1811.1200 ;
        RECT 693.8800 1816.0800 695.4800 1816.5600 ;
        RECT 682.1200 1805.2000 685.1200 1805.6800 ;
        RECT 682.1200 1810.6400 685.1200 1811.1200 ;
        RECT 682.1200 1816.0800 685.1200 1816.5600 ;
        RECT 693.8800 1794.3200 695.4800 1794.8000 ;
        RECT 693.8800 1799.7600 695.4800 1800.2400 ;
        RECT 682.1200 1794.3200 685.1200 1794.8000 ;
        RECT 682.1200 1799.7600 685.1200 1800.2400 ;
        RECT 886.2200 1778.0000 889.2200 1778.4800 ;
        RECT 886.2200 1783.4400 889.2200 1783.9200 ;
        RECT 886.2200 1788.8800 889.2200 1789.3600 ;
        RECT 873.8800 1778.0000 875.4800 1778.4800 ;
        RECT 873.8800 1783.4400 875.4800 1783.9200 ;
        RECT 873.8800 1788.8800 875.4800 1789.3600 ;
        RECT 886.2200 1767.1200 889.2200 1767.6000 ;
        RECT 886.2200 1772.5600 889.2200 1773.0400 ;
        RECT 873.8800 1767.1200 875.4800 1767.6000 ;
        RECT 873.8800 1772.5600 875.4800 1773.0400 ;
        RECT 886.2200 1750.8000 889.2200 1751.2800 ;
        RECT 886.2200 1756.2400 889.2200 1756.7200 ;
        RECT 886.2200 1761.6800 889.2200 1762.1600 ;
        RECT 873.8800 1750.8000 875.4800 1751.2800 ;
        RECT 873.8800 1756.2400 875.4800 1756.7200 ;
        RECT 873.8800 1761.6800 875.4800 1762.1600 ;
        RECT 886.2200 1739.9200 889.2200 1740.4000 ;
        RECT 886.2200 1745.3600 889.2200 1745.8400 ;
        RECT 873.8800 1739.9200 875.4800 1740.4000 ;
        RECT 873.8800 1745.3600 875.4800 1745.8400 ;
        RECT 828.8800 1778.0000 830.4800 1778.4800 ;
        RECT 828.8800 1783.4400 830.4800 1783.9200 ;
        RECT 828.8800 1788.8800 830.4800 1789.3600 ;
        RECT 828.8800 1767.1200 830.4800 1767.6000 ;
        RECT 828.8800 1772.5600 830.4800 1773.0400 ;
        RECT 828.8800 1750.8000 830.4800 1751.2800 ;
        RECT 828.8800 1756.2400 830.4800 1756.7200 ;
        RECT 828.8800 1761.6800 830.4800 1762.1600 ;
        RECT 828.8800 1739.9200 830.4800 1740.4000 ;
        RECT 828.8800 1745.3600 830.4800 1745.8400 ;
        RECT 886.2200 1723.6000 889.2200 1724.0800 ;
        RECT 886.2200 1729.0400 889.2200 1729.5200 ;
        RECT 886.2200 1734.4800 889.2200 1734.9600 ;
        RECT 873.8800 1723.6000 875.4800 1724.0800 ;
        RECT 873.8800 1729.0400 875.4800 1729.5200 ;
        RECT 873.8800 1734.4800 875.4800 1734.9600 ;
        RECT 886.2200 1712.7200 889.2200 1713.2000 ;
        RECT 886.2200 1718.1600 889.2200 1718.6400 ;
        RECT 873.8800 1712.7200 875.4800 1713.2000 ;
        RECT 873.8800 1718.1600 875.4800 1718.6400 ;
        RECT 886.2200 1696.4000 889.2200 1696.8800 ;
        RECT 886.2200 1701.8400 889.2200 1702.3200 ;
        RECT 886.2200 1707.2800 889.2200 1707.7600 ;
        RECT 873.8800 1696.4000 875.4800 1696.8800 ;
        RECT 873.8800 1701.8400 875.4800 1702.3200 ;
        RECT 873.8800 1707.2800 875.4800 1707.7600 ;
        RECT 886.2200 1690.9600 889.2200 1691.4400 ;
        RECT 873.8800 1690.9600 875.4800 1691.4400 ;
        RECT 828.8800 1723.6000 830.4800 1724.0800 ;
        RECT 828.8800 1729.0400 830.4800 1729.5200 ;
        RECT 828.8800 1734.4800 830.4800 1734.9600 ;
        RECT 828.8800 1712.7200 830.4800 1713.2000 ;
        RECT 828.8800 1718.1600 830.4800 1718.6400 ;
        RECT 828.8800 1696.4000 830.4800 1696.8800 ;
        RECT 828.8800 1701.8400 830.4800 1702.3200 ;
        RECT 828.8800 1707.2800 830.4800 1707.7600 ;
        RECT 828.8800 1690.9600 830.4800 1691.4400 ;
        RECT 783.8800 1778.0000 785.4800 1778.4800 ;
        RECT 783.8800 1783.4400 785.4800 1783.9200 ;
        RECT 783.8800 1788.8800 785.4800 1789.3600 ;
        RECT 783.8800 1767.1200 785.4800 1767.6000 ;
        RECT 783.8800 1772.5600 785.4800 1773.0400 ;
        RECT 738.8800 1778.0000 740.4800 1778.4800 ;
        RECT 738.8800 1783.4400 740.4800 1783.9200 ;
        RECT 738.8800 1788.8800 740.4800 1789.3600 ;
        RECT 738.8800 1767.1200 740.4800 1767.6000 ;
        RECT 738.8800 1772.5600 740.4800 1773.0400 ;
        RECT 783.8800 1750.8000 785.4800 1751.2800 ;
        RECT 783.8800 1756.2400 785.4800 1756.7200 ;
        RECT 783.8800 1761.6800 785.4800 1762.1600 ;
        RECT 783.8800 1739.9200 785.4800 1740.4000 ;
        RECT 783.8800 1745.3600 785.4800 1745.8400 ;
        RECT 738.8800 1750.8000 740.4800 1751.2800 ;
        RECT 738.8800 1756.2400 740.4800 1756.7200 ;
        RECT 738.8800 1761.6800 740.4800 1762.1600 ;
        RECT 738.8800 1739.9200 740.4800 1740.4000 ;
        RECT 738.8800 1745.3600 740.4800 1745.8400 ;
        RECT 693.8800 1778.0000 695.4800 1778.4800 ;
        RECT 693.8800 1783.4400 695.4800 1783.9200 ;
        RECT 693.8800 1788.8800 695.4800 1789.3600 ;
        RECT 682.1200 1778.0000 685.1200 1778.4800 ;
        RECT 682.1200 1783.4400 685.1200 1783.9200 ;
        RECT 682.1200 1788.8800 685.1200 1789.3600 ;
        RECT 693.8800 1767.1200 695.4800 1767.6000 ;
        RECT 693.8800 1772.5600 695.4800 1773.0400 ;
        RECT 682.1200 1767.1200 685.1200 1767.6000 ;
        RECT 682.1200 1772.5600 685.1200 1773.0400 ;
        RECT 693.8800 1750.8000 695.4800 1751.2800 ;
        RECT 693.8800 1756.2400 695.4800 1756.7200 ;
        RECT 693.8800 1761.6800 695.4800 1762.1600 ;
        RECT 682.1200 1750.8000 685.1200 1751.2800 ;
        RECT 682.1200 1756.2400 685.1200 1756.7200 ;
        RECT 682.1200 1761.6800 685.1200 1762.1600 ;
        RECT 693.8800 1739.9200 695.4800 1740.4000 ;
        RECT 693.8800 1745.3600 695.4800 1745.8400 ;
        RECT 682.1200 1739.9200 685.1200 1740.4000 ;
        RECT 682.1200 1745.3600 685.1200 1745.8400 ;
        RECT 783.8800 1723.6000 785.4800 1724.0800 ;
        RECT 783.8800 1729.0400 785.4800 1729.5200 ;
        RECT 783.8800 1734.4800 785.4800 1734.9600 ;
        RECT 783.8800 1712.7200 785.4800 1713.2000 ;
        RECT 783.8800 1718.1600 785.4800 1718.6400 ;
        RECT 738.8800 1723.6000 740.4800 1724.0800 ;
        RECT 738.8800 1729.0400 740.4800 1729.5200 ;
        RECT 738.8800 1734.4800 740.4800 1734.9600 ;
        RECT 738.8800 1712.7200 740.4800 1713.2000 ;
        RECT 738.8800 1718.1600 740.4800 1718.6400 ;
        RECT 783.8800 1696.4000 785.4800 1696.8800 ;
        RECT 783.8800 1701.8400 785.4800 1702.3200 ;
        RECT 783.8800 1707.2800 785.4800 1707.7600 ;
        RECT 783.8800 1690.9600 785.4800 1691.4400 ;
        RECT 738.8800 1696.4000 740.4800 1696.8800 ;
        RECT 738.8800 1701.8400 740.4800 1702.3200 ;
        RECT 738.8800 1707.2800 740.4800 1707.7600 ;
        RECT 738.8800 1690.9600 740.4800 1691.4400 ;
        RECT 693.8800 1723.6000 695.4800 1724.0800 ;
        RECT 693.8800 1729.0400 695.4800 1729.5200 ;
        RECT 693.8800 1734.4800 695.4800 1734.9600 ;
        RECT 682.1200 1723.6000 685.1200 1724.0800 ;
        RECT 682.1200 1729.0400 685.1200 1729.5200 ;
        RECT 682.1200 1734.4800 685.1200 1734.9600 ;
        RECT 693.8800 1712.7200 695.4800 1713.2000 ;
        RECT 693.8800 1718.1600 695.4800 1718.6400 ;
        RECT 682.1200 1712.7200 685.1200 1713.2000 ;
        RECT 682.1200 1718.1600 685.1200 1718.6400 ;
        RECT 693.8800 1696.4000 695.4800 1696.8800 ;
        RECT 693.8800 1701.8400 695.4800 1702.3200 ;
        RECT 693.8800 1707.2800 695.4800 1707.7600 ;
        RECT 682.1200 1696.4000 685.1200 1696.8800 ;
        RECT 682.1200 1701.8400 685.1200 1702.3200 ;
        RECT 682.1200 1707.2800 685.1200 1707.7600 ;
        RECT 682.1200 1690.9600 685.1200 1691.4400 ;
        RECT 693.8800 1690.9600 695.4800 1691.4400 ;
        RECT 682.1200 1895.8700 889.2200 1898.8700 ;
        RECT 682.1200 1682.7700 889.2200 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 1453.1300 875.4800 1669.2300 ;
        RECT 828.8800 1453.1300 830.4800 1669.2300 ;
        RECT 783.8800 1453.1300 785.4800 1669.2300 ;
        RECT 738.8800 1453.1300 740.4800 1669.2300 ;
        RECT 693.8800 1453.1300 695.4800 1669.2300 ;
        RECT 886.2200 1453.1300 889.2200 1669.2300 ;
        RECT 682.1200 1453.1300 685.1200 1669.2300 ;
      LAYER met3 ;
        RECT 886.2200 1646.2800 889.2200 1646.7600 ;
        RECT 886.2200 1651.7200 889.2200 1652.2000 ;
        RECT 873.8800 1646.2800 875.4800 1646.7600 ;
        RECT 873.8800 1651.7200 875.4800 1652.2000 ;
        RECT 886.2200 1657.1600 889.2200 1657.6400 ;
        RECT 873.8800 1657.1600 875.4800 1657.6400 ;
        RECT 886.2200 1635.4000 889.2200 1635.8800 ;
        RECT 886.2200 1640.8400 889.2200 1641.3200 ;
        RECT 873.8800 1635.4000 875.4800 1635.8800 ;
        RECT 873.8800 1640.8400 875.4800 1641.3200 ;
        RECT 886.2200 1619.0800 889.2200 1619.5600 ;
        RECT 886.2200 1624.5200 889.2200 1625.0000 ;
        RECT 873.8800 1619.0800 875.4800 1619.5600 ;
        RECT 873.8800 1624.5200 875.4800 1625.0000 ;
        RECT 886.2200 1629.9600 889.2200 1630.4400 ;
        RECT 873.8800 1629.9600 875.4800 1630.4400 ;
        RECT 828.8800 1646.2800 830.4800 1646.7600 ;
        RECT 828.8800 1651.7200 830.4800 1652.2000 ;
        RECT 828.8800 1657.1600 830.4800 1657.6400 ;
        RECT 828.8800 1635.4000 830.4800 1635.8800 ;
        RECT 828.8800 1640.8400 830.4800 1641.3200 ;
        RECT 828.8800 1619.0800 830.4800 1619.5600 ;
        RECT 828.8800 1624.5200 830.4800 1625.0000 ;
        RECT 828.8800 1629.9600 830.4800 1630.4400 ;
        RECT 886.2200 1602.7600 889.2200 1603.2400 ;
        RECT 886.2200 1608.2000 889.2200 1608.6800 ;
        RECT 886.2200 1613.6400 889.2200 1614.1200 ;
        RECT 873.8800 1602.7600 875.4800 1603.2400 ;
        RECT 873.8800 1608.2000 875.4800 1608.6800 ;
        RECT 873.8800 1613.6400 875.4800 1614.1200 ;
        RECT 886.2200 1591.8800 889.2200 1592.3600 ;
        RECT 886.2200 1597.3200 889.2200 1597.8000 ;
        RECT 873.8800 1591.8800 875.4800 1592.3600 ;
        RECT 873.8800 1597.3200 875.4800 1597.8000 ;
        RECT 886.2200 1575.5600 889.2200 1576.0400 ;
        RECT 886.2200 1581.0000 889.2200 1581.4800 ;
        RECT 886.2200 1586.4400 889.2200 1586.9200 ;
        RECT 873.8800 1575.5600 875.4800 1576.0400 ;
        RECT 873.8800 1581.0000 875.4800 1581.4800 ;
        RECT 873.8800 1586.4400 875.4800 1586.9200 ;
        RECT 886.2200 1564.6800 889.2200 1565.1600 ;
        RECT 886.2200 1570.1200 889.2200 1570.6000 ;
        RECT 873.8800 1564.6800 875.4800 1565.1600 ;
        RECT 873.8800 1570.1200 875.4800 1570.6000 ;
        RECT 828.8800 1602.7600 830.4800 1603.2400 ;
        RECT 828.8800 1608.2000 830.4800 1608.6800 ;
        RECT 828.8800 1613.6400 830.4800 1614.1200 ;
        RECT 828.8800 1591.8800 830.4800 1592.3600 ;
        RECT 828.8800 1597.3200 830.4800 1597.8000 ;
        RECT 828.8800 1575.5600 830.4800 1576.0400 ;
        RECT 828.8800 1581.0000 830.4800 1581.4800 ;
        RECT 828.8800 1586.4400 830.4800 1586.9200 ;
        RECT 828.8800 1564.6800 830.4800 1565.1600 ;
        RECT 828.8800 1570.1200 830.4800 1570.6000 ;
        RECT 783.8800 1646.2800 785.4800 1646.7600 ;
        RECT 783.8800 1651.7200 785.4800 1652.2000 ;
        RECT 783.8800 1657.1600 785.4800 1657.6400 ;
        RECT 738.8800 1646.2800 740.4800 1646.7600 ;
        RECT 738.8800 1651.7200 740.4800 1652.2000 ;
        RECT 738.8800 1657.1600 740.4800 1657.6400 ;
        RECT 783.8800 1635.4000 785.4800 1635.8800 ;
        RECT 783.8800 1640.8400 785.4800 1641.3200 ;
        RECT 783.8800 1619.0800 785.4800 1619.5600 ;
        RECT 783.8800 1624.5200 785.4800 1625.0000 ;
        RECT 783.8800 1629.9600 785.4800 1630.4400 ;
        RECT 738.8800 1635.4000 740.4800 1635.8800 ;
        RECT 738.8800 1640.8400 740.4800 1641.3200 ;
        RECT 738.8800 1619.0800 740.4800 1619.5600 ;
        RECT 738.8800 1624.5200 740.4800 1625.0000 ;
        RECT 738.8800 1629.9600 740.4800 1630.4400 ;
        RECT 693.8800 1646.2800 695.4800 1646.7600 ;
        RECT 693.8800 1651.7200 695.4800 1652.2000 ;
        RECT 682.1200 1651.7200 685.1200 1652.2000 ;
        RECT 682.1200 1646.2800 685.1200 1646.7600 ;
        RECT 682.1200 1657.1600 685.1200 1657.6400 ;
        RECT 693.8800 1657.1600 695.4800 1657.6400 ;
        RECT 693.8800 1635.4000 695.4800 1635.8800 ;
        RECT 693.8800 1640.8400 695.4800 1641.3200 ;
        RECT 682.1200 1640.8400 685.1200 1641.3200 ;
        RECT 682.1200 1635.4000 685.1200 1635.8800 ;
        RECT 693.8800 1619.0800 695.4800 1619.5600 ;
        RECT 693.8800 1624.5200 695.4800 1625.0000 ;
        RECT 682.1200 1624.5200 685.1200 1625.0000 ;
        RECT 682.1200 1619.0800 685.1200 1619.5600 ;
        RECT 682.1200 1629.9600 685.1200 1630.4400 ;
        RECT 693.8800 1629.9600 695.4800 1630.4400 ;
        RECT 783.8800 1602.7600 785.4800 1603.2400 ;
        RECT 783.8800 1608.2000 785.4800 1608.6800 ;
        RECT 783.8800 1613.6400 785.4800 1614.1200 ;
        RECT 783.8800 1591.8800 785.4800 1592.3600 ;
        RECT 783.8800 1597.3200 785.4800 1597.8000 ;
        RECT 738.8800 1602.7600 740.4800 1603.2400 ;
        RECT 738.8800 1608.2000 740.4800 1608.6800 ;
        RECT 738.8800 1613.6400 740.4800 1614.1200 ;
        RECT 738.8800 1591.8800 740.4800 1592.3600 ;
        RECT 738.8800 1597.3200 740.4800 1597.8000 ;
        RECT 783.8800 1575.5600 785.4800 1576.0400 ;
        RECT 783.8800 1581.0000 785.4800 1581.4800 ;
        RECT 783.8800 1586.4400 785.4800 1586.9200 ;
        RECT 783.8800 1564.6800 785.4800 1565.1600 ;
        RECT 783.8800 1570.1200 785.4800 1570.6000 ;
        RECT 738.8800 1575.5600 740.4800 1576.0400 ;
        RECT 738.8800 1581.0000 740.4800 1581.4800 ;
        RECT 738.8800 1586.4400 740.4800 1586.9200 ;
        RECT 738.8800 1564.6800 740.4800 1565.1600 ;
        RECT 738.8800 1570.1200 740.4800 1570.6000 ;
        RECT 693.8800 1602.7600 695.4800 1603.2400 ;
        RECT 693.8800 1608.2000 695.4800 1608.6800 ;
        RECT 693.8800 1613.6400 695.4800 1614.1200 ;
        RECT 682.1200 1602.7600 685.1200 1603.2400 ;
        RECT 682.1200 1608.2000 685.1200 1608.6800 ;
        RECT 682.1200 1613.6400 685.1200 1614.1200 ;
        RECT 693.8800 1591.8800 695.4800 1592.3600 ;
        RECT 693.8800 1597.3200 695.4800 1597.8000 ;
        RECT 682.1200 1591.8800 685.1200 1592.3600 ;
        RECT 682.1200 1597.3200 685.1200 1597.8000 ;
        RECT 693.8800 1575.5600 695.4800 1576.0400 ;
        RECT 693.8800 1581.0000 695.4800 1581.4800 ;
        RECT 693.8800 1586.4400 695.4800 1586.9200 ;
        RECT 682.1200 1575.5600 685.1200 1576.0400 ;
        RECT 682.1200 1581.0000 685.1200 1581.4800 ;
        RECT 682.1200 1586.4400 685.1200 1586.9200 ;
        RECT 693.8800 1564.6800 695.4800 1565.1600 ;
        RECT 693.8800 1570.1200 695.4800 1570.6000 ;
        RECT 682.1200 1564.6800 685.1200 1565.1600 ;
        RECT 682.1200 1570.1200 685.1200 1570.6000 ;
        RECT 886.2200 1548.3600 889.2200 1548.8400 ;
        RECT 886.2200 1553.8000 889.2200 1554.2800 ;
        RECT 886.2200 1559.2400 889.2200 1559.7200 ;
        RECT 873.8800 1548.3600 875.4800 1548.8400 ;
        RECT 873.8800 1553.8000 875.4800 1554.2800 ;
        RECT 873.8800 1559.2400 875.4800 1559.7200 ;
        RECT 886.2200 1537.4800 889.2200 1537.9600 ;
        RECT 886.2200 1542.9200 889.2200 1543.4000 ;
        RECT 873.8800 1537.4800 875.4800 1537.9600 ;
        RECT 873.8800 1542.9200 875.4800 1543.4000 ;
        RECT 886.2200 1521.1600 889.2200 1521.6400 ;
        RECT 886.2200 1526.6000 889.2200 1527.0800 ;
        RECT 886.2200 1532.0400 889.2200 1532.5200 ;
        RECT 873.8800 1521.1600 875.4800 1521.6400 ;
        RECT 873.8800 1526.6000 875.4800 1527.0800 ;
        RECT 873.8800 1532.0400 875.4800 1532.5200 ;
        RECT 886.2200 1510.2800 889.2200 1510.7600 ;
        RECT 886.2200 1515.7200 889.2200 1516.2000 ;
        RECT 873.8800 1510.2800 875.4800 1510.7600 ;
        RECT 873.8800 1515.7200 875.4800 1516.2000 ;
        RECT 828.8800 1548.3600 830.4800 1548.8400 ;
        RECT 828.8800 1553.8000 830.4800 1554.2800 ;
        RECT 828.8800 1559.2400 830.4800 1559.7200 ;
        RECT 828.8800 1537.4800 830.4800 1537.9600 ;
        RECT 828.8800 1542.9200 830.4800 1543.4000 ;
        RECT 828.8800 1521.1600 830.4800 1521.6400 ;
        RECT 828.8800 1526.6000 830.4800 1527.0800 ;
        RECT 828.8800 1532.0400 830.4800 1532.5200 ;
        RECT 828.8800 1510.2800 830.4800 1510.7600 ;
        RECT 828.8800 1515.7200 830.4800 1516.2000 ;
        RECT 886.2200 1493.9600 889.2200 1494.4400 ;
        RECT 886.2200 1499.4000 889.2200 1499.8800 ;
        RECT 886.2200 1504.8400 889.2200 1505.3200 ;
        RECT 873.8800 1493.9600 875.4800 1494.4400 ;
        RECT 873.8800 1499.4000 875.4800 1499.8800 ;
        RECT 873.8800 1504.8400 875.4800 1505.3200 ;
        RECT 886.2200 1483.0800 889.2200 1483.5600 ;
        RECT 886.2200 1488.5200 889.2200 1489.0000 ;
        RECT 873.8800 1483.0800 875.4800 1483.5600 ;
        RECT 873.8800 1488.5200 875.4800 1489.0000 ;
        RECT 886.2200 1466.7600 889.2200 1467.2400 ;
        RECT 886.2200 1472.2000 889.2200 1472.6800 ;
        RECT 886.2200 1477.6400 889.2200 1478.1200 ;
        RECT 873.8800 1466.7600 875.4800 1467.2400 ;
        RECT 873.8800 1472.2000 875.4800 1472.6800 ;
        RECT 873.8800 1477.6400 875.4800 1478.1200 ;
        RECT 886.2200 1461.3200 889.2200 1461.8000 ;
        RECT 873.8800 1461.3200 875.4800 1461.8000 ;
        RECT 828.8800 1493.9600 830.4800 1494.4400 ;
        RECT 828.8800 1499.4000 830.4800 1499.8800 ;
        RECT 828.8800 1504.8400 830.4800 1505.3200 ;
        RECT 828.8800 1483.0800 830.4800 1483.5600 ;
        RECT 828.8800 1488.5200 830.4800 1489.0000 ;
        RECT 828.8800 1466.7600 830.4800 1467.2400 ;
        RECT 828.8800 1472.2000 830.4800 1472.6800 ;
        RECT 828.8800 1477.6400 830.4800 1478.1200 ;
        RECT 828.8800 1461.3200 830.4800 1461.8000 ;
        RECT 783.8800 1548.3600 785.4800 1548.8400 ;
        RECT 783.8800 1553.8000 785.4800 1554.2800 ;
        RECT 783.8800 1559.2400 785.4800 1559.7200 ;
        RECT 783.8800 1537.4800 785.4800 1537.9600 ;
        RECT 783.8800 1542.9200 785.4800 1543.4000 ;
        RECT 738.8800 1548.3600 740.4800 1548.8400 ;
        RECT 738.8800 1553.8000 740.4800 1554.2800 ;
        RECT 738.8800 1559.2400 740.4800 1559.7200 ;
        RECT 738.8800 1537.4800 740.4800 1537.9600 ;
        RECT 738.8800 1542.9200 740.4800 1543.4000 ;
        RECT 783.8800 1521.1600 785.4800 1521.6400 ;
        RECT 783.8800 1526.6000 785.4800 1527.0800 ;
        RECT 783.8800 1532.0400 785.4800 1532.5200 ;
        RECT 783.8800 1510.2800 785.4800 1510.7600 ;
        RECT 783.8800 1515.7200 785.4800 1516.2000 ;
        RECT 738.8800 1521.1600 740.4800 1521.6400 ;
        RECT 738.8800 1526.6000 740.4800 1527.0800 ;
        RECT 738.8800 1532.0400 740.4800 1532.5200 ;
        RECT 738.8800 1510.2800 740.4800 1510.7600 ;
        RECT 738.8800 1515.7200 740.4800 1516.2000 ;
        RECT 693.8800 1548.3600 695.4800 1548.8400 ;
        RECT 693.8800 1553.8000 695.4800 1554.2800 ;
        RECT 693.8800 1559.2400 695.4800 1559.7200 ;
        RECT 682.1200 1548.3600 685.1200 1548.8400 ;
        RECT 682.1200 1553.8000 685.1200 1554.2800 ;
        RECT 682.1200 1559.2400 685.1200 1559.7200 ;
        RECT 693.8800 1537.4800 695.4800 1537.9600 ;
        RECT 693.8800 1542.9200 695.4800 1543.4000 ;
        RECT 682.1200 1537.4800 685.1200 1537.9600 ;
        RECT 682.1200 1542.9200 685.1200 1543.4000 ;
        RECT 693.8800 1521.1600 695.4800 1521.6400 ;
        RECT 693.8800 1526.6000 695.4800 1527.0800 ;
        RECT 693.8800 1532.0400 695.4800 1532.5200 ;
        RECT 682.1200 1521.1600 685.1200 1521.6400 ;
        RECT 682.1200 1526.6000 685.1200 1527.0800 ;
        RECT 682.1200 1532.0400 685.1200 1532.5200 ;
        RECT 693.8800 1510.2800 695.4800 1510.7600 ;
        RECT 693.8800 1515.7200 695.4800 1516.2000 ;
        RECT 682.1200 1510.2800 685.1200 1510.7600 ;
        RECT 682.1200 1515.7200 685.1200 1516.2000 ;
        RECT 783.8800 1493.9600 785.4800 1494.4400 ;
        RECT 783.8800 1499.4000 785.4800 1499.8800 ;
        RECT 783.8800 1504.8400 785.4800 1505.3200 ;
        RECT 783.8800 1483.0800 785.4800 1483.5600 ;
        RECT 783.8800 1488.5200 785.4800 1489.0000 ;
        RECT 738.8800 1493.9600 740.4800 1494.4400 ;
        RECT 738.8800 1499.4000 740.4800 1499.8800 ;
        RECT 738.8800 1504.8400 740.4800 1505.3200 ;
        RECT 738.8800 1483.0800 740.4800 1483.5600 ;
        RECT 738.8800 1488.5200 740.4800 1489.0000 ;
        RECT 783.8800 1466.7600 785.4800 1467.2400 ;
        RECT 783.8800 1472.2000 785.4800 1472.6800 ;
        RECT 783.8800 1477.6400 785.4800 1478.1200 ;
        RECT 783.8800 1461.3200 785.4800 1461.8000 ;
        RECT 738.8800 1466.7600 740.4800 1467.2400 ;
        RECT 738.8800 1472.2000 740.4800 1472.6800 ;
        RECT 738.8800 1477.6400 740.4800 1478.1200 ;
        RECT 738.8800 1461.3200 740.4800 1461.8000 ;
        RECT 693.8800 1493.9600 695.4800 1494.4400 ;
        RECT 693.8800 1499.4000 695.4800 1499.8800 ;
        RECT 693.8800 1504.8400 695.4800 1505.3200 ;
        RECT 682.1200 1493.9600 685.1200 1494.4400 ;
        RECT 682.1200 1499.4000 685.1200 1499.8800 ;
        RECT 682.1200 1504.8400 685.1200 1505.3200 ;
        RECT 693.8800 1483.0800 695.4800 1483.5600 ;
        RECT 693.8800 1488.5200 695.4800 1489.0000 ;
        RECT 682.1200 1483.0800 685.1200 1483.5600 ;
        RECT 682.1200 1488.5200 685.1200 1489.0000 ;
        RECT 693.8800 1466.7600 695.4800 1467.2400 ;
        RECT 693.8800 1472.2000 695.4800 1472.6800 ;
        RECT 693.8800 1477.6400 695.4800 1478.1200 ;
        RECT 682.1200 1466.7600 685.1200 1467.2400 ;
        RECT 682.1200 1472.2000 685.1200 1472.6800 ;
        RECT 682.1200 1477.6400 685.1200 1478.1200 ;
        RECT 682.1200 1461.3200 685.1200 1461.8000 ;
        RECT 693.8800 1461.3200 695.4800 1461.8000 ;
        RECT 682.1200 1666.2300 889.2200 1669.2300 ;
        RECT 682.1200 1453.1300 889.2200 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 1223.4900 875.4800 1439.5900 ;
        RECT 828.8800 1223.4900 830.4800 1439.5900 ;
        RECT 783.8800 1223.4900 785.4800 1439.5900 ;
        RECT 738.8800 1223.4900 740.4800 1439.5900 ;
        RECT 693.8800 1223.4900 695.4800 1439.5900 ;
        RECT 886.2200 1223.4900 889.2200 1439.5900 ;
        RECT 682.1200 1223.4900 685.1200 1439.5900 ;
      LAYER met3 ;
        RECT 886.2200 1416.6400 889.2200 1417.1200 ;
        RECT 886.2200 1422.0800 889.2200 1422.5600 ;
        RECT 873.8800 1416.6400 875.4800 1417.1200 ;
        RECT 873.8800 1422.0800 875.4800 1422.5600 ;
        RECT 886.2200 1427.5200 889.2200 1428.0000 ;
        RECT 873.8800 1427.5200 875.4800 1428.0000 ;
        RECT 886.2200 1405.7600 889.2200 1406.2400 ;
        RECT 886.2200 1411.2000 889.2200 1411.6800 ;
        RECT 873.8800 1405.7600 875.4800 1406.2400 ;
        RECT 873.8800 1411.2000 875.4800 1411.6800 ;
        RECT 886.2200 1389.4400 889.2200 1389.9200 ;
        RECT 886.2200 1394.8800 889.2200 1395.3600 ;
        RECT 873.8800 1389.4400 875.4800 1389.9200 ;
        RECT 873.8800 1394.8800 875.4800 1395.3600 ;
        RECT 886.2200 1400.3200 889.2200 1400.8000 ;
        RECT 873.8800 1400.3200 875.4800 1400.8000 ;
        RECT 828.8800 1416.6400 830.4800 1417.1200 ;
        RECT 828.8800 1422.0800 830.4800 1422.5600 ;
        RECT 828.8800 1427.5200 830.4800 1428.0000 ;
        RECT 828.8800 1405.7600 830.4800 1406.2400 ;
        RECT 828.8800 1411.2000 830.4800 1411.6800 ;
        RECT 828.8800 1389.4400 830.4800 1389.9200 ;
        RECT 828.8800 1394.8800 830.4800 1395.3600 ;
        RECT 828.8800 1400.3200 830.4800 1400.8000 ;
        RECT 886.2200 1373.1200 889.2200 1373.6000 ;
        RECT 886.2200 1378.5600 889.2200 1379.0400 ;
        RECT 886.2200 1384.0000 889.2200 1384.4800 ;
        RECT 873.8800 1373.1200 875.4800 1373.6000 ;
        RECT 873.8800 1378.5600 875.4800 1379.0400 ;
        RECT 873.8800 1384.0000 875.4800 1384.4800 ;
        RECT 886.2200 1362.2400 889.2200 1362.7200 ;
        RECT 886.2200 1367.6800 889.2200 1368.1600 ;
        RECT 873.8800 1362.2400 875.4800 1362.7200 ;
        RECT 873.8800 1367.6800 875.4800 1368.1600 ;
        RECT 886.2200 1345.9200 889.2200 1346.4000 ;
        RECT 886.2200 1351.3600 889.2200 1351.8400 ;
        RECT 886.2200 1356.8000 889.2200 1357.2800 ;
        RECT 873.8800 1345.9200 875.4800 1346.4000 ;
        RECT 873.8800 1351.3600 875.4800 1351.8400 ;
        RECT 873.8800 1356.8000 875.4800 1357.2800 ;
        RECT 886.2200 1335.0400 889.2200 1335.5200 ;
        RECT 886.2200 1340.4800 889.2200 1340.9600 ;
        RECT 873.8800 1335.0400 875.4800 1335.5200 ;
        RECT 873.8800 1340.4800 875.4800 1340.9600 ;
        RECT 828.8800 1373.1200 830.4800 1373.6000 ;
        RECT 828.8800 1378.5600 830.4800 1379.0400 ;
        RECT 828.8800 1384.0000 830.4800 1384.4800 ;
        RECT 828.8800 1362.2400 830.4800 1362.7200 ;
        RECT 828.8800 1367.6800 830.4800 1368.1600 ;
        RECT 828.8800 1345.9200 830.4800 1346.4000 ;
        RECT 828.8800 1351.3600 830.4800 1351.8400 ;
        RECT 828.8800 1356.8000 830.4800 1357.2800 ;
        RECT 828.8800 1335.0400 830.4800 1335.5200 ;
        RECT 828.8800 1340.4800 830.4800 1340.9600 ;
        RECT 783.8800 1416.6400 785.4800 1417.1200 ;
        RECT 783.8800 1422.0800 785.4800 1422.5600 ;
        RECT 783.8800 1427.5200 785.4800 1428.0000 ;
        RECT 738.8800 1416.6400 740.4800 1417.1200 ;
        RECT 738.8800 1422.0800 740.4800 1422.5600 ;
        RECT 738.8800 1427.5200 740.4800 1428.0000 ;
        RECT 783.8800 1405.7600 785.4800 1406.2400 ;
        RECT 783.8800 1411.2000 785.4800 1411.6800 ;
        RECT 783.8800 1389.4400 785.4800 1389.9200 ;
        RECT 783.8800 1394.8800 785.4800 1395.3600 ;
        RECT 783.8800 1400.3200 785.4800 1400.8000 ;
        RECT 738.8800 1405.7600 740.4800 1406.2400 ;
        RECT 738.8800 1411.2000 740.4800 1411.6800 ;
        RECT 738.8800 1389.4400 740.4800 1389.9200 ;
        RECT 738.8800 1394.8800 740.4800 1395.3600 ;
        RECT 738.8800 1400.3200 740.4800 1400.8000 ;
        RECT 693.8800 1416.6400 695.4800 1417.1200 ;
        RECT 693.8800 1422.0800 695.4800 1422.5600 ;
        RECT 682.1200 1422.0800 685.1200 1422.5600 ;
        RECT 682.1200 1416.6400 685.1200 1417.1200 ;
        RECT 682.1200 1427.5200 685.1200 1428.0000 ;
        RECT 693.8800 1427.5200 695.4800 1428.0000 ;
        RECT 693.8800 1405.7600 695.4800 1406.2400 ;
        RECT 693.8800 1411.2000 695.4800 1411.6800 ;
        RECT 682.1200 1411.2000 685.1200 1411.6800 ;
        RECT 682.1200 1405.7600 685.1200 1406.2400 ;
        RECT 693.8800 1389.4400 695.4800 1389.9200 ;
        RECT 693.8800 1394.8800 695.4800 1395.3600 ;
        RECT 682.1200 1394.8800 685.1200 1395.3600 ;
        RECT 682.1200 1389.4400 685.1200 1389.9200 ;
        RECT 682.1200 1400.3200 685.1200 1400.8000 ;
        RECT 693.8800 1400.3200 695.4800 1400.8000 ;
        RECT 783.8800 1373.1200 785.4800 1373.6000 ;
        RECT 783.8800 1378.5600 785.4800 1379.0400 ;
        RECT 783.8800 1384.0000 785.4800 1384.4800 ;
        RECT 783.8800 1362.2400 785.4800 1362.7200 ;
        RECT 783.8800 1367.6800 785.4800 1368.1600 ;
        RECT 738.8800 1373.1200 740.4800 1373.6000 ;
        RECT 738.8800 1378.5600 740.4800 1379.0400 ;
        RECT 738.8800 1384.0000 740.4800 1384.4800 ;
        RECT 738.8800 1362.2400 740.4800 1362.7200 ;
        RECT 738.8800 1367.6800 740.4800 1368.1600 ;
        RECT 783.8800 1345.9200 785.4800 1346.4000 ;
        RECT 783.8800 1351.3600 785.4800 1351.8400 ;
        RECT 783.8800 1356.8000 785.4800 1357.2800 ;
        RECT 783.8800 1335.0400 785.4800 1335.5200 ;
        RECT 783.8800 1340.4800 785.4800 1340.9600 ;
        RECT 738.8800 1345.9200 740.4800 1346.4000 ;
        RECT 738.8800 1351.3600 740.4800 1351.8400 ;
        RECT 738.8800 1356.8000 740.4800 1357.2800 ;
        RECT 738.8800 1335.0400 740.4800 1335.5200 ;
        RECT 738.8800 1340.4800 740.4800 1340.9600 ;
        RECT 693.8800 1373.1200 695.4800 1373.6000 ;
        RECT 693.8800 1378.5600 695.4800 1379.0400 ;
        RECT 693.8800 1384.0000 695.4800 1384.4800 ;
        RECT 682.1200 1373.1200 685.1200 1373.6000 ;
        RECT 682.1200 1378.5600 685.1200 1379.0400 ;
        RECT 682.1200 1384.0000 685.1200 1384.4800 ;
        RECT 693.8800 1362.2400 695.4800 1362.7200 ;
        RECT 693.8800 1367.6800 695.4800 1368.1600 ;
        RECT 682.1200 1362.2400 685.1200 1362.7200 ;
        RECT 682.1200 1367.6800 685.1200 1368.1600 ;
        RECT 693.8800 1345.9200 695.4800 1346.4000 ;
        RECT 693.8800 1351.3600 695.4800 1351.8400 ;
        RECT 693.8800 1356.8000 695.4800 1357.2800 ;
        RECT 682.1200 1345.9200 685.1200 1346.4000 ;
        RECT 682.1200 1351.3600 685.1200 1351.8400 ;
        RECT 682.1200 1356.8000 685.1200 1357.2800 ;
        RECT 693.8800 1335.0400 695.4800 1335.5200 ;
        RECT 693.8800 1340.4800 695.4800 1340.9600 ;
        RECT 682.1200 1335.0400 685.1200 1335.5200 ;
        RECT 682.1200 1340.4800 685.1200 1340.9600 ;
        RECT 886.2200 1318.7200 889.2200 1319.2000 ;
        RECT 886.2200 1324.1600 889.2200 1324.6400 ;
        RECT 886.2200 1329.6000 889.2200 1330.0800 ;
        RECT 873.8800 1318.7200 875.4800 1319.2000 ;
        RECT 873.8800 1324.1600 875.4800 1324.6400 ;
        RECT 873.8800 1329.6000 875.4800 1330.0800 ;
        RECT 886.2200 1307.8400 889.2200 1308.3200 ;
        RECT 886.2200 1313.2800 889.2200 1313.7600 ;
        RECT 873.8800 1307.8400 875.4800 1308.3200 ;
        RECT 873.8800 1313.2800 875.4800 1313.7600 ;
        RECT 886.2200 1291.5200 889.2200 1292.0000 ;
        RECT 886.2200 1296.9600 889.2200 1297.4400 ;
        RECT 886.2200 1302.4000 889.2200 1302.8800 ;
        RECT 873.8800 1291.5200 875.4800 1292.0000 ;
        RECT 873.8800 1296.9600 875.4800 1297.4400 ;
        RECT 873.8800 1302.4000 875.4800 1302.8800 ;
        RECT 886.2200 1280.6400 889.2200 1281.1200 ;
        RECT 886.2200 1286.0800 889.2200 1286.5600 ;
        RECT 873.8800 1280.6400 875.4800 1281.1200 ;
        RECT 873.8800 1286.0800 875.4800 1286.5600 ;
        RECT 828.8800 1318.7200 830.4800 1319.2000 ;
        RECT 828.8800 1324.1600 830.4800 1324.6400 ;
        RECT 828.8800 1329.6000 830.4800 1330.0800 ;
        RECT 828.8800 1307.8400 830.4800 1308.3200 ;
        RECT 828.8800 1313.2800 830.4800 1313.7600 ;
        RECT 828.8800 1291.5200 830.4800 1292.0000 ;
        RECT 828.8800 1296.9600 830.4800 1297.4400 ;
        RECT 828.8800 1302.4000 830.4800 1302.8800 ;
        RECT 828.8800 1280.6400 830.4800 1281.1200 ;
        RECT 828.8800 1286.0800 830.4800 1286.5600 ;
        RECT 886.2200 1264.3200 889.2200 1264.8000 ;
        RECT 886.2200 1269.7600 889.2200 1270.2400 ;
        RECT 886.2200 1275.2000 889.2200 1275.6800 ;
        RECT 873.8800 1264.3200 875.4800 1264.8000 ;
        RECT 873.8800 1269.7600 875.4800 1270.2400 ;
        RECT 873.8800 1275.2000 875.4800 1275.6800 ;
        RECT 886.2200 1253.4400 889.2200 1253.9200 ;
        RECT 886.2200 1258.8800 889.2200 1259.3600 ;
        RECT 873.8800 1253.4400 875.4800 1253.9200 ;
        RECT 873.8800 1258.8800 875.4800 1259.3600 ;
        RECT 886.2200 1237.1200 889.2200 1237.6000 ;
        RECT 886.2200 1242.5600 889.2200 1243.0400 ;
        RECT 886.2200 1248.0000 889.2200 1248.4800 ;
        RECT 873.8800 1237.1200 875.4800 1237.6000 ;
        RECT 873.8800 1242.5600 875.4800 1243.0400 ;
        RECT 873.8800 1248.0000 875.4800 1248.4800 ;
        RECT 886.2200 1231.6800 889.2200 1232.1600 ;
        RECT 873.8800 1231.6800 875.4800 1232.1600 ;
        RECT 828.8800 1264.3200 830.4800 1264.8000 ;
        RECT 828.8800 1269.7600 830.4800 1270.2400 ;
        RECT 828.8800 1275.2000 830.4800 1275.6800 ;
        RECT 828.8800 1253.4400 830.4800 1253.9200 ;
        RECT 828.8800 1258.8800 830.4800 1259.3600 ;
        RECT 828.8800 1237.1200 830.4800 1237.6000 ;
        RECT 828.8800 1242.5600 830.4800 1243.0400 ;
        RECT 828.8800 1248.0000 830.4800 1248.4800 ;
        RECT 828.8800 1231.6800 830.4800 1232.1600 ;
        RECT 783.8800 1318.7200 785.4800 1319.2000 ;
        RECT 783.8800 1324.1600 785.4800 1324.6400 ;
        RECT 783.8800 1329.6000 785.4800 1330.0800 ;
        RECT 783.8800 1307.8400 785.4800 1308.3200 ;
        RECT 783.8800 1313.2800 785.4800 1313.7600 ;
        RECT 738.8800 1318.7200 740.4800 1319.2000 ;
        RECT 738.8800 1324.1600 740.4800 1324.6400 ;
        RECT 738.8800 1329.6000 740.4800 1330.0800 ;
        RECT 738.8800 1307.8400 740.4800 1308.3200 ;
        RECT 738.8800 1313.2800 740.4800 1313.7600 ;
        RECT 783.8800 1291.5200 785.4800 1292.0000 ;
        RECT 783.8800 1296.9600 785.4800 1297.4400 ;
        RECT 783.8800 1302.4000 785.4800 1302.8800 ;
        RECT 783.8800 1280.6400 785.4800 1281.1200 ;
        RECT 783.8800 1286.0800 785.4800 1286.5600 ;
        RECT 738.8800 1291.5200 740.4800 1292.0000 ;
        RECT 738.8800 1296.9600 740.4800 1297.4400 ;
        RECT 738.8800 1302.4000 740.4800 1302.8800 ;
        RECT 738.8800 1280.6400 740.4800 1281.1200 ;
        RECT 738.8800 1286.0800 740.4800 1286.5600 ;
        RECT 693.8800 1318.7200 695.4800 1319.2000 ;
        RECT 693.8800 1324.1600 695.4800 1324.6400 ;
        RECT 693.8800 1329.6000 695.4800 1330.0800 ;
        RECT 682.1200 1318.7200 685.1200 1319.2000 ;
        RECT 682.1200 1324.1600 685.1200 1324.6400 ;
        RECT 682.1200 1329.6000 685.1200 1330.0800 ;
        RECT 693.8800 1307.8400 695.4800 1308.3200 ;
        RECT 693.8800 1313.2800 695.4800 1313.7600 ;
        RECT 682.1200 1307.8400 685.1200 1308.3200 ;
        RECT 682.1200 1313.2800 685.1200 1313.7600 ;
        RECT 693.8800 1291.5200 695.4800 1292.0000 ;
        RECT 693.8800 1296.9600 695.4800 1297.4400 ;
        RECT 693.8800 1302.4000 695.4800 1302.8800 ;
        RECT 682.1200 1291.5200 685.1200 1292.0000 ;
        RECT 682.1200 1296.9600 685.1200 1297.4400 ;
        RECT 682.1200 1302.4000 685.1200 1302.8800 ;
        RECT 693.8800 1280.6400 695.4800 1281.1200 ;
        RECT 693.8800 1286.0800 695.4800 1286.5600 ;
        RECT 682.1200 1280.6400 685.1200 1281.1200 ;
        RECT 682.1200 1286.0800 685.1200 1286.5600 ;
        RECT 783.8800 1264.3200 785.4800 1264.8000 ;
        RECT 783.8800 1269.7600 785.4800 1270.2400 ;
        RECT 783.8800 1275.2000 785.4800 1275.6800 ;
        RECT 783.8800 1253.4400 785.4800 1253.9200 ;
        RECT 783.8800 1258.8800 785.4800 1259.3600 ;
        RECT 738.8800 1264.3200 740.4800 1264.8000 ;
        RECT 738.8800 1269.7600 740.4800 1270.2400 ;
        RECT 738.8800 1275.2000 740.4800 1275.6800 ;
        RECT 738.8800 1253.4400 740.4800 1253.9200 ;
        RECT 738.8800 1258.8800 740.4800 1259.3600 ;
        RECT 783.8800 1237.1200 785.4800 1237.6000 ;
        RECT 783.8800 1242.5600 785.4800 1243.0400 ;
        RECT 783.8800 1248.0000 785.4800 1248.4800 ;
        RECT 783.8800 1231.6800 785.4800 1232.1600 ;
        RECT 738.8800 1237.1200 740.4800 1237.6000 ;
        RECT 738.8800 1242.5600 740.4800 1243.0400 ;
        RECT 738.8800 1248.0000 740.4800 1248.4800 ;
        RECT 738.8800 1231.6800 740.4800 1232.1600 ;
        RECT 693.8800 1264.3200 695.4800 1264.8000 ;
        RECT 693.8800 1269.7600 695.4800 1270.2400 ;
        RECT 693.8800 1275.2000 695.4800 1275.6800 ;
        RECT 682.1200 1264.3200 685.1200 1264.8000 ;
        RECT 682.1200 1269.7600 685.1200 1270.2400 ;
        RECT 682.1200 1275.2000 685.1200 1275.6800 ;
        RECT 693.8800 1253.4400 695.4800 1253.9200 ;
        RECT 693.8800 1258.8800 695.4800 1259.3600 ;
        RECT 682.1200 1253.4400 685.1200 1253.9200 ;
        RECT 682.1200 1258.8800 685.1200 1259.3600 ;
        RECT 693.8800 1237.1200 695.4800 1237.6000 ;
        RECT 693.8800 1242.5600 695.4800 1243.0400 ;
        RECT 693.8800 1248.0000 695.4800 1248.4800 ;
        RECT 682.1200 1237.1200 685.1200 1237.6000 ;
        RECT 682.1200 1242.5600 685.1200 1243.0400 ;
        RECT 682.1200 1248.0000 685.1200 1248.4800 ;
        RECT 682.1200 1231.6800 685.1200 1232.1600 ;
        RECT 693.8800 1231.6800 695.4800 1232.1600 ;
        RECT 682.1200 1436.5900 889.2200 1439.5900 ;
        RECT 682.1200 1223.4900 889.2200 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 993.8500 875.4800 1209.9500 ;
        RECT 828.8800 993.8500 830.4800 1209.9500 ;
        RECT 783.8800 993.8500 785.4800 1209.9500 ;
        RECT 738.8800 993.8500 740.4800 1209.9500 ;
        RECT 693.8800 993.8500 695.4800 1209.9500 ;
        RECT 886.2200 993.8500 889.2200 1209.9500 ;
        RECT 682.1200 993.8500 685.1200 1209.9500 ;
      LAYER met3 ;
        RECT 886.2200 1187.0000 889.2200 1187.4800 ;
        RECT 886.2200 1192.4400 889.2200 1192.9200 ;
        RECT 873.8800 1187.0000 875.4800 1187.4800 ;
        RECT 873.8800 1192.4400 875.4800 1192.9200 ;
        RECT 886.2200 1197.8800 889.2200 1198.3600 ;
        RECT 873.8800 1197.8800 875.4800 1198.3600 ;
        RECT 886.2200 1176.1200 889.2200 1176.6000 ;
        RECT 886.2200 1181.5600 889.2200 1182.0400 ;
        RECT 873.8800 1176.1200 875.4800 1176.6000 ;
        RECT 873.8800 1181.5600 875.4800 1182.0400 ;
        RECT 886.2200 1159.8000 889.2200 1160.2800 ;
        RECT 886.2200 1165.2400 889.2200 1165.7200 ;
        RECT 873.8800 1159.8000 875.4800 1160.2800 ;
        RECT 873.8800 1165.2400 875.4800 1165.7200 ;
        RECT 886.2200 1170.6800 889.2200 1171.1600 ;
        RECT 873.8800 1170.6800 875.4800 1171.1600 ;
        RECT 828.8800 1187.0000 830.4800 1187.4800 ;
        RECT 828.8800 1192.4400 830.4800 1192.9200 ;
        RECT 828.8800 1197.8800 830.4800 1198.3600 ;
        RECT 828.8800 1176.1200 830.4800 1176.6000 ;
        RECT 828.8800 1181.5600 830.4800 1182.0400 ;
        RECT 828.8800 1159.8000 830.4800 1160.2800 ;
        RECT 828.8800 1165.2400 830.4800 1165.7200 ;
        RECT 828.8800 1170.6800 830.4800 1171.1600 ;
        RECT 886.2200 1143.4800 889.2200 1143.9600 ;
        RECT 886.2200 1148.9200 889.2200 1149.4000 ;
        RECT 886.2200 1154.3600 889.2200 1154.8400 ;
        RECT 873.8800 1143.4800 875.4800 1143.9600 ;
        RECT 873.8800 1148.9200 875.4800 1149.4000 ;
        RECT 873.8800 1154.3600 875.4800 1154.8400 ;
        RECT 886.2200 1132.6000 889.2200 1133.0800 ;
        RECT 886.2200 1138.0400 889.2200 1138.5200 ;
        RECT 873.8800 1132.6000 875.4800 1133.0800 ;
        RECT 873.8800 1138.0400 875.4800 1138.5200 ;
        RECT 886.2200 1116.2800 889.2200 1116.7600 ;
        RECT 886.2200 1121.7200 889.2200 1122.2000 ;
        RECT 886.2200 1127.1600 889.2200 1127.6400 ;
        RECT 873.8800 1116.2800 875.4800 1116.7600 ;
        RECT 873.8800 1121.7200 875.4800 1122.2000 ;
        RECT 873.8800 1127.1600 875.4800 1127.6400 ;
        RECT 886.2200 1105.4000 889.2200 1105.8800 ;
        RECT 886.2200 1110.8400 889.2200 1111.3200 ;
        RECT 873.8800 1105.4000 875.4800 1105.8800 ;
        RECT 873.8800 1110.8400 875.4800 1111.3200 ;
        RECT 828.8800 1143.4800 830.4800 1143.9600 ;
        RECT 828.8800 1148.9200 830.4800 1149.4000 ;
        RECT 828.8800 1154.3600 830.4800 1154.8400 ;
        RECT 828.8800 1132.6000 830.4800 1133.0800 ;
        RECT 828.8800 1138.0400 830.4800 1138.5200 ;
        RECT 828.8800 1116.2800 830.4800 1116.7600 ;
        RECT 828.8800 1121.7200 830.4800 1122.2000 ;
        RECT 828.8800 1127.1600 830.4800 1127.6400 ;
        RECT 828.8800 1105.4000 830.4800 1105.8800 ;
        RECT 828.8800 1110.8400 830.4800 1111.3200 ;
        RECT 783.8800 1187.0000 785.4800 1187.4800 ;
        RECT 783.8800 1192.4400 785.4800 1192.9200 ;
        RECT 783.8800 1197.8800 785.4800 1198.3600 ;
        RECT 738.8800 1187.0000 740.4800 1187.4800 ;
        RECT 738.8800 1192.4400 740.4800 1192.9200 ;
        RECT 738.8800 1197.8800 740.4800 1198.3600 ;
        RECT 783.8800 1176.1200 785.4800 1176.6000 ;
        RECT 783.8800 1181.5600 785.4800 1182.0400 ;
        RECT 783.8800 1159.8000 785.4800 1160.2800 ;
        RECT 783.8800 1165.2400 785.4800 1165.7200 ;
        RECT 783.8800 1170.6800 785.4800 1171.1600 ;
        RECT 738.8800 1176.1200 740.4800 1176.6000 ;
        RECT 738.8800 1181.5600 740.4800 1182.0400 ;
        RECT 738.8800 1159.8000 740.4800 1160.2800 ;
        RECT 738.8800 1165.2400 740.4800 1165.7200 ;
        RECT 738.8800 1170.6800 740.4800 1171.1600 ;
        RECT 693.8800 1187.0000 695.4800 1187.4800 ;
        RECT 693.8800 1192.4400 695.4800 1192.9200 ;
        RECT 682.1200 1192.4400 685.1200 1192.9200 ;
        RECT 682.1200 1187.0000 685.1200 1187.4800 ;
        RECT 682.1200 1197.8800 685.1200 1198.3600 ;
        RECT 693.8800 1197.8800 695.4800 1198.3600 ;
        RECT 693.8800 1176.1200 695.4800 1176.6000 ;
        RECT 693.8800 1181.5600 695.4800 1182.0400 ;
        RECT 682.1200 1181.5600 685.1200 1182.0400 ;
        RECT 682.1200 1176.1200 685.1200 1176.6000 ;
        RECT 693.8800 1159.8000 695.4800 1160.2800 ;
        RECT 693.8800 1165.2400 695.4800 1165.7200 ;
        RECT 682.1200 1165.2400 685.1200 1165.7200 ;
        RECT 682.1200 1159.8000 685.1200 1160.2800 ;
        RECT 682.1200 1170.6800 685.1200 1171.1600 ;
        RECT 693.8800 1170.6800 695.4800 1171.1600 ;
        RECT 783.8800 1143.4800 785.4800 1143.9600 ;
        RECT 783.8800 1148.9200 785.4800 1149.4000 ;
        RECT 783.8800 1154.3600 785.4800 1154.8400 ;
        RECT 783.8800 1132.6000 785.4800 1133.0800 ;
        RECT 783.8800 1138.0400 785.4800 1138.5200 ;
        RECT 738.8800 1143.4800 740.4800 1143.9600 ;
        RECT 738.8800 1148.9200 740.4800 1149.4000 ;
        RECT 738.8800 1154.3600 740.4800 1154.8400 ;
        RECT 738.8800 1132.6000 740.4800 1133.0800 ;
        RECT 738.8800 1138.0400 740.4800 1138.5200 ;
        RECT 783.8800 1116.2800 785.4800 1116.7600 ;
        RECT 783.8800 1121.7200 785.4800 1122.2000 ;
        RECT 783.8800 1127.1600 785.4800 1127.6400 ;
        RECT 783.8800 1105.4000 785.4800 1105.8800 ;
        RECT 783.8800 1110.8400 785.4800 1111.3200 ;
        RECT 738.8800 1116.2800 740.4800 1116.7600 ;
        RECT 738.8800 1121.7200 740.4800 1122.2000 ;
        RECT 738.8800 1127.1600 740.4800 1127.6400 ;
        RECT 738.8800 1105.4000 740.4800 1105.8800 ;
        RECT 738.8800 1110.8400 740.4800 1111.3200 ;
        RECT 693.8800 1143.4800 695.4800 1143.9600 ;
        RECT 693.8800 1148.9200 695.4800 1149.4000 ;
        RECT 693.8800 1154.3600 695.4800 1154.8400 ;
        RECT 682.1200 1143.4800 685.1200 1143.9600 ;
        RECT 682.1200 1148.9200 685.1200 1149.4000 ;
        RECT 682.1200 1154.3600 685.1200 1154.8400 ;
        RECT 693.8800 1132.6000 695.4800 1133.0800 ;
        RECT 693.8800 1138.0400 695.4800 1138.5200 ;
        RECT 682.1200 1132.6000 685.1200 1133.0800 ;
        RECT 682.1200 1138.0400 685.1200 1138.5200 ;
        RECT 693.8800 1116.2800 695.4800 1116.7600 ;
        RECT 693.8800 1121.7200 695.4800 1122.2000 ;
        RECT 693.8800 1127.1600 695.4800 1127.6400 ;
        RECT 682.1200 1116.2800 685.1200 1116.7600 ;
        RECT 682.1200 1121.7200 685.1200 1122.2000 ;
        RECT 682.1200 1127.1600 685.1200 1127.6400 ;
        RECT 693.8800 1105.4000 695.4800 1105.8800 ;
        RECT 693.8800 1110.8400 695.4800 1111.3200 ;
        RECT 682.1200 1105.4000 685.1200 1105.8800 ;
        RECT 682.1200 1110.8400 685.1200 1111.3200 ;
        RECT 886.2200 1089.0800 889.2200 1089.5600 ;
        RECT 886.2200 1094.5200 889.2200 1095.0000 ;
        RECT 886.2200 1099.9600 889.2200 1100.4400 ;
        RECT 873.8800 1089.0800 875.4800 1089.5600 ;
        RECT 873.8800 1094.5200 875.4800 1095.0000 ;
        RECT 873.8800 1099.9600 875.4800 1100.4400 ;
        RECT 886.2200 1078.2000 889.2200 1078.6800 ;
        RECT 886.2200 1083.6400 889.2200 1084.1200 ;
        RECT 873.8800 1078.2000 875.4800 1078.6800 ;
        RECT 873.8800 1083.6400 875.4800 1084.1200 ;
        RECT 886.2200 1061.8800 889.2200 1062.3600 ;
        RECT 886.2200 1067.3200 889.2200 1067.8000 ;
        RECT 886.2200 1072.7600 889.2200 1073.2400 ;
        RECT 873.8800 1061.8800 875.4800 1062.3600 ;
        RECT 873.8800 1067.3200 875.4800 1067.8000 ;
        RECT 873.8800 1072.7600 875.4800 1073.2400 ;
        RECT 886.2200 1051.0000 889.2200 1051.4800 ;
        RECT 886.2200 1056.4400 889.2200 1056.9200 ;
        RECT 873.8800 1051.0000 875.4800 1051.4800 ;
        RECT 873.8800 1056.4400 875.4800 1056.9200 ;
        RECT 828.8800 1089.0800 830.4800 1089.5600 ;
        RECT 828.8800 1094.5200 830.4800 1095.0000 ;
        RECT 828.8800 1099.9600 830.4800 1100.4400 ;
        RECT 828.8800 1078.2000 830.4800 1078.6800 ;
        RECT 828.8800 1083.6400 830.4800 1084.1200 ;
        RECT 828.8800 1061.8800 830.4800 1062.3600 ;
        RECT 828.8800 1067.3200 830.4800 1067.8000 ;
        RECT 828.8800 1072.7600 830.4800 1073.2400 ;
        RECT 828.8800 1051.0000 830.4800 1051.4800 ;
        RECT 828.8800 1056.4400 830.4800 1056.9200 ;
        RECT 886.2200 1034.6800 889.2200 1035.1600 ;
        RECT 886.2200 1040.1200 889.2200 1040.6000 ;
        RECT 886.2200 1045.5600 889.2200 1046.0400 ;
        RECT 873.8800 1034.6800 875.4800 1035.1600 ;
        RECT 873.8800 1040.1200 875.4800 1040.6000 ;
        RECT 873.8800 1045.5600 875.4800 1046.0400 ;
        RECT 886.2200 1023.8000 889.2200 1024.2800 ;
        RECT 886.2200 1029.2400 889.2200 1029.7200 ;
        RECT 873.8800 1023.8000 875.4800 1024.2800 ;
        RECT 873.8800 1029.2400 875.4800 1029.7200 ;
        RECT 886.2200 1007.4800 889.2200 1007.9600 ;
        RECT 886.2200 1012.9200 889.2200 1013.4000 ;
        RECT 886.2200 1018.3600 889.2200 1018.8400 ;
        RECT 873.8800 1007.4800 875.4800 1007.9600 ;
        RECT 873.8800 1012.9200 875.4800 1013.4000 ;
        RECT 873.8800 1018.3600 875.4800 1018.8400 ;
        RECT 886.2200 1002.0400 889.2200 1002.5200 ;
        RECT 873.8800 1002.0400 875.4800 1002.5200 ;
        RECT 828.8800 1034.6800 830.4800 1035.1600 ;
        RECT 828.8800 1040.1200 830.4800 1040.6000 ;
        RECT 828.8800 1045.5600 830.4800 1046.0400 ;
        RECT 828.8800 1023.8000 830.4800 1024.2800 ;
        RECT 828.8800 1029.2400 830.4800 1029.7200 ;
        RECT 828.8800 1007.4800 830.4800 1007.9600 ;
        RECT 828.8800 1012.9200 830.4800 1013.4000 ;
        RECT 828.8800 1018.3600 830.4800 1018.8400 ;
        RECT 828.8800 1002.0400 830.4800 1002.5200 ;
        RECT 783.8800 1089.0800 785.4800 1089.5600 ;
        RECT 783.8800 1094.5200 785.4800 1095.0000 ;
        RECT 783.8800 1099.9600 785.4800 1100.4400 ;
        RECT 783.8800 1078.2000 785.4800 1078.6800 ;
        RECT 783.8800 1083.6400 785.4800 1084.1200 ;
        RECT 738.8800 1089.0800 740.4800 1089.5600 ;
        RECT 738.8800 1094.5200 740.4800 1095.0000 ;
        RECT 738.8800 1099.9600 740.4800 1100.4400 ;
        RECT 738.8800 1078.2000 740.4800 1078.6800 ;
        RECT 738.8800 1083.6400 740.4800 1084.1200 ;
        RECT 783.8800 1061.8800 785.4800 1062.3600 ;
        RECT 783.8800 1067.3200 785.4800 1067.8000 ;
        RECT 783.8800 1072.7600 785.4800 1073.2400 ;
        RECT 783.8800 1051.0000 785.4800 1051.4800 ;
        RECT 783.8800 1056.4400 785.4800 1056.9200 ;
        RECT 738.8800 1061.8800 740.4800 1062.3600 ;
        RECT 738.8800 1067.3200 740.4800 1067.8000 ;
        RECT 738.8800 1072.7600 740.4800 1073.2400 ;
        RECT 738.8800 1051.0000 740.4800 1051.4800 ;
        RECT 738.8800 1056.4400 740.4800 1056.9200 ;
        RECT 693.8800 1089.0800 695.4800 1089.5600 ;
        RECT 693.8800 1094.5200 695.4800 1095.0000 ;
        RECT 693.8800 1099.9600 695.4800 1100.4400 ;
        RECT 682.1200 1089.0800 685.1200 1089.5600 ;
        RECT 682.1200 1094.5200 685.1200 1095.0000 ;
        RECT 682.1200 1099.9600 685.1200 1100.4400 ;
        RECT 693.8800 1078.2000 695.4800 1078.6800 ;
        RECT 693.8800 1083.6400 695.4800 1084.1200 ;
        RECT 682.1200 1078.2000 685.1200 1078.6800 ;
        RECT 682.1200 1083.6400 685.1200 1084.1200 ;
        RECT 693.8800 1061.8800 695.4800 1062.3600 ;
        RECT 693.8800 1067.3200 695.4800 1067.8000 ;
        RECT 693.8800 1072.7600 695.4800 1073.2400 ;
        RECT 682.1200 1061.8800 685.1200 1062.3600 ;
        RECT 682.1200 1067.3200 685.1200 1067.8000 ;
        RECT 682.1200 1072.7600 685.1200 1073.2400 ;
        RECT 693.8800 1051.0000 695.4800 1051.4800 ;
        RECT 693.8800 1056.4400 695.4800 1056.9200 ;
        RECT 682.1200 1051.0000 685.1200 1051.4800 ;
        RECT 682.1200 1056.4400 685.1200 1056.9200 ;
        RECT 783.8800 1034.6800 785.4800 1035.1600 ;
        RECT 783.8800 1040.1200 785.4800 1040.6000 ;
        RECT 783.8800 1045.5600 785.4800 1046.0400 ;
        RECT 783.8800 1023.8000 785.4800 1024.2800 ;
        RECT 783.8800 1029.2400 785.4800 1029.7200 ;
        RECT 738.8800 1034.6800 740.4800 1035.1600 ;
        RECT 738.8800 1040.1200 740.4800 1040.6000 ;
        RECT 738.8800 1045.5600 740.4800 1046.0400 ;
        RECT 738.8800 1023.8000 740.4800 1024.2800 ;
        RECT 738.8800 1029.2400 740.4800 1029.7200 ;
        RECT 783.8800 1007.4800 785.4800 1007.9600 ;
        RECT 783.8800 1012.9200 785.4800 1013.4000 ;
        RECT 783.8800 1018.3600 785.4800 1018.8400 ;
        RECT 783.8800 1002.0400 785.4800 1002.5200 ;
        RECT 738.8800 1007.4800 740.4800 1007.9600 ;
        RECT 738.8800 1012.9200 740.4800 1013.4000 ;
        RECT 738.8800 1018.3600 740.4800 1018.8400 ;
        RECT 738.8800 1002.0400 740.4800 1002.5200 ;
        RECT 693.8800 1034.6800 695.4800 1035.1600 ;
        RECT 693.8800 1040.1200 695.4800 1040.6000 ;
        RECT 693.8800 1045.5600 695.4800 1046.0400 ;
        RECT 682.1200 1034.6800 685.1200 1035.1600 ;
        RECT 682.1200 1040.1200 685.1200 1040.6000 ;
        RECT 682.1200 1045.5600 685.1200 1046.0400 ;
        RECT 693.8800 1023.8000 695.4800 1024.2800 ;
        RECT 693.8800 1029.2400 695.4800 1029.7200 ;
        RECT 682.1200 1023.8000 685.1200 1024.2800 ;
        RECT 682.1200 1029.2400 685.1200 1029.7200 ;
        RECT 693.8800 1007.4800 695.4800 1007.9600 ;
        RECT 693.8800 1012.9200 695.4800 1013.4000 ;
        RECT 693.8800 1018.3600 695.4800 1018.8400 ;
        RECT 682.1200 1007.4800 685.1200 1007.9600 ;
        RECT 682.1200 1012.9200 685.1200 1013.4000 ;
        RECT 682.1200 1018.3600 685.1200 1018.8400 ;
        RECT 682.1200 1002.0400 685.1200 1002.5200 ;
        RECT 693.8800 1002.0400 695.4800 1002.5200 ;
        RECT 682.1200 1206.9500 889.2200 1209.9500 ;
        RECT 682.1200 993.8500 889.2200 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 873.8800 764.2100 875.4800 980.3100 ;
        RECT 828.8800 764.2100 830.4800 980.3100 ;
        RECT 783.8800 764.2100 785.4800 980.3100 ;
        RECT 738.8800 764.2100 740.4800 980.3100 ;
        RECT 693.8800 764.2100 695.4800 980.3100 ;
        RECT 886.2200 764.2100 889.2200 980.3100 ;
        RECT 682.1200 764.2100 685.1200 980.3100 ;
      LAYER met3 ;
        RECT 886.2200 957.3600 889.2200 957.8400 ;
        RECT 886.2200 962.8000 889.2200 963.2800 ;
        RECT 873.8800 957.3600 875.4800 957.8400 ;
        RECT 873.8800 962.8000 875.4800 963.2800 ;
        RECT 886.2200 968.2400 889.2200 968.7200 ;
        RECT 873.8800 968.2400 875.4800 968.7200 ;
        RECT 886.2200 946.4800 889.2200 946.9600 ;
        RECT 886.2200 951.9200 889.2200 952.4000 ;
        RECT 873.8800 946.4800 875.4800 946.9600 ;
        RECT 873.8800 951.9200 875.4800 952.4000 ;
        RECT 886.2200 930.1600 889.2200 930.6400 ;
        RECT 886.2200 935.6000 889.2200 936.0800 ;
        RECT 873.8800 930.1600 875.4800 930.6400 ;
        RECT 873.8800 935.6000 875.4800 936.0800 ;
        RECT 886.2200 941.0400 889.2200 941.5200 ;
        RECT 873.8800 941.0400 875.4800 941.5200 ;
        RECT 828.8800 957.3600 830.4800 957.8400 ;
        RECT 828.8800 962.8000 830.4800 963.2800 ;
        RECT 828.8800 968.2400 830.4800 968.7200 ;
        RECT 828.8800 946.4800 830.4800 946.9600 ;
        RECT 828.8800 951.9200 830.4800 952.4000 ;
        RECT 828.8800 930.1600 830.4800 930.6400 ;
        RECT 828.8800 935.6000 830.4800 936.0800 ;
        RECT 828.8800 941.0400 830.4800 941.5200 ;
        RECT 886.2200 913.8400 889.2200 914.3200 ;
        RECT 886.2200 919.2800 889.2200 919.7600 ;
        RECT 886.2200 924.7200 889.2200 925.2000 ;
        RECT 873.8800 913.8400 875.4800 914.3200 ;
        RECT 873.8800 919.2800 875.4800 919.7600 ;
        RECT 873.8800 924.7200 875.4800 925.2000 ;
        RECT 886.2200 902.9600 889.2200 903.4400 ;
        RECT 886.2200 908.4000 889.2200 908.8800 ;
        RECT 873.8800 902.9600 875.4800 903.4400 ;
        RECT 873.8800 908.4000 875.4800 908.8800 ;
        RECT 886.2200 886.6400 889.2200 887.1200 ;
        RECT 886.2200 892.0800 889.2200 892.5600 ;
        RECT 886.2200 897.5200 889.2200 898.0000 ;
        RECT 873.8800 886.6400 875.4800 887.1200 ;
        RECT 873.8800 892.0800 875.4800 892.5600 ;
        RECT 873.8800 897.5200 875.4800 898.0000 ;
        RECT 886.2200 875.7600 889.2200 876.2400 ;
        RECT 886.2200 881.2000 889.2200 881.6800 ;
        RECT 873.8800 875.7600 875.4800 876.2400 ;
        RECT 873.8800 881.2000 875.4800 881.6800 ;
        RECT 828.8800 913.8400 830.4800 914.3200 ;
        RECT 828.8800 919.2800 830.4800 919.7600 ;
        RECT 828.8800 924.7200 830.4800 925.2000 ;
        RECT 828.8800 902.9600 830.4800 903.4400 ;
        RECT 828.8800 908.4000 830.4800 908.8800 ;
        RECT 828.8800 886.6400 830.4800 887.1200 ;
        RECT 828.8800 892.0800 830.4800 892.5600 ;
        RECT 828.8800 897.5200 830.4800 898.0000 ;
        RECT 828.8800 875.7600 830.4800 876.2400 ;
        RECT 828.8800 881.2000 830.4800 881.6800 ;
        RECT 783.8800 957.3600 785.4800 957.8400 ;
        RECT 783.8800 962.8000 785.4800 963.2800 ;
        RECT 783.8800 968.2400 785.4800 968.7200 ;
        RECT 738.8800 957.3600 740.4800 957.8400 ;
        RECT 738.8800 962.8000 740.4800 963.2800 ;
        RECT 738.8800 968.2400 740.4800 968.7200 ;
        RECT 783.8800 946.4800 785.4800 946.9600 ;
        RECT 783.8800 951.9200 785.4800 952.4000 ;
        RECT 783.8800 930.1600 785.4800 930.6400 ;
        RECT 783.8800 935.6000 785.4800 936.0800 ;
        RECT 783.8800 941.0400 785.4800 941.5200 ;
        RECT 738.8800 946.4800 740.4800 946.9600 ;
        RECT 738.8800 951.9200 740.4800 952.4000 ;
        RECT 738.8800 930.1600 740.4800 930.6400 ;
        RECT 738.8800 935.6000 740.4800 936.0800 ;
        RECT 738.8800 941.0400 740.4800 941.5200 ;
        RECT 693.8800 957.3600 695.4800 957.8400 ;
        RECT 693.8800 962.8000 695.4800 963.2800 ;
        RECT 682.1200 962.8000 685.1200 963.2800 ;
        RECT 682.1200 957.3600 685.1200 957.8400 ;
        RECT 682.1200 968.2400 685.1200 968.7200 ;
        RECT 693.8800 968.2400 695.4800 968.7200 ;
        RECT 693.8800 946.4800 695.4800 946.9600 ;
        RECT 693.8800 951.9200 695.4800 952.4000 ;
        RECT 682.1200 951.9200 685.1200 952.4000 ;
        RECT 682.1200 946.4800 685.1200 946.9600 ;
        RECT 693.8800 930.1600 695.4800 930.6400 ;
        RECT 693.8800 935.6000 695.4800 936.0800 ;
        RECT 682.1200 935.6000 685.1200 936.0800 ;
        RECT 682.1200 930.1600 685.1200 930.6400 ;
        RECT 682.1200 941.0400 685.1200 941.5200 ;
        RECT 693.8800 941.0400 695.4800 941.5200 ;
        RECT 783.8800 913.8400 785.4800 914.3200 ;
        RECT 783.8800 919.2800 785.4800 919.7600 ;
        RECT 783.8800 924.7200 785.4800 925.2000 ;
        RECT 783.8800 902.9600 785.4800 903.4400 ;
        RECT 783.8800 908.4000 785.4800 908.8800 ;
        RECT 738.8800 913.8400 740.4800 914.3200 ;
        RECT 738.8800 919.2800 740.4800 919.7600 ;
        RECT 738.8800 924.7200 740.4800 925.2000 ;
        RECT 738.8800 902.9600 740.4800 903.4400 ;
        RECT 738.8800 908.4000 740.4800 908.8800 ;
        RECT 783.8800 886.6400 785.4800 887.1200 ;
        RECT 783.8800 892.0800 785.4800 892.5600 ;
        RECT 783.8800 897.5200 785.4800 898.0000 ;
        RECT 783.8800 875.7600 785.4800 876.2400 ;
        RECT 783.8800 881.2000 785.4800 881.6800 ;
        RECT 738.8800 886.6400 740.4800 887.1200 ;
        RECT 738.8800 892.0800 740.4800 892.5600 ;
        RECT 738.8800 897.5200 740.4800 898.0000 ;
        RECT 738.8800 875.7600 740.4800 876.2400 ;
        RECT 738.8800 881.2000 740.4800 881.6800 ;
        RECT 693.8800 913.8400 695.4800 914.3200 ;
        RECT 693.8800 919.2800 695.4800 919.7600 ;
        RECT 693.8800 924.7200 695.4800 925.2000 ;
        RECT 682.1200 913.8400 685.1200 914.3200 ;
        RECT 682.1200 919.2800 685.1200 919.7600 ;
        RECT 682.1200 924.7200 685.1200 925.2000 ;
        RECT 693.8800 902.9600 695.4800 903.4400 ;
        RECT 693.8800 908.4000 695.4800 908.8800 ;
        RECT 682.1200 902.9600 685.1200 903.4400 ;
        RECT 682.1200 908.4000 685.1200 908.8800 ;
        RECT 693.8800 886.6400 695.4800 887.1200 ;
        RECT 693.8800 892.0800 695.4800 892.5600 ;
        RECT 693.8800 897.5200 695.4800 898.0000 ;
        RECT 682.1200 886.6400 685.1200 887.1200 ;
        RECT 682.1200 892.0800 685.1200 892.5600 ;
        RECT 682.1200 897.5200 685.1200 898.0000 ;
        RECT 693.8800 875.7600 695.4800 876.2400 ;
        RECT 693.8800 881.2000 695.4800 881.6800 ;
        RECT 682.1200 875.7600 685.1200 876.2400 ;
        RECT 682.1200 881.2000 685.1200 881.6800 ;
        RECT 886.2200 859.4400 889.2200 859.9200 ;
        RECT 886.2200 864.8800 889.2200 865.3600 ;
        RECT 886.2200 870.3200 889.2200 870.8000 ;
        RECT 873.8800 859.4400 875.4800 859.9200 ;
        RECT 873.8800 864.8800 875.4800 865.3600 ;
        RECT 873.8800 870.3200 875.4800 870.8000 ;
        RECT 886.2200 848.5600 889.2200 849.0400 ;
        RECT 886.2200 854.0000 889.2200 854.4800 ;
        RECT 873.8800 848.5600 875.4800 849.0400 ;
        RECT 873.8800 854.0000 875.4800 854.4800 ;
        RECT 886.2200 832.2400 889.2200 832.7200 ;
        RECT 886.2200 837.6800 889.2200 838.1600 ;
        RECT 886.2200 843.1200 889.2200 843.6000 ;
        RECT 873.8800 832.2400 875.4800 832.7200 ;
        RECT 873.8800 837.6800 875.4800 838.1600 ;
        RECT 873.8800 843.1200 875.4800 843.6000 ;
        RECT 886.2200 821.3600 889.2200 821.8400 ;
        RECT 886.2200 826.8000 889.2200 827.2800 ;
        RECT 873.8800 821.3600 875.4800 821.8400 ;
        RECT 873.8800 826.8000 875.4800 827.2800 ;
        RECT 828.8800 859.4400 830.4800 859.9200 ;
        RECT 828.8800 864.8800 830.4800 865.3600 ;
        RECT 828.8800 870.3200 830.4800 870.8000 ;
        RECT 828.8800 848.5600 830.4800 849.0400 ;
        RECT 828.8800 854.0000 830.4800 854.4800 ;
        RECT 828.8800 832.2400 830.4800 832.7200 ;
        RECT 828.8800 837.6800 830.4800 838.1600 ;
        RECT 828.8800 843.1200 830.4800 843.6000 ;
        RECT 828.8800 821.3600 830.4800 821.8400 ;
        RECT 828.8800 826.8000 830.4800 827.2800 ;
        RECT 886.2200 805.0400 889.2200 805.5200 ;
        RECT 886.2200 810.4800 889.2200 810.9600 ;
        RECT 886.2200 815.9200 889.2200 816.4000 ;
        RECT 873.8800 805.0400 875.4800 805.5200 ;
        RECT 873.8800 810.4800 875.4800 810.9600 ;
        RECT 873.8800 815.9200 875.4800 816.4000 ;
        RECT 886.2200 794.1600 889.2200 794.6400 ;
        RECT 886.2200 799.6000 889.2200 800.0800 ;
        RECT 873.8800 794.1600 875.4800 794.6400 ;
        RECT 873.8800 799.6000 875.4800 800.0800 ;
        RECT 886.2200 777.8400 889.2200 778.3200 ;
        RECT 886.2200 783.2800 889.2200 783.7600 ;
        RECT 886.2200 788.7200 889.2200 789.2000 ;
        RECT 873.8800 777.8400 875.4800 778.3200 ;
        RECT 873.8800 783.2800 875.4800 783.7600 ;
        RECT 873.8800 788.7200 875.4800 789.2000 ;
        RECT 886.2200 772.4000 889.2200 772.8800 ;
        RECT 873.8800 772.4000 875.4800 772.8800 ;
        RECT 828.8800 805.0400 830.4800 805.5200 ;
        RECT 828.8800 810.4800 830.4800 810.9600 ;
        RECT 828.8800 815.9200 830.4800 816.4000 ;
        RECT 828.8800 794.1600 830.4800 794.6400 ;
        RECT 828.8800 799.6000 830.4800 800.0800 ;
        RECT 828.8800 777.8400 830.4800 778.3200 ;
        RECT 828.8800 783.2800 830.4800 783.7600 ;
        RECT 828.8800 788.7200 830.4800 789.2000 ;
        RECT 828.8800 772.4000 830.4800 772.8800 ;
        RECT 783.8800 859.4400 785.4800 859.9200 ;
        RECT 783.8800 864.8800 785.4800 865.3600 ;
        RECT 783.8800 870.3200 785.4800 870.8000 ;
        RECT 783.8800 848.5600 785.4800 849.0400 ;
        RECT 783.8800 854.0000 785.4800 854.4800 ;
        RECT 738.8800 859.4400 740.4800 859.9200 ;
        RECT 738.8800 864.8800 740.4800 865.3600 ;
        RECT 738.8800 870.3200 740.4800 870.8000 ;
        RECT 738.8800 848.5600 740.4800 849.0400 ;
        RECT 738.8800 854.0000 740.4800 854.4800 ;
        RECT 783.8800 832.2400 785.4800 832.7200 ;
        RECT 783.8800 837.6800 785.4800 838.1600 ;
        RECT 783.8800 843.1200 785.4800 843.6000 ;
        RECT 783.8800 821.3600 785.4800 821.8400 ;
        RECT 783.8800 826.8000 785.4800 827.2800 ;
        RECT 738.8800 832.2400 740.4800 832.7200 ;
        RECT 738.8800 837.6800 740.4800 838.1600 ;
        RECT 738.8800 843.1200 740.4800 843.6000 ;
        RECT 738.8800 821.3600 740.4800 821.8400 ;
        RECT 738.8800 826.8000 740.4800 827.2800 ;
        RECT 693.8800 859.4400 695.4800 859.9200 ;
        RECT 693.8800 864.8800 695.4800 865.3600 ;
        RECT 693.8800 870.3200 695.4800 870.8000 ;
        RECT 682.1200 859.4400 685.1200 859.9200 ;
        RECT 682.1200 864.8800 685.1200 865.3600 ;
        RECT 682.1200 870.3200 685.1200 870.8000 ;
        RECT 693.8800 848.5600 695.4800 849.0400 ;
        RECT 693.8800 854.0000 695.4800 854.4800 ;
        RECT 682.1200 848.5600 685.1200 849.0400 ;
        RECT 682.1200 854.0000 685.1200 854.4800 ;
        RECT 693.8800 832.2400 695.4800 832.7200 ;
        RECT 693.8800 837.6800 695.4800 838.1600 ;
        RECT 693.8800 843.1200 695.4800 843.6000 ;
        RECT 682.1200 832.2400 685.1200 832.7200 ;
        RECT 682.1200 837.6800 685.1200 838.1600 ;
        RECT 682.1200 843.1200 685.1200 843.6000 ;
        RECT 693.8800 821.3600 695.4800 821.8400 ;
        RECT 693.8800 826.8000 695.4800 827.2800 ;
        RECT 682.1200 821.3600 685.1200 821.8400 ;
        RECT 682.1200 826.8000 685.1200 827.2800 ;
        RECT 783.8800 805.0400 785.4800 805.5200 ;
        RECT 783.8800 810.4800 785.4800 810.9600 ;
        RECT 783.8800 815.9200 785.4800 816.4000 ;
        RECT 783.8800 794.1600 785.4800 794.6400 ;
        RECT 783.8800 799.6000 785.4800 800.0800 ;
        RECT 738.8800 805.0400 740.4800 805.5200 ;
        RECT 738.8800 810.4800 740.4800 810.9600 ;
        RECT 738.8800 815.9200 740.4800 816.4000 ;
        RECT 738.8800 794.1600 740.4800 794.6400 ;
        RECT 738.8800 799.6000 740.4800 800.0800 ;
        RECT 783.8800 777.8400 785.4800 778.3200 ;
        RECT 783.8800 783.2800 785.4800 783.7600 ;
        RECT 783.8800 788.7200 785.4800 789.2000 ;
        RECT 783.8800 772.4000 785.4800 772.8800 ;
        RECT 738.8800 777.8400 740.4800 778.3200 ;
        RECT 738.8800 783.2800 740.4800 783.7600 ;
        RECT 738.8800 788.7200 740.4800 789.2000 ;
        RECT 738.8800 772.4000 740.4800 772.8800 ;
        RECT 693.8800 805.0400 695.4800 805.5200 ;
        RECT 693.8800 810.4800 695.4800 810.9600 ;
        RECT 693.8800 815.9200 695.4800 816.4000 ;
        RECT 682.1200 805.0400 685.1200 805.5200 ;
        RECT 682.1200 810.4800 685.1200 810.9600 ;
        RECT 682.1200 815.9200 685.1200 816.4000 ;
        RECT 693.8800 794.1600 695.4800 794.6400 ;
        RECT 693.8800 799.6000 695.4800 800.0800 ;
        RECT 682.1200 794.1600 685.1200 794.6400 ;
        RECT 682.1200 799.6000 685.1200 800.0800 ;
        RECT 693.8800 777.8400 695.4800 778.3200 ;
        RECT 693.8800 783.2800 695.4800 783.7600 ;
        RECT 693.8800 788.7200 695.4800 789.2000 ;
        RECT 682.1200 777.8400 685.1200 778.3200 ;
        RECT 682.1200 783.2800 685.1200 783.7600 ;
        RECT 682.1200 788.7200 685.1200 789.2000 ;
        RECT 682.1200 772.4000 685.1200 772.8800 ;
        RECT 693.8800 772.4000 695.4800 772.8800 ;
        RECT 682.1200 977.3100 889.2200 980.3100 ;
        RECT 682.1200 764.2100 889.2200 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single2'
    PORT
      LAYER met4 ;
        RECT 1136.3400 2830.6100 1138.3400 2857.5400 ;
        RECT 903.3400 2830.6100 905.3400 2857.5400 ;
      LAYER met3 ;
        RECT 1136.3400 2847.3200 1138.3400 2847.8000 ;
        RECT 903.3400 2847.3200 905.3400 2847.8000 ;
        RECT 1136.3400 2836.4400 1138.3400 2836.9200 ;
        RECT 1136.3400 2841.8800 1138.3400 2842.3600 ;
        RECT 903.3400 2836.4400 905.3400 2836.9200 ;
        RECT 903.3400 2841.8800 905.3400 2842.3600 ;
        RECT 903.3400 2855.5400 1138.3400 2857.5400 ;
        RECT 903.3400 2830.6100 1138.3400 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single2'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 534.5700 1094.1000 750.6700 ;
        RECT 1048.1000 534.5700 1049.1000 750.6700 ;
        RECT 1003.1000 534.5700 1004.1000 750.6700 ;
        RECT 958.1000 534.5700 959.1000 750.6700 ;
        RECT 913.1000 534.5700 914.1000 750.6700 ;
        RECT 1136.3400 534.5700 1139.3400 750.6700 ;
        RECT 902.3400 534.5700 905.3400 750.6700 ;
      LAYER met3 ;
        RECT 1136.3400 733.1600 1139.3400 733.6400 ;
        RECT 1136.3400 738.6000 1139.3400 739.0800 ;
        RECT 1093.1000 733.1600 1094.1000 733.6400 ;
        RECT 1093.1000 738.6000 1094.1000 739.0800 ;
        RECT 1136.3400 722.2800 1139.3400 722.7600 ;
        RECT 1136.3400 727.7200 1139.3400 728.2000 ;
        RECT 1136.3400 711.4000 1139.3400 711.8800 ;
        RECT 1136.3400 716.8400 1139.3400 717.3200 ;
        RECT 1136.3400 705.9600 1139.3400 706.4400 ;
        RECT 1093.1000 722.2800 1094.1000 722.7600 ;
        RECT 1093.1000 727.7200 1094.1000 728.2000 ;
        RECT 1093.1000 705.9600 1094.1000 706.4400 ;
        RECT 1093.1000 711.4000 1094.1000 711.8800 ;
        RECT 1093.1000 716.8400 1094.1000 717.3200 ;
        RECT 1048.1000 733.1600 1049.1000 733.6400 ;
        RECT 1048.1000 738.6000 1049.1000 739.0800 ;
        RECT 1048.1000 722.2800 1049.1000 722.7600 ;
        RECT 1048.1000 727.7200 1049.1000 728.2000 ;
        RECT 1048.1000 705.9600 1049.1000 706.4400 ;
        RECT 1048.1000 711.4000 1049.1000 711.8800 ;
        RECT 1048.1000 716.8400 1049.1000 717.3200 ;
        RECT 1136.3400 689.6400 1139.3400 690.1200 ;
        RECT 1136.3400 695.0800 1139.3400 695.5600 ;
        RECT 1136.3400 700.5200 1139.3400 701.0000 ;
        RECT 1136.3400 684.2000 1139.3400 684.6800 ;
        RECT 1136.3400 673.3200 1139.3400 673.8000 ;
        RECT 1136.3400 678.7600 1139.3400 679.2400 ;
        RECT 1093.1000 689.6400 1094.1000 690.1200 ;
        RECT 1093.1000 695.0800 1094.1000 695.5600 ;
        RECT 1093.1000 700.5200 1094.1000 701.0000 ;
        RECT 1093.1000 673.3200 1094.1000 673.8000 ;
        RECT 1093.1000 678.7600 1094.1000 679.2400 ;
        RECT 1093.1000 684.2000 1094.1000 684.6800 ;
        RECT 1136.3400 662.4400 1139.3400 662.9200 ;
        RECT 1136.3400 667.8800 1139.3400 668.3600 ;
        RECT 1136.3400 651.5600 1139.3400 652.0400 ;
        RECT 1136.3400 657.0000 1139.3400 657.4800 ;
        RECT 1136.3400 646.1200 1139.3400 646.6000 ;
        RECT 1093.1000 662.4400 1094.1000 662.9200 ;
        RECT 1093.1000 667.8800 1094.1000 668.3600 ;
        RECT 1093.1000 646.1200 1094.1000 646.6000 ;
        RECT 1093.1000 651.5600 1094.1000 652.0400 ;
        RECT 1093.1000 657.0000 1094.1000 657.4800 ;
        RECT 1048.1000 689.6400 1049.1000 690.1200 ;
        RECT 1048.1000 695.0800 1049.1000 695.5600 ;
        RECT 1048.1000 700.5200 1049.1000 701.0000 ;
        RECT 1048.1000 673.3200 1049.1000 673.8000 ;
        RECT 1048.1000 678.7600 1049.1000 679.2400 ;
        RECT 1048.1000 684.2000 1049.1000 684.6800 ;
        RECT 1048.1000 662.4400 1049.1000 662.9200 ;
        RECT 1048.1000 667.8800 1049.1000 668.3600 ;
        RECT 1048.1000 646.1200 1049.1000 646.6000 ;
        RECT 1048.1000 651.5600 1049.1000 652.0400 ;
        RECT 1048.1000 657.0000 1049.1000 657.4800 ;
        RECT 1003.1000 733.1600 1004.1000 733.6400 ;
        RECT 1003.1000 738.6000 1004.1000 739.0800 ;
        RECT 1003.1000 722.2800 1004.1000 722.7600 ;
        RECT 1003.1000 727.7200 1004.1000 728.2000 ;
        RECT 1003.1000 705.9600 1004.1000 706.4400 ;
        RECT 1003.1000 711.4000 1004.1000 711.8800 ;
        RECT 1003.1000 716.8400 1004.1000 717.3200 ;
        RECT 958.1000 733.1600 959.1000 733.6400 ;
        RECT 958.1000 738.6000 959.1000 739.0800 ;
        RECT 913.1000 738.6000 914.1000 739.0800 ;
        RECT 913.1000 733.1600 914.1000 733.6400 ;
        RECT 902.3400 738.6000 905.3400 739.0800 ;
        RECT 902.3400 733.1600 905.3400 733.6400 ;
        RECT 958.1000 722.2800 959.1000 722.7600 ;
        RECT 958.1000 727.7200 959.1000 728.2000 ;
        RECT 958.1000 705.9600 959.1000 706.4400 ;
        RECT 958.1000 711.4000 959.1000 711.8800 ;
        RECT 958.1000 716.8400 959.1000 717.3200 ;
        RECT 902.3400 727.7200 905.3400 728.2000 ;
        RECT 913.1000 727.7200 914.1000 728.2000 ;
        RECT 902.3400 722.2800 905.3400 722.7600 ;
        RECT 913.1000 722.2800 914.1000 722.7600 ;
        RECT 913.1000 716.8400 914.1000 717.3200 ;
        RECT 913.1000 711.4000 914.1000 711.8800 ;
        RECT 902.3400 716.8400 905.3400 717.3200 ;
        RECT 902.3400 711.4000 905.3400 711.8800 ;
        RECT 902.3400 705.9600 905.3400 706.4400 ;
        RECT 913.1000 705.9600 914.1000 706.4400 ;
        RECT 1003.1000 689.6400 1004.1000 690.1200 ;
        RECT 1003.1000 695.0800 1004.1000 695.5600 ;
        RECT 1003.1000 700.5200 1004.1000 701.0000 ;
        RECT 1003.1000 673.3200 1004.1000 673.8000 ;
        RECT 1003.1000 678.7600 1004.1000 679.2400 ;
        RECT 1003.1000 684.2000 1004.1000 684.6800 ;
        RECT 1003.1000 662.4400 1004.1000 662.9200 ;
        RECT 1003.1000 667.8800 1004.1000 668.3600 ;
        RECT 1003.1000 646.1200 1004.1000 646.6000 ;
        RECT 1003.1000 651.5600 1004.1000 652.0400 ;
        RECT 1003.1000 657.0000 1004.1000 657.4800 ;
        RECT 958.1000 689.6400 959.1000 690.1200 ;
        RECT 958.1000 695.0800 959.1000 695.5600 ;
        RECT 958.1000 700.5200 959.1000 701.0000 ;
        RECT 958.1000 673.3200 959.1000 673.8000 ;
        RECT 958.1000 678.7600 959.1000 679.2400 ;
        RECT 958.1000 684.2000 959.1000 684.6800 ;
        RECT 902.3400 700.5200 905.3400 701.0000 ;
        RECT 913.1000 700.5200 914.1000 701.0000 ;
        RECT 902.3400 689.6400 905.3400 690.1200 ;
        RECT 913.1000 689.6400 914.1000 690.1200 ;
        RECT 902.3400 695.0800 905.3400 695.5600 ;
        RECT 913.1000 695.0800 914.1000 695.5600 ;
        RECT 902.3400 684.2000 905.3400 684.6800 ;
        RECT 913.1000 684.2000 914.1000 684.6800 ;
        RECT 913.1000 678.7600 914.1000 679.2400 ;
        RECT 913.1000 673.3200 914.1000 673.8000 ;
        RECT 902.3400 678.7600 905.3400 679.2400 ;
        RECT 902.3400 673.3200 905.3400 673.8000 ;
        RECT 958.1000 662.4400 959.1000 662.9200 ;
        RECT 958.1000 667.8800 959.1000 668.3600 ;
        RECT 958.1000 646.1200 959.1000 646.6000 ;
        RECT 958.1000 651.5600 959.1000 652.0400 ;
        RECT 958.1000 657.0000 959.1000 657.4800 ;
        RECT 902.3400 667.8800 905.3400 668.3600 ;
        RECT 913.1000 667.8800 914.1000 668.3600 ;
        RECT 902.3400 662.4400 905.3400 662.9200 ;
        RECT 913.1000 662.4400 914.1000 662.9200 ;
        RECT 913.1000 657.0000 914.1000 657.4800 ;
        RECT 913.1000 651.5600 914.1000 652.0400 ;
        RECT 902.3400 657.0000 905.3400 657.4800 ;
        RECT 902.3400 651.5600 905.3400 652.0400 ;
        RECT 902.3400 646.1200 905.3400 646.6000 ;
        RECT 913.1000 646.1200 914.1000 646.6000 ;
        RECT 1136.3400 629.8000 1139.3400 630.2800 ;
        RECT 1136.3400 635.2400 1139.3400 635.7200 ;
        RECT 1136.3400 640.6800 1139.3400 641.1600 ;
        RECT 1136.3400 624.3600 1139.3400 624.8400 ;
        RECT 1136.3400 613.4800 1139.3400 613.9600 ;
        RECT 1136.3400 618.9200 1139.3400 619.4000 ;
        RECT 1093.1000 629.8000 1094.1000 630.2800 ;
        RECT 1093.1000 635.2400 1094.1000 635.7200 ;
        RECT 1093.1000 640.6800 1094.1000 641.1600 ;
        RECT 1093.1000 613.4800 1094.1000 613.9600 ;
        RECT 1093.1000 618.9200 1094.1000 619.4000 ;
        RECT 1093.1000 624.3600 1094.1000 624.8400 ;
        RECT 1136.3400 602.6000 1139.3400 603.0800 ;
        RECT 1136.3400 608.0400 1139.3400 608.5200 ;
        RECT 1136.3400 591.7200 1139.3400 592.2000 ;
        RECT 1136.3400 597.1600 1139.3400 597.6400 ;
        RECT 1136.3400 586.2800 1139.3400 586.7600 ;
        RECT 1093.1000 602.6000 1094.1000 603.0800 ;
        RECT 1093.1000 608.0400 1094.1000 608.5200 ;
        RECT 1093.1000 586.2800 1094.1000 586.7600 ;
        RECT 1093.1000 591.7200 1094.1000 592.2000 ;
        RECT 1093.1000 597.1600 1094.1000 597.6400 ;
        RECT 1048.1000 629.8000 1049.1000 630.2800 ;
        RECT 1048.1000 635.2400 1049.1000 635.7200 ;
        RECT 1048.1000 640.6800 1049.1000 641.1600 ;
        RECT 1048.1000 613.4800 1049.1000 613.9600 ;
        RECT 1048.1000 618.9200 1049.1000 619.4000 ;
        RECT 1048.1000 624.3600 1049.1000 624.8400 ;
        RECT 1048.1000 602.6000 1049.1000 603.0800 ;
        RECT 1048.1000 608.0400 1049.1000 608.5200 ;
        RECT 1048.1000 586.2800 1049.1000 586.7600 ;
        RECT 1048.1000 591.7200 1049.1000 592.2000 ;
        RECT 1048.1000 597.1600 1049.1000 597.6400 ;
        RECT 1136.3400 569.9600 1139.3400 570.4400 ;
        RECT 1136.3400 575.4000 1139.3400 575.8800 ;
        RECT 1136.3400 580.8400 1139.3400 581.3200 ;
        RECT 1136.3400 564.5200 1139.3400 565.0000 ;
        RECT 1136.3400 553.6400 1139.3400 554.1200 ;
        RECT 1136.3400 559.0800 1139.3400 559.5600 ;
        RECT 1093.1000 569.9600 1094.1000 570.4400 ;
        RECT 1093.1000 575.4000 1094.1000 575.8800 ;
        RECT 1093.1000 580.8400 1094.1000 581.3200 ;
        RECT 1093.1000 553.6400 1094.1000 554.1200 ;
        RECT 1093.1000 559.0800 1094.1000 559.5600 ;
        RECT 1093.1000 564.5200 1094.1000 565.0000 ;
        RECT 1136.3400 542.7600 1139.3400 543.2400 ;
        RECT 1136.3400 548.2000 1139.3400 548.6800 ;
        RECT 1093.1000 542.7600 1094.1000 543.2400 ;
        RECT 1093.1000 548.2000 1094.1000 548.6800 ;
        RECT 1048.1000 569.9600 1049.1000 570.4400 ;
        RECT 1048.1000 575.4000 1049.1000 575.8800 ;
        RECT 1048.1000 580.8400 1049.1000 581.3200 ;
        RECT 1048.1000 553.6400 1049.1000 554.1200 ;
        RECT 1048.1000 559.0800 1049.1000 559.5600 ;
        RECT 1048.1000 564.5200 1049.1000 565.0000 ;
        RECT 1048.1000 542.7600 1049.1000 543.2400 ;
        RECT 1048.1000 548.2000 1049.1000 548.6800 ;
        RECT 1003.1000 629.8000 1004.1000 630.2800 ;
        RECT 1003.1000 635.2400 1004.1000 635.7200 ;
        RECT 1003.1000 640.6800 1004.1000 641.1600 ;
        RECT 1003.1000 613.4800 1004.1000 613.9600 ;
        RECT 1003.1000 618.9200 1004.1000 619.4000 ;
        RECT 1003.1000 624.3600 1004.1000 624.8400 ;
        RECT 1003.1000 602.6000 1004.1000 603.0800 ;
        RECT 1003.1000 608.0400 1004.1000 608.5200 ;
        RECT 1003.1000 586.2800 1004.1000 586.7600 ;
        RECT 1003.1000 591.7200 1004.1000 592.2000 ;
        RECT 1003.1000 597.1600 1004.1000 597.6400 ;
        RECT 958.1000 629.8000 959.1000 630.2800 ;
        RECT 958.1000 635.2400 959.1000 635.7200 ;
        RECT 958.1000 640.6800 959.1000 641.1600 ;
        RECT 958.1000 613.4800 959.1000 613.9600 ;
        RECT 958.1000 618.9200 959.1000 619.4000 ;
        RECT 958.1000 624.3600 959.1000 624.8400 ;
        RECT 902.3400 640.6800 905.3400 641.1600 ;
        RECT 913.1000 640.6800 914.1000 641.1600 ;
        RECT 902.3400 629.8000 905.3400 630.2800 ;
        RECT 913.1000 629.8000 914.1000 630.2800 ;
        RECT 902.3400 635.2400 905.3400 635.7200 ;
        RECT 913.1000 635.2400 914.1000 635.7200 ;
        RECT 902.3400 624.3600 905.3400 624.8400 ;
        RECT 913.1000 624.3600 914.1000 624.8400 ;
        RECT 913.1000 618.9200 914.1000 619.4000 ;
        RECT 913.1000 613.4800 914.1000 613.9600 ;
        RECT 902.3400 618.9200 905.3400 619.4000 ;
        RECT 902.3400 613.4800 905.3400 613.9600 ;
        RECT 958.1000 602.6000 959.1000 603.0800 ;
        RECT 958.1000 608.0400 959.1000 608.5200 ;
        RECT 958.1000 586.2800 959.1000 586.7600 ;
        RECT 958.1000 591.7200 959.1000 592.2000 ;
        RECT 958.1000 597.1600 959.1000 597.6400 ;
        RECT 902.3400 608.0400 905.3400 608.5200 ;
        RECT 913.1000 608.0400 914.1000 608.5200 ;
        RECT 902.3400 602.6000 905.3400 603.0800 ;
        RECT 913.1000 602.6000 914.1000 603.0800 ;
        RECT 913.1000 597.1600 914.1000 597.6400 ;
        RECT 913.1000 591.7200 914.1000 592.2000 ;
        RECT 902.3400 597.1600 905.3400 597.6400 ;
        RECT 902.3400 591.7200 905.3400 592.2000 ;
        RECT 902.3400 586.2800 905.3400 586.7600 ;
        RECT 913.1000 586.2800 914.1000 586.7600 ;
        RECT 1003.1000 569.9600 1004.1000 570.4400 ;
        RECT 1003.1000 575.4000 1004.1000 575.8800 ;
        RECT 1003.1000 580.8400 1004.1000 581.3200 ;
        RECT 1003.1000 553.6400 1004.1000 554.1200 ;
        RECT 1003.1000 559.0800 1004.1000 559.5600 ;
        RECT 1003.1000 564.5200 1004.1000 565.0000 ;
        RECT 1003.1000 542.7600 1004.1000 543.2400 ;
        RECT 1003.1000 548.2000 1004.1000 548.6800 ;
        RECT 958.1000 569.9600 959.1000 570.4400 ;
        RECT 958.1000 575.4000 959.1000 575.8800 ;
        RECT 958.1000 580.8400 959.1000 581.3200 ;
        RECT 958.1000 553.6400 959.1000 554.1200 ;
        RECT 958.1000 559.0800 959.1000 559.5600 ;
        RECT 958.1000 564.5200 959.1000 565.0000 ;
        RECT 902.3400 580.8400 905.3400 581.3200 ;
        RECT 913.1000 580.8400 914.1000 581.3200 ;
        RECT 902.3400 569.9600 905.3400 570.4400 ;
        RECT 913.1000 569.9600 914.1000 570.4400 ;
        RECT 902.3400 575.4000 905.3400 575.8800 ;
        RECT 913.1000 575.4000 914.1000 575.8800 ;
        RECT 902.3400 564.5200 905.3400 565.0000 ;
        RECT 913.1000 564.5200 914.1000 565.0000 ;
        RECT 913.1000 559.0800 914.1000 559.5600 ;
        RECT 913.1000 553.6400 914.1000 554.1200 ;
        RECT 902.3400 559.0800 905.3400 559.5600 ;
        RECT 902.3400 553.6400 905.3400 554.1200 ;
        RECT 958.1000 542.7600 959.1000 543.2400 ;
        RECT 958.1000 548.2000 959.1000 548.6800 ;
        RECT 902.3400 548.2000 905.3400 548.6800 ;
        RECT 913.1000 548.2000 914.1000 548.6800 ;
        RECT 902.3400 542.7600 905.3400 543.2400 ;
        RECT 913.1000 542.7600 914.1000 543.2400 ;
        RECT 902.3400 747.6700 1139.3400 750.6700 ;
        RECT 902.3400 534.5700 1139.3400 537.5700 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 304.9300 1094.1000 521.0300 ;
        RECT 1048.1000 304.9300 1049.1000 521.0300 ;
        RECT 1003.1000 304.9300 1004.1000 521.0300 ;
        RECT 958.1000 304.9300 959.1000 521.0300 ;
        RECT 913.1000 304.9300 914.1000 521.0300 ;
        RECT 1136.3400 304.9300 1139.3400 521.0300 ;
        RECT 902.3400 304.9300 905.3400 521.0300 ;
      LAYER met3 ;
        RECT 1136.3400 503.5200 1139.3400 504.0000 ;
        RECT 1136.3400 508.9600 1139.3400 509.4400 ;
        RECT 1093.1000 503.5200 1094.1000 504.0000 ;
        RECT 1093.1000 508.9600 1094.1000 509.4400 ;
        RECT 1136.3400 492.6400 1139.3400 493.1200 ;
        RECT 1136.3400 498.0800 1139.3400 498.5600 ;
        RECT 1136.3400 481.7600 1139.3400 482.2400 ;
        RECT 1136.3400 487.2000 1139.3400 487.6800 ;
        RECT 1136.3400 476.3200 1139.3400 476.8000 ;
        RECT 1093.1000 492.6400 1094.1000 493.1200 ;
        RECT 1093.1000 498.0800 1094.1000 498.5600 ;
        RECT 1093.1000 476.3200 1094.1000 476.8000 ;
        RECT 1093.1000 481.7600 1094.1000 482.2400 ;
        RECT 1093.1000 487.2000 1094.1000 487.6800 ;
        RECT 1048.1000 503.5200 1049.1000 504.0000 ;
        RECT 1048.1000 508.9600 1049.1000 509.4400 ;
        RECT 1048.1000 492.6400 1049.1000 493.1200 ;
        RECT 1048.1000 498.0800 1049.1000 498.5600 ;
        RECT 1048.1000 476.3200 1049.1000 476.8000 ;
        RECT 1048.1000 481.7600 1049.1000 482.2400 ;
        RECT 1048.1000 487.2000 1049.1000 487.6800 ;
        RECT 1136.3400 460.0000 1139.3400 460.4800 ;
        RECT 1136.3400 465.4400 1139.3400 465.9200 ;
        RECT 1136.3400 470.8800 1139.3400 471.3600 ;
        RECT 1136.3400 454.5600 1139.3400 455.0400 ;
        RECT 1136.3400 443.6800 1139.3400 444.1600 ;
        RECT 1136.3400 449.1200 1139.3400 449.6000 ;
        RECT 1093.1000 460.0000 1094.1000 460.4800 ;
        RECT 1093.1000 465.4400 1094.1000 465.9200 ;
        RECT 1093.1000 470.8800 1094.1000 471.3600 ;
        RECT 1093.1000 443.6800 1094.1000 444.1600 ;
        RECT 1093.1000 449.1200 1094.1000 449.6000 ;
        RECT 1093.1000 454.5600 1094.1000 455.0400 ;
        RECT 1136.3400 432.8000 1139.3400 433.2800 ;
        RECT 1136.3400 438.2400 1139.3400 438.7200 ;
        RECT 1136.3400 421.9200 1139.3400 422.4000 ;
        RECT 1136.3400 427.3600 1139.3400 427.8400 ;
        RECT 1136.3400 416.4800 1139.3400 416.9600 ;
        RECT 1093.1000 432.8000 1094.1000 433.2800 ;
        RECT 1093.1000 438.2400 1094.1000 438.7200 ;
        RECT 1093.1000 416.4800 1094.1000 416.9600 ;
        RECT 1093.1000 421.9200 1094.1000 422.4000 ;
        RECT 1093.1000 427.3600 1094.1000 427.8400 ;
        RECT 1048.1000 460.0000 1049.1000 460.4800 ;
        RECT 1048.1000 465.4400 1049.1000 465.9200 ;
        RECT 1048.1000 470.8800 1049.1000 471.3600 ;
        RECT 1048.1000 443.6800 1049.1000 444.1600 ;
        RECT 1048.1000 449.1200 1049.1000 449.6000 ;
        RECT 1048.1000 454.5600 1049.1000 455.0400 ;
        RECT 1048.1000 432.8000 1049.1000 433.2800 ;
        RECT 1048.1000 438.2400 1049.1000 438.7200 ;
        RECT 1048.1000 416.4800 1049.1000 416.9600 ;
        RECT 1048.1000 421.9200 1049.1000 422.4000 ;
        RECT 1048.1000 427.3600 1049.1000 427.8400 ;
        RECT 1003.1000 503.5200 1004.1000 504.0000 ;
        RECT 1003.1000 508.9600 1004.1000 509.4400 ;
        RECT 1003.1000 492.6400 1004.1000 493.1200 ;
        RECT 1003.1000 498.0800 1004.1000 498.5600 ;
        RECT 1003.1000 476.3200 1004.1000 476.8000 ;
        RECT 1003.1000 481.7600 1004.1000 482.2400 ;
        RECT 1003.1000 487.2000 1004.1000 487.6800 ;
        RECT 958.1000 503.5200 959.1000 504.0000 ;
        RECT 958.1000 508.9600 959.1000 509.4400 ;
        RECT 913.1000 508.9600 914.1000 509.4400 ;
        RECT 913.1000 503.5200 914.1000 504.0000 ;
        RECT 902.3400 508.9600 905.3400 509.4400 ;
        RECT 902.3400 503.5200 905.3400 504.0000 ;
        RECT 958.1000 492.6400 959.1000 493.1200 ;
        RECT 958.1000 498.0800 959.1000 498.5600 ;
        RECT 958.1000 476.3200 959.1000 476.8000 ;
        RECT 958.1000 481.7600 959.1000 482.2400 ;
        RECT 958.1000 487.2000 959.1000 487.6800 ;
        RECT 902.3400 498.0800 905.3400 498.5600 ;
        RECT 913.1000 498.0800 914.1000 498.5600 ;
        RECT 902.3400 492.6400 905.3400 493.1200 ;
        RECT 913.1000 492.6400 914.1000 493.1200 ;
        RECT 913.1000 487.2000 914.1000 487.6800 ;
        RECT 913.1000 481.7600 914.1000 482.2400 ;
        RECT 902.3400 487.2000 905.3400 487.6800 ;
        RECT 902.3400 481.7600 905.3400 482.2400 ;
        RECT 902.3400 476.3200 905.3400 476.8000 ;
        RECT 913.1000 476.3200 914.1000 476.8000 ;
        RECT 1003.1000 460.0000 1004.1000 460.4800 ;
        RECT 1003.1000 465.4400 1004.1000 465.9200 ;
        RECT 1003.1000 470.8800 1004.1000 471.3600 ;
        RECT 1003.1000 443.6800 1004.1000 444.1600 ;
        RECT 1003.1000 449.1200 1004.1000 449.6000 ;
        RECT 1003.1000 454.5600 1004.1000 455.0400 ;
        RECT 1003.1000 432.8000 1004.1000 433.2800 ;
        RECT 1003.1000 438.2400 1004.1000 438.7200 ;
        RECT 1003.1000 416.4800 1004.1000 416.9600 ;
        RECT 1003.1000 421.9200 1004.1000 422.4000 ;
        RECT 1003.1000 427.3600 1004.1000 427.8400 ;
        RECT 958.1000 460.0000 959.1000 460.4800 ;
        RECT 958.1000 465.4400 959.1000 465.9200 ;
        RECT 958.1000 470.8800 959.1000 471.3600 ;
        RECT 958.1000 443.6800 959.1000 444.1600 ;
        RECT 958.1000 449.1200 959.1000 449.6000 ;
        RECT 958.1000 454.5600 959.1000 455.0400 ;
        RECT 902.3400 470.8800 905.3400 471.3600 ;
        RECT 913.1000 470.8800 914.1000 471.3600 ;
        RECT 902.3400 460.0000 905.3400 460.4800 ;
        RECT 913.1000 460.0000 914.1000 460.4800 ;
        RECT 902.3400 465.4400 905.3400 465.9200 ;
        RECT 913.1000 465.4400 914.1000 465.9200 ;
        RECT 902.3400 454.5600 905.3400 455.0400 ;
        RECT 913.1000 454.5600 914.1000 455.0400 ;
        RECT 913.1000 449.1200 914.1000 449.6000 ;
        RECT 913.1000 443.6800 914.1000 444.1600 ;
        RECT 902.3400 449.1200 905.3400 449.6000 ;
        RECT 902.3400 443.6800 905.3400 444.1600 ;
        RECT 958.1000 432.8000 959.1000 433.2800 ;
        RECT 958.1000 438.2400 959.1000 438.7200 ;
        RECT 958.1000 416.4800 959.1000 416.9600 ;
        RECT 958.1000 421.9200 959.1000 422.4000 ;
        RECT 958.1000 427.3600 959.1000 427.8400 ;
        RECT 902.3400 438.2400 905.3400 438.7200 ;
        RECT 913.1000 438.2400 914.1000 438.7200 ;
        RECT 902.3400 432.8000 905.3400 433.2800 ;
        RECT 913.1000 432.8000 914.1000 433.2800 ;
        RECT 913.1000 427.3600 914.1000 427.8400 ;
        RECT 913.1000 421.9200 914.1000 422.4000 ;
        RECT 902.3400 427.3600 905.3400 427.8400 ;
        RECT 902.3400 421.9200 905.3400 422.4000 ;
        RECT 902.3400 416.4800 905.3400 416.9600 ;
        RECT 913.1000 416.4800 914.1000 416.9600 ;
        RECT 1136.3400 400.1600 1139.3400 400.6400 ;
        RECT 1136.3400 405.6000 1139.3400 406.0800 ;
        RECT 1136.3400 411.0400 1139.3400 411.5200 ;
        RECT 1136.3400 394.7200 1139.3400 395.2000 ;
        RECT 1136.3400 383.8400 1139.3400 384.3200 ;
        RECT 1136.3400 389.2800 1139.3400 389.7600 ;
        RECT 1093.1000 400.1600 1094.1000 400.6400 ;
        RECT 1093.1000 405.6000 1094.1000 406.0800 ;
        RECT 1093.1000 411.0400 1094.1000 411.5200 ;
        RECT 1093.1000 383.8400 1094.1000 384.3200 ;
        RECT 1093.1000 389.2800 1094.1000 389.7600 ;
        RECT 1093.1000 394.7200 1094.1000 395.2000 ;
        RECT 1136.3400 372.9600 1139.3400 373.4400 ;
        RECT 1136.3400 378.4000 1139.3400 378.8800 ;
        RECT 1136.3400 362.0800 1139.3400 362.5600 ;
        RECT 1136.3400 367.5200 1139.3400 368.0000 ;
        RECT 1136.3400 356.6400 1139.3400 357.1200 ;
        RECT 1093.1000 372.9600 1094.1000 373.4400 ;
        RECT 1093.1000 378.4000 1094.1000 378.8800 ;
        RECT 1093.1000 356.6400 1094.1000 357.1200 ;
        RECT 1093.1000 362.0800 1094.1000 362.5600 ;
        RECT 1093.1000 367.5200 1094.1000 368.0000 ;
        RECT 1048.1000 400.1600 1049.1000 400.6400 ;
        RECT 1048.1000 405.6000 1049.1000 406.0800 ;
        RECT 1048.1000 411.0400 1049.1000 411.5200 ;
        RECT 1048.1000 383.8400 1049.1000 384.3200 ;
        RECT 1048.1000 389.2800 1049.1000 389.7600 ;
        RECT 1048.1000 394.7200 1049.1000 395.2000 ;
        RECT 1048.1000 372.9600 1049.1000 373.4400 ;
        RECT 1048.1000 378.4000 1049.1000 378.8800 ;
        RECT 1048.1000 356.6400 1049.1000 357.1200 ;
        RECT 1048.1000 362.0800 1049.1000 362.5600 ;
        RECT 1048.1000 367.5200 1049.1000 368.0000 ;
        RECT 1136.3400 340.3200 1139.3400 340.8000 ;
        RECT 1136.3400 345.7600 1139.3400 346.2400 ;
        RECT 1136.3400 351.2000 1139.3400 351.6800 ;
        RECT 1136.3400 334.8800 1139.3400 335.3600 ;
        RECT 1136.3400 324.0000 1139.3400 324.4800 ;
        RECT 1136.3400 329.4400 1139.3400 329.9200 ;
        RECT 1093.1000 340.3200 1094.1000 340.8000 ;
        RECT 1093.1000 345.7600 1094.1000 346.2400 ;
        RECT 1093.1000 351.2000 1094.1000 351.6800 ;
        RECT 1093.1000 324.0000 1094.1000 324.4800 ;
        RECT 1093.1000 329.4400 1094.1000 329.9200 ;
        RECT 1093.1000 334.8800 1094.1000 335.3600 ;
        RECT 1136.3400 313.1200 1139.3400 313.6000 ;
        RECT 1136.3400 318.5600 1139.3400 319.0400 ;
        RECT 1093.1000 313.1200 1094.1000 313.6000 ;
        RECT 1093.1000 318.5600 1094.1000 319.0400 ;
        RECT 1048.1000 340.3200 1049.1000 340.8000 ;
        RECT 1048.1000 345.7600 1049.1000 346.2400 ;
        RECT 1048.1000 351.2000 1049.1000 351.6800 ;
        RECT 1048.1000 324.0000 1049.1000 324.4800 ;
        RECT 1048.1000 329.4400 1049.1000 329.9200 ;
        RECT 1048.1000 334.8800 1049.1000 335.3600 ;
        RECT 1048.1000 313.1200 1049.1000 313.6000 ;
        RECT 1048.1000 318.5600 1049.1000 319.0400 ;
        RECT 1003.1000 400.1600 1004.1000 400.6400 ;
        RECT 1003.1000 405.6000 1004.1000 406.0800 ;
        RECT 1003.1000 411.0400 1004.1000 411.5200 ;
        RECT 1003.1000 383.8400 1004.1000 384.3200 ;
        RECT 1003.1000 389.2800 1004.1000 389.7600 ;
        RECT 1003.1000 394.7200 1004.1000 395.2000 ;
        RECT 1003.1000 372.9600 1004.1000 373.4400 ;
        RECT 1003.1000 378.4000 1004.1000 378.8800 ;
        RECT 1003.1000 356.6400 1004.1000 357.1200 ;
        RECT 1003.1000 362.0800 1004.1000 362.5600 ;
        RECT 1003.1000 367.5200 1004.1000 368.0000 ;
        RECT 958.1000 400.1600 959.1000 400.6400 ;
        RECT 958.1000 405.6000 959.1000 406.0800 ;
        RECT 958.1000 411.0400 959.1000 411.5200 ;
        RECT 958.1000 383.8400 959.1000 384.3200 ;
        RECT 958.1000 389.2800 959.1000 389.7600 ;
        RECT 958.1000 394.7200 959.1000 395.2000 ;
        RECT 902.3400 411.0400 905.3400 411.5200 ;
        RECT 913.1000 411.0400 914.1000 411.5200 ;
        RECT 902.3400 400.1600 905.3400 400.6400 ;
        RECT 913.1000 400.1600 914.1000 400.6400 ;
        RECT 902.3400 405.6000 905.3400 406.0800 ;
        RECT 913.1000 405.6000 914.1000 406.0800 ;
        RECT 902.3400 394.7200 905.3400 395.2000 ;
        RECT 913.1000 394.7200 914.1000 395.2000 ;
        RECT 913.1000 389.2800 914.1000 389.7600 ;
        RECT 913.1000 383.8400 914.1000 384.3200 ;
        RECT 902.3400 389.2800 905.3400 389.7600 ;
        RECT 902.3400 383.8400 905.3400 384.3200 ;
        RECT 958.1000 372.9600 959.1000 373.4400 ;
        RECT 958.1000 378.4000 959.1000 378.8800 ;
        RECT 958.1000 356.6400 959.1000 357.1200 ;
        RECT 958.1000 362.0800 959.1000 362.5600 ;
        RECT 958.1000 367.5200 959.1000 368.0000 ;
        RECT 902.3400 378.4000 905.3400 378.8800 ;
        RECT 913.1000 378.4000 914.1000 378.8800 ;
        RECT 902.3400 372.9600 905.3400 373.4400 ;
        RECT 913.1000 372.9600 914.1000 373.4400 ;
        RECT 913.1000 367.5200 914.1000 368.0000 ;
        RECT 913.1000 362.0800 914.1000 362.5600 ;
        RECT 902.3400 367.5200 905.3400 368.0000 ;
        RECT 902.3400 362.0800 905.3400 362.5600 ;
        RECT 902.3400 356.6400 905.3400 357.1200 ;
        RECT 913.1000 356.6400 914.1000 357.1200 ;
        RECT 1003.1000 340.3200 1004.1000 340.8000 ;
        RECT 1003.1000 345.7600 1004.1000 346.2400 ;
        RECT 1003.1000 351.2000 1004.1000 351.6800 ;
        RECT 1003.1000 324.0000 1004.1000 324.4800 ;
        RECT 1003.1000 329.4400 1004.1000 329.9200 ;
        RECT 1003.1000 334.8800 1004.1000 335.3600 ;
        RECT 1003.1000 313.1200 1004.1000 313.6000 ;
        RECT 1003.1000 318.5600 1004.1000 319.0400 ;
        RECT 958.1000 340.3200 959.1000 340.8000 ;
        RECT 958.1000 345.7600 959.1000 346.2400 ;
        RECT 958.1000 351.2000 959.1000 351.6800 ;
        RECT 958.1000 324.0000 959.1000 324.4800 ;
        RECT 958.1000 329.4400 959.1000 329.9200 ;
        RECT 958.1000 334.8800 959.1000 335.3600 ;
        RECT 902.3400 351.2000 905.3400 351.6800 ;
        RECT 913.1000 351.2000 914.1000 351.6800 ;
        RECT 902.3400 340.3200 905.3400 340.8000 ;
        RECT 913.1000 340.3200 914.1000 340.8000 ;
        RECT 902.3400 345.7600 905.3400 346.2400 ;
        RECT 913.1000 345.7600 914.1000 346.2400 ;
        RECT 902.3400 334.8800 905.3400 335.3600 ;
        RECT 913.1000 334.8800 914.1000 335.3600 ;
        RECT 913.1000 329.4400 914.1000 329.9200 ;
        RECT 913.1000 324.0000 914.1000 324.4800 ;
        RECT 902.3400 329.4400 905.3400 329.9200 ;
        RECT 902.3400 324.0000 905.3400 324.4800 ;
        RECT 958.1000 313.1200 959.1000 313.6000 ;
        RECT 958.1000 318.5600 959.1000 319.0400 ;
        RECT 902.3400 318.5600 905.3400 319.0400 ;
        RECT 913.1000 318.5600 914.1000 319.0400 ;
        RECT 902.3400 313.1200 905.3400 313.6000 ;
        RECT 913.1000 313.1200 914.1000 313.6000 ;
        RECT 902.3400 518.0300 1139.3400 521.0300 ;
        RECT 902.3400 304.9300 1139.3400 307.9300 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 75.2900 1094.1000 291.3900 ;
        RECT 1048.1000 75.2900 1049.1000 291.3900 ;
        RECT 1003.1000 75.2900 1004.1000 291.3900 ;
        RECT 958.1000 75.2900 959.1000 291.3900 ;
        RECT 913.1000 75.2900 914.1000 291.3900 ;
        RECT 1136.3400 75.2900 1139.3400 291.3900 ;
        RECT 902.3400 75.2900 905.3400 291.3900 ;
      LAYER met3 ;
        RECT 1136.3400 273.8800 1139.3400 274.3600 ;
        RECT 1136.3400 279.3200 1139.3400 279.8000 ;
        RECT 1093.1000 273.8800 1094.1000 274.3600 ;
        RECT 1093.1000 279.3200 1094.1000 279.8000 ;
        RECT 1136.3400 263.0000 1139.3400 263.4800 ;
        RECT 1136.3400 268.4400 1139.3400 268.9200 ;
        RECT 1136.3400 252.1200 1139.3400 252.6000 ;
        RECT 1136.3400 257.5600 1139.3400 258.0400 ;
        RECT 1136.3400 246.6800 1139.3400 247.1600 ;
        RECT 1093.1000 263.0000 1094.1000 263.4800 ;
        RECT 1093.1000 268.4400 1094.1000 268.9200 ;
        RECT 1093.1000 246.6800 1094.1000 247.1600 ;
        RECT 1093.1000 252.1200 1094.1000 252.6000 ;
        RECT 1093.1000 257.5600 1094.1000 258.0400 ;
        RECT 1048.1000 273.8800 1049.1000 274.3600 ;
        RECT 1048.1000 279.3200 1049.1000 279.8000 ;
        RECT 1048.1000 263.0000 1049.1000 263.4800 ;
        RECT 1048.1000 268.4400 1049.1000 268.9200 ;
        RECT 1048.1000 246.6800 1049.1000 247.1600 ;
        RECT 1048.1000 252.1200 1049.1000 252.6000 ;
        RECT 1048.1000 257.5600 1049.1000 258.0400 ;
        RECT 1136.3400 230.3600 1139.3400 230.8400 ;
        RECT 1136.3400 235.8000 1139.3400 236.2800 ;
        RECT 1136.3400 241.2400 1139.3400 241.7200 ;
        RECT 1136.3400 224.9200 1139.3400 225.4000 ;
        RECT 1136.3400 214.0400 1139.3400 214.5200 ;
        RECT 1136.3400 219.4800 1139.3400 219.9600 ;
        RECT 1093.1000 230.3600 1094.1000 230.8400 ;
        RECT 1093.1000 235.8000 1094.1000 236.2800 ;
        RECT 1093.1000 241.2400 1094.1000 241.7200 ;
        RECT 1093.1000 214.0400 1094.1000 214.5200 ;
        RECT 1093.1000 219.4800 1094.1000 219.9600 ;
        RECT 1093.1000 224.9200 1094.1000 225.4000 ;
        RECT 1136.3400 203.1600 1139.3400 203.6400 ;
        RECT 1136.3400 208.6000 1139.3400 209.0800 ;
        RECT 1136.3400 192.2800 1139.3400 192.7600 ;
        RECT 1136.3400 197.7200 1139.3400 198.2000 ;
        RECT 1136.3400 186.8400 1139.3400 187.3200 ;
        RECT 1093.1000 203.1600 1094.1000 203.6400 ;
        RECT 1093.1000 208.6000 1094.1000 209.0800 ;
        RECT 1093.1000 186.8400 1094.1000 187.3200 ;
        RECT 1093.1000 192.2800 1094.1000 192.7600 ;
        RECT 1093.1000 197.7200 1094.1000 198.2000 ;
        RECT 1048.1000 230.3600 1049.1000 230.8400 ;
        RECT 1048.1000 235.8000 1049.1000 236.2800 ;
        RECT 1048.1000 241.2400 1049.1000 241.7200 ;
        RECT 1048.1000 214.0400 1049.1000 214.5200 ;
        RECT 1048.1000 219.4800 1049.1000 219.9600 ;
        RECT 1048.1000 224.9200 1049.1000 225.4000 ;
        RECT 1048.1000 203.1600 1049.1000 203.6400 ;
        RECT 1048.1000 208.6000 1049.1000 209.0800 ;
        RECT 1048.1000 186.8400 1049.1000 187.3200 ;
        RECT 1048.1000 192.2800 1049.1000 192.7600 ;
        RECT 1048.1000 197.7200 1049.1000 198.2000 ;
        RECT 1003.1000 273.8800 1004.1000 274.3600 ;
        RECT 1003.1000 279.3200 1004.1000 279.8000 ;
        RECT 1003.1000 263.0000 1004.1000 263.4800 ;
        RECT 1003.1000 268.4400 1004.1000 268.9200 ;
        RECT 1003.1000 246.6800 1004.1000 247.1600 ;
        RECT 1003.1000 252.1200 1004.1000 252.6000 ;
        RECT 1003.1000 257.5600 1004.1000 258.0400 ;
        RECT 958.1000 273.8800 959.1000 274.3600 ;
        RECT 958.1000 279.3200 959.1000 279.8000 ;
        RECT 913.1000 279.3200 914.1000 279.8000 ;
        RECT 913.1000 273.8800 914.1000 274.3600 ;
        RECT 902.3400 279.3200 905.3400 279.8000 ;
        RECT 902.3400 273.8800 905.3400 274.3600 ;
        RECT 958.1000 263.0000 959.1000 263.4800 ;
        RECT 958.1000 268.4400 959.1000 268.9200 ;
        RECT 958.1000 246.6800 959.1000 247.1600 ;
        RECT 958.1000 252.1200 959.1000 252.6000 ;
        RECT 958.1000 257.5600 959.1000 258.0400 ;
        RECT 902.3400 268.4400 905.3400 268.9200 ;
        RECT 913.1000 268.4400 914.1000 268.9200 ;
        RECT 902.3400 263.0000 905.3400 263.4800 ;
        RECT 913.1000 263.0000 914.1000 263.4800 ;
        RECT 913.1000 257.5600 914.1000 258.0400 ;
        RECT 913.1000 252.1200 914.1000 252.6000 ;
        RECT 902.3400 257.5600 905.3400 258.0400 ;
        RECT 902.3400 252.1200 905.3400 252.6000 ;
        RECT 902.3400 246.6800 905.3400 247.1600 ;
        RECT 913.1000 246.6800 914.1000 247.1600 ;
        RECT 1003.1000 230.3600 1004.1000 230.8400 ;
        RECT 1003.1000 235.8000 1004.1000 236.2800 ;
        RECT 1003.1000 241.2400 1004.1000 241.7200 ;
        RECT 1003.1000 214.0400 1004.1000 214.5200 ;
        RECT 1003.1000 219.4800 1004.1000 219.9600 ;
        RECT 1003.1000 224.9200 1004.1000 225.4000 ;
        RECT 1003.1000 203.1600 1004.1000 203.6400 ;
        RECT 1003.1000 208.6000 1004.1000 209.0800 ;
        RECT 1003.1000 186.8400 1004.1000 187.3200 ;
        RECT 1003.1000 192.2800 1004.1000 192.7600 ;
        RECT 1003.1000 197.7200 1004.1000 198.2000 ;
        RECT 958.1000 230.3600 959.1000 230.8400 ;
        RECT 958.1000 235.8000 959.1000 236.2800 ;
        RECT 958.1000 241.2400 959.1000 241.7200 ;
        RECT 958.1000 214.0400 959.1000 214.5200 ;
        RECT 958.1000 219.4800 959.1000 219.9600 ;
        RECT 958.1000 224.9200 959.1000 225.4000 ;
        RECT 902.3400 241.2400 905.3400 241.7200 ;
        RECT 913.1000 241.2400 914.1000 241.7200 ;
        RECT 902.3400 230.3600 905.3400 230.8400 ;
        RECT 913.1000 230.3600 914.1000 230.8400 ;
        RECT 902.3400 235.8000 905.3400 236.2800 ;
        RECT 913.1000 235.8000 914.1000 236.2800 ;
        RECT 902.3400 224.9200 905.3400 225.4000 ;
        RECT 913.1000 224.9200 914.1000 225.4000 ;
        RECT 913.1000 219.4800 914.1000 219.9600 ;
        RECT 913.1000 214.0400 914.1000 214.5200 ;
        RECT 902.3400 219.4800 905.3400 219.9600 ;
        RECT 902.3400 214.0400 905.3400 214.5200 ;
        RECT 958.1000 203.1600 959.1000 203.6400 ;
        RECT 958.1000 208.6000 959.1000 209.0800 ;
        RECT 958.1000 186.8400 959.1000 187.3200 ;
        RECT 958.1000 192.2800 959.1000 192.7600 ;
        RECT 958.1000 197.7200 959.1000 198.2000 ;
        RECT 902.3400 208.6000 905.3400 209.0800 ;
        RECT 913.1000 208.6000 914.1000 209.0800 ;
        RECT 902.3400 203.1600 905.3400 203.6400 ;
        RECT 913.1000 203.1600 914.1000 203.6400 ;
        RECT 913.1000 197.7200 914.1000 198.2000 ;
        RECT 913.1000 192.2800 914.1000 192.7600 ;
        RECT 902.3400 197.7200 905.3400 198.2000 ;
        RECT 902.3400 192.2800 905.3400 192.7600 ;
        RECT 902.3400 186.8400 905.3400 187.3200 ;
        RECT 913.1000 186.8400 914.1000 187.3200 ;
        RECT 1136.3400 170.5200 1139.3400 171.0000 ;
        RECT 1136.3400 175.9600 1139.3400 176.4400 ;
        RECT 1136.3400 181.4000 1139.3400 181.8800 ;
        RECT 1136.3400 165.0800 1139.3400 165.5600 ;
        RECT 1136.3400 154.2000 1139.3400 154.6800 ;
        RECT 1136.3400 159.6400 1139.3400 160.1200 ;
        RECT 1093.1000 170.5200 1094.1000 171.0000 ;
        RECT 1093.1000 175.9600 1094.1000 176.4400 ;
        RECT 1093.1000 181.4000 1094.1000 181.8800 ;
        RECT 1093.1000 154.2000 1094.1000 154.6800 ;
        RECT 1093.1000 159.6400 1094.1000 160.1200 ;
        RECT 1093.1000 165.0800 1094.1000 165.5600 ;
        RECT 1136.3400 143.3200 1139.3400 143.8000 ;
        RECT 1136.3400 148.7600 1139.3400 149.2400 ;
        RECT 1136.3400 132.4400 1139.3400 132.9200 ;
        RECT 1136.3400 137.8800 1139.3400 138.3600 ;
        RECT 1136.3400 127.0000 1139.3400 127.4800 ;
        RECT 1093.1000 143.3200 1094.1000 143.8000 ;
        RECT 1093.1000 148.7600 1094.1000 149.2400 ;
        RECT 1093.1000 127.0000 1094.1000 127.4800 ;
        RECT 1093.1000 132.4400 1094.1000 132.9200 ;
        RECT 1093.1000 137.8800 1094.1000 138.3600 ;
        RECT 1048.1000 170.5200 1049.1000 171.0000 ;
        RECT 1048.1000 175.9600 1049.1000 176.4400 ;
        RECT 1048.1000 181.4000 1049.1000 181.8800 ;
        RECT 1048.1000 154.2000 1049.1000 154.6800 ;
        RECT 1048.1000 159.6400 1049.1000 160.1200 ;
        RECT 1048.1000 165.0800 1049.1000 165.5600 ;
        RECT 1048.1000 143.3200 1049.1000 143.8000 ;
        RECT 1048.1000 148.7600 1049.1000 149.2400 ;
        RECT 1048.1000 127.0000 1049.1000 127.4800 ;
        RECT 1048.1000 132.4400 1049.1000 132.9200 ;
        RECT 1048.1000 137.8800 1049.1000 138.3600 ;
        RECT 1136.3400 110.6800 1139.3400 111.1600 ;
        RECT 1136.3400 116.1200 1139.3400 116.6000 ;
        RECT 1136.3400 121.5600 1139.3400 122.0400 ;
        RECT 1136.3400 105.2400 1139.3400 105.7200 ;
        RECT 1136.3400 94.3600 1139.3400 94.8400 ;
        RECT 1136.3400 99.8000 1139.3400 100.2800 ;
        RECT 1093.1000 110.6800 1094.1000 111.1600 ;
        RECT 1093.1000 116.1200 1094.1000 116.6000 ;
        RECT 1093.1000 121.5600 1094.1000 122.0400 ;
        RECT 1093.1000 94.3600 1094.1000 94.8400 ;
        RECT 1093.1000 99.8000 1094.1000 100.2800 ;
        RECT 1093.1000 105.2400 1094.1000 105.7200 ;
        RECT 1136.3400 83.4800 1139.3400 83.9600 ;
        RECT 1136.3400 88.9200 1139.3400 89.4000 ;
        RECT 1093.1000 83.4800 1094.1000 83.9600 ;
        RECT 1093.1000 88.9200 1094.1000 89.4000 ;
        RECT 1048.1000 110.6800 1049.1000 111.1600 ;
        RECT 1048.1000 116.1200 1049.1000 116.6000 ;
        RECT 1048.1000 121.5600 1049.1000 122.0400 ;
        RECT 1048.1000 94.3600 1049.1000 94.8400 ;
        RECT 1048.1000 99.8000 1049.1000 100.2800 ;
        RECT 1048.1000 105.2400 1049.1000 105.7200 ;
        RECT 1048.1000 83.4800 1049.1000 83.9600 ;
        RECT 1048.1000 88.9200 1049.1000 89.4000 ;
        RECT 1003.1000 170.5200 1004.1000 171.0000 ;
        RECT 1003.1000 175.9600 1004.1000 176.4400 ;
        RECT 1003.1000 181.4000 1004.1000 181.8800 ;
        RECT 1003.1000 154.2000 1004.1000 154.6800 ;
        RECT 1003.1000 159.6400 1004.1000 160.1200 ;
        RECT 1003.1000 165.0800 1004.1000 165.5600 ;
        RECT 1003.1000 143.3200 1004.1000 143.8000 ;
        RECT 1003.1000 148.7600 1004.1000 149.2400 ;
        RECT 1003.1000 127.0000 1004.1000 127.4800 ;
        RECT 1003.1000 132.4400 1004.1000 132.9200 ;
        RECT 1003.1000 137.8800 1004.1000 138.3600 ;
        RECT 958.1000 170.5200 959.1000 171.0000 ;
        RECT 958.1000 175.9600 959.1000 176.4400 ;
        RECT 958.1000 181.4000 959.1000 181.8800 ;
        RECT 958.1000 154.2000 959.1000 154.6800 ;
        RECT 958.1000 159.6400 959.1000 160.1200 ;
        RECT 958.1000 165.0800 959.1000 165.5600 ;
        RECT 902.3400 181.4000 905.3400 181.8800 ;
        RECT 913.1000 181.4000 914.1000 181.8800 ;
        RECT 902.3400 170.5200 905.3400 171.0000 ;
        RECT 913.1000 170.5200 914.1000 171.0000 ;
        RECT 902.3400 175.9600 905.3400 176.4400 ;
        RECT 913.1000 175.9600 914.1000 176.4400 ;
        RECT 902.3400 165.0800 905.3400 165.5600 ;
        RECT 913.1000 165.0800 914.1000 165.5600 ;
        RECT 913.1000 159.6400 914.1000 160.1200 ;
        RECT 913.1000 154.2000 914.1000 154.6800 ;
        RECT 902.3400 159.6400 905.3400 160.1200 ;
        RECT 902.3400 154.2000 905.3400 154.6800 ;
        RECT 958.1000 143.3200 959.1000 143.8000 ;
        RECT 958.1000 148.7600 959.1000 149.2400 ;
        RECT 958.1000 127.0000 959.1000 127.4800 ;
        RECT 958.1000 132.4400 959.1000 132.9200 ;
        RECT 958.1000 137.8800 959.1000 138.3600 ;
        RECT 902.3400 148.7600 905.3400 149.2400 ;
        RECT 913.1000 148.7600 914.1000 149.2400 ;
        RECT 902.3400 143.3200 905.3400 143.8000 ;
        RECT 913.1000 143.3200 914.1000 143.8000 ;
        RECT 913.1000 137.8800 914.1000 138.3600 ;
        RECT 913.1000 132.4400 914.1000 132.9200 ;
        RECT 902.3400 137.8800 905.3400 138.3600 ;
        RECT 902.3400 132.4400 905.3400 132.9200 ;
        RECT 902.3400 127.0000 905.3400 127.4800 ;
        RECT 913.1000 127.0000 914.1000 127.4800 ;
        RECT 1003.1000 110.6800 1004.1000 111.1600 ;
        RECT 1003.1000 116.1200 1004.1000 116.6000 ;
        RECT 1003.1000 121.5600 1004.1000 122.0400 ;
        RECT 1003.1000 94.3600 1004.1000 94.8400 ;
        RECT 1003.1000 99.8000 1004.1000 100.2800 ;
        RECT 1003.1000 105.2400 1004.1000 105.7200 ;
        RECT 1003.1000 83.4800 1004.1000 83.9600 ;
        RECT 1003.1000 88.9200 1004.1000 89.4000 ;
        RECT 958.1000 110.6800 959.1000 111.1600 ;
        RECT 958.1000 116.1200 959.1000 116.6000 ;
        RECT 958.1000 121.5600 959.1000 122.0400 ;
        RECT 958.1000 94.3600 959.1000 94.8400 ;
        RECT 958.1000 99.8000 959.1000 100.2800 ;
        RECT 958.1000 105.2400 959.1000 105.7200 ;
        RECT 902.3400 121.5600 905.3400 122.0400 ;
        RECT 913.1000 121.5600 914.1000 122.0400 ;
        RECT 902.3400 110.6800 905.3400 111.1600 ;
        RECT 913.1000 110.6800 914.1000 111.1600 ;
        RECT 902.3400 116.1200 905.3400 116.6000 ;
        RECT 913.1000 116.1200 914.1000 116.6000 ;
        RECT 902.3400 105.2400 905.3400 105.7200 ;
        RECT 913.1000 105.2400 914.1000 105.7200 ;
        RECT 913.1000 99.8000 914.1000 100.2800 ;
        RECT 913.1000 94.3600 914.1000 94.8400 ;
        RECT 902.3400 99.8000 905.3400 100.2800 ;
        RECT 902.3400 94.3600 905.3400 94.8400 ;
        RECT 958.1000 83.4800 959.1000 83.9600 ;
        RECT 958.1000 88.9200 959.1000 89.4000 ;
        RECT 902.3400 88.9200 905.3400 89.4000 ;
        RECT 913.1000 88.9200 914.1000 89.4000 ;
        RECT 902.3400 83.4800 905.3400 83.9600 ;
        RECT 913.1000 83.4800 914.1000 83.9600 ;
        RECT 902.3400 288.3900 1139.3400 291.3900 ;
        RECT 902.3400 75.2900 1139.3400 78.2900 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'S_term_single2'
    PORT
      LAYER met4 ;
        RECT 903.3400 34.6700 905.3400 61.6000 ;
        RECT 1136.3400 34.6700 1138.3400 61.6000 ;
      LAYER met3 ;
        RECT 1136.3400 51.3800 1138.3400 51.8600 ;
        RECT 903.3400 51.3800 905.3400 51.8600 ;
        RECT 1136.3400 45.9400 1138.3400 46.4200 ;
        RECT 1136.3400 40.5000 1138.3400 40.9800 ;
        RECT 903.3400 45.9400 905.3400 46.4200 ;
        RECT 903.3400 40.5000 905.3400 40.9800 ;
        RECT 903.3400 59.6000 1138.3400 61.6000 ;
        RECT 903.3400 34.6700 1138.3400 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single2'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 2601.3300 1094.1000 2817.4300 ;
        RECT 1048.1000 2601.3300 1049.1000 2817.4300 ;
        RECT 1003.1000 2601.3300 1004.1000 2817.4300 ;
        RECT 958.1000 2601.3300 959.1000 2817.4300 ;
        RECT 913.1000 2601.3300 914.1000 2817.4300 ;
        RECT 1136.3400 2601.3300 1139.3400 2817.4300 ;
        RECT 902.3400 2601.3300 905.3400 2817.4300 ;
      LAYER met3 ;
        RECT 1136.3400 2799.9200 1139.3400 2800.4000 ;
        RECT 1136.3400 2805.3600 1139.3400 2805.8400 ;
        RECT 1093.1000 2799.9200 1094.1000 2800.4000 ;
        RECT 1093.1000 2805.3600 1094.1000 2805.8400 ;
        RECT 1136.3400 2789.0400 1139.3400 2789.5200 ;
        RECT 1136.3400 2794.4800 1139.3400 2794.9600 ;
        RECT 1136.3400 2778.1600 1139.3400 2778.6400 ;
        RECT 1136.3400 2783.6000 1139.3400 2784.0800 ;
        RECT 1136.3400 2772.7200 1139.3400 2773.2000 ;
        RECT 1093.1000 2789.0400 1094.1000 2789.5200 ;
        RECT 1093.1000 2794.4800 1094.1000 2794.9600 ;
        RECT 1093.1000 2772.7200 1094.1000 2773.2000 ;
        RECT 1093.1000 2778.1600 1094.1000 2778.6400 ;
        RECT 1093.1000 2783.6000 1094.1000 2784.0800 ;
        RECT 1048.1000 2799.9200 1049.1000 2800.4000 ;
        RECT 1048.1000 2805.3600 1049.1000 2805.8400 ;
        RECT 1048.1000 2789.0400 1049.1000 2789.5200 ;
        RECT 1048.1000 2794.4800 1049.1000 2794.9600 ;
        RECT 1048.1000 2772.7200 1049.1000 2773.2000 ;
        RECT 1048.1000 2778.1600 1049.1000 2778.6400 ;
        RECT 1048.1000 2783.6000 1049.1000 2784.0800 ;
        RECT 1136.3400 2756.4000 1139.3400 2756.8800 ;
        RECT 1136.3400 2761.8400 1139.3400 2762.3200 ;
        RECT 1136.3400 2767.2800 1139.3400 2767.7600 ;
        RECT 1136.3400 2750.9600 1139.3400 2751.4400 ;
        RECT 1136.3400 2740.0800 1139.3400 2740.5600 ;
        RECT 1136.3400 2745.5200 1139.3400 2746.0000 ;
        RECT 1093.1000 2756.4000 1094.1000 2756.8800 ;
        RECT 1093.1000 2761.8400 1094.1000 2762.3200 ;
        RECT 1093.1000 2767.2800 1094.1000 2767.7600 ;
        RECT 1093.1000 2740.0800 1094.1000 2740.5600 ;
        RECT 1093.1000 2745.5200 1094.1000 2746.0000 ;
        RECT 1093.1000 2750.9600 1094.1000 2751.4400 ;
        RECT 1136.3400 2729.2000 1139.3400 2729.6800 ;
        RECT 1136.3400 2734.6400 1139.3400 2735.1200 ;
        RECT 1136.3400 2718.3200 1139.3400 2718.8000 ;
        RECT 1136.3400 2723.7600 1139.3400 2724.2400 ;
        RECT 1136.3400 2712.8800 1139.3400 2713.3600 ;
        RECT 1093.1000 2729.2000 1094.1000 2729.6800 ;
        RECT 1093.1000 2734.6400 1094.1000 2735.1200 ;
        RECT 1093.1000 2712.8800 1094.1000 2713.3600 ;
        RECT 1093.1000 2718.3200 1094.1000 2718.8000 ;
        RECT 1093.1000 2723.7600 1094.1000 2724.2400 ;
        RECT 1048.1000 2756.4000 1049.1000 2756.8800 ;
        RECT 1048.1000 2761.8400 1049.1000 2762.3200 ;
        RECT 1048.1000 2767.2800 1049.1000 2767.7600 ;
        RECT 1048.1000 2740.0800 1049.1000 2740.5600 ;
        RECT 1048.1000 2745.5200 1049.1000 2746.0000 ;
        RECT 1048.1000 2750.9600 1049.1000 2751.4400 ;
        RECT 1048.1000 2729.2000 1049.1000 2729.6800 ;
        RECT 1048.1000 2734.6400 1049.1000 2735.1200 ;
        RECT 1048.1000 2712.8800 1049.1000 2713.3600 ;
        RECT 1048.1000 2718.3200 1049.1000 2718.8000 ;
        RECT 1048.1000 2723.7600 1049.1000 2724.2400 ;
        RECT 1003.1000 2799.9200 1004.1000 2800.4000 ;
        RECT 1003.1000 2805.3600 1004.1000 2805.8400 ;
        RECT 1003.1000 2789.0400 1004.1000 2789.5200 ;
        RECT 1003.1000 2794.4800 1004.1000 2794.9600 ;
        RECT 1003.1000 2772.7200 1004.1000 2773.2000 ;
        RECT 1003.1000 2778.1600 1004.1000 2778.6400 ;
        RECT 1003.1000 2783.6000 1004.1000 2784.0800 ;
        RECT 958.1000 2799.9200 959.1000 2800.4000 ;
        RECT 958.1000 2805.3600 959.1000 2805.8400 ;
        RECT 913.1000 2805.3600 914.1000 2805.8400 ;
        RECT 913.1000 2799.9200 914.1000 2800.4000 ;
        RECT 902.3400 2805.3600 905.3400 2805.8400 ;
        RECT 902.3400 2799.9200 905.3400 2800.4000 ;
        RECT 958.1000 2789.0400 959.1000 2789.5200 ;
        RECT 958.1000 2794.4800 959.1000 2794.9600 ;
        RECT 958.1000 2772.7200 959.1000 2773.2000 ;
        RECT 958.1000 2778.1600 959.1000 2778.6400 ;
        RECT 958.1000 2783.6000 959.1000 2784.0800 ;
        RECT 902.3400 2794.4800 905.3400 2794.9600 ;
        RECT 913.1000 2794.4800 914.1000 2794.9600 ;
        RECT 902.3400 2789.0400 905.3400 2789.5200 ;
        RECT 913.1000 2789.0400 914.1000 2789.5200 ;
        RECT 913.1000 2783.6000 914.1000 2784.0800 ;
        RECT 913.1000 2778.1600 914.1000 2778.6400 ;
        RECT 902.3400 2783.6000 905.3400 2784.0800 ;
        RECT 902.3400 2778.1600 905.3400 2778.6400 ;
        RECT 902.3400 2772.7200 905.3400 2773.2000 ;
        RECT 913.1000 2772.7200 914.1000 2773.2000 ;
        RECT 1003.1000 2756.4000 1004.1000 2756.8800 ;
        RECT 1003.1000 2761.8400 1004.1000 2762.3200 ;
        RECT 1003.1000 2767.2800 1004.1000 2767.7600 ;
        RECT 1003.1000 2740.0800 1004.1000 2740.5600 ;
        RECT 1003.1000 2745.5200 1004.1000 2746.0000 ;
        RECT 1003.1000 2750.9600 1004.1000 2751.4400 ;
        RECT 1003.1000 2729.2000 1004.1000 2729.6800 ;
        RECT 1003.1000 2734.6400 1004.1000 2735.1200 ;
        RECT 1003.1000 2712.8800 1004.1000 2713.3600 ;
        RECT 1003.1000 2718.3200 1004.1000 2718.8000 ;
        RECT 1003.1000 2723.7600 1004.1000 2724.2400 ;
        RECT 958.1000 2756.4000 959.1000 2756.8800 ;
        RECT 958.1000 2761.8400 959.1000 2762.3200 ;
        RECT 958.1000 2767.2800 959.1000 2767.7600 ;
        RECT 958.1000 2740.0800 959.1000 2740.5600 ;
        RECT 958.1000 2745.5200 959.1000 2746.0000 ;
        RECT 958.1000 2750.9600 959.1000 2751.4400 ;
        RECT 902.3400 2767.2800 905.3400 2767.7600 ;
        RECT 913.1000 2767.2800 914.1000 2767.7600 ;
        RECT 902.3400 2756.4000 905.3400 2756.8800 ;
        RECT 913.1000 2756.4000 914.1000 2756.8800 ;
        RECT 902.3400 2761.8400 905.3400 2762.3200 ;
        RECT 913.1000 2761.8400 914.1000 2762.3200 ;
        RECT 902.3400 2750.9600 905.3400 2751.4400 ;
        RECT 913.1000 2750.9600 914.1000 2751.4400 ;
        RECT 913.1000 2745.5200 914.1000 2746.0000 ;
        RECT 913.1000 2740.0800 914.1000 2740.5600 ;
        RECT 902.3400 2745.5200 905.3400 2746.0000 ;
        RECT 902.3400 2740.0800 905.3400 2740.5600 ;
        RECT 958.1000 2729.2000 959.1000 2729.6800 ;
        RECT 958.1000 2734.6400 959.1000 2735.1200 ;
        RECT 958.1000 2712.8800 959.1000 2713.3600 ;
        RECT 958.1000 2718.3200 959.1000 2718.8000 ;
        RECT 958.1000 2723.7600 959.1000 2724.2400 ;
        RECT 902.3400 2734.6400 905.3400 2735.1200 ;
        RECT 913.1000 2734.6400 914.1000 2735.1200 ;
        RECT 902.3400 2729.2000 905.3400 2729.6800 ;
        RECT 913.1000 2729.2000 914.1000 2729.6800 ;
        RECT 913.1000 2723.7600 914.1000 2724.2400 ;
        RECT 913.1000 2718.3200 914.1000 2718.8000 ;
        RECT 902.3400 2723.7600 905.3400 2724.2400 ;
        RECT 902.3400 2718.3200 905.3400 2718.8000 ;
        RECT 902.3400 2712.8800 905.3400 2713.3600 ;
        RECT 913.1000 2712.8800 914.1000 2713.3600 ;
        RECT 1136.3400 2696.5600 1139.3400 2697.0400 ;
        RECT 1136.3400 2702.0000 1139.3400 2702.4800 ;
        RECT 1136.3400 2707.4400 1139.3400 2707.9200 ;
        RECT 1136.3400 2691.1200 1139.3400 2691.6000 ;
        RECT 1136.3400 2680.2400 1139.3400 2680.7200 ;
        RECT 1136.3400 2685.6800 1139.3400 2686.1600 ;
        RECT 1093.1000 2696.5600 1094.1000 2697.0400 ;
        RECT 1093.1000 2702.0000 1094.1000 2702.4800 ;
        RECT 1093.1000 2707.4400 1094.1000 2707.9200 ;
        RECT 1093.1000 2680.2400 1094.1000 2680.7200 ;
        RECT 1093.1000 2685.6800 1094.1000 2686.1600 ;
        RECT 1093.1000 2691.1200 1094.1000 2691.6000 ;
        RECT 1136.3400 2669.3600 1139.3400 2669.8400 ;
        RECT 1136.3400 2674.8000 1139.3400 2675.2800 ;
        RECT 1136.3400 2658.4800 1139.3400 2658.9600 ;
        RECT 1136.3400 2663.9200 1139.3400 2664.4000 ;
        RECT 1136.3400 2653.0400 1139.3400 2653.5200 ;
        RECT 1093.1000 2669.3600 1094.1000 2669.8400 ;
        RECT 1093.1000 2674.8000 1094.1000 2675.2800 ;
        RECT 1093.1000 2653.0400 1094.1000 2653.5200 ;
        RECT 1093.1000 2658.4800 1094.1000 2658.9600 ;
        RECT 1093.1000 2663.9200 1094.1000 2664.4000 ;
        RECT 1048.1000 2696.5600 1049.1000 2697.0400 ;
        RECT 1048.1000 2702.0000 1049.1000 2702.4800 ;
        RECT 1048.1000 2707.4400 1049.1000 2707.9200 ;
        RECT 1048.1000 2680.2400 1049.1000 2680.7200 ;
        RECT 1048.1000 2685.6800 1049.1000 2686.1600 ;
        RECT 1048.1000 2691.1200 1049.1000 2691.6000 ;
        RECT 1048.1000 2669.3600 1049.1000 2669.8400 ;
        RECT 1048.1000 2674.8000 1049.1000 2675.2800 ;
        RECT 1048.1000 2653.0400 1049.1000 2653.5200 ;
        RECT 1048.1000 2658.4800 1049.1000 2658.9600 ;
        RECT 1048.1000 2663.9200 1049.1000 2664.4000 ;
        RECT 1136.3400 2636.7200 1139.3400 2637.2000 ;
        RECT 1136.3400 2642.1600 1139.3400 2642.6400 ;
        RECT 1136.3400 2647.6000 1139.3400 2648.0800 ;
        RECT 1136.3400 2631.2800 1139.3400 2631.7600 ;
        RECT 1136.3400 2620.4000 1139.3400 2620.8800 ;
        RECT 1136.3400 2625.8400 1139.3400 2626.3200 ;
        RECT 1093.1000 2636.7200 1094.1000 2637.2000 ;
        RECT 1093.1000 2642.1600 1094.1000 2642.6400 ;
        RECT 1093.1000 2647.6000 1094.1000 2648.0800 ;
        RECT 1093.1000 2620.4000 1094.1000 2620.8800 ;
        RECT 1093.1000 2625.8400 1094.1000 2626.3200 ;
        RECT 1093.1000 2631.2800 1094.1000 2631.7600 ;
        RECT 1136.3400 2609.5200 1139.3400 2610.0000 ;
        RECT 1136.3400 2614.9600 1139.3400 2615.4400 ;
        RECT 1093.1000 2609.5200 1094.1000 2610.0000 ;
        RECT 1093.1000 2614.9600 1094.1000 2615.4400 ;
        RECT 1048.1000 2636.7200 1049.1000 2637.2000 ;
        RECT 1048.1000 2642.1600 1049.1000 2642.6400 ;
        RECT 1048.1000 2647.6000 1049.1000 2648.0800 ;
        RECT 1048.1000 2620.4000 1049.1000 2620.8800 ;
        RECT 1048.1000 2625.8400 1049.1000 2626.3200 ;
        RECT 1048.1000 2631.2800 1049.1000 2631.7600 ;
        RECT 1048.1000 2609.5200 1049.1000 2610.0000 ;
        RECT 1048.1000 2614.9600 1049.1000 2615.4400 ;
        RECT 1003.1000 2696.5600 1004.1000 2697.0400 ;
        RECT 1003.1000 2702.0000 1004.1000 2702.4800 ;
        RECT 1003.1000 2707.4400 1004.1000 2707.9200 ;
        RECT 1003.1000 2680.2400 1004.1000 2680.7200 ;
        RECT 1003.1000 2685.6800 1004.1000 2686.1600 ;
        RECT 1003.1000 2691.1200 1004.1000 2691.6000 ;
        RECT 1003.1000 2669.3600 1004.1000 2669.8400 ;
        RECT 1003.1000 2674.8000 1004.1000 2675.2800 ;
        RECT 1003.1000 2653.0400 1004.1000 2653.5200 ;
        RECT 1003.1000 2658.4800 1004.1000 2658.9600 ;
        RECT 1003.1000 2663.9200 1004.1000 2664.4000 ;
        RECT 958.1000 2696.5600 959.1000 2697.0400 ;
        RECT 958.1000 2702.0000 959.1000 2702.4800 ;
        RECT 958.1000 2707.4400 959.1000 2707.9200 ;
        RECT 958.1000 2680.2400 959.1000 2680.7200 ;
        RECT 958.1000 2685.6800 959.1000 2686.1600 ;
        RECT 958.1000 2691.1200 959.1000 2691.6000 ;
        RECT 902.3400 2707.4400 905.3400 2707.9200 ;
        RECT 913.1000 2707.4400 914.1000 2707.9200 ;
        RECT 902.3400 2696.5600 905.3400 2697.0400 ;
        RECT 913.1000 2696.5600 914.1000 2697.0400 ;
        RECT 902.3400 2702.0000 905.3400 2702.4800 ;
        RECT 913.1000 2702.0000 914.1000 2702.4800 ;
        RECT 902.3400 2691.1200 905.3400 2691.6000 ;
        RECT 913.1000 2691.1200 914.1000 2691.6000 ;
        RECT 913.1000 2685.6800 914.1000 2686.1600 ;
        RECT 913.1000 2680.2400 914.1000 2680.7200 ;
        RECT 902.3400 2685.6800 905.3400 2686.1600 ;
        RECT 902.3400 2680.2400 905.3400 2680.7200 ;
        RECT 958.1000 2669.3600 959.1000 2669.8400 ;
        RECT 958.1000 2674.8000 959.1000 2675.2800 ;
        RECT 958.1000 2653.0400 959.1000 2653.5200 ;
        RECT 958.1000 2658.4800 959.1000 2658.9600 ;
        RECT 958.1000 2663.9200 959.1000 2664.4000 ;
        RECT 902.3400 2674.8000 905.3400 2675.2800 ;
        RECT 913.1000 2674.8000 914.1000 2675.2800 ;
        RECT 902.3400 2669.3600 905.3400 2669.8400 ;
        RECT 913.1000 2669.3600 914.1000 2669.8400 ;
        RECT 913.1000 2663.9200 914.1000 2664.4000 ;
        RECT 913.1000 2658.4800 914.1000 2658.9600 ;
        RECT 902.3400 2663.9200 905.3400 2664.4000 ;
        RECT 902.3400 2658.4800 905.3400 2658.9600 ;
        RECT 902.3400 2653.0400 905.3400 2653.5200 ;
        RECT 913.1000 2653.0400 914.1000 2653.5200 ;
        RECT 1003.1000 2636.7200 1004.1000 2637.2000 ;
        RECT 1003.1000 2642.1600 1004.1000 2642.6400 ;
        RECT 1003.1000 2647.6000 1004.1000 2648.0800 ;
        RECT 1003.1000 2620.4000 1004.1000 2620.8800 ;
        RECT 1003.1000 2625.8400 1004.1000 2626.3200 ;
        RECT 1003.1000 2631.2800 1004.1000 2631.7600 ;
        RECT 1003.1000 2609.5200 1004.1000 2610.0000 ;
        RECT 1003.1000 2614.9600 1004.1000 2615.4400 ;
        RECT 958.1000 2636.7200 959.1000 2637.2000 ;
        RECT 958.1000 2642.1600 959.1000 2642.6400 ;
        RECT 958.1000 2647.6000 959.1000 2648.0800 ;
        RECT 958.1000 2620.4000 959.1000 2620.8800 ;
        RECT 958.1000 2625.8400 959.1000 2626.3200 ;
        RECT 958.1000 2631.2800 959.1000 2631.7600 ;
        RECT 902.3400 2647.6000 905.3400 2648.0800 ;
        RECT 913.1000 2647.6000 914.1000 2648.0800 ;
        RECT 902.3400 2636.7200 905.3400 2637.2000 ;
        RECT 913.1000 2636.7200 914.1000 2637.2000 ;
        RECT 902.3400 2642.1600 905.3400 2642.6400 ;
        RECT 913.1000 2642.1600 914.1000 2642.6400 ;
        RECT 902.3400 2631.2800 905.3400 2631.7600 ;
        RECT 913.1000 2631.2800 914.1000 2631.7600 ;
        RECT 913.1000 2625.8400 914.1000 2626.3200 ;
        RECT 913.1000 2620.4000 914.1000 2620.8800 ;
        RECT 902.3400 2625.8400 905.3400 2626.3200 ;
        RECT 902.3400 2620.4000 905.3400 2620.8800 ;
        RECT 958.1000 2609.5200 959.1000 2610.0000 ;
        RECT 958.1000 2614.9600 959.1000 2615.4400 ;
        RECT 902.3400 2614.9600 905.3400 2615.4400 ;
        RECT 913.1000 2614.9600 914.1000 2615.4400 ;
        RECT 902.3400 2609.5200 905.3400 2610.0000 ;
        RECT 913.1000 2609.5200 914.1000 2610.0000 ;
        RECT 902.3400 2814.4300 1139.3400 2817.4300 ;
        RECT 902.3400 2601.3300 1139.3400 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 2371.6900 1094.1000 2587.7900 ;
        RECT 1048.1000 2371.6900 1049.1000 2587.7900 ;
        RECT 1003.1000 2371.6900 1004.1000 2587.7900 ;
        RECT 958.1000 2371.6900 959.1000 2587.7900 ;
        RECT 913.1000 2371.6900 914.1000 2587.7900 ;
        RECT 1136.3400 2371.6900 1139.3400 2587.7900 ;
        RECT 902.3400 2371.6900 905.3400 2587.7900 ;
      LAYER met3 ;
        RECT 1136.3400 2570.2800 1139.3400 2570.7600 ;
        RECT 1136.3400 2575.7200 1139.3400 2576.2000 ;
        RECT 1093.1000 2570.2800 1094.1000 2570.7600 ;
        RECT 1093.1000 2575.7200 1094.1000 2576.2000 ;
        RECT 1136.3400 2559.4000 1139.3400 2559.8800 ;
        RECT 1136.3400 2564.8400 1139.3400 2565.3200 ;
        RECT 1136.3400 2548.5200 1139.3400 2549.0000 ;
        RECT 1136.3400 2553.9600 1139.3400 2554.4400 ;
        RECT 1136.3400 2543.0800 1139.3400 2543.5600 ;
        RECT 1093.1000 2559.4000 1094.1000 2559.8800 ;
        RECT 1093.1000 2564.8400 1094.1000 2565.3200 ;
        RECT 1093.1000 2543.0800 1094.1000 2543.5600 ;
        RECT 1093.1000 2548.5200 1094.1000 2549.0000 ;
        RECT 1093.1000 2553.9600 1094.1000 2554.4400 ;
        RECT 1048.1000 2570.2800 1049.1000 2570.7600 ;
        RECT 1048.1000 2575.7200 1049.1000 2576.2000 ;
        RECT 1048.1000 2559.4000 1049.1000 2559.8800 ;
        RECT 1048.1000 2564.8400 1049.1000 2565.3200 ;
        RECT 1048.1000 2543.0800 1049.1000 2543.5600 ;
        RECT 1048.1000 2548.5200 1049.1000 2549.0000 ;
        RECT 1048.1000 2553.9600 1049.1000 2554.4400 ;
        RECT 1136.3400 2526.7600 1139.3400 2527.2400 ;
        RECT 1136.3400 2532.2000 1139.3400 2532.6800 ;
        RECT 1136.3400 2537.6400 1139.3400 2538.1200 ;
        RECT 1136.3400 2521.3200 1139.3400 2521.8000 ;
        RECT 1136.3400 2510.4400 1139.3400 2510.9200 ;
        RECT 1136.3400 2515.8800 1139.3400 2516.3600 ;
        RECT 1093.1000 2526.7600 1094.1000 2527.2400 ;
        RECT 1093.1000 2532.2000 1094.1000 2532.6800 ;
        RECT 1093.1000 2537.6400 1094.1000 2538.1200 ;
        RECT 1093.1000 2510.4400 1094.1000 2510.9200 ;
        RECT 1093.1000 2515.8800 1094.1000 2516.3600 ;
        RECT 1093.1000 2521.3200 1094.1000 2521.8000 ;
        RECT 1136.3400 2499.5600 1139.3400 2500.0400 ;
        RECT 1136.3400 2505.0000 1139.3400 2505.4800 ;
        RECT 1136.3400 2488.6800 1139.3400 2489.1600 ;
        RECT 1136.3400 2494.1200 1139.3400 2494.6000 ;
        RECT 1136.3400 2483.2400 1139.3400 2483.7200 ;
        RECT 1093.1000 2499.5600 1094.1000 2500.0400 ;
        RECT 1093.1000 2505.0000 1094.1000 2505.4800 ;
        RECT 1093.1000 2483.2400 1094.1000 2483.7200 ;
        RECT 1093.1000 2488.6800 1094.1000 2489.1600 ;
        RECT 1093.1000 2494.1200 1094.1000 2494.6000 ;
        RECT 1048.1000 2526.7600 1049.1000 2527.2400 ;
        RECT 1048.1000 2532.2000 1049.1000 2532.6800 ;
        RECT 1048.1000 2537.6400 1049.1000 2538.1200 ;
        RECT 1048.1000 2510.4400 1049.1000 2510.9200 ;
        RECT 1048.1000 2515.8800 1049.1000 2516.3600 ;
        RECT 1048.1000 2521.3200 1049.1000 2521.8000 ;
        RECT 1048.1000 2499.5600 1049.1000 2500.0400 ;
        RECT 1048.1000 2505.0000 1049.1000 2505.4800 ;
        RECT 1048.1000 2483.2400 1049.1000 2483.7200 ;
        RECT 1048.1000 2488.6800 1049.1000 2489.1600 ;
        RECT 1048.1000 2494.1200 1049.1000 2494.6000 ;
        RECT 1003.1000 2570.2800 1004.1000 2570.7600 ;
        RECT 1003.1000 2575.7200 1004.1000 2576.2000 ;
        RECT 1003.1000 2559.4000 1004.1000 2559.8800 ;
        RECT 1003.1000 2564.8400 1004.1000 2565.3200 ;
        RECT 1003.1000 2543.0800 1004.1000 2543.5600 ;
        RECT 1003.1000 2548.5200 1004.1000 2549.0000 ;
        RECT 1003.1000 2553.9600 1004.1000 2554.4400 ;
        RECT 958.1000 2570.2800 959.1000 2570.7600 ;
        RECT 958.1000 2575.7200 959.1000 2576.2000 ;
        RECT 913.1000 2575.7200 914.1000 2576.2000 ;
        RECT 913.1000 2570.2800 914.1000 2570.7600 ;
        RECT 902.3400 2575.7200 905.3400 2576.2000 ;
        RECT 902.3400 2570.2800 905.3400 2570.7600 ;
        RECT 958.1000 2559.4000 959.1000 2559.8800 ;
        RECT 958.1000 2564.8400 959.1000 2565.3200 ;
        RECT 958.1000 2543.0800 959.1000 2543.5600 ;
        RECT 958.1000 2548.5200 959.1000 2549.0000 ;
        RECT 958.1000 2553.9600 959.1000 2554.4400 ;
        RECT 902.3400 2564.8400 905.3400 2565.3200 ;
        RECT 913.1000 2564.8400 914.1000 2565.3200 ;
        RECT 902.3400 2559.4000 905.3400 2559.8800 ;
        RECT 913.1000 2559.4000 914.1000 2559.8800 ;
        RECT 913.1000 2553.9600 914.1000 2554.4400 ;
        RECT 913.1000 2548.5200 914.1000 2549.0000 ;
        RECT 902.3400 2553.9600 905.3400 2554.4400 ;
        RECT 902.3400 2548.5200 905.3400 2549.0000 ;
        RECT 902.3400 2543.0800 905.3400 2543.5600 ;
        RECT 913.1000 2543.0800 914.1000 2543.5600 ;
        RECT 1003.1000 2526.7600 1004.1000 2527.2400 ;
        RECT 1003.1000 2532.2000 1004.1000 2532.6800 ;
        RECT 1003.1000 2537.6400 1004.1000 2538.1200 ;
        RECT 1003.1000 2510.4400 1004.1000 2510.9200 ;
        RECT 1003.1000 2515.8800 1004.1000 2516.3600 ;
        RECT 1003.1000 2521.3200 1004.1000 2521.8000 ;
        RECT 1003.1000 2499.5600 1004.1000 2500.0400 ;
        RECT 1003.1000 2505.0000 1004.1000 2505.4800 ;
        RECT 1003.1000 2483.2400 1004.1000 2483.7200 ;
        RECT 1003.1000 2488.6800 1004.1000 2489.1600 ;
        RECT 1003.1000 2494.1200 1004.1000 2494.6000 ;
        RECT 958.1000 2526.7600 959.1000 2527.2400 ;
        RECT 958.1000 2532.2000 959.1000 2532.6800 ;
        RECT 958.1000 2537.6400 959.1000 2538.1200 ;
        RECT 958.1000 2510.4400 959.1000 2510.9200 ;
        RECT 958.1000 2515.8800 959.1000 2516.3600 ;
        RECT 958.1000 2521.3200 959.1000 2521.8000 ;
        RECT 902.3400 2537.6400 905.3400 2538.1200 ;
        RECT 913.1000 2537.6400 914.1000 2538.1200 ;
        RECT 902.3400 2526.7600 905.3400 2527.2400 ;
        RECT 913.1000 2526.7600 914.1000 2527.2400 ;
        RECT 902.3400 2532.2000 905.3400 2532.6800 ;
        RECT 913.1000 2532.2000 914.1000 2532.6800 ;
        RECT 902.3400 2521.3200 905.3400 2521.8000 ;
        RECT 913.1000 2521.3200 914.1000 2521.8000 ;
        RECT 913.1000 2515.8800 914.1000 2516.3600 ;
        RECT 913.1000 2510.4400 914.1000 2510.9200 ;
        RECT 902.3400 2515.8800 905.3400 2516.3600 ;
        RECT 902.3400 2510.4400 905.3400 2510.9200 ;
        RECT 958.1000 2499.5600 959.1000 2500.0400 ;
        RECT 958.1000 2505.0000 959.1000 2505.4800 ;
        RECT 958.1000 2483.2400 959.1000 2483.7200 ;
        RECT 958.1000 2488.6800 959.1000 2489.1600 ;
        RECT 958.1000 2494.1200 959.1000 2494.6000 ;
        RECT 902.3400 2505.0000 905.3400 2505.4800 ;
        RECT 913.1000 2505.0000 914.1000 2505.4800 ;
        RECT 902.3400 2499.5600 905.3400 2500.0400 ;
        RECT 913.1000 2499.5600 914.1000 2500.0400 ;
        RECT 913.1000 2494.1200 914.1000 2494.6000 ;
        RECT 913.1000 2488.6800 914.1000 2489.1600 ;
        RECT 902.3400 2494.1200 905.3400 2494.6000 ;
        RECT 902.3400 2488.6800 905.3400 2489.1600 ;
        RECT 902.3400 2483.2400 905.3400 2483.7200 ;
        RECT 913.1000 2483.2400 914.1000 2483.7200 ;
        RECT 1136.3400 2466.9200 1139.3400 2467.4000 ;
        RECT 1136.3400 2472.3600 1139.3400 2472.8400 ;
        RECT 1136.3400 2477.8000 1139.3400 2478.2800 ;
        RECT 1136.3400 2461.4800 1139.3400 2461.9600 ;
        RECT 1136.3400 2450.6000 1139.3400 2451.0800 ;
        RECT 1136.3400 2456.0400 1139.3400 2456.5200 ;
        RECT 1093.1000 2466.9200 1094.1000 2467.4000 ;
        RECT 1093.1000 2472.3600 1094.1000 2472.8400 ;
        RECT 1093.1000 2477.8000 1094.1000 2478.2800 ;
        RECT 1093.1000 2450.6000 1094.1000 2451.0800 ;
        RECT 1093.1000 2456.0400 1094.1000 2456.5200 ;
        RECT 1093.1000 2461.4800 1094.1000 2461.9600 ;
        RECT 1136.3400 2439.7200 1139.3400 2440.2000 ;
        RECT 1136.3400 2445.1600 1139.3400 2445.6400 ;
        RECT 1136.3400 2428.8400 1139.3400 2429.3200 ;
        RECT 1136.3400 2434.2800 1139.3400 2434.7600 ;
        RECT 1136.3400 2423.4000 1139.3400 2423.8800 ;
        RECT 1093.1000 2439.7200 1094.1000 2440.2000 ;
        RECT 1093.1000 2445.1600 1094.1000 2445.6400 ;
        RECT 1093.1000 2423.4000 1094.1000 2423.8800 ;
        RECT 1093.1000 2428.8400 1094.1000 2429.3200 ;
        RECT 1093.1000 2434.2800 1094.1000 2434.7600 ;
        RECT 1048.1000 2466.9200 1049.1000 2467.4000 ;
        RECT 1048.1000 2472.3600 1049.1000 2472.8400 ;
        RECT 1048.1000 2477.8000 1049.1000 2478.2800 ;
        RECT 1048.1000 2450.6000 1049.1000 2451.0800 ;
        RECT 1048.1000 2456.0400 1049.1000 2456.5200 ;
        RECT 1048.1000 2461.4800 1049.1000 2461.9600 ;
        RECT 1048.1000 2439.7200 1049.1000 2440.2000 ;
        RECT 1048.1000 2445.1600 1049.1000 2445.6400 ;
        RECT 1048.1000 2423.4000 1049.1000 2423.8800 ;
        RECT 1048.1000 2428.8400 1049.1000 2429.3200 ;
        RECT 1048.1000 2434.2800 1049.1000 2434.7600 ;
        RECT 1136.3400 2407.0800 1139.3400 2407.5600 ;
        RECT 1136.3400 2412.5200 1139.3400 2413.0000 ;
        RECT 1136.3400 2417.9600 1139.3400 2418.4400 ;
        RECT 1136.3400 2401.6400 1139.3400 2402.1200 ;
        RECT 1136.3400 2390.7600 1139.3400 2391.2400 ;
        RECT 1136.3400 2396.2000 1139.3400 2396.6800 ;
        RECT 1093.1000 2407.0800 1094.1000 2407.5600 ;
        RECT 1093.1000 2412.5200 1094.1000 2413.0000 ;
        RECT 1093.1000 2417.9600 1094.1000 2418.4400 ;
        RECT 1093.1000 2390.7600 1094.1000 2391.2400 ;
        RECT 1093.1000 2396.2000 1094.1000 2396.6800 ;
        RECT 1093.1000 2401.6400 1094.1000 2402.1200 ;
        RECT 1136.3400 2379.8800 1139.3400 2380.3600 ;
        RECT 1136.3400 2385.3200 1139.3400 2385.8000 ;
        RECT 1093.1000 2379.8800 1094.1000 2380.3600 ;
        RECT 1093.1000 2385.3200 1094.1000 2385.8000 ;
        RECT 1048.1000 2407.0800 1049.1000 2407.5600 ;
        RECT 1048.1000 2412.5200 1049.1000 2413.0000 ;
        RECT 1048.1000 2417.9600 1049.1000 2418.4400 ;
        RECT 1048.1000 2390.7600 1049.1000 2391.2400 ;
        RECT 1048.1000 2396.2000 1049.1000 2396.6800 ;
        RECT 1048.1000 2401.6400 1049.1000 2402.1200 ;
        RECT 1048.1000 2379.8800 1049.1000 2380.3600 ;
        RECT 1048.1000 2385.3200 1049.1000 2385.8000 ;
        RECT 1003.1000 2466.9200 1004.1000 2467.4000 ;
        RECT 1003.1000 2472.3600 1004.1000 2472.8400 ;
        RECT 1003.1000 2477.8000 1004.1000 2478.2800 ;
        RECT 1003.1000 2450.6000 1004.1000 2451.0800 ;
        RECT 1003.1000 2456.0400 1004.1000 2456.5200 ;
        RECT 1003.1000 2461.4800 1004.1000 2461.9600 ;
        RECT 1003.1000 2439.7200 1004.1000 2440.2000 ;
        RECT 1003.1000 2445.1600 1004.1000 2445.6400 ;
        RECT 1003.1000 2423.4000 1004.1000 2423.8800 ;
        RECT 1003.1000 2428.8400 1004.1000 2429.3200 ;
        RECT 1003.1000 2434.2800 1004.1000 2434.7600 ;
        RECT 958.1000 2466.9200 959.1000 2467.4000 ;
        RECT 958.1000 2472.3600 959.1000 2472.8400 ;
        RECT 958.1000 2477.8000 959.1000 2478.2800 ;
        RECT 958.1000 2450.6000 959.1000 2451.0800 ;
        RECT 958.1000 2456.0400 959.1000 2456.5200 ;
        RECT 958.1000 2461.4800 959.1000 2461.9600 ;
        RECT 902.3400 2477.8000 905.3400 2478.2800 ;
        RECT 913.1000 2477.8000 914.1000 2478.2800 ;
        RECT 902.3400 2466.9200 905.3400 2467.4000 ;
        RECT 913.1000 2466.9200 914.1000 2467.4000 ;
        RECT 902.3400 2472.3600 905.3400 2472.8400 ;
        RECT 913.1000 2472.3600 914.1000 2472.8400 ;
        RECT 902.3400 2461.4800 905.3400 2461.9600 ;
        RECT 913.1000 2461.4800 914.1000 2461.9600 ;
        RECT 913.1000 2456.0400 914.1000 2456.5200 ;
        RECT 913.1000 2450.6000 914.1000 2451.0800 ;
        RECT 902.3400 2456.0400 905.3400 2456.5200 ;
        RECT 902.3400 2450.6000 905.3400 2451.0800 ;
        RECT 958.1000 2439.7200 959.1000 2440.2000 ;
        RECT 958.1000 2445.1600 959.1000 2445.6400 ;
        RECT 958.1000 2423.4000 959.1000 2423.8800 ;
        RECT 958.1000 2428.8400 959.1000 2429.3200 ;
        RECT 958.1000 2434.2800 959.1000 2434.7600 ;
        RECT 902.3400 2445.1600 905.3400 2445.6400 ;
        RECT 913.1000 2445.1600 914.1000 2445.6400 ;
        RECT 902.3400 2439.7200 905.3400 2440.2000 ;
        RECT 913.1000 2439.7200 914.1000 2440.2000 ;
        RECT 913.1000 2434.2800 914.1000 2434.7600 ;
        RECT 913.1000 2428.8400 914.1000 2429.3200 ;
        RECT 902.3400 2434.2800 905.3400 2434.7600 ;
        RECT 902.3400 2428.8400 905.3400 2429.3200 ;
        RECT 902.3400 2423.4000 905.3400 2423.8800 ;
        RECT 913.1000 2423.4000 914.1000 2423.8800 ;
        RECT 1003.1000 2407.0800 1004.1000 2407.5600 ;
        RECT 1003.1000 2412.5200 1004.1000 2413.0000 ;
        RECT 1003.1000 2417.9600 1004.1000 2418.4400 ;
        RECT 1003.1000 2390.7600 1004.1000 2391.2400 ;
        RECT 1003.1000 2396.2000 1004.1000 2396.6800 ;
        RECT 1003.1000 2401.6400 1004.1000 2402.1200 ;
        RECT 1003.1000 2379.8800 1004.1000 2380.3600 ;
        RECT 1003.1000 2385.3200 1004.1000 2385.8000 ;
        RECT 958.1000 2407.0800 959.1000 2407.5600 ;
        RECT 958.1000 2412.5200 959.1000 2413.0000 ;
        RECT 958.1000 2417.9600 959.1000 2418.4400 ;
        RECT 958.1000 2390.7600 959.1000 2391.2400 ;
        RECT 958.1000 2396.2000 959.1000 2396.6800 ;
        RECT 958.1000 2401.6400 959.1000 2402.1200 ;
        RECT 902.3400 2417.9600 905.3400 2418.4400 ;
        RECT 913.1000 2417.9600 914.1000 2418.4400 ;
        RECT 902.3400 2407.0800 905.3400 2407.5600 ;
        RECT 913.1000 2407.0800 914.1000 2407.5600 ;
        RECT 902.3400 2412.5200 905.3400 2413.0000 ;
        RECT 913.1000 2412.5200 914.1000 2413.0000 ;
        RECT 902.3400 2401.6400 905.3400 2402.1200 ;
        RECT 913.1000 2401.6400 914.1000 2402.1200 ;
        RECT 913.1000 2396.2000 914.1000 2396.6800 ;
        RECT 913.1000 2390.7600 914.1000 2391.2400 ;
        RECT 902.3400 2396.2000 905.3400 2396.6800 ;
        RECT 902.3400 2390.7600 905.3400 2391.2400 ;
        RECT 958.1000 2379.8800 959.1000 2380.3600 ;
        RECT 958.1000 2385.3200 959.1000 2385.8000 ;
        RECT 902.3400 2385.3200 905.3400 2385.8000 ;
        RECT 913.1000 2385.3200 914.1000 2385.8000 ;
        RECT 902.3400 2379.8800 905.3400 2380.3600 ;
        RECT 913.1000 2379.8800 914.1000 2380.3600 ;
        RECT 902.3400 2584.7900 1139.3400 2587.7900 ;
        RECT 902.3400 2371.6900 1139.3400 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 2142.0500 1094.1000 2358.1500 ;
        RECT 1048.1000 2142.0500 1049.1000 2358.1500 ;
        RECT 1003.1000 2142.0500 1004.1000 2358.1500 ;
        RECT 958.1000 2142.0500 959.1000 2358.1500 ;
        RECT 913.1000 2142.0500 914.1000 2358.1500 ;
        RECT 1136.3400 2142.0500 1139.3400 2358.1500 ;
        RECT 902.3400 2142.0500 905.3400 2358.1500 ;
      LAYER met3 ;
        RECT 1136.3400 2340.6400 1139.3400 2341.1200 ;
        RECT 1136.3400 2346.0800 1139.3400 2346.5600 ;
        RECT 1093.1000 2340.6400 1094.1000 2341.1200 ;
        RECT 1093.1000 2346.0800 1094.1000 2346.5600 ;
        RECT 1136.3400 2329.7600 1139.3400 2330.2400 ;
        RECT 1136.3400 2335.2000 1139.3400 2335.6800 ;
        RECT 1136.3400 2318.8800 1139.3400 2319.3600 ;
        RECT 1136.3400 2324.3200 1139.3400 2324.8000 ;
        RECT 1136.3400 2313.4400 1139.3400 2313.9200 ;
        RECT 1093.1000 2329.7600 1094.1000 2330.2400 ;
        RECT 1093.1000 2335.2000 1094.1000 2335.6800 ;
        RECT 1093.1000 2313.4400 1094.1000 2313.9200 ;
        RECT 1093.1000 2318.8800 1094.1000 2319.3600 ;
        RECT 1093.1000 2324.3200 1094.1000 2324.8000 ;
        RECT 1048.1000 2340.6400 1049.1000 2341.1200 ;
        RECT 1048.1000 2346.0800 1049.1000 2346.5600 ;
        RECT 1048.1000 2329.7600 1049.1000 2330.2400 ;
        RECT 1048.1000 2335.2000 1049.1000 2335.6800 ;
        RECT 1048.1000 2313.4400 1049.1000 2313.9200 ;
        RECT 1048.1000 2318.8800 1049.1000 2319.3600 ;
        RECT 1048.1000 2324.3200 1049.1000 2324.8000 ;
        RECT 1136.3400 2297.1200 1139.3400 2297.6000 ;
        RECT 1136.3400 2302.5600 1139.3400 2303.0400 ;
        RECT 1136.3400 2308.0000 1139.3400 2308.4800 ;
        RECT 1136.3400 2291.6800 1139.3400 2292.1600 ;
        RECT 1136.3400 2280.8000 1139.3400 2281.2800 ;
        RECT 1136.3400 2286.2400 1139.3400 2286.7200 ;
        RECT 1093.1000 2297.1200 1094.1000 2297.6000 ;
        RECT 1093.1000 2302.5600 1094.1000 2303.0400 ;
        RECT 1093.1000 2308.0000 1094.1000 2308.4800 ;
        RECT 1093.1000 2280.8000 1094.1000 2281.2800 ;
        RECT 1093.1000 2286.2400 1094.1000 2286.7200 ;
        RECT 1093.1000 2291.6800 1094.1000 2292.1600 ;
        RECT 1136.3400 2269.9200 1139.3400 2270.4000 ;
        RECT 1136.3400 2275.3600 1139.3400 2275.8400 ;
        RECT 1136.3400 2259.0400 1139.3400 2259.5200 ;
        RECT 1136.3400 2264.4800 1139.3400 2264.9600 ;
        RECT 1136.3400 2253.6000 1139.3400 2254.0800 ;
        RECT 1093.1000 2269.9200 1094.1000 2270.4000 ;
        RECT 1093.1000 2275.3600 1094.1000 2275.8400 ;
        RECT 1093.1000 2253.6000 1094.1000 2254.0800 ;
        RECT 1093.1000 2259.0400 1094.1000 2259.5200 ;
        RECT 1093.1000 2264.4800 1094.1000 2264.9600 ;
        RECT 1048.1000 2297.1200 1049.1000 2297.6000 ;
        RECT 1048.1000 2302.5600 1049.1000 2303.0400 ;
        RECT 1048.1000 2308.0000 1049.1000 2308.4800 ;
        RECT 1048.1000 2280.8000 1049.1000 2281.2800 ;
        RECT 1048.1000 2286.2400 1049.1000 2286.7200 ;
        RECT 1048.1000 2291.6800 1049.1000 2292.1600 ;
        RECT 1048.1000 2269.9200 1049.1000 2270.4000 ;
        RECT 1048.1000 2275.3600 1049.1000 2275.8400 ;
        RECT 1048.1000 2253.6000 1049.1000 2254.0800 ;
        RECT 1048.1000 2259.0400 1049.1000 2259.5200 ;
        RECT 1048.1000 2264.4800 1049.1000 2264.9600 ;
        RECT 1003.1000 2340.6400 1004.1000 2341.1200 ;
        RECT 1003.1000 2346.0800 1004.1000 2346.5600 ;
        RECT 1003.1000 2329.7600 1004.1000 2330.2400 ;
        RECT 1003.1000 2335.2000 1004.1000 2335.6800 ;
        RECT 1003.1000 2313.4400 1004.1000 2313.9200 ;
        RECT 1003.1000 2318.8800 1004.1000 2319.3600 ;
        RECT 1003.1000 2324.3200 1004.1000 2324.8000 ;
        RECT 958.1000 2340.6400 959.1000 2341.1200 ;
        RECT 958.1000 2346.0800 959.1000 2346.5600 ;
        RECT 913.1000 2346.0800 914.1000 2346.5600 ;
        RECT 913.1000 2340.6400 914.1000 2341.1200 ;
        RECT 902.3400 2346.0800 905.3400 2346.5600 ;
        RECT 902.3400 2340.6400 905.3400 2341.1200 ;
        RECT 958.1000 2329.7600 959.1000 2330.2400 ;
        RECT 958.1000 2335.2000 959.1000 2335.6800 ;
        RECT 958.1000 2313.4400 959.1000 2313.9200 ;
        RECT 958.1000 2318.8800 959.1000 2319.3600 ;
        RECT 958.1000 2324.3200 959.1000 2324.8000 ;
        RECT 902.3400 2335.2000 905.3400 2335.6800 ;
        RECT 913.1000 2335.2000 914.1000 2335.6800 ;
        RECT 902.3400 2329.7600 905.3400 2330.2400 ;
        RECT 913.1000 2329.7600 914.1000 2330.2400 ;
        RECT 913.1000 2324.3200 914.1000 2324.8000 ;
        RECT 913.1000 2318.8800 914.1000 2319.3600 ;
        RECT 902.3400 2324.3200 905.3400 2324.8000 ;
        RECT 902.3400 2318.8800 905.3400 2319.3600 ;
        RECT 902.3400 2313.4400 905.3400 2313.9200 ;
        RECT 913.1000 2313.4400 914.1000 2313.9200 ;
        RECT 1003.1000 2297.1200 1004.1000 2297.6000 ;
        RECT 1003.1000 2302.5600 1004.1000 2303.0400 ;
        RECT 1003.1000 2308.0000 1004.1000 2308.4800 ;
        RECT 1003.1000 2280.8000 1004.1000 2281.2800 ;
        RECT 1003.1000 2286.2400 1004.1000 2286.7200 ;
        RECT 1003.1000 2291.6800 1004.1000 2292.1600 ;
        RECT 1003.1000 2269.9200 1004.1000 2270.4000 ;
        RECT 1003.1000 2275.3600 1004.1000 2275.8400 ;
        RECT 1003.1000 2253.6000 1004.1000 2254.0800 ;
        RECT 1003.1000 2259.0400 1004.1000 2259.5200 ;
        RECT 1003.1000 2264.4800 1004.1000 2264.9600 ;
        RECT 958.1000 2297.1200 959.1000 2297.6000 ;
        RECT 958.1000 2302.5600 959.1000 2303.0400 ;
        RECT 958.1000 2308.0000 959.1000 2308.4800 ;
        RECT 958.1000 2280.8000 959.1000 2281.2800 ;
        RECT 958.1000 2286.2400 959.1000 2286.7200 ;
        RECT 958.1000 2291.6800 959.1000 2292.1600 ;
        RECT 902.3400 2308.0000 905.3400 2308.4800 ;
        RECT 913.1000 2308.0000 914.1000 2308.4800 ;
        RECT 902.3400 2297.1200 905.3400 2297.6000 ;
        RECT 913.1000 2297.1200 914.1000 2297.6000 ;
        RECT 902.3400 2302.5600 905.3400 2303.0400 ;
        RECT 913.1000 2302.5600 914.1000 2303.0400 ;
        RECT 902.3400 2291.6800 905.3400 2292.1600 ;
        RECT 913.1000 2291.6800 914.1000 2292.1600 ;
        RECT 913.1000 2286.2400 914.1000 2286.7200 ;
        RECT 913.1000 2280.8000 914.1000 2281.2800 ;
        RECT 902.3400 2286.2400 905.3400 2286.7200 ;
        RECT 902.3400 2280.8000 905.3400 2281.2800 ;
        RECT 958.1000 2269.9200 959.1000 2270.4000 ;
        RECT 958.1000 2275.3600 959.1000 2275.8400 ;
        RECT 958.1000 2253.6000 959.1000 2254.0800 ;
        RECT 958.1000 2259.0400 959.1000 2259.5200 ;
        RECT 958.1000 2264.4800 959.1000 2264.9600 ;
        RECT 902.3400 2275.3600 905.3400 2275.8400 ;
        RECT 913.1000 2275.3600 914.1000 2275.8400 ;
        RECT 902.3400 2269.9200 905.3400 2270.4000 ;
        RECT 913.1000 2269.9200 914.1000 2270.4000 ;
        RECT 913.1000 2264.4800 914.1000 2264.9600 ;
        RECT 913.1000 2259.0400 914.1000 2259.5200 ;
        RECT 902.3400 2264.4800 905.3400 2264.9600 ;
        RECT 902.3400 2259.0400 905.3400 2259.5200 ;
        RECT 902.3400 2253.6000 905.3400 2254.0800 ;
        RECT 913.1000 2253.6000 914.1000 2254.0800 ;
        RECT 1136.3400 2237.2800 1139.3400 2237.7600 ;
        RECT 1136.3400 2242.7200 1139.3400 2243.2000 ;
        RECT 1136.3400 2248.1600 1139.3400 2248.6400 ;
        RECT 1136.3400 2231.8400 1139.3400 2232.3200 ;
        RECT 1136.3400 2220.9600 1139.3400 2221.4400 ;
        RECT 1136.3400 2226.4000 1139.3400 2226.8800 ;
        RECT 1093.1000 2237.2800 1094.1000 2237.7600 ;
        RECT 1093.1000 2242.7200 1094.1000 2243.2000 ;
        RECT 1093.1000 2248.1600 1094.1000 2248.6400 ;
        RECT 1093.1000 2220.9600 1094.1000 2221.4400 ;
        RECT 1093.1000 2226.4000 1094.1000 2226.8800 ;
        RECT 1093.1000 2231.8400 1094.1000 2232.3200 ;
        RECT 1136.3400 2210.0800 1139.3400 2210.5600 ;
        RECT 1136.3400 2215.5200 1139.3400 2216.0000 ;
        RECT 1136.3400 2199.2000 1139.3400 2199.6800 ;
        RECT 1136.3400 2204.6400 1139.3400 2205.1200 ;
        RECT 1136.3400 2193.7600 1139.3400 2194.2400 ;
        RECT 1093.1000 2210.0800 1094.1000 2210.5600 ;
        RECT 1093.1000 2215.5200 1094.1000 2216.0000 ;
        RECT 1093.1000 2193.7600 1094.1000 2194.2400 ;
        RECT 1093.1000 2199.2000 1094.1000 2199.6800 ;
        RECT 1093.1000 2204.6400 1094.1000 2205.1200 ;
        RECT 1048.1000 2237.2800 1049.1000 2237.7600 ;
        RECT 1048.1000 2242.7200 1049.1000 2243.2000 ;
        RECT 1048.1000 2248.1600 1049.1000 2248.6400 ;
        RECT 1048.1000 2220.9600 1049.1000 2221.4400 ;
        RECT 1048.1000 2226.4000 1049.1000 2226.8800 ;
        RECT 1048.1000 2231.8400 1049.1000 2232.3200 ;
        RECT 1048.1000 2210.0800 1049.1000 2210.5600 ;
        RECT 1048.1000 2215.5200 1049.1000 2216.0000 ;
        RECT 1048.1000 2193.7600 1049.1000 2194.2400 ;
        RECT 1048.1000 2199.2000 1049.1000 2199.6800 ;
        RECT 1048.1000 2204.6400 1049.1000 2205.1200 ;
        RECT 1136.3400 2177.4400 1139.3400 2177.9200 ;
        RECT 1136.3400 2182.8800 1139.3400 2183.3600 ;
        RECT 1136.3400 2188.3200 1139.3400 2188.8000 ;
        RECT 1136.3400 2172.0000 1139.3400 2172.4800 ;
        RECT 1136.3400 2161.1200 1139.3400 2161.6000 ;
        RECT 1136.3400 2166.5600 1139.3400 2167.0400 ;
        RECT 1093.1000 2177.4400 1094.1000 2177.9200 ;
        RECT 1093.1000 2182.8800 1094.1000 2183.3600 ;
        RECT 1093.1000 2188.3200 1094.1000 2188.8000 ;
        RECT 1093.1000 2161.1200 1094.1000 2161.6000 ;
        RECT 1093.1000 2166.5600 1094.1000 2167.0400 ;
        RECT 1093.1000 2172.0000 1094.1000 2172.4800 ;
        RECT 1136.3400 2150.2400 1139.3400 2150.7200 ;
        RECT 1136.3400 2155.6800 1139.3400 2156.1600 ;
        RECT 1093.1000 2150.2400 1094.1000 2150.7200 ;
        RECT 1093.1000 2155.6800 1094.1000 2156.1600 ;
        RECT 1048.1000 2177.4400 1049.1000 2177.9200 ;
        RECT 1048.1000 2182.8800 1049.1000 2183.3600 ;
        RECT 1048.1000 2188.3200 1049.1000 2188.8000 ;
        RECT 1048.1000 2161.1200 1049.1000 2161.6000 ;
        RECT 1048.1000 2166.5600 1049.1000 2167.0400 ;
        RECT 1048.1000 2172.0000 1049.1000 2172.4800 ;
        RECT 1048.1000 2150.2400 1049.1000 2150.7200 ;
        RECT 1048.1000 2155.6800 1049.1000 2156.1600 ;
        RECT 1003.1000 2237.2800 1004.1000 2237.7600 ;
        RECT 1003.1000 2242.7200 1004.1000 2243.2000 ;
        RECT 1003.1000 2248.1600 1004.1000 2248.6400 ;
        RECT 1003.1000 2220.9600 1004.1000 2221.4400 ;
        RECT 1003.1000 2226.4000 1004.1000 2226.8800 ;
        RECT 1003.1000 2231.8400 1004.1000 2232.3200 ;
        RECT 1003.1000 2210.0800 1004.1000 2210.5600 ;
        RECT 1003.1000 2215.5200 1004.1000 2216.0000 ;
        RECT 1003.1000 2193.7600 1004.1000 2194.2400 ;
        RECT 1003.1000 2199.2000 1004.1000 2199.6800 ;
        RECT 1003.1000 2204.6400 1004.1000 2205.1200 ;
        RECT 958.1000 2237.2800 959.1000 2237.7600 ;
        RECT 958.1000 2242.7200 959.1000 2243.2000 ;
        RECT 958.1000 2248.1600 959.1000 2248.6400 ;
        RECT 958.1000 2220.9600 959.1000 2221.4400 ;
        RECT 958.1000 2226.4000 959.1000 2226.8800 ;
        RECT 958.1000 2231.8400 959.1000 2232.3200 ;
        RECT 902.3400 2248.1600 905.3400 2248.6400 ;
        RECT 913.1000 2248.1600 914.1000 2248.6400 ;
        RECT 902.3400 2237.2800 905.3400 2237.7600 ;
        RECT 913.1000 2237.2800 914.1000 2237.7600 ;
        RECT 902.3400 2242.7200 905.3400 2243.2000 ;
        RECT 913.1000 2242.7200 914.1000 2243.2000 ;
        RECT 902.3400 2231.8400 905.3400 2232.3200 ;
        RECT 913.1000 2231.8400 914.1000 2232.3200 ;
        RECT 913.1000 2226.4000 914.1000 2226.8800 ;
        RECT 913.1000 2220.9600 914.1000 2221.4400 ;
        RECT 902.3400 2226.4000 905.3400 2226.8800 ;
        RECT 902.3400 2220.9600 905.3400 2221.4400 ;
        RECT 958.1000 2210.0800 959.1000 2210.5600 ;
        RECT 958.1000 2215.5200 959.1000 2216.0000 ;
        RECT 958.1000 2193.7600 959.1000 2194.2400 ;
        RECT 958.1000 2199.2000 959.1000 2199.6800 ;
        RECT 958.1000 2204.6400 959.1000 2205.1200 ;
        RECT 902.3400 2215.5200 905.3400 2216.0000 ;
        RECT 913.1000 2215.5200 914.1000 2216.0000 ;
        RECT 902.3400 2210.0800 905.3400 2210.5600 ;
        RECT 913.1000 2210.0800 914.1000 2210.5600 ;
        RECT 913.1000 2204.6400 914.1000 2205.1200 ;
        RECT 913.1000 2199.2000 914.1000 2199.6800 ;
        RECT 902.3400 2204.6400 905.3400 2205.1200 ;
        RECT 902.3400 2199.2000 905.3400 2199.6800 ;
        RECT 902.3400 2193.7600 905.3400 2194.2400 ;
        RECT 913.1000 2193.7600 914.1000 2194.2400 ;
        RECT 1003.1000 2177.4400 1004.1000 2177.9200 ;
        RECT 1003.1000 2182.8800 1004.1000 2183.3600 ;
        RECT 1003.1000 2188.3200 1004.1000 2188.8000 ;
        RECT 1003.1000 2161.1200 1004.1000 2161.6000 ;
        RECT 1003.1000 2166.5600 1004.1000 2167.0400 ;
        RECT 1003.1000 2172.0000 1004.1000 2172.4800 ;
        RECT 1003.1000 2150.2400 1004.1000 2150.7200 ;
        RECT 1003.1000 2155.6800 1004.1000 2156.1600 ;
        RECT 958.1000 2177.4400 959.1000 2177.9200 ;
        RECT 958.1000 2182.8800 959.1000 2183.3600 ;
        RECT 958.1000 2188.3200 959.1000 2188.8000 ;
        RECT 958.1000 2161.1200 959.1000 2161.6000 ;
        RECT 958.1000 2166.5600 959.1000 2167.0400 ;
        RECT 958.1000 2172.0000 959.1000 2172.4800 ;
        RECT 902.3400 2188.3200 905.3400 2188.8000 ;
        RECT 913.1000 2188.3200 914.1000 2188.8000 ;
        RECT 902.3400 2177.4400 905.3400 2177.9200 ;
        RECT 913.1000 2177.4400 914.1000 2177.9200 ;
        RECT 902.3400 2182.8800 905.3400 2183.3600 ;
        RECT 913.1000 2182.8800 914.1000 2183.3600 ;
        RECT 902.3400 2172.0000 905.3400 2172.4800 ;
        RECT 913.1000 2172.0000 914.1000 2172.4800 ;
        RECT 913.1000 2166.5600 914.1000 2167.0400 ;
        RECT 913.1000 2161.1200 914.1000 2161.6000 ;
        RECT 902.3400 2166.5600 905.3400 2167.0400 ;
        RECT 902.3400 2161.1200 905.3400 2161.6000 ;
        RECT 958.1000 2150.2400 959.1000 2150.7200 ;
        RECT 958.1000 2155.6800 959.1000 2156.1600 ;
        RECT 902.3400 2155.6800 905.3400 2156.1600 ;
        RECT 913.1000 2155.6800 914.1000 2156.1600 ;
        RECT 902.3400 2150.2400 905.3400 2150.7200 ;
        RECT 913.1000 2150.2400 914.1000 2150.7200 ;
        RECT 902.3400 2355.1500 1139.3400 2358.1500 ;
        RECT 902.3400 2142.0500 1139.3400 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 1912.4100 1094.1000 2128.5100 ;
        RECT 1048.1000 1912.4100 1049.1000 2128.5100 ;
        RECT 1003.1000 1912.4100 1004.1000 2128.5100 ;
        RECT 958.1000 1912.4100 959.1000 2128.5100 ;
        RECT 913.1000 1912.4100 914.1000 2128.5100 ;
        RECT 1136.3400 1912.4100 1139.3400 2128.5100 ;
        RECT 902.3400 1912.4100 905.3400 2128.5100 ;
      LAYER met3 ;
        RECT 1136.3400 2111.0000 1139.3400 2111.4800 ;
        RECT 1136.3400 2116.4400 1139.3400 2116.9200 ;
        RECT 1093.1000 2111.0000 1094.1000 2111.4800 ;
        RECT 1093.1000 2116.4400 1094.1000 2116.9200 ;
        RECT 1136.3400 2100.1200 1139.3400 2100.6000 ;
        RECT 1136.3400 2105.5600 1139.3400 2106.0400 ;
        RECT 1136.3400 2089.2400 1139.3400 2089.7200 ;
        RECT 1136.3400 2094.6800 1139.3400 2095.1600 ;
        RECT 1136.3400 2083.8000 1139.3400 2084.2800 ;
        RECT 1093.1000 2100.1200 1094.1000 2100.6000 ;
        RECT 1093.1000 2105.5600 1094.1000 2106.0400 ;
        RECT 1093.1000 2083.8000 1094.1000 2084.2800 ;
        RECT 1093.1000 2089.2400 1094.1000 2089.7200 ;
        RECT 1093.1000 2094.6800 1094.1000 2095.1600 ;
        RECT 1048.1000 2111.0000 1049.1000 2111.4800 ;
        RECT 1048.1000 2116.4400 1049.1000 2116.9200 ;
        RECT 1048.1000 2100.1200 1049.1000 2100.6000 ;
        RECT 1048.1000 2105.5600 1049.1000 2106.0400 ;
        RECT 1048.1000 2083.8000 1049.1000 2084.2800 ;
        RECT 1048.1000 2089.2400 1049.1000 2089.7200 ;
        RECT 1048.1000 2094.6800 1049.1000 2095.1600 ;
        RECT 1136.3400 2067.4800 1139.3400 2067.9600 ;
        RECT 1136.3400 2072.9200 1139.3400 2073.4000 ;
        RECT 1136.3400 2078.3600 1139.3400 2078.8400 ;
        RECT 1136.3400 2062.0400 1139.3400 2062.5200 ;
        RECT 1136.3400 2051.1600 1139.3400 2051.6400 ;
        RECT 1136.3400 2056.6000 1139.3400 2057.0800 ;
        RECT 1093.1000 2067.4800 1094.1000 2067.9600 ;
        RECT 1093.1000 2072.9200 1094.1000 2073.4000 ;
        RECT 1093.1000 2078.3600 1094.1000 2078.8400 ;
        RECT 1093.1000 2051.1600 1094.1000 2051.6400 ;
        RECT 1093.1000 2056.6000 1094.1000 2057.0800 ;
        RECT 1093.1000 2062.0400 1094.1000 2062.5200 ;
        RECT 1136.3400 2040.2800 1139.3400 2040.7600 ;
        RECT 1136.3400 2045.7200 1139.3400 2046.2000 ;
        RECT 1136.3400 2029.4000 1139.3400 2029.8800 ;
        RECT 1136.3400 2034.8400 1139.3400 2035.3200 ;
        RECT 1136.3400 2023.9600 1139.3400 2024.4400 ;
        RECT 1093.1000 2040.2800 1094.1000 2040.7600 ;
        RECT 1093.1000 2045.7200 1094.1000 2046.2000 ;
        RECT 1093.1000 2023.9600 1094.1000 2024.4400 ;
        RECT 1093.1000 2029.4000 1094.1000 2029.8800 ;
        RECT 1093.1000 2034.8400 1094.1000 2035.3200 ;
        RECT 1048.1000 2067.4800 1049.1000 2067.9600 ;
        RECT 1048.1000 2072.9200 1049.1000 2073.4000 ;
        RECT 1048.1000 2078.3600 1049.1000 2078.8400 ;
        RECT 1048.1000 2051.1600 1049.1000 2051.6400 ;
        RECT 1048.1000 2056.6000 1049.1000 2057.0800 ;
        RECT 1048.1000 2062.0400 1049.1000 2062.5200 ;
        RECT 1048.1000 2040.2800 1049.1000 2040.7600 ;
        RECT 1048.1000 2045.7200 1049.1000 2046.2000 ;
        RECT 1048.1000 2023.9600 1049.1000 2024.4400 ;
        RECT 1048.1000 2029.4000 1049.1000 2029.8800 ;
        RECT 1048.1000 2034.8400 1049.1000 2035.3200 ;
        RECT 1003.1000 2111.0000 1004.1000 2111.4800 ;
        RECT 1003.1000 2116.4400 1004.1000 2116.9200 ;
        RECT 1003.1000 2100.1200 1004.1000 2100.6000 ;
        RECT 1003.1000 2105.5600 1004.1000 2106.0400 ;
        RECT 1003.1000 2083.8000 1004.1000 2084.2800 ;
        RECT 1003.1000 2089.2400 1004.1000 2089.7200 ;
        RECT 1003.1000 2094.6800 1004.1000 2095.1600 ;
        RECT 958.1000 2111.0000 959.1000 2111.4800 ;
        RECT 958.1000 2116.4400 959.1000 2116.9200 ;
        RECT 913.1000 2116.4400 914.1000 2116.9200 ;
        RECT 913.1000 2111.0000 914.1000 2111.4800 ;
        RECT 902.3400 2116.4400 905.3400 2116.9200 ;
        RECT 902.3400 2111.0000 905.3400 2111.4800 ;
        RECT 958.1000 2100.1200 959.1000 2100.6000 ;
        RECT 958.1000 2105.5600 959.1000 2106.0400 ;
        RECT 958.1000 2083.8000 959.1000 2084.2800 ;
        RECT 958.1000 2089.2400 959.1000 2089.7200 ;
        RECT 958.1000 2094.6800 959.1000 2095.1600 ;
        RECT 902.3400 2105.5600 905.3400 2106.0400 ;
        RECT 913.1000 2105.5600 914.1000 2106.0400 ;
        RECT 902.3400 2100.1200 905.3400 2100.6000 ;
        RECT 913.1000 2100.1200 914.1000 2100.6000 ;
        RECT 913.1000 2094.6800 914.1000 2095.1600 ;
        RECT 913.1000 2089.2400 914.1000 2089.7200 ;
        RECT 902.3400 2094.6800 905.3400 2095.1600 ;
        RECT 902.3400 2089.2400 905.3400 2089.7200 ;
        RECT 902.3400 2083.8000 905.3400 2084.2800 ;
        RECT 913.1000 2083.8000 914.1000 2084.2800 ;
        RECT 1003.1000 2067.4800 1004.1000 2067.9600 ;
        RECT 1003.1000 2072.9200 1004.1000 2073.4000 ;
        RECT 1003.1000 2078.3600 1004.1000 2078.8400 ;
        RECT 1003.1000 2051.1600 1004.1000 2051.6400 ;
        RECT 1003.1000 2056.6000 1004.1000 2057.0800 ;
        RECT 1003.1000 2062.0400 1004.1000 2062.5200 ;
        RECT 1003.1000 2040.2800 1004.1000 2040.7600 ;
        RECT 1003.1000 2045.7200 1004.1000 2046.2000 ;
        RECT 1003.1000 2023.9600 1004.1000 2024.4400 ;
        RECT 1003.1000 2029.4000 1004.1000 2029.8800 ;
        RECT 1003.1000 2034.8400 1004.1000 2035.3200 ;
        RECT 958.1000 2067.4800 959.1000 2067.9600 ;
        RECT 958.1000 2072.9200 959.1000 2073.4000 ;
        RECT 958.1000 2078.3600 959.1000 2078.8400 ;
        RECT 958.1000 2051.1600 959.1000 2051.6400 ;
        RECT 958.1000 2056.6000 959.1000 2057.0800 ;
        RECT 958.1000 2062.0400 959.1000 2062.5200 ;
        RECT 902.3400 2078.3600 905.3400 2078.8400 ;
        RECT 913.1000 2078.3600 914.1000 2078.8400 ;
        RECT 902.3400 2067.4800 905.3400 2067.9600 ;
        RECT 913.1000 2067.4800 914.1000 2067.9600 ;
        RECT 902.3400 2072.9200 905.3400 2073.4000 ;
        RECT 913.1000 2072.9200 914.1000 2073.4000 ;
        RECT 902.3400 2062.0400 905.3400 2062.5200 ;
        RECT 913.1000 2062.0400 914.1000 2062.5200 ;
        RECT 913.1000 2056.6000 914.1000 2057.0800 ;
        RECT 913.1000 2051.1600 914.1000 2051.6400 ;
        RECT 902.3400 2056.6000 905.3400 2057.0800 ;
        RECT 902.3400 2051.1600 905.3400 2051.6400 ;
        RECT 958.1000 2040.2800 959.1000 2040.7600 ;
        RECT 958.1000 2045.7200 959.1000 2046.2000 ;
        RECT 958.1000 2023.9600 959.1000 2024.4400 ;
        RECT 958.1000 2029.4000 959.1000 2029.8800 ;
        RECT 958.1000 2034.8400 959.1000 2035.3200 ;
        RECT 902.3400 2045.7200 905.3400 2046.2000 ;
        RECT 913.1000 2045.7200 914.1000 2046.2000 ;
        RECT 902.3400 2040.2800 905.3400 2040.7600 ;
        RECT 913.1000 2040.2800 914.1000 2040.7600 ;
        RECT 913.1000 2034.8400 914.1000 2035.3200 ;
        RECT 913.1000 2029.4000 914.1000 2029.8800 ;
        RECT 902.3400 2034.8400 905.3400 2035.3200 ;
        RECT 902.3400 2029.4000 905.3400 2029.8800 ;
        RECT 902.3400 2023.9600 905.3400 2024.4400 ;
        RECT 913.1000 2023.9600 914.1000 2024.4400 ;
        RECT 1136.3400 2007.6400 1139.3400 2008.1200 ;
        RECT 1136.3400 2013.0800 1139.3400 2013.5600 ;
        RECT 1136.3400 2018.5200 1139.3400 2019.0000 ;
        RECT 1136.3400 2002.2000 1139.3400 2002.6800 ;
        RECT 1136.3400 1991.3200 1139.3400 1991.8000 ;
        RECT 1136.3400 1996.7600 1139.3400 1997.2400 ;
        RECT 1093.1000 2007.6400 1094.1000 2008.1200 ;
        RECT 1093.1000 2013.0800 1094.1000 2013.5600 ;
        RECT 1093.1000 2018.5200 1094.1000 2019.0000 ;
        RECT 1093.1000 1991.3200 1094.1000 1991.8000 ;
        RECT 1093.1000 1996.7600 1094.1000 1997.2400 ;
        RECT 1093.1000 2002.2000 1094.1000 2002.6800 ;
        RECT 1136.3400 1980.4400 1139.3400 1980.9200 ;
        RECT 1136.3400 1985.8800 1139.3400 1986.3600 ;
        RECT 1136.3400 1969.5600 1139.3400 1970.0400 ;
        RECT 1136.3400 1975.0000 1139.3400 1975.4800 ;
        RECT 1136.3400 1964.1200 1139.3400 1964.6000 ;
        RECT 1093.1000 1980.4400 1094.1000 1980.9200 ;
        RECT 1093.1000 1985.8800 1094.1000 1986.3600 ;
        RECT 1093.1000 1964.1200 1094.1000 1964.6000 ;
        RECT 1093.1000 1969.5600 1094.1000 1970.0400 ;
        RECT 1093.1000 1975.0000 1094.1000 1975.4800 ;
        RECT 1048.1000 2007.6400 1049.1000 2008.1200 ;
        RECT 1048.1000 2013.0800 1049.1000 2013.5600 ;
        RECT 1048.1000 2018.5200 1049.1000 2019.0000 ;
        RECT 1048.1000 1991.3200 1049.1000 1991.8000 ;
        RECT 1048.1000 1996.7600 1049.1000 1997.2400 ;
        RECT 1048.1000 2002.2000 1049.1000 2002.6800 ;
        RECT 1048.1000 1980.4400 1049.1000 1980.9200 ;
        RECT 1048.1000 1985.8800 1049.1000 1986.3600 ;
        RECT 1048.1000 1964.1200 1049.1000 1964.6000 ;
        RECT 1048.1000 1969.5600 1049.1000 1970.0400 ;
        RECT 1048.1000 1975.0000 1049.1000 1975.4800 ;
        RECT 1136.3400 1947.8000 1139.3400 1948.2800 ;
        RECT 1136.3400 1953.2400 1139.3400 1953.7200 ;
        RECT 1136.3400 1958.6800 1139.3400 1959.1600 ;
        RECT 1136.3400 1942.3600 1139.3400 1942.8400 ;
        RECT 1136.3400 1931.4800 1139.3400 1931.9600 ;
        RECT 1136.3400 1936.9200 1139.3400 1937.4000 ;
        RECT 1093.1000 1947.8000 1094.1000 1948.2800 ;
        RECT 1093.1000 1953.2400 1094.1000 1953.7200 ;
        RECT 1093.1000 1958.6800 1094.1000 1959.1600 ;
        RECT 1093.1000 1931.4800 1094.1000 1931.9600 ;
        RECT 1093.1000 1936.9200 1094.1000 1937.4000 ;
        RECT 1093.1000 1942.3600 1094.1000 1942.8400 ;
        RECT 1136.3400 1920.6000 1139.3400 1921.0800 ;
        RECT 1136.3400 1926.0400 1139.3400 1926.5200 ;
        RECT 1093.1000 1920.6000 1094.1000 1921.0800 ;
        RECT 1093.1000 1926.0400 1094.1000 1926.5200 ;
        RECT 1048.1000 1947.8000 1049.1000 1948.2800 ;
        RECT 1048.1000 1953.2400 1049.1000 1953.7200 ;
        RECT 1048.1000 1958.6800 1049.1000 1959.1600 ;
        RECT 1048.1000 1931.4800 1049.1000 1931.9600 ;
        RECT 1048.1000 1936.9200 1049.1000 1937.4000 ;
        RECT 1048.1000 1942.3600 1049.1000 1942.8400 ;
        RECT 1048.1000 1920.6000 1049.1000 1921.0800 ;
        RECT 1048.1000 1926.0400 1049.1000 1926.5200 ;
        RECT 1003.1000 2007.6400 1004.1000 2008.1200 ;
        RECT 1003.1000 2013.0800 1004.1000 2013.5600 ;
        RECT 1003.1000 2018.5200 1004.1000 2019.0000 ;
        RECT 1003.1000 1991.3200 1004.1000 1991.8000 ;
        RECT 1003.1000 1996.7600 1004.1000 1997.2400 ;
        RECT 1003.1000 2002.2000 1004.1000 2002.6800 ;
        RECT 1003.1000 1980.4400 1004.1000 1980.9200 ;
        RECT 1003.1000 1985.8800 1004.1000 1986.3600 ;
        RECT 1003.1000 1964.1200 1004.1000 1964.6000 ;
        RECT 1003.1000 1969.5600 1004.1000 1970.0400 ;
        RECT 1003.1000 1975.0000 1004.1000 1975.4800 ;
        RECT 958.1000 2007.6400 959.1000 2008.1200 ;
        RECT 958.1000 2013.0800 959.1000 2013.5600 ;
        RECT 958.1000 2018.5200 959.1000 2019.0000 ;
        RECT 958.1000 1991.3200 959.1000 1991.8000 ;
        RECT 958.1000 1996.7600 959.1000 1997.2400 ;
        RECT 958.1000 2002.2000 959.1000 2002.6800 ;
        RECT 902.3400 2018.5200 905.3400 2019.0000 ;
        RECT 913.1000 2018.5200 914.1000 2019.0000 ;
        RECT 902.3400 2007.6400 905.3400 2008.1200 ;
        RECT 913.1000 2007.6400 914.1000 2008.1200 ;
        RECT 902.3400 2013.0800 905.3400 2013.5600 ;
        RECT 913.1000 2013.0800 914.1000 2013.5600 ;
        RECT 902.3400 2002.2000 905.3400 2002.6800 ;
        RECT 913.1000 2002.2000 914.1000 2002.6800 ;
        RECT 913.1000 1996.7600 914.1000 1997.2400 ;
        RECT 913.1000 1991.3200 914.1000 1991.8000 ;
        RECT 902.3400 1996.7600 905.3400 1997.2400 ;
        RECT 902.3400 1991.3200 905.3400 1991.8000 ;
        RECT 958.1000 1980.4400 959.1000 1980.9200 ;
        RECT 958.1000 1985.8800 959.1000 1986.3600 ;
        RECT 958.1000 1964.1200 959.1000 1964.6000 ;
        RECT 958.1000 1969.5600 959.1000 1970.0400 ;
        RECT 958.1000 1975.0000 959.1000 1975.4800 ;
        RECT 902.3400 1985.8800 905.3400 1986.3600 ;
        RECT 913.1000 1985.8800 914.1000 1986.3600 ;
        RECT 902.3400 1980.4400 905.3400 1980.9200 ;
        RECT 913.1000 1980.4400 914.1000 1980.9200 ;
        RECT 913.1000 1975.0000 914.1000 1975.4800 ;
        RECT 913.1000 1969.5600 914.1000 1970.0400 ;
        RECT 902.3400 1975.0000 905.3400 1975.4800 ;
        RECT 902.3400 1969.5600 905.3400 1970.0400 ;
        RECT 902.3400 1964.1200 905.3400 1964.6000 ;
        RECT 913.1000 1964.1200 914.1000 1964.6000 ;
        RECT 1003.1000 1947.8000 1004.1000 1948.2800 ;
        RECT 1003.1000 1953.2400 1004.1000 1953.7200 ;
        RECT 1003.1000 1958.6800 1004.1000 1959.1600 ;
        RECT 1003.1000 1931.4800 1004.1000 1931.9600 ;
        RECT 1003.1000 1936.9200 1004.1000 1937.4000 ;
        RECT 1003.1000 1942.3600 1004.1000 1942.8400 ;
        RECT 1003.1000 1920.6000 1004.1000 1921.0800 ;
        RECT 1003.1000 1926.0400 1004.1000 1926.5200 ;
        RECT 958.1000 1947.8000 959.1000 1948.2800 ;
        RECT 958.1000 1953.2400 959.1000 1953.7200 ;
        RECT 958.1000 1958.6800 959.1000 1959.1600 ;
        RECT 958.1000 1931.4800 959.1000 1931.9600 ;
        RECT 958.1000 1936.9200 959.1000 1937.4000 ;
        RECT 958.1000 1942.3600 959.1000 1942.8400 ;
        RECT 902.3400 1958.6800 905.3400 1959.1600 ;
        RECT 913.1000 1958.6800 914.1000 1959.1600 ;
        RECT 902.3400 1947.8000 905.3400 1948.2800 ;
        RECT 913.1000 1947.8000 914.1000 1948.2800 ;
        RECT 902.3400 1953.2400 905.3400 1953.7200 ;
        RECT 913.1000 1953.2400 914.1000 1953.7200 ;
        RECT 902.3400 1942.3600 905.3400 1942.8400 ;
        RECT 913.1000 1942.3600 914.1000 1942.8400 ;
        RECT 913.1000 1936.9200 914.1000 1937.4000 ;
        RECT 913.1000 1931.4800 914.1000 1931.9600 ;
        RECT 902.3400 1936.9200 905.3400 1937.4000 ;
        RECT 902.3400 1931.4800 905.3400 1931.9600 ;
        RECT 958.1000 1920.6000 959.1000 1921.0800 ;
        RECT 958.1000 1926.0400 959.1000 1926.5200 ;
        RECT 902.3400 1926.0400 905.3400 1926.5200 ;
        RECT 913.1000 1926.0400 914.1000 1926.5200 ;
        RECT 902.3400 1920.6000 905.3400 1921.0800 ;
        RECT 913.1000 1920.6000 914.1000 1921.0800 ;
        RECT 902.3400 2125.5100 1139.3400 2128.5100 ;
        RECT 902.3400 1912.4100 1139.3400 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 1682.7700 1094.1000 1898.8700 ;
        RECT 1048.1000 1682.7700 1049.1000 1898.8700 ;
        RECT 1003.1000 1682.7700 1004.1000 1898.8700 ;
        RECT 958.1000 1682.7700 959.1000 1898.8700 ;
        RECT 913.1000 1682.7700 914.1000 1898.8700 ;
        RECT 1136.3400 1682.7700 1139.3400 1898.8700 ;
        RECT 902.3400 1682.7700 905.3400 1898.8700 ;
      LAYER met3 ;
        RECT 1136.3400 1881.3600 1139.3400 1881.8400 ;
        RECT 1136.3400 1886.8000 1139.3400 1887.2800 ;
        RECT 1093.1000 1881.3600 1094.1000 1881.8400 ;
        RECT 1093.1000 1886.8000 1094.1000 1887.2800 ;
        RECT 1136.3400 1870.4800 1139.3400 1870.9600 ;
        RECT 1136.3400 1875.9200 1139.3400 1876.4000 ;
        RECT 1136.3400 1859.6000 1139.3400 1860.0800 ;
        RECT 1136.3400 1865.0400 1139.3400 1865.5200 ;
        RECT 1136.3400 1854.1600 1139.3400 1854.6400 ;
        RECT 1093.1000 1870.4800 1094.1000 1870.9600 ;
        RECT 1093.1000 1875.9200 1094.1000 1876.4000 ;
        RECT 1093.1000 1854.1600 1094.1000 1854.6400 ;
        RECT 1093.1000 1859.6000 1094.1000 1860.0800 ;
        RECT 1093.1000 1865.0400 1094.1000 1865.5200 ;
        RECT 1048.1000 1881.3600 1049.1000 1881.8400 ;
        RECT 1048.1000 1886.8000 1049.1000 1887.2800 ;
        RECT 1048.1000 1870.4800 1049.1000 1870.9600 ;
        RECT 1048.1000 1875.9200 1049.1000 1876.4000 ;
        RECT 1048.1000 1854.1600 1049.1000 1854.6400 ;
        RECT 1048.1000 1859.6000 1049.1000 1860.0800 ;
        RECT 1048.1000 1865.0400 1049.1000 1865.5200 ;
        RECT 1136.3400 1837.8400 1139.3400 1838.3200 ;
        RECT 1136.3400 1843.2800 1139.3400 1843.7600 ;
        RECT 1136.3400 1848.7200 1139.3400 1849.2000 ;
        RECT 1136.3400 1832.4000 1139.3400 1832.8800 ;
        RECT 1136.3400 1821.5200 1139.3400 1822.0000 ;
        RECT 1136.3400 1826.9600 1139.3400 1827.4400 ;
        RECT 1093.1000 1837.8400 1094.1000 1838.3200 ;
        RECT 1093.1000 1843.2800 1094.1000 1843.7600 ;
        RECT 1093.1000 1848.7200 1094.1000 1849.2000 ;
        RECT 1093.1000 1821.5200 1094.1000 1822.0000 ;
        RECT 1093.1000 1826.9600 1094.1000 1827.4400 ;
        RECT 1093.1000 1832.4000 1094.1000 1832.8800 ;
        RECT 1136.3400 1810.6400 1139.3400 1811.1200 ;
        RECT 1136.3400 1816.0800 1139.3400 1816.5600 ;
        RECT 1136.3400 1799.7600 1139.3400 1800.2400 ;
        RECT 1136.3400 1805.2000 1139.3400 1805.6800 ;
        RECT 1136.3400 1794.3200 1139.3400 1794.8000 ;
        RECT 1093.1000 1810.6400 1094.1000 1811.1200 ;
        RECT 1093.1000 1816.0800 1094.1000 1816.5600 ;
        RECT 1093.1000 1794.3200 1094.1000 1794.8000 ;
        RECT 1093.1000 1799.7600 1094.1000 1800.2400 ;
        RECT 1093.1000 1805.2000 1094.1000 1805.6800 ;
        RECT 1048.1000 1837.8400 1049.1000 1838.3200 ;
        RECT 1048.1000 1843.2800 1049.1000 1843.7600 ;
        RECT 1048.1000 1848.7200 1049.1000 1849.2000 ;
        RECT 1048.1000 1821.5200 1049.1000 1822.0000 ;
        RECT 1048.1000 1826.9600 1049.1000 1827.4400 ;
        RECT 1048.1000 1832.4000 1049.1000 1832.8800 ;
        RECT 1048.1000 1810.6400 1049.1000 1811.1200 ;
        RECT 1048.1000 1816.0800 1049.1000 1816.5600 ;
        RECT 1048.1000 1794.3200 1049.1000 1794.8000 ;
        RECT 1048.1000 1799.7600 1049.1000 1800.2400 ;
        RECT 1048.1000 1805.2000 1049.1000 1805.6800 ;
        RECT 1003.1000 1881.3600 1004.1000 1881.8400 ;
        RECT 1003.1000 1886.8000 1004.1000 1887.2800 ;
        RECT 1003.1000 1870.4800 1004.1000 1870.9600 ;
        RECT 1003.1000 1875.9200 1004.1000 1876.4000 ;
        RECT 1003.1000 1854.1600 1004.1000 1854.6400 ;
        RECT 1003.1000 1859.6000 1004.1000 1860.0800 ;
        RECT 1003.1000 1865.0400 1004.1000 1865.5200 ;
        RECT 958.1000 1881.3600 959.1000 1881.8400 ;
        RECT 958.1000 1886.8000 959.1000 1887.2800 ;
        RECT 913.1000 1886.8000 914.1000 1887.2800 ;
        RECT 913.1000 1881.3600 914.1000 1881.8400 ;
        RECT 902.3400 1886.8000 905.3400 1887.2800 ;
        RECT 902.3400 1881.3600 905.3400 1881.8400 ;
        RECT 958.1000 1870.4800 959.1000 1870.9600 ;
        RECT 958.1000 1875.9200 959.1000 1876.4000 ;
        RECT 958.1000 1854.1600 959.1000 1854.6400 ;
        RECT 958.1000 1859.6000 959.1000 1860.0800 ;
        RECT 958.1000 1865.0400 959.1000 1865.5200 ;
        RECT 902.3400 1875.9200 905.3400 1876.4000 ;
        RECT 913.1000 1875.9200 914.1000 1876.4000 ;
        RECT 902.3400 1870.4800 905.3400 1870.9600 ;
        RECT 913.1000 1870.4800 914.1000 1870.9600 ;
        RECT 913.1000 1865.0400 914.1000 1865.5200 ;
        RECT 913.1000 1859.6000 914.1000 1860.0800 ;
        RECT 902.3400 1865.0400 905.3400 1865.5200 ;
        RECT 902.3400 1859.6000 905.3400 1860.0800 ;
        RECT 902.3400 1854.1600 905.3400 1854.6400 ;
        RECT 913.1000 1854.1600 914.1000 1854.6400 ;
        RECT 1003.1000 1837.8400 1004.1000 1838.3200 ;
        RECT 1003.1000 1843.2800 1004.1000 1843.7600 ;
        RECT 1003.1000 1848.7200 1004.1000 1849.2000 ;
        RECT 1003.1000 1821.5200 1004.1000 1822.0000 ;
        RECT 1003.1000 1826.9600 1004.1000 1827.4400 ;
        RECT 1003.1000 1832.4000 1004.1000 1832.8800 ;
        RECT 1003.1000 1810.6400 1004.1000 1811.1200 ;
        RECT 1003.1000 1816.0800 1004.1000 1816.5600 ;
        RECT 1003.1000 1794.3200 1004.1000 1794.8000 ;
        RECT 1003.1000 1799.7600 1004.1000 1800.2400 ;
        RECT 1003.1000 1805.2000 1004.1000 1805.6800 ;
        RECT 958.1000 1837.8400 959.1000 1838.3200 ;
        RECT 958.1000 1843.2800 959.1000 1843.7600 ;
        RECT 958.1000 1848.7200 959.1000 1849.2000 ;
        RECT 958.1000 1821.5200 959.1000 1822.0000 ;
        RECT 958.1000 1826.9600 959.1000 1827.4400 ;
        RECT 958.1000 1832.4000 959.1000 1832.8800 ;
        RECT 902.3400 1848.7200 905.3400 1849.2000 ;
        RECT 913.1000 1848.7200 914.1000 1849.2000 ;
        RECT 902.3400 1837.8400 905.3400 1838.3200 ;
        RECT 913.1000 1837.8400 914.1000 1838.3200 ;
        RECT 902.3400 1843.2800 905.3400 1843.7600 ;
        RECT 913.1000 1843.2800 914.1000 1843.7600 ;
        RECT 902.3400 1832.4000 905.3400 1832.8800 ;
        RECT 913.1000 1832.4000 914.1000 1832.8800 ;
        RECT 913.1000 1826.9600 914.1000 1827.4400 ;
        RECT 913.1000 1821.5200 914.1000 1822.0000 ;
        RECT 902.3400 1826.9600 905.3400 1827.4400 ;
        RECT 902.3400 1821.5200 905.3400 1822.0000 ;
        RECT 958.1000 1810.6400 959.1000 1811.1200 ;
        RECT 958.1000 1816.0800 959.1000 1816.5600 ;
        RECT 958.1000 1794.3200 959.1000 1794.8000 ;
        RECT 958.1000 1799.7600 959.1000 1800.2400 ;
        RECT 958.1000 1805.2000 959.1000 1805.6800 ;
        RECT 902.3400 1816.0800 905.3400 1816.5600 ;
        RECT 913.1000 1816.0800 914.1000 1816.5600 ;
        RECT 902.3400 1810.6400 905.3400 1811.1200 ;
        RECT 913.1000 1810.6400 914.1000 1811.1200 ;
        RECT 913.1000 1805.2000 914.1000 1805.6800 ;
        RECT 913.1000 1799.7600 914.1000 1800.2400 ;
        RECT 902.3400 1805.2000 905.3400 1805.6800 ;
        RECT 902.3400 1799.7600 905.3400 1800.2400 ;
        RECT 902.3400 1794.3200 905.3400 1794.8000 ;
        RECT 913.1000 1794.3200 914.1000 1794.8000 ;
        RECT 1136.3400 1778.0000 1139.3400 1778.4800 ;
        RECT 1136.3400 1783.4400 1139.3400 1783.9200 ;
        RECT 1136.3400 1788.8800 1139.3400 1789.3600 ;
        RECT 1136.3400 1772.5600 1139.3400 1773.0400 ;
        RECT 1136.3400 1761.6800 1139.3400 1762.1600 ;
        RECT 1136.3400 1767.1200 1139.3400 1767.6000 ;
        RECT 1093.1000 1778.0000 1094.1000 1778.4800 ;
        RECT 1093.1000 1783.4400 1094.1000 1783.9200 ;
        RECT 1093.1000 1788.8800 1094.1000 1789.3600 ;
        RECT 1093.1000 1761.6800 1094.1000 1762.1600 ;
        RECT 1093.1000 1767.1200 1094.1000 1767.6000 ;
        RECT 1093.1000 1772.5600 1094.1000 1773.0400 ;
        RECT 1136.3400 1750.8000 1139.3400 1751.2800 ;
        RECT 1136.3400 1756.2400 1139.3400 1756.7200 ;
        RECT 1136.3400 1739.9200 1139.3400 1740.4000 ;
        RECT 1136.3400 1745.3600 1139.3400 1745.8400 ;
        RECT 1136.3400 1734.4800 1139.3400 1734.9600 ;
        RECT 1093.1000 1750.8000 1094.1000 1751.2800 ;
        RECT 1093.1000 1756.2400 1094.1000 1756.7200 ;
        RECT 1093.1000 1734.4800 1094.1000 1734.9600 ;
        RECT 1093.1000 1739.9200 1094.1000 1740.4000 ;
        RECT 1093.1000 1745.3600 1094.1000 1745.8400 ;
        RECT 1048.1000 1778.0000 1049.1000 1778.4800 ;
        RECT 1048.1000 1783.4400 1049.1000 1783.9200 ;
        RECT 1048.1000 1788.8800 1049.1000 1789.3600 ;
        RECT 1048.1000 1761.6800 1049.1000 1762.1600 ;
        RECT 1048.1000 1767.1200 1049.1000 1767.6000 ;
        RECT 1048.1000 1772.5600 1049.1000 1773.0400 ;
        RECT 1048.1000 1750.8000 1049.1000 1751.2800 ;
        RECT 1048.1000 1756.2400 1049.1000 1756.7200 ;
        RECT 1048.1000 1734.4800 1049.1000 1734.9600 ;
        RECT 1048.1000 1739.9200 1049.1000 1740.4000 ;
        RECT 1048.1000 1745.3600 1049.1000 1745.8400 ;
        RECT 1136.3400 1718.1600 1139.3400 1718.6400 ;
        RECT 1136.3400 1723.6000 1139.3400 1724.0800 ;
        RECT 1136.3400 1729.0400 1139.3400 1729.5200 ;
        RECT 1136.3400 1712.7200 1139.3400 1713.2000 ;
        RECT 1136.3400 1701.8400 1139.3400 1702.3200 ;
        RECT 1136.3400 1707.2800 1139.3400 1707.7600 ;
        RECT 1093.1000 1718.1600 1094.1000 1718.6400 ;
        RECT 1093.1000 1723.6000 1094.1000 1724.0800 ;
        RECT 1093.1000 1729.0400 1094.1000 1729.5200 ;
        RECT 1093.1000 1701.8400 1094.1000 1702.3200 ;
        RECT 1093.1000 1707.2800 1094.1000 1707.7600 ;
        RECT 1093.1000 1712.7200 1094.1000 1713.2000 ;
        RECT 1136.3400 1690.9600 1139.3400 1691.4400 ;
        RECT 1136.3400 1696.4000 1139.3400 1696.8800 ;
        RECT 1093.1000 1690.9600 1094.1000 1691.4400 ;
        RECT 1093.1000 1696.4000 1094.1000 1696.8800 ;
        RECT 1048.1000 1718.1600 1049.1000 1718.6400 ;
        RECT 1048.1000 1723.6000 1049.1000 1724.0800 ;
        RECT 1048.1000 1729.0400 1049.1000 1729.5200 ;
        RECT 1048.1000 1701.8400 1049.1000 1702.3200 ;
        RECT 1048.1000 1707.2800 1049.1000 1707.7600 ;
        RECT 1048.1000 1712.7200 1049.1000 1713.2000 ;
        RECT 1048.1000 1690.9600 1049.1000 1691.4400 ;
        RECT 1048.1000 1696.4000 1049.1000 1696.8800 ;
        RECT 1003.1000 1778.0000 1004.1000 1778.4800 ;
        RECT 1003.1000 1783.4400 1004.1000 1783.9200 ;
        RECT 1003.1000 1788.8800 1004.1000 1789.3600 ;
        RECT 1003.1000 1761.6800 1004.1000 1762.1600 ;
        RECT 1003.1000 1767.1200 1004.1000 1767.6000 ;
        RECT 1003.1000 1772.5600 1004.1000 1773.0400 ;
        RECT 1003.1000 1750.8000 1004.1000 1751.2800 ;
        RECT 1003.1000 1756.2400 1004.1000 1756.7200 ;
        RECT 1003.1000 1734.4800 1004.1000 1734.9600 ;
        RECT 1003.1000 1739.9200 1004.1000 1740.4000 ;
        RECT 1003.1000 1745.3600 1004.1000 1745.8400 ;
        RECT 958.1000 1778.0000 959.1000 1778.4800 ;
        RECT 958.1000 1783.4400 959.1000 1783.9200 ;
        RECT 958.1000 1788.8800 959.1000 1789.3600 ;
        RECT 958.1000 1761.6800 959.1000 1762.1600 ;
        RECT 958.1000 1767.1200 959.1000 1767.6000 ;
        RECT 958.1000 1772.5600 959.1000 1773.0400 ;
        RECT 902.3400 1788.8800 905.3400 1789.3600 ;
        RECT 913.1000 1788.8800 914.1000 1789.3600 ;
        RECT 902.3400 1778.0000 905.3400 1778.4800 ;
        RECT 913.1000 1778.0000 914.1000 1778.4800 ;
        RECT 902.3400 1783.4400 905.3400 1783.9200 ;
        RECT 913.1000 1783.4400 914.1000 1783.9200 ;
        RECT 902.3400 1772.5600 905.3400 1773.0400 ;
        RECT 913.1000 1772.5600 914.1000 1773.0400 ;
        RECT 913.1000 1767.1200 914.1000 1767.6000 ;
        RECT 913.1000 1761.6800 914.1000 1762.1600 ;
        RECT 902.3400 1767.1200 905.3400 1767.6000 ;
        RECT 902.3400 1761.6800 905.3400 1762.1600 ;
        RECT 958.1000 1750.8000 959.1000 1751.2800 ;
        RECT 958.1000 1756.2400 959.1000 1756.7200 ;
        RECT 958.1000 1734.4800 959.1000 1734.9600 ;
        RECT 958.1000 1739.9200 959.1000 1740.4000 ;
        RECT 958.1000 1745.3600 959.1000 1745.8400 ;
        RECT 902.3400 1756.2400 905.3400 1756.7200 ;
        RECT 913.1000 1756.2400 914.1000 1756.7200 ;
        RECT 902.3400 1750.8000 905.3400 1751.2800 ;
        RECT 913.1000 1750.8000 914.1000 1751.2800 ;
        RECT 913.1000 1745.3600 914.1000 1745.8400 ;
        RECT 913.1000 1739.9200 914.1000 1740.4000 ;
        RECT 902.3400 1745.3600 905.3400 1745.8400 ;
        RECT 902.3400 1739.9200 905.3400 1740.4000 ;
        RECT 902.3400 1734.4800 905.3400 1734.9600 ;
        RECT 913.1000 1734.4800 914.1000 1734.9600 ;
        RECT 1003.1000 1718.1600 1004.1000 1718.6400 ;
        RECT 1003.1000 1723.6000 1004.1000 1724.0800 ;
        RECT 1003.1000 1729.0400 1004.1000 1729.5200 ;
        RECT 1003.1000 1701.8400 1004.1000 1702.3200 ;
        RECT 1003.1000 1707.2800 1004.1000 1707.7600 ;
        RECT 1003.1000 1712.7200 1004.1000 1713.2000 ;
        RECT 1003.1000 1690.9600 1004.1000 1691.4400 ;
        RECT 1003.1000 1696.4000 1004.1000 1696.8800 ;
        RECT 958.1000 1718.1600 959.1000 1718.6400 ;
        RECT 958.1000 1723.6000 959.1000 1724.0800 ;
        RECT 958.1000 1729.0400 959.1000 1729.5200 ;
        RECT 958.1000 1701.8400 959.1000 1702.3200 ;
        RECT 958.1000 1707.2800 959.1000 1707.7600 ;
        RECT 958.1000 1712.7200 959.1000 1713.2000 ;
        RECT 902.3400 1729.0400 905.3400 1729.5200 ;
        RECT 913.1000 1729.0400 914.1000 1729.5200 ;
        RECT 902.3400 1718.1600 905.3400 1718.6400 ;
        RECT 913.1000 1718.1600 914.1000 1718.6400 ;
        RECT 902.3400 1723.6000 905.3400 1724.0800 ;
        RECT 913.1000 1723.6000 914.1000 1724.0800 ;
        RECT 902.3400 1712.7200 905.3400 1713.2000 ;
        RECT 913.1000 1712.7200 914.1000 1713.2000 ;
        RECT 913.1000 1707.2800 914.1000 1707.7600 ;
        RECT 913.1000 1701.8400 914.1000 1702.3200 ;
        RECT 902.3400 1707.2800 905.3400 1707.7600 ;
        RECT 902.3400 1701.8400 905.3400 1702.3200 ;
        RECT 958.1000 1690.9600 959.1000 1691.4400 ;
        RECT 958.1000 1696.4000 959.1000 1696.8800 ;
        RECT 902.3400 1696.4000 905.3400 1696.8800 ;
        RECT 913.1000 1696.4000 914.1000 1696.8800 ;
        RECT 902.3400 1690.9600 905.3400 1691.4400 ;
        RECT 913.1000 1690.9600 914.1000 1691.4400 ;
        RECT 902.3400 1895.8700 1139.3400 1898.8700 ;
        RECT 902.3400 1682.7700 1139.3400 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 1453.1300 1094.1000 1669.2300 ;
        RECT 1048.1000 1453.1300 1049.1000 1669.2300 ;
        RECT 1003.1000 1453.1300 1004.1000 1669.2300 ;
        RECT 958.1000 1453.1300 959.1000 1669.2300 ;
        RECT 913.1000 1453.1300 914.1000 1669.2300 ;
        RECT 1136.3400 1453.1300 1139.3400 1669.2300 ;
        RECT 902.3400 1453.1300 905.3400 1669.2300 ;
      LAYER met3 ;
        RECT 1136.3400 1651.7200 1139.3400 1652.2000 ;
        RECT 1136.3400 1657.1600 1139.3400 1657.6400 ;
        RECT 1093.1000 1651.7200 1094.1000 1652.2000 ;
        RECT 1093.1000 1657.1600 1094.1000 1657.6400 ;
        RECT 1136.3400 1640.8400 1139.3400 1641.3200 ;
        RECT 1136.3400 1646.2800 1139.3400 1646.7600 ;
        RECT 1136.3400 1629.9600 1139.3400 1630.4400 ;
        RECT 1136.3400 1635.4000 1139.3400 1635.8800 ;
        RECT 1136.3400 1624.5200 1139.3400 1625.0000 ;
        RECT 1093.1000 1640.8400 1094.1000 1641.3200 ;
        RECT 1093.1000 1646.2800 1094.1000 1646.7600 ;
        RECT 1093.1000 1624.5200 1094.1000 1625.0000 ;
        RECT 1093.1000 1629.9600 1094.1000 1630.4400 ;
        RECT 1093.1000 1635.4000 1094.1000 1635.8800 ;
        RECT 1048.1000 1651.7200 1049.1000 1652.2000 ;
        RECT 1048.1000 1657.1600 1049.1000 1657.6400 ;
        RECT 1048.1000 1640.8400 1049.1000 1641.3200 ;
        RECT 1048.1000 1646.2800 1049.1000 1646.7600 ;
        RECT 1048.1000 1624.5200 1049.1000 1625.0000 ;
        RECT 1048.1000 1629.9600 1049.1000 1630.4400 ;
        RECT 1048.1000 1635.4000 1049.1000 1635.8800 ;
        RECT 1136.3400 1608.2000 1139.3400 1608.6800 ;
        RECT 1136.3400 1613.6400 1139.3400 1614.1200 ;
        RECT 1136.3400 1619.0800 1139.3400 1619.5600 ;
        RECT 1136.3400 1602.7600 1139.3400 1603.2400 ;
        RECT 1136.3400 1591.8800 1139.3400 1592.3600 ;
        RECT 1136.3400 1597.3200 1139.3400 1597.8000 ;
        RECT 1093.1000 1608.2000 1094.1000 1608.6800 ;
        RECT 1093.1000 1613.6400 1094.1000 1614.1200 ;
        RECT 1093.1000 1619.0800 1094.1000 1619.5600 ;
        RECT 1093.1000 1591.8800 1094.1000 1592.3600 ;
        RECT 1093.1000 1597.3200 1094.1000 1597.8000 ;
        RECT 1093.1000 1602.7600 1094.1000 1603.2400 ;
        RECT 1136.3400 1581.0000 1139.3400 1581.4800 ;
        RECT 1136.3400 1586.4400 1139.3400 1586.9200 ;
        RECT 1136.3400 1570.1200 1139.3400 1570.6000 ;
        RECT 1136.3400 1575.5600 1139.3400 1576.0400 ;
        RECT 1136.3400 1564.6800 1139.3400 1565.1600 ;
        RECT 1093.1000 1581.0000 1094.1000 1581.4800 ;
        RECT 1093.1000 1586.4400 1094.1000 1586.9200 ;
        RECT 1093.1000 1564.6800 1094.1000 1565.1600 ;
        RECT 1093.1000 1570.1200 1094.1000 1570.6000 ;
        RECT 1093.1000 1575.5600 1094.1000 1576.0400 ;
        RECT 1048.1000 1608.2000 1049.1000 1608.6800 ;
        RECT 1048.1000 1613.6400 1049.1000 1614.1200 ;
        RECT 1048.1000 1619.0800 1049.1000 1619.5600 ;
        RECT 1048.1000 1591.8800 1049.1000 1592.3600 ;
        RECT 1048.1000 1597.3200 1049.1000 1597.8000 ;
        RECT 1048.1000 1602.7600 1049.1000 1603.2400 ;
        RECT 1048.1000 1581.0000 1049.1000 1581.4800 ;
        RECT 1048.1000 1586.4400 1049.1000 1586.9200 ;
        RECT 1048.1000 1564.6800 1049.1000 1565.1600 ;
        RECT 1048.1000 1570.1200 1049.1000 1570.6000 ;
        RECT 1048.1000 1575.5600 1049.1000 1576.0400 ;
        RECT 1003.1000 1651.7200 1004.1000 1652.2000 ;
        RECT 1003.1000 1657.1600 1004.1000 1657.6400 ;
        RECT 1003.1000 1640.8400 1004.1000 1641.3200 ;
        RECT 1003.1000 1646.2800 1004.1000 1646.7600 ;
        RECT 1003.1000 1624.5200 1004.1000 1625.0000 ;
        RECT 1003.1000 1629.9600 1004.1000 1630.4400 ;
        RECT 1003.1000 1635.4000 1004.1000 1635.8800 ;
        RECT 958.1000 1651.7200 959.1000 1652.2000 ;
        RECT 958.1000 1657.1600 959.1000 1657.6400 ;
        RECT 913.1000 1657.1600 914.1000 1657.6400 ;
        RECT 913.1000 1651.7200 914.1000 1652.2000 ;
        RECT 902.3400 1657.1600 905.3400 1657.6400 ;
        RECT 902.3400 1651.7200 905.3400 1652.2000 ;
        RECT 958.1000 1640.8400 959.1000 1641.3200 ;
        RECT 958.1000 1646.2800 959.1000 1646.7600 ;
        RECT 958.1000 1624.5200 959.1000 1625.0000 ;
        RECT 958.1000 1629.9600 959.1000 1630.4400 ;
        RECT 958.1000 1635.4000 959.1000 1635.8800 ;
        RECT 902.3400 1646.2800 905.3400 1646.7600 ;
        RECT 913.1000 1646.2800 914.1000 1646.7600 ;
        RECT 902.3400 1640.8400 905.3400 1641.3200 ;
        RECT 913.1000 1640.8400 914.1000 1641.3200 ;
        RECT 913.1000 1635.4000 914.1000 1635.8800 ;
        RECT 913.1000 1629.9600 914.1000 1630.4400 ;
        RECT 902.3400 1635.4000 905.3400 1635.8800 ;
        RECT 902.3400 1629.9600 905.3400 1630.4400 ;
        RECT 902.3400 1624.5200 905.3400 1625.0000 ;
        RECT 913.1000 1624.5200 914.1000 1625.0000 ;
        RECT 1003.1000 1608.2000 1004.1000 1608.6800 ;
        RECT 1003.1000 1613.6400 1004.1000 1614.1200 ;
        RECT 1003.1000 1619.0800 1004.1000 1619.5600 ;
        RECT 1003.1000 1591.8800 1004.1000 1592.3600 ;
        RECT 1003.1000 1597.3200 1004.1000 1597.8000 ;
        RECT 1003.1000 1602.7600 1004.1000 1603.2400 ;
        RECT 1003.1000 1581.0000 1004.1000 1581.4800 ;
        RECT 1003.1000 1586.4400 1004.1000 1586.9200 ;
        RECT 1003.1000 1564.6800 1004.1000 1565.1600 ;
        RECT 1003.1000 1570.1200 1004.1000 1570.6000 ;
        RECT 1003.1000 1575.5600 1004.1000 1576.0400 ;
        RECT 958.1000 1608.2000 959.1000 1608.6800 ;
        RECT 958.1000 1613.6400 959.1000 1614.1200 ;
        RECT 958.1000 1619.0800 959.1000 1619.5600 ;
        RECT 958.1000 1591.8800 959.1000 1592.3600 ;
        RECT 958.1000 1597.3200 959.1000 1597.8000 ;
        RECT 958.1000 1602.7600 959.1000 1603.2400 ;
        RECT 902.3400 1619.0800 905.3400 1619.5600 ;
        RECT 913.1000 1619.0800 914.1000 1619.5600 ;
        RECT 902.3400 1608.2000 905.3400 1608.6800 ;
        RECT 913.1000 1608.2000 914.1000 1608.6800 ;
        RECT 902.3400 1613.6400 905.3400 1614.1200 ;
        RECT 913.1000 1613.6400 914.1000 1614.1200 ;
        RECT 902.3400 1602.7600 905.3400 1603.2400 ;
        RECT 913.1000 1602.7600 914.1000 1603.2400 ;
        RECT 913.1000 1597.3200 914.1000 1597.8000 ;
        RECT 913.1000 1591.8800 914.1000 1592.3600 ;
        RECT 902.3400 1597.3200 905.3400 1597.8000 ;
        RECT 902.3400 1591.8800 905.3400 1592.3600 ;
        RECT 958.1000 1581.0000 959.1000 1581.4800 ;
        RECT 958.1000 1586.4400 959.1000 1586.9200 ;
        RECT 958.1000 1564.6800 959.1000 1565.1600 ;
        RECT 958.1000 1570.1200 959.1000 1570.6000 ;
        RECT 958.1000 1575.5600 959.1000 1576.0400 ;
        RECT 902.3400 1586.4400 905.3400 1586.9200 ;
        RECT 913.1000 1586.4400 914.1000 1586.9200 ;
        RECT 902.3400 1581.0000 905.3400 1581.4800 ;
        RECT 913.1000 1581.0000 914.1000 1581.4800 ;
        RECT 913.1000 1575.5600 914.1000 1576.0400 ;
        RECT 913.1000 1570.1200 914.1000 1570.6000 ;
        RECT 902.3400 1575.5600 905.3400 1576.0400 ;
        RECT 902.3400 1570.1200 905.3400 1570.6000 ;
        RECT 902.3400 1564.6800 905.3400 1565.1600 ;
        RECT 913.1000 1564.6800 914.1000 1565.1600 ;
        RECT 1136.3400 1548.3600 1139.3400 1548.8400 ;
        RECT 1136.3400 1553.8000 1139.3400 1554.2800 ;
        RECT 1136.3400 1559.2400 1139.3400 1559.7200 ;
        RECT 1136.3400 1542.9200 1139.3400 1543.4000 ;
        RECT 1136.3400 1532.0400 1139.3400 1532.5200 ;
        RECT 1136.3400 1537.4800 1139.3400 1537.9600 ;
        RECT 1093.1000 1548.3600 1094.1000 1548.8400 ;
        RECT 1093.1000 1553.8000 1094.1000 1554.2800 ;
        RECT 1093.1000 1559.2400 1094.1000 1559.7200 ;
        RECT 1093.1000 1532.0400 1094.1000 1532.5200 ;
        RECT 1093.1000 1537.4800 1094.1000 1537.9600 ;
        RECT 1093.1000 1542.9200 1094.1000 1543.4000 ;
        RECT 1136.3400 1521.1600 1139.3400 1521.6400 ;
        RECT 1136.3400 1526.6000 1139.3400 1527.0800 ;
        RECT 1136.3400 1510.2800 1139.3400 1510.7600 ;
        RECT 1136.3400 1515.7200 1139.3400 1516.2000 ;
        RECT 1136.3400 1504.8400 1139.3400 1505.3200 ;
        RECT 1093.1000 1521.1600 1094.1000 1521.6400 ;
        RECT 1093.1000 1526.6000 1094.1000 1527.0800 ;
        RECT 1093.1000 1504.8400 1094.1000 1505.3200 ;
        RECT 1093.1000 1510.2800 1094.1000 1510.7600 ;
        RECT 1093.1000 1515.7200 1094.1000 1516.2000 ;
        RECT 1048.1000 1548.3600 1049.1000 1548.8400 ;
        RECT 1048.1000 1553.8000 1049.1000 1554.2800 ;
        RECT 1048.1000 1559.2400 1049.1000 1559.7200 ;
        RECT 1048.1000 1532.0400 1049.1000 1532.5200 ;
        RECT 1048.1000 1537.4800 1049.1000 1537.9600 ;
        RECT 1048.1000 1542.9200 1049.1000 1543.4000 ;
        RECT 1048.1000 1521.1600 1049.1000 1521.6400 ;
        RECT 1048.1000 1526.6000 1049.1000 1527.0800 ;
        RECT 1048.1000 1504.8400 1049.1000 1505.3200 ;
        RECT 1048.1000 1510.2800 1049.1000 1510.7600 ;
        RECT 1048.1000 1515.7200 1049.1000 1516.2000 ;
        RECT 1136.3400 1488.5200 1139.3400 1489.0000 ;
        RECT 1136.3400 1493.9600 1139.3400 1494.4400 ;
        RECT 1136.3400 1499.4000 1139.3400 1499.8800 ;
        RECT 1136.3400 1483.0800 1139.3400 1483.5600 ;
        RECT 1136.3400 1472.2000 1139.3400 1472.6800 ;
        RECT 1136.3400 1477.6400 1139.3400 1478.1200 ;
        RECT 1093.1000 1488.5200 1094.1000 1489.0000 ;
        RECT 1093.1000 1493.9600 1094.1000 1494.4400 ;
        RECT 1093.1000 1499.4000 1094.1000 1499.8800 ;
        RECT 1093.1000 1472.2000 1094.1000 1472.6800 ;
        RECT 1093.1000 1477.6400 1094.1000 1478.1200 ;
        RECT 1093.1000 1483.0800 1094.1000 1483.5600 ;
        RECT 1136.3400 1461.3200 1139.3400 1461.8000 ;
        RECT 1136.3400 1466.7600 1139.3400 1467.2400 ;
        RECT 1093.1000 1461.3200 1094.1000 1461.8000 ;
        RECT 1093.1000 1466.7600 1094.1000 1467.2400 ;
        RECT 1048.1000 1488.5200 1049.1000 1489.0000 ;
        RECT 1048.1000 1493.9600 1049.1000 1494.4400 ;
        RECT 1048.1000 1499.4000 1049.1000 1499.8800 ;
        RECT 1048.1000 1472.2000 1049.1000 1472.6800 ;
        RECT 1048.1000 1477.6400 1049.1000 1478.1200 ;
        RECT 1048.1000 1483.0800 1049.1000 1483.5600 ;
        RECT 1048.1000 1461.3200 1049.1000 1461.8000 ;
        RECT 1048.1000 1466.7600 1049.1000 1467.2400 ;
        RECT 1003.1000 1548.3600 1004.1000 1548.8400 ;
        RECT 1003.1000 1553.8000 1004.1000 1554.2800 ;
        RECT 1003.1000 1559.2400 1004.1000 1559.7200 ;
        RECT 1003.1000 1532.0400 1004.1000 1532.5200 ;
        RECT 1003.1000 1537.4800 1004.1000 1537.9600 ;
        RECT 1003.1000 1542.9200 1004.1000 1543.4000 ;
        RECT 1003.1000 1521.1600 1004.1000 1521.6400 ;
        RECT 1003.1000 1526.6000 1004.1000 1527.0800 ;
        RECT 1003.1000 1504.8400 1004.1000 1505.3200 ;
        RECT 1003.1000 1510.2800 1004.1000 1510.7600 ;
        RECT 1003.1000 1515.7200 1004.1000 1516.2000 ;
        RECT 958.1000 1548.3600 959.1000 1548.8400 ;
        RECT 958.1000 1553.8000 959.1000 1554.2800 ;
        RECT 958.1000 1559.2400 959.1000 1559.7200 ;
        RECT 958.1000 1532.0400 959.1000 1532.5200 ;
        RECT 958.1000 1537.4800 959.1000 1537.9600 ;
        RECT 958.1000 1542.9200 959.1000 1543.4000 ;
        RECT 902.3400 1559.2400 905.3400 1559.7200 ;
        RECT 913.1000 1559.2400 914.1000 1559.7200 ;
        RECT 902.3400 1548.3600 905.3400 1548.8400 ;
        RECT 913.1000 1548.3600 914.1000 1548.8400 ;
        RECT 902.3400 1553.8000 905.3400 1554.2800 ;
        RECT 913.1000 1553.8000 914.1000 1554.2800 ;
        RECT 902.3400 1542.9200 905.3400 1543.4000 ;
        RECT 913.1000 1542.9200 914.1000 1543.4000 ;
        RECT 913.1000 1537.4800 914.1000 1537.9600 ;
        RECT 913.1000 1532.0400 914.1000 1532.5200 ;
        RECT 902.3400 1537.4800 905.3400 1537.9600 ;
        RECT 902.3400 1532.0400 905.3400 1532.5200 ;
        RECT 958.1000 1521.1600 959.1000 1521.6400 ;
        RECT 958.1000 1526.6000 959.1000 1527.0800 ;
        RECT 958.1000 1504.8400 959.1000 1505.3200 ;
        RECT 958.1000 1510.2800 959.1000 1510.7600 ;
        RECT 958.1000 1515.7200 959.1000 1516.2000 ;
        RECT 902.3400 1526.6000 905.3400 1527.0800 ;
        RECT 913.1000 1526.6000 914.1000 1527.0800 ;
        RECT 902.3400 1521.1600 905.3400 1521.6400 ;
        RECT 913.1000 1521.1600 914.1000 1521.6400 ;
        RECT 913.1000 1515.7200 914.1000 1516.2000 ;
        RECT 913.1000 1510.2800 914.1000 1510.7600 ;
        RECT 902.3400 1515.7200 905.3400 1516.2000 ;
        RECT 902.3400 1510.2800 905.3400 1510.7600 ;
        RECT 902.3400 1504.8400 905.3400 1505.3200 ;
        RECT 913.1000 1504.8400 914.1000 1505.3200 ;
        RECT 1003.1000 1488.5200 1004.1000 1489.0000 ;
        RECT 1003.1000 1493.9600 1004.1000 1494.4400 ;
        RECT 1003.1000 1499.4000 1004.1000 1499.8800 ;
        RECT 1003.1000 1472.2000 1004.1000 1472.6800 ;
        RECT 1003.1000 1477.6400 1004.1000 1478.1200 ;
        RECT 1003.1000 1483.0800 1004.1000 1483.5600 ;
        RECT 1003.1000 1461.3200 1004.1000 1461.8000 ;
        RECT 1003.1000 1466.7600 1004.1000 1467.2400 ;
        RECT 958.1000 1488.5200 959.1000 1489.0000 ;
        RECT 958.1000 1493.9600 959.1000 1494.4400 ;
        RECT 958.1000 1499.4000 959.1000 1499.8800 ;
        RECT 958.1000 1472.2000 959.1000 1472.6800 ;
        RECT 958.1000 1477.6400 959.1000 1478.1200 ;
        RECT 958.1000 1483.0800 959.1000 1483.5600 ;
        RECT 902.3400 1499.4000 905.3400 1499.8800 ;
        RECT 913.1000 1499.4000 914.1000 1499.8800 ;
        RECT 902.3400 1488.5200 905.3400 1489.0000 ;
        RECT 913.1000 1488.5200 914.1000 1489.0000 ;
        RECT 902.3400 1493.9600 905.3400 1494.4400 ;
        RECT 913.1000 1493.9600 914.1000 1494.4400 ;
        RECT 902.3400 1483.0800 905.3400 1483.5600 ;
        RECT 913.1000 1483.0800 914.1000 1483.5600 ;
        RECT 913.1000 1477.6400 914.1000 1478.1200 ;
        RECT 913.1000 1472.2000 914.1000 1472.6800 ;
        RECT 902.3400 1477.6400 905.3400 1478.1200 ;
        RECT 902.3400 1472.2000 905.3400 1472.6800 ;
        RECT 958.1000 1461.3200 959.1000 1461.8000 ;
        RECT 958.1000 1466.7600 959.1000 1467.2400 ;
        RECT 902.3400 1466.7600 905.3400 1467.2400 ;
        RECT 913.1000 1466.7600 914.1000 1467.2400 ;
        RECT 902.3400 1461.3200 905.3400 1461.8000 ;
        RECT 913.1000 1461.3200 914.1000 1461.8000 ;
        RECT 902.3400 1666.2300 1139.3400 1669.2300 ;
        RECT 902.3400 1453.1300 1139.3400 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 1223.4900 1094.1000 1439.5900 ;
        RECT 1048.1000 1223.4900 1049.1000 1439.5900 ;
        RECT 1003.1000 1223.4900 1004.1000 1439.5900 ;
        RECT 958.1000 1223.4900 959.1000 1439.5900 ;
        RECT 913.1000 1223.4900 914.1000 1439.5900 ;
        RECT 1136.3400 1223.4900 1139.3400 1439.5900 ;
        RECT 902.3400 1223.4900 905.3400 1439.5900 ;
      LAYER met3 ;
        RECT 1136.3400 1422.0800 1139.3400 1422.5600 ;
        RECT 1136.3400 1427.5200 1139.3400 1428.0000 ;
        RECT 1093.1000 1422.0800 1094.1000 1422.5600 ;
        RECT 1093.1000 1427.5200 1094.1000 1428.0000 ;
        RECT 1136.3400 1411.2000 1139.3400 1411.6800 ;
        RECT 1136.3400 1416.6400 1139.3400 1417.1200 ;
        RECT 1136.3400 1400.3200 1139.3400 1400.8000 ;
        RECT 1136.3400 1405.7600 1139.3400 1406.2400 ;
        RECT 1136.3400 1394.8800 1139.3400 1395.3600 ;
        RECT 1093.1000 1411.2000 1094.1000 1411.6800 ;
        RECT 1093.1000 1416.6400 1094.1000 1417.1200 ;
        RECT 1093.1000 1394.8800 1094.1000 1395.3600 ;
        RECT 1093.1000 1400.3200 1094.1000 1400.8000 ;
        RECT 1093.1000 1405.7600 1094.1000 1406.2400 ;
        RECT 1048.1000 1422.0800 1049.1000 1422.5600 ;
        RECT 1048.1000 1427.5200 1049.1000 1428.0000 ;
        RECT 1048.1000 1411.2000 1049.1000 1411.6800 ;
        RECT 1048.1000 1416.6400 1049.1000 1417.1200 ;
        RECT 1048.1000 1394.8800 1049.1000 1395.3600 ;
        RECT 1048.1000 1400.3200 1049.1000 1400.8000 ;
        RECT 1048.1000 1405.7600 1049.1000 1406.2400 ;
        RECT 1136.3400 1378.5600 1139.3400 1379.0400 ;
        RECT 1136.3400 1384.0000 1139.3400 1384.4800 ;
        RECT 1136.3400 1389.4400 1139.3400 1389.9200 ;
        RECT 1136.3400 1373.1200 1139.3400 1373.6000 ;
        RECT 1136.3400 1362.2400 1139.3400 1362.7200 ;
        RECT 1136.3400 1367.6800 1139.3400 1368.1600 ;
        RECT 1093.1000 1378.5600 1094.1000 1379.0400 ;
        RECT 1093.1000 1384.0000 1094.1000 1384.4800 ;
        RECT 1093.1000 1389.4400 1094.1000 1389.9200 ;
        RECT 1093.1000 1362.2400 1094.1000 1362.7200 ;
        RECT 1093.1000 1367.6800 1094.1000 1368.1600 ;
        RECT 1093.1000 1373.1200 1094.1000 1373.6000 ;
        RECT 1136.3400 1351.3600 1139.3400 1351.8400 ;
        RECT 1136.3400 1356.8000 1139.3400 1357.2800 ;
        RECT 1136.3400 1340.4800 1139.3400 1340.9600 ;
        RECT 1136.3400 1345.9200 1139.3400 1346.4000 ;
        RECT 1136.3400 1335.0400 1139.3400 1335.5200 ;
        RECT 1093.1000 1351.3600 1094.1000 1351.8400 ;
        RECT 1093.1000 1356.8000 1094.1000 1357.2800 ;
        RECT 1093.1000 1335.0400 1094.1000 1335.5200 ;
        RECT 1093.1000 1340.4800 1094.1000 1340.9600 ;
        RECT 1093.1000 1345.9200 1094.1000 1346.4000 ;
        RECT 1048.1000 1378.5600 1049.1000 1379.0400 ;
        RECT 1048.1000 1384.0000 1049.1000 1384.4800 ;
        RECT 1048.1000 1389.4400 1049.1000 1389.9200 ;
        RECT 1048.1000 1362.2400 1049.1000 1362.7200 ;
        RECT 1048.1000 1367.6800 1049.1000 1368.1600 ;
        RECT 1048.1000 1373.1200 1049.1000 1373.6000 ;
        RECT 1048.1000 1351.3600 1049.1000 1351.8400 ;
        RECT 1048.1000 1356.8000 1049.1000 1357.2800 ;
        RECT 1048.1000 1335.0400 1049.1000 1335.5200 ;
        RECT 1048.1000 1340.4800 1049.1000 1340.9600 ;
        RECT 1048.1000 1345.9200 1049.1000 1346.4000 ;
        RECT 1003.1000 1422.0800 1004.1000 1422.5600 ;
        RECT 1003.1000 1427.5200 1004.1000 1428.0000 ;
        RECT 1003.1000 1411.2000 1004.1000 1411.6800 ;
        RECT 1003.1000 1416.6400 1004.1000 1417.1200 ;
        RECT 1003.1000 1394.8800 1004.1000 1395.3600 ;
        RECT 1003.1000 1400.3200 1004.1000 1400.8000 ;
        RECT 1003.1000 1405.7600 1004.1000 1406.2400 ;
        RECT 958.1000 1422.0800 959.1000 1422.5600 ;
        RECT 958.1000 1427.5200 959.1000 1428.0000 ;
        RECT 913.1000 1427.5200 914.1000 1428.0000 ;
        RECT 913.1000 1422.0800 914.1000 1422.5600 ;
        RECT 902.3400 1427.5200 905.3400 1428.0000 ;
        RECT 902.3400 1422.0800 905.3400 1422.5600 ;
        RECT 958.1000 1411.2000 959.1000 1411.6800 ;
        RECT 958.1000 1416.6400 959.1000 1417.1200 ;
        RECT 958.1000 1394.8800 959.1000 1395.3600 ;
        RECT 958.1000 1400.3200 959.1000 1400.8000 ;
        RECT 958.1000 1405.7600 959.1000 1406.2400 ;
        RECT 902.3400 1416.6400 905.3400 1417.1200 ;
        RECT 913.1000 1416.6400 914.1000 1417.1200 ;
        RECT 902.3400 1411.2000 905.3400 1411.6800 ;
        RECT 913.1000 1411.2000 914.1000 1411.6800 ;
        RECT 913.1000 1405.7600 914.1000 1406.2400 ;
        RECT 913.1000 1400.3200 914.1000 1400.8000 ;
        RECT 902.3400 1405.7600 905.3400 1406.2400 ;
        RECT 902.3400 1400.3200 905.3400 1400.8000 ;
        RECT 902.3400 1394.8800 905.3400 1395.3600 ;
        RECT 913.1000 1394.8800 914.1000 1395.3600 ;
        RECT 1003.1000 1378.5600 1004.1000 1379.0400 ;
        RECT 1003.1000 1384.0000 1004.1000 1384.4800 ;
        RECT 1003.1000 1389.4400 1004.1000 1389.9200 ;
        RECT 1003.1000 1362.2400 1004.1000 1362.7200 ;
        RECT 1003.1000 1367.6800 1004.1000 1368.1600 ;
        RECT 1003.1000 1373.1200 1004.1000 1373.6000 ;
        RECT 1003.1000 1351.3600 1004.1000 1351.8400 ;
        RECT 1003.1000 1356.8000 1004.1000 1357.2800 ;
        RECT 1003.1000 1335.0400 1004.1000 1335.5200 ;
        RECT 1003.1000 1340.4800 1004.1000 1340.9600 ;
        RECT 1003.1000 1345.9200 1004.1000 1346.4000 ;
        RECT 958.1000 1378.5600 959.1000 1379.0400 ;
        RECT 958.1000 1384.0000 959.1000 1384.4800 ;
        RECT 958.1000 1389.4400 959.1000 1389.9200 ;
        RECT 958.1000 1362.2400 959.1000 1362.7200 ;
        RECT 958.1000 1367.6800 959.1000 1368.1600 ;
        RECT 958.1000 1373.1200 959.1000 1373.6000 ;
        RECT 902.3400 1389.4400 905.3400 1389.9200 ;
        RECT 913.1000 1389.4400 914.1000 1389.9200 ;
        RECT 902.3400 1378.5600 905.3400 1379.0400 ;
        RECT 913.1000 1378.5600 914.1000 1379.0400 ;
        RECT 902.3400 1384.0000 905.3400 1384.4800 ;
        RECT 913.1000 1384.0000 914.1000 1384.4800 ;
        RECT 902.3400 1373.1200 905.3400 1373.6000 ;
        RECT 913.1000 1373.1200 914.1000 1373.6000 ;
        RECT 913.1000 1367.6800 914.1000 1368.1600 ;
        RECT 913.1000 1362.2400 914.1000 1362.7200 ;
        RECT 902.3400 1367.6800 905.3400 1368.1600 ;
        RECT 902.3400 1362.2400 905.3400 1362.7200 ;
        RECT 958.1000 1351.3600 959.1000 1351.8400 ;
        RECT 958.1000 1356.8000 959.1000 1357.2800 ;
        RECT 958.1000 1335.0400 959.1000 1335.5200 ;
        RECT 958.1000 1340.4800 959.1000 1340.9600 ;
        RECT 958.1000 1345.9200 959.1000 1346.4000 ;
        RECT 902.3400 1356.8000 905.3400 1357.2800 ;
        RECT 913.1000 1356.8000 914.1000 1357.2800 ;
        RECT 902.3400 1351.3600 905.3400 1351.8400 ;
        RECT 913.1000 1351.3600 914.1000 1351.8400 ;
        RECT 913.1000 1345.9200 914.1000 1346.4000 ;
        RECT 913.1000 1340.4800 914.1000 1340.9600 ;
        RECT 902.3400 1345.9200 905.3400 1346.4000 ;
        RECT 902.3400 1340.4800 905.3400 1340.9600 ;
        RECT 902.3400 1335.0400 905.3400 1335.5200 ;
        RECT 913.1000 1335.0400 914.1000 1335.5200 ;
        RECT 1136.3400 1318.7200 1139.3400 1319.2000 ;
        RECT 1136.3400 1324.1600 1139.3400 1324.6400 ;
        RECT 1136.3400 1329.6000 1139.3400 1330.0800 ;
        RECT 1136.3400 1313.2800 1139.3400 1313.7600 ;
        RECT 1136.3400 1302.4000 1139.3400 1302.8800 ;
        RECT 1136.3400 1307.8400 1139.3400 1308.3200 ;
        RECT 1093.1000 1318.7200 1094.1000 1319.2000 ;
        RECT 1093.1000 1324.1600 1094.1000 1324.6400 ;
        RECT 1093.1000 1329.6000 1094.1000 1330.0800 ;
        RECT 1093.1000 1302.4000 1094.1000 1302.8800 ;
        RECT 1093.1000 1307.8400 1094.1000 1308.3200 ;
        RECT 1093.1000 1313.2800 1094.1000 1313.7600 ;
        RECT 1136.3400 1291.5200 1139.3400 1292.0000 ;
        RECT 1136.3400 1296.9600 1139.3400 1297.4400 ;
        RECT 1136.3400 1280.6400 1139.3400 1281.1200 ;
        RECT 1136.3400 1286.0800 1139.3400 1286.5600 ;
        RECT 1136.3400 1275.2000 1139.3400 1275.6800 ;
        RECT 1093.1000 1291.5200 1094.1000 1292.0000 ;
        RECT 1093.1000 1296.9600 1094.1000 1297.4400 ;
        RECT 1093.1000 1275.2000 1094.1000 1275.6800 ;
        RECT 1093.1000 1280.6400 1094.1000 1281.1200 ;
        RECT 1093.1000 1286.0800 1094.1000 1286.5600 ;
        RECT 1048.1000 1318.7200 1049.1000 1319.2000 ;
        RECT 1048.1000 1324.1600 1049.1000 1324.6400 ;
        RECT 1048.1000 1329.6000 1049.1000 1330.0800 ;
        RECT 1048.1000 1302.4000 1049.1000 1302.8800 ;
        RECT 1048.1000 1307.8400 1049.1000 1308.3200 ;
        RECT 1048.1000 1313.2800 1049.1000 1313.7600 ;
        RECT 1048.1000 1291.5200 1049.1000 1292.0000 ;
        RECT 1048.1000 1296.9600 1049.1000 1297.4400 ;
        RECT 1048.1000 1275.2000 1049.1000 1275.6800 ;
        RECT 1048.1000 1280.6400 1049.1000 1281.1200 ;
        RECT 1048.1000 1286.0800 1049.1000 1286.5600 ;
        RECT 1136.3400 1258.8800 1139.3400 1259.3600 ;
        RECT 1136.3400 1264.3200 1139.3400 1264.8000 ;
        RECT 1136.3400 1269.7600 1139.3400 1270.2400 ;
        RECT 1136.3400 1253.4400 1139.3400 1253.9200 ;
        RECT 1136.3400 1242.5600 1139.3400 1243.0400 ;
        RECT 1136.3400 1248.0000 1139.3400 1248.4800 ;
        RECT 1093.1000 1258.8800 1094.1000 1259.3600 ;
        RECT 1093.1000 1264.3200 1094.1000 1264.8000 ;
        RECT 1093.1000 1269.7600 1094.1000 1270.2400 ;
        RECT 1093.1000 1242.5600 1094.1000 1243.0400 ;
        RECT 1093.1000 1248.0000 1094.1000 1248.4800 ;
        RECT 1093.1000 1253.4400 1094.1000 1253.9200 ;
        RECT 1136.3400 1231.6800 1139.3400 1232.1600 ;
        RECT 1136.3400 1237.1200 1139.3400 1237.6000 ;
        RECT 1093.1000 1231.6800 1094.1000 1232.1600 ;
        RECT 1093.1000 1237.1200 1094.1000 1237.6000 ;
        RECT 1048.1000 1258.8800 1049.1000 1259.3600 ;
        RECT 1048.1000 1264.3200 1049.1000 1264.8000 ;
        RECT 1048.1000 1269.7600 1049.1000 1270.2400 ;
        RECT 1048.1000 1242.5600 1049.1000 1243.0400 ;
        RECT 1048.1000 1248.0000 1049.1000 1248.4800 ;
        RECT 1048.1000 1253.4400 1049.1000 1253.9200 ;
        RECT 1048.1000 1231.6800 1049.1000 1232.1600 ;
        RECT 1048.1000 1237.1200 1049.1000 1237.6000 ;
        RECT 1003.1000 1318.7200 1004.1000 1319.2000 ;
        RECT 1003.1000 1324.1600 1004.1000 1324.6400 ;
        RECT 1003.1000 1329.6000 1004.1000 1330.0800 ;
        RECT 1003.1000 1302.4000 1004.1000 1302.8800 ;
        RECT 1003.1000 1307.8400 1004.1000 1308.3200 ;
        RECT 1003.1000 1313.2800 1004.1000 1313.7600 ;
        RECT 1003.1000 1291.5200 1004.1000 1292.0000 ;
        RECT 1003.1000 1296.9600 1004.1000 1297.4400 ;
        RECT 1003.1000 1275.2000 1004.1000 1275.6800 ;
        RECT 1003.1000 1280.6400 1004.1000 1281.1200 ;
        RECT 1003.1000 1286.0800 1004.1000 1286.5600 ;
        RECT 958.1000 1318.7200 959.1000 1319.2000 ;
        RECT 958.1000 1324.1600 959.1000 1324.6400 ;
        RECT 958.1000 1329.6000 959.1000 1330.0800 ;
        RECT 958.1000 1302.4000 959.1000 1302.8800 ;
        RECT 958.1000 1307.8400 959.1000 1308.3200 ;
        RECT 958.1000 1313.2800 959.1000 1313.7600 ;
        RECT 902.3400 1329.6000 905.3400 1330.0800 ;
        RECT 913.1000 1329.6000 914.1000 1330.0800 ;
        RECT 902.3400 1318.7200 905.3400 1319.2000 ;
        RECT 913.1000 1318.7200 914.1000 1319.2000 ;
        RECT 902.3400 1324.1600 905.3400 1324.6400 ;
        RECT 913.1000 1324.1600 914.1000 1324.6400 ;
        RECT 902.3400 1313.2800 905.3400 1313.7600 ;
        RECT 913.1000 1313.2800 914.1000 1313.7600 ;
        RECT 913.1000 1307.8400 914.1000 1308.3200 ;
        RECT 913.1000 1302.4000 914.1000 1302.8800 ;
        RECT 902.3400 1307.8400 905.3400 1308.3200 ;
        RECT 902.3400 1302.4000 905.3400 1302.8800 ;
        RECT 958.1000 1291.5200 959.1000 1292.0000 ;
        RECT 958.1000 1296.9600 959.1000 1297.4400 ;
        RECT 958.1000 1275.2000 959.1000 1275.6800 ;
        RECT 958.1000 1280.6400 959.1000 1281.1200 ;
        RECT 958.1000 1286.0800 959.1000 1286.5600 ;
        RECT 902.3400 1296.9600 905.3400 1297.4400 ;
        RECT 913.1000 1296.9600 914.1000 1297.4400 ;
        RECT 902.3400 1291.5200 905.3400 1292.0000 ;
        RECT 913.1000 1291.5200 914.1000 1292.0000 ;
        RECT 913.1000 1286.0800 914.1000 1286.5600 ;
        RECT 913.1000 1280.6400 914.1000 1281.1200 ;
        RECT 902.3400 1286.0800 905.3400 1286.5600 ;
        RECT 902.3400 1280.6400 905.3400 1281.1200 ;
        RECT 902.3400 1275.2000 905.3400 1275.6800 ;
        RECT 913.1000 1275.2000 914.1000 1275.6800 ;
        RECT 1003.1000 1258.8800 1004.1000 1259.3600 ;
        RECT 1003.1000 1264.3200 1004.1000 1264.8000 ;
        RECT 1003.1000 1269.7600 1004.1000 1270.2400 ;
        RECT 1003.1000 1242.5600 1004.1000 1243.0400 ;
        RECT 1003.1000 1248.0000 1004.1000 1248.4800 ;
        RECT 1003.1000 1253.4400 1004.1000 1253.9200 ;
        RECT 1003.1000 1231.6800 1004.1000 1232.1600 ;
        RECT 1003.1000 1237.1200 1004.1000 1237.6000 ;
        RECT 958.1000 1258.8800 959.1000 1259.3600 ;
        RECT 958.1000 1264.3200 959.1000 1264.8000 ;
        RECT 958.1000 1269.7600 959.1000 1270.2400 ;
        RECT 958.1000 1242.5600 959.1000 1243.0400 ;
        RECT 958.1000 1248.0000 959.1000 1248.4800 ;
        RECT 958.1000 1253.4400 959.1000 1253.9200 ;
        RECT 902.3400 1269.7600 905.3400 1270.2400 ;
        RECT 913.1000 1269.7600 914.1000 1270.2400 ;
        RECT 902.3400 1258.8800 905.3400 1259.3600 ;
        RECT 913.1000 1258.8800 914.1000 1259.3600 ;
        RECT 902.3400 1264.3200 905.3400 1264.8000 ;
        RECT 913.1000 1264.3200 914.1000 1264.8000 ;
        RECT 902.3400 1253.4400 905.3400 1253.9200 ;
        RECT 913.1000 1253.4400 914.1000 1253.9200 ;
        RECT 913.1000 1248.0000 914.1000 1248.4800 ;
        RECT 913.1000 1242.5600 914.1000 1243.0400 ;
        RECT 902.3400 1248.0000 905.3400 1248.4800 ;
        RECT 902.3400 1242.5600 905.3400 1243.0400 ;
        RECT 958.1000 1231.6800 959.1000 1232.1600 ;
        RECT 958.1000 1237.1200 959.1000 1237.6000 ;
        RECT 902.3400 1237.1200 905.3400 1237.6000 ;
        RECT 913.1000 1237.1200 914.1000 1237.6000 ;
        RECT 902.3400 1231.6800 905.3400 1232.1600 ;
        RECT 913.1000 1231.6800 914.1000 1232.1600 ;
        RECT 902.3400 1436.5900 1139.3400 1439.5900 ;
        RECT 902.3400 1223.4900 1139.3400 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 993.8500 1094.1000 1209.9500 ;
        RECT 1048.1000 993.8500 1049.1000 1209.9500 ;
        RECT 1003.1000 993.8500 1004.1000 1209.9500 ;
        RECT 958.1000 993.8500 959.1000 1209.9500 ;
        RECT 913.1000 993.8500 914.1000 1209.9500 ;
        RECT 1136.3400 993.8500 1139.3400 1209.9500 ;
        RECT 902.3400 993.8500 905.3400 1209.9500 ;
      LAYER met3 ;
        RECT 1136.3400 1192.4400 1139.3400 1192.9200 ;
        RECT 1136.3400 1197.8800 1139.3400 1198.3600 ;
        RECT 1093.1000 1192.4400 1094.1000 1192.9200 ;
        RECT 1093.1000 1197.8800 1094.1000 1198.3600 ;
        RECT 1136.3400 1181.5600 1139.3400 1182.0400 ;
        RECT 1136.3400 1187.0000 1139.3400 1187.4800 ;
        RECT 1136.3400 1170.6800 1139.3400 1171.1600 ;
        RECT 1136.3400 1176.1200 1139.3400 1176.6000 ;
        RECT 1136.3400 1165.2400 1139.3400 1165.7200 ;
        RECT 1093.1000 1181.5600 1094.1000 1182.0400 ;
        RECT 1093.1000 1187.0000 1094.1000 1187.4800 ;
        RECT 1093.1000 1165.2400 1094.1000 1165.7200 ;
        RECT 1093.1000 1170.6800 1094.1000 1171.1600 ;
        RECT 1093.1000 1176.1200 1094.1000 1176.6000 ;
        RECT 1048.1000 1192.4400 1049.1000 1192.9200 ;
        RECT 1048.1000 1197.8800 1049.1000 1198.3600 ;
        RECT 1048.1000 1181.5600 1049.1000 1182.0400 ;
        RECT 1048.1000 1187.0000 1049.1000 1187.4800 ;
        RECT 1048.1000 1165.2400 1049.1000 1165.7200 ;
        RECT 1048.1000 1170.6800 1049.1000 1171.1600 ;
        RECT 1048.1000 1176.1200 1049.1000 1176.6000 ;
        RECT 1136.3400 1148.9200 1139.3400 1149.4000 ;
        RECT 1136.3400 1154.3600 1139.3400 1154.8400 ;
        RECT 1136.3400 1159.8000 1139.3400 1160.2800 ;
        RECT 1136.3400 1143.4800 1139.3400 1143.9600 ;
        RECT 1136.3400 1132.6000 1139.3400 1133.0800 ;
        RECT 1136.3400 1138.0400 1139.3400 1138.5200 ;
        RECT 1093.1000 1148.9200 1094.1000 1149.4000 ;
        RECT 1093.1000 1154.3600 1094.1000 1154.8400 ;
        RECT 1093.1000 1159.8000 1094.1000 1160.2800 ;
        RECT 1093.1000 1132.6000 1094.1000 1133.0800 ;
        RECT 1093.1000 1138.0400 1094.1000 1138.5200 ;
        RECT 1093.1000 1143.4800 1094.1000 1143.9600 ;
        RECT 1136.3400 1121.7200 1139.3400 1122.2000 ;
        RECT 1136.3400 1127.1600 1139.3400 1127.6400 ;
        RECT 1136.3400 1110.8400 1139.3400 1111.3200 ;
        RECT 1136.3400 1116.2800 1139.3400 1116.7600 ;
        RECT 1136.3400 1105.4000 1139.3400 1105.8800 ;
        RECT 1093.1000 1121.7200 1094.1000 1122.2000 ;
        RECT 1093.1000 1127.1600 1094.1000 1127.6400 ;
        RECT 1093.1000 1105.4000 1094.1000 1105.8800 ;
        RECT 1093.1000 1110.8400 1094.1000 1111.3200 ;
        RECT 1093.1000 1116.2800 1094.1000 1116.7600 ;
        RECT 1048.1000 1148.9200 1049.1000 1149.4000 ;
        RECT 1048.1000 1154.3600 1049.1000 1154.8400 ;
        RECT 1048.1000 1159.8000 1049.1000 1160.2800 ;
        RECT 1048.1000 1132.6000 1049.1000 1133.0800 ;
        RECT 1048.1000 1138.0400 1049.1000 1138.5200 ;
        RECT 1048.1000 1143.4800 1049.1000 1143.9600 ;
        RECT 1048.1000 1121.7200 1049.1000 1122.2000 ;
        RECT 1048.1000 1127.1600 1049.1000 1127.6400 ;
        RECT 1048.1000 1105.4000 1049.1000 1105.8800 ;
        RECT 1048.1000 1110.8400 1049.1000 1111.3200 ;
        RECT 1048.1000 1116.2800 1049.1000 1116.7600 ;
        RECT 1003.1000 1192.4400 1004.1000 1192.9200 ;
        RECT 1003.1000 1197.8800 1004.1000 1198.3600 ;
        RECT 1003.1000 1181.5600 1004.1000 1182.0400 ;
        RECT 1003.1000 1187.0000 1004.1000 1187.4800 ;
        RECT 1003.1000 1165.2400 1004.1000 1165.7200 ;
        RECT 1003.1000 1170.6800 1004.1000 1171.1600 ;
        RECT 1003.1000 1176.1200 1004.1000 1176.6000 ;
        RECT 958.1000 1192.4400 959.1000 1192.9200 ;
        RECT 958.1000 1197.8800 959.1000 1198.3600 ;
        RECT 913.1000 1197.8800 914.1000 1198.3600 ;
        RECT 913.1000 1192.4400 914.1000 1192.9200 ;
        RECT 902.3400 1197.8800 905.3400 1198.3600 ;
        RECT 902.3400 1192.4400 905.3400 1192.9200 ;
        RECT 958.1000 1181.5600 959.1000 1182.0400 ;
        RECT 958.1000 1187.0000 959.1000 1187.4800 ;
        RECT 958.1000 1165.2400 959.1000 1165.7200 ;
        RECT 958.1000 1170.6800 959.1000 1171.1600 ;
        RECT 958.1000 1176.1200 959.1000 1176.6000 ;
        RECT 902.3400 1187.0000 905.3400 1187.4800 ;
        RECT 913.1000 1187.0000 914.1000 1187.4800 ;
        RECT 902.3400 1181.5600 905.3400 1182.0400 ;
        RECT 913.1000 1181.5600 914.1000 1182.0400 ;
        RECT 913.1000 1176.1200 914.1000 1176.6000 ;
        RECT 913.1000 1170.6800 914.1000 1171.1600 ;
        RECT 902.3400 1176.1200 905.3400 1176.6000 ;
        RECT 902.3400 1170.6800 905.3400 1171.1600 ;
        RECT 902.3400 1165.2400 905.3400 1165.7200 ;
        RECT 913.1000 1165.2400 914.1000 1165.7200 ;
        RECT 1003.1000 1148.9200 1004.1000 1149.4000 ;
        RECT 1003.1000 1154.3600 1004.1000 1154.8400 ;
        RECT 1003.1000 1159.8000 1004.1000 1160.2800 ;
        RECT 1003.1000 1132.6000 1004.1000 1133.0800 ;
        RECT 1003.1000 1138.0400 1004.1000 1138.5200 ;
        RECT 1003.1000 1143.4800 1004.1000 1143.9600 ;
        RECT 1003.1000 1121.7200 1004.1000 1122.2000 ;
        RECT 1003.1000 1127.1600 1004.1000 1127.6400 ;
        RECT 1003.1000 1105.4000 1004.1000 1105.8800 ;
        RECT 1003.1000 1110.8400 1004.1000 1111.3200 ;
        RECT 1003.1000 1116.2800 1004.1000 1116.7600 ;
        RECT 958.1000 1148.9200 959.1000 1149.4000 ;
        RECT 958.1000 1154.3600 959.1000 1154.8400 ;
        RECT 958.1000 1159.8000 959.1000 1160.2800 ;
        RECT 958.1000 1132.6000 959.1000 1133.0800 ;
        RECT 958.1000 1138.0400 959.1000 1138.5200 ;
        RECT 958.1000 1143.4800 959.1000 1143.9600 ;
        RECT 902.3400 1159.8000 905.3400 1160.2800 ;
        RECT 913.1000 1159.8000 914.1000 1160.2800 ;
        RECT 902.3400 1148.9200 905.3400 1149.4000 ;
        RECT 913.1000 1148.9200 914.1000 1149.4000 ;
        RECT 902.3400 1154.3600 905.3400 1154.8400 ;
        RECT 913.1000 1154.3600 914.1000 1154.8400 ;
        RECT 902.3400 1143.4800 905.3400 1143.9600 ;
        RECT 913.1000 1143.4800 914.1000 1143.9600 ;
        RECT 913.1000 1138.0400 914.1000 1138.5200 ;
        RECT 913.1000 1132.6000 914.1000 1133.0800 ;
        RECT 902.3400 1138.0400 905.3400 1138.5200 ;
        RECT 902.3400 1132.6000 905.3400 1133.0800 ;
        RECT 958.1000 1121.7200 959.1000 1122.2000 ;
        RECT 958.1000 1127.1600 959.1000 1127.6400 ;
        RECT 958.1000 1105.4000 959.1000 1105.8800 ;
        RECT 958.1000 1110.8400 959.1000 1111.3200 ;
        RECT 958.1000 1116.2800 959.1000 1116.7600 ;
        RECT 902.3400 1127.1600 905.3400 1127.6400 ;
        RECT 913.1000 1127.1600 914.1000 1127.6400 ;
        RECT 902.3400 1121.7200 905.3400 1122.2000 ;
        RECT 913.1000 1121.7200 914.1000 1122.2000 ;
        RECT 913.1000 1116.2800 914.1000 1116.7600 ;
        RECT 913.1000 1110.8400 914.1000 1111.3200 ;
        RECT 902.3400 1116.2800 905.3400 1116.7600 ;
        RECT 902.3400 1110.8400 905.3400 1111.3200 ;
        RECT 902.3400 1105.4000 905.3400 1105.8800 ;
        RECT 913.1000 1105.4000 914.1000 1105.8800 ;
        RECT 1136.3400 1089.0800 1139.3400 1089.5600 ;
        RECT 1136.3400 1094.5200 1139.3400 1095.0000 ;
        RECT 1136.3400 1099.9600 1139.3400 1100.4400 ;
        RECT 1136.3400 1083.6400 1139.3400 1084.1200 ;
        RECT 1136.3400 1072.7600 1139.3400 1073.2400 ;
        RECT 1136.3400 1078.2000 1139.3400 1078.6800 ;
        RECT 1093.1000 1089.0800 1094.1000 1089.5600 ;
        RECT 1093.1000 1094.5200 1094.1000 1095.0000 ;
        RECT 1093.1000 1099.9600 1094.1000 1100.4400 ;
        RECT 1093.1000 1072.7600 1094.1000 1073.2400 ;
        RECT 1093.1000 1078.2000 1094.1000 1078.6800 ;
        RECT 1093.1000 1083.6400 1094.1000 1084.1200 ;
        RECT 1136.3400 1061.8800 1139.3400 1062.3600 ;
        RECT 1136.3400 1067.3200 1139.3400 1067.8000 ;
        RECT 1136.3400 1051.0000 1139.3400 1051.4800 ;
        RECT 1136.3400 1056.4400 1139.3400 1056.9200 ;
        RECT 1136.3400 1045.5600 1139.3400 1046.0400 ;
        RECT 1093.1000 1061.8800 1094.1000 1062.3600 ;
        RECT 1093.1000 1067.3200 1094.1000 1067.8000 ;
        RECT 1093.1000 1045.5600 1094.1000 1046.0400 ;
        RECT 1093.1000 1051.0000 1094.1000 1051.4800 ;
        RECT 1093.1000 1056.4400 1094.1000 1056.9200 ;
        RECT 1048.1000 1089.0800 1049.1000 1089.5600 ;
        RECT 1048.1000 1094.5200 1049.1000 1095.0000 ;
        RECT 1048.1000 1099.9600 1049.1000 1100.4400 ;
        RECT 1048.1000 1072.7600 1049.1000 1073.2400 ;
        RECT 1048.1000 1078.2000 1049.1000 1078.6800 ;
        RECT 1048.1000 1083.6400 1049.1000 1084.1200 ;
        RECT 1048.1000 1061.8800 1049.1000 1062.3600 ;
        RECT 1048.1000 1067.3200 1049.1000 1067.8000 ;
        RECT 1048.1000 1045.5600 1049.1000 1046.0400 ;
        RECT 1048.1000 1051.0000 1049.1000 1051.4800 ;
        RECT 1048.1000 1056.4400 1049.1000 1056.9200 ;
        RECT 1136.3400 1029.2400 1139.3400 1029.7200 ;
        RECT 1136.3400 1034.6800 1139.3400 1035.1600 ;
        RECT 1136.3400 1040.1200 1139.3400 1040.6000 ;
        RECT 1136.3400 1023.8000 1139.3400 1024.2800 ;
        RECT 1136.3400 1012.9200 1139.3400 1013.4000 ;
        RECT 1136.3400 1018.3600 1139.3400 1018.8400 ;
        RECT 1093.1000 1029.2400 1094.1000 1029.7200 ;
        RECT 1093.1000 1034.6800 1094.1000 1035.1600 ;
        RECT 1093.1000 1040.1200 1094.1000 1040.6000 ;
        RECT 1093.1000 1012.9200 1094.1000 1013.4000 ;
        RECT 1093.1000 1018.3600 1094.1000 1018.8400 ;
        RECT 1093.1000 1023.8000 1094.1000 1024.2800 ;
        RECT 1136.3400 1002.0400 1139.3400 1002.5200 ;
        RECT 1136.3400 1007.4800 1139.3400 1007.9600 ;
        RECT 1093.1000 1002.0400 1094.1000 1002.5200 ;
        RECT 1093.1000 1007.4800 1094.1000 1007.9600 ;
        RECT 1048.1000 1029.2400 1049.1000 1029.7200 ;
        RECT 1048.1000 1034.6800 1049.1000 1035.1600 ;
        RECT 1048.1000 1040.1200 1049.1000 1040.6000 ;
        RECT 1048.1000 1012.9200 1049.1000 1013.4000 ;
        RECT 1048.1000 1018.3600 1049.1000 1018.8400 ;
        RECT 1048.1000 1023.8000 1049.1000 1024.2800 ;
        RECT 1048.1000 1002.0400 1049.1000 1002.5200 ;
        RECT 1048.1000 1007.4800 1049.1000 1007.9600 ;
        RECT 1003.1000 1089.0800 1004.1000 1089.5600 ;
        RECT 1003.1000 1094.5200 1004.1000 1095.0000 ;
        RECT 1003.1000 1099.9600 1004.1000 1100.4400 ;
        RECT 1003.1000 1072.7600 1004.1000 1073.2400 ;
        RECT 1003.1000 1078.2000 1004.1000 1078.6800 ;
        RECT 1003.1000 1083.6400 1004.1000 1084.1200 ;
        RECT 1003.1000 1061.8800 1004.1000 1062.3600 ;
        RECT 1003.1000 1067.3200 1004.1000 1067.8000 ;
        RECT 1003.1000 1045.5600 1004.1000 1046.0400 ;
        RECT 1003.1000 1051.0000 1004.1000 1051.4800 ;
        RECT 1003.1000 1056.4400 1004.1000 1056.9200 ;
        RECT 958.1000 1089.0800 959.1000 1089.5600 ;
        RECT 958.1000 1094.5200 959.1000 1095.0000 ;
        RECT 958.1000 1099.9600 959.1000 1100.4400 ;
        RECT 958.1000 1072.7600 959.1000 1073.2400 ;
        RECT 958.1000 1078.2000 959.1000 1078.6800 ;
        RECT 958.1000 1083.6400 959.1000 1084.1200 ;
        RECT 902.3400 1099.9600 905.3400 1100.4400 ;
        RECT 913.1000 1099.9600 914.1000 1100.4400 ;
        RECT 902.3400 1089.0800 905.3400 1089.5600 ;
        RECT 913.1000 1089.0800 914.1000 1089.5600 ;
        RECT 902.3400 1094.5200 905.3400 1095.0000 ;
        RECT 913.1000 1094.5200 914.1000 1095.0000 ;
        RECT 902.3400 1083.6400 905.3400 1084.1200 ;
        RECT 913.1000 1083.6400 914.1000 1084.1200 ;
        RECT 913.1000 1078.2000 914.1000 1078.6800 ;
        RECT 913.1000 1072.7600 914.1000 1073.2400 ;
        RECT 902.3400 1078.2000 905.3400 1078.6800 ;
        RECT 902.3400 1072.7600 905.3400 1073.2400 ;
        RECT 958.1000 1061.8800 959.1000 1062.3600 ;
        RECT 958.1000 1067.3200 959.1000 1067.8000 ;
        RECT 958.1000 1045.5600 959.1000 1046.0400 ;
        RECT 958.1000 1051.0000 959.1000 1051.4800 ;
        RECT 958.1000 1056.4400 959.1000 1056.9200 ;
        RECT 902.3400 1067.3200 905.3400 1067.8000 ;
        RECT 913.1000 1067.3200 914.1000 1067.8000 ;
        RECT 902.3400 1061.8800 905.3400 1062.3600 ;
        RECT 913.1000 1061.8800 914.1000 1062.3600 ;
        RECT 913.1000 1056.4400 914.1000 1056.9200 ;
        RECT 913.1000 1051.0000 914.1000 1051.4800 ;
        RECT 902.3400 1056.4400 905.3400 1056.9200 ;
        RECT 902.3400 1051.0000 905.3400 1051.4800 ;
        RECT 902.3400 1045.5600 905.3400 1046.0400 ;
        RECT 913.1000 1045.5600 914.1000 1046.0400 ;
        RECT 1003.1000 1029.2400 1004.1000 1029.7200 ;
        RECT 1003.1000 1034.6800 1004.1000 1035.1600 ;
        RECT 1003.1000 1040.1200 1004.1000 1040.6000 ;
        RECT 1003.1000 1012.9200 1004.1000 1013.4000 ;
        RECT 1003.1000 1018.3600 1004.1000 1018.8400 ;
        RECT 1003.1000 1023.8000 1004.1000 1024.2800 ;
        RECT 1003.1000 1002.0400 1004.1000 1002.5200 ;
        RECT 1003.1000 1007.4800 1004.1000 1007.9600 ;
        RECT 958.1000 1029.2400 959.1000 1029.7200 ;
        RECT 958.1000 1034.6800 959.1000 1035.1600 ;
        RECT 958.1000 1040.1200 959.1000 1040.6000 ;
        RECT 958.1000 1012.9200 959.1000 1013.4000 ;
        RECT 958.1000 1018.3600 959.1000 1018.8400 ;
        RECT 958.1000 1023.8000 959.1000 1024.2800 ;
        RECT 902.3400 1040.1200 905.3400 1040.6000 ;
        RECT 913.1000 1040.1200 914.1000 1040.6000 ;
        RECT 902.3400 1029.2400 905.3400 1029.7200 ;
        RECT 913.1000 1029.2400 914.1000 1029.7200 ;
        RECT 902.3400 1034.6800 905.3400 1035.1600 ;
        RECT 913.1000 1034.6800 914.1000 1035.1600 ;
        RECT 902.3400 1023.8000 905.3400 1024.2800 ;
        RECT 913.1000 1023.8000 914.1000 1024.2800 ;
        RECT 913.1000 1018.3600 914.1000 1018.8400 ;
        RECT 913.1000 1012.9200 914.1000 1013.4000 ;
        RECT 902.3400 1018.3600 905.3400 1018.8400 ;
        RECT 902.3400 1012.9200 905.3400 1013.4000 ;
        RECT 958.1000 1002.0400 959.1000 1002.5200 ;
        RECT 958.1000 1007.4800 959.1000 1007.9600 ;
        RECT 902.3400 1007.4800 905.3400 1007.9600 ;
        RECT 913.1000 1007.4800 914.1000 1007.9600 ;
        RECT 902.3400 1002.0400 905.3400 1002.5200 ;
        RECT 913.1000 1002.0400 914.1000 1002.5200 ;
        RECT 902.3400 1206.9500 1139.3400 1209.9500 ;
        RECT 902.3400 993.8500 1139.3400 996.8500 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'RegFile'
    PORT
      LAYER met4 ;
        RECT 1093.1000 764.2100 1094.1000 980.3100 ;
        RECT 1048.1000 764.2100 1049.1000 980.3100 ;
        RECT 1003.1000 764.2100 1004.1000 980.3100 ;
        RECT 958.1000 764.2100 959.1000 980.3100 ;
        RECT 913.1000 764.2100 914.1000 980.3100 ;
        RECT 1136.3400 764.2100 1139.3400 980.3100 ;
        RECT 902.3400 764.2100 905.3400 980.3100 ;
      LAYER met3 ;
        RECT 1136.3400 962.8000 1139.3400 963.2800 ;
        RECT 1136.3400 968.2400 1139.3400 968.7200 ;
        RECT 1093.1000 962.8000 1094.1000 963.2800 ;
        RECT 1093.1000 968.2400 1094.1000 968.7200 ;
        RECT 1136.3400 951.9200 1139.3400 952.4000 ;
        RECT 1136.3400 957.3600 1139.3400 957.8400 ;
        RECT 1136.3400 941.0400 1139.3400 941.5200 ;
        RECT 1136.3400 946.4800 1139.3400 946.9600 ;
        RECT 1136.3400 935.6000 1139.3400 936.0800 ;
        RECT 1093.1000 951.9200 1094.1000 952.4000 ;
        RECT 1093.1000 957.3600 1094.1000 957.8400 ;
        RECT 1093.1000 935.6000 1094.1000 936.0800 ;
        RECT 1093.1000 941.0400 1094.1000 941.5200 ;
        RECT 1093.1000 946.4800 1094.1000 946.9600 ;
        RECT 1048.1000 962.8000 1049.1000 963.2800 ;
        RECT 1048.1000 968.2400 1049.1000 968.7200 ;
        RECT 1048.1000 951.9200 1049.1000 952.4000 ;
        RECT 1048.1000 957.3600 1049.1000 957.8400 ;
        RECT 1048.1000 935.6000 1049.1000 936.0800 ;
        RECT 1048.1000 941.0400 1049.1000 941.5200 ;
        RECT 1048.1000 946.4800 1049.1000 946.9600 ;
        RECT 1136.3400 919.2800 1139.3400 919.7600 ;
        RECT 1136.3400 924.7200 1139.3400 925.2000 ;
        RECT 1136.3400 930.1600 1139.3400 930.6400 ;
        RECT 1136.3400 913.8400 1139.3400 914.3200 ;
        RECT 1136.3400 902.9600 1139.3400 903.4400 ;
        RECT 1136.3400 908.4000 1139.3400 908.8800 ;
        RECT 1093.1000 919.2800 1094.1000 919.7600 ;
        RECT 1093.1000 924.7200 1094.1000 925.2000 ;
        RECT 1093.1000 930.1600 1094.1000 930.6400 ;
        RECT 1093.1000 902.9600 1094.1000 903.4400 ;
        RECT 1093.1000 908.4000 1094.1000 908.8800 ;
        RECT 1093.1000 913.8400 1094.1000 914.3200 ;
        RECT 1136.3400 892.0800 1139.3400 892.5600 ;
        RECT 1136.3400 897.5200 1139.3400 898.0000 ;
        RECT 1136.3400 881.2000 1139.3400 881.6800 ;
        RECT 1136.3400 886.6400 1139.3400 887.1200 ;
        RECT 1136.3400 875.7600 1139.3400 876.2400 ;
        RECT 1093.1000 892.0800 1094.1000 892.5600 ;
        RECT 1093.1000 897.5200 1094.1000 898.0000 ;
        RECT 1093.1000 875.7600 1094.1000 876.2400 ;
        RECT 1093.1000 881.2000 1094.1000 881.6800 ;
        RECT 1093.1000 886.6400 1094.1000 887.1200 ;
        RECT 1048.1000 919.2800 1049.1000 919.7600 ;
        RECT 1048.1000 924.7200 1049.1000 925.2000 ;
        RECT 1048.1000 930.1600 1049.1000 930.6400 ;
        RECT 1048.1000 902.9600 1049.1000 903.4400 ;
        RECT 1048.1000 908.4000 1049.1000 908.8800 ;
        RECT 1048.1000 913.8400 1049.1000 914.3200 ;
        RECT 1048.1000 892.0800 1049.1000 892.5600 ;
        RECT 1048.1000 897.5200 1049.1000 898.0000 ;
        RECT 1048.1000 875.7600 1049.1000 876.2400 ;
        RECT 1048.1000 881.2000 1049.1000 881.6800 ;
        RECT 1048.1000 886.6400 1049.1000 887.1200 ;
        RECT 1003.1000 962.8000 1004.1000 963.2800 ;
        RECT 1003.1000 968.2400 1004.1000 968.7200 ;
        RECT 1003.1000 951.9200 1004.1000 952.4000 ;
        RECT 1003.1000 957.3600 1004.1000 957.8400 ;
        RECT 1003.1000 935.6000 1004.1000 936.0800 ;
        RECT 1003.1000 941.0400 1004.1000 941.5200 ;
        RECT 1003.1000 946.4800 1004.1000 946.9600 ;
        RECT 958.1000 962.8000 959.1000 963.2800 ;
        RECT 958.1000 968.2400 959.1000 968.7200 ;
        RECT 913.1000 968.2400 914.1000 968.7200 ;
        RECT 913.1000 962.8000 914.1000 963.2800 ;
        RECT 902.3400 968.2400 905.3400 968.7200 ;
        RECT 902.3400 962.8000 905.3400 963.2800 ;
        RECT 958.1000 951.9200 959.1000 952.4000 ;
        RECT 958.1000 957.3600 959.1000 957.8400 ;
        RECT 958.1000 935.6000 959.1000 936.0800 ;
        RECT 958.1000 941.0400 959.1000 941.5200 ;
        RECT 958.1000 946.4800 959.1000 946.9600 ;
        RECT 902.3400 957.3600 905.3400 957.8400 ;
        RECT 913.1000 957.3600 914.1000 957.8400 ;
        RECT 902.3400 951.9200 905.3400 952.4000 ;
        RECT 913.1000 951.9200 914.1000 952.4000 ;
        RECT 913.1000 946.4800 914.1000 946.9600 ;
        RECT 913.1000 941.0400 914.1000 941.5200 ;
        RECT 902.3400 946.4800 905.3400 946.9600 ;
        RECT 902.3400 941.0400 905.3400 941.5200 ;
        RECT 902.3400 935.6000 905.3400 936.0800 ;
        RECT 913.1000 935.6000 914.1000 936.0800 ;
        RECT 1003.1000 919.2800 1004.1000 919.7600 ;
        RECT 1003.1000 924.7200 1004.1000 925.2000 ;
        RECT 1003.1000 930.1600 1004.1000 930.6400 ;
        RECT 1003.1000 902.9600 1004.1000 903.4400 ;
        RECT 1003.1000 908.4000 1004.1000 908.8800 ;
        RECT 1003.1000 913.8400 1004.1000 914.3200 ;
        RECT 1003.1000 892.0800 1004.1000 892.5600 ;
        RECT 1003.1000 897.5200 1004.1000 898.0000 ;
        RECT 1003.1000 875.7600 1004.1000 876.2400 ;
        RECT 1003.1000 881.2000 1004.1000 881.6800 ;
        RECT 1003.1000 886.6400 1004.1000 887.1200 ;
        RECT 958.1000 919.2800 959.1000 919.7600 ;
        RECT 958.1000 924.7200 959.1000 925.2000 ;
        RECT 958.1000 930.1600 959.1000 930.6400 ;
        RECT 958.1000 902.9600 959.1000 903.4400 ;
        RECT 958.1000 908.4000 959.1000 908.8800 ;
        RECT 958.1000 913.8400 959.1000 914.3200 ;
        RECT 902.3400 930.1600 905.3400 930.6400 ;
        RECT 913.1000 930.1600 914.1000 930.6400 ;
        RECT 902.3400 919.2800 905.3400 919.7600 ;
        RECT 913.1000 919.2800 914.1000 919.7600 ;
        RECT 902.3400 924.7200 905.3400 925.2000 ;
        RECT 913.1000 924.7200 914.1000 925.2000 ;
        RECT 902.3400 913.8400 905.3400 914.3200 ;
        RECT 913.1000 913.8400 914.1000 914.3200 ;
        RECT 913.1000 908.4000 914.1000 908.8800 ;
        RECT 913.1000 902.9600 914.1000 903.4400 ;
        RECT 902.3400 908.4000 905.3400 908.8800 ;
        RECT 902.3400 902.9600 905.3400 903.4400 ;
        RECT 958.1000 892.0800 959.1000 892.5600 ;
        RECT 958.1000 897.5200 959.1000 898.0000 ;
        RECT 958.1000 875.7600 959.1000 876.2400 ;
        RECT 958.1000 881.2000 959.1000 881.6800 ;
        RECT 958.1000 886.6400 959.1000 887.1200 ;
        RECT 902.3400 897.5200 905.3400 898.0000 ;
        RECT 913.1000 897.5200 914.1000 898.0000 ;
        RECT 902.3400 892.0800 905.3400 892.5600 ;
        RECT 913.1000 892.0800 914.1000 892.5600 ;
        RECT 913.1000 886.6400 914.1000 887.1200 ;
        RECT 913.1000 881.2000 914.1000 881.6800 ;
        RECT 902.3400 886.6400 905.3400 887.1200 ;
        RECT 902.3400 881.2000 905.3400 881.6800 ;
        RECT 902.3400 875.7600 905.3400 876.2400 ;
        RECT 913.1000 875.7600 914.1000 876.2400 ;
        RECT 1136.3400 859.4400 1139.3400 859.9200 ;
        RECT 1136.3400 864.8800 1139.3400 865.3600 ;
        RECT 1136.3400 870.3200 1139.3400 870.8000 ;
        RECT 1136.3400 854.0000 1139.3400 854.4800 ;
        RECT 1136.3400 843.1200 1139.3400 843.6000 ;
        RECT 1136.3400 848.5600 1139.3400 849.0400 ;
        RECT 1093.1000 859.4400 1094.1000 859.9200 ;
        RECT 1093.1000 864.8800 1094.1000 865.3600 ;
        RECT 1093.1000 870.3200 1094.1000 870.8000 ;
        RECT 1093.1000 843.1200 1094.1000 843.6000 ;
        RECT 1093.1000 848.5600 1094.1000 849.0400 ;
        RECT 1093.1000 854.0000 1094.1000 854.4800 ;
        RECT 1136.3400 832.2400 1139.3400 832.7200 ;
        RECT 1136.3400 837.6800 1139.3400 838.1600 ;
        RECT 1136.3400 821.3600 1139.3400 821.8400 ;
        RECT 1136.3400 826.8000 1139.3400 827.2800 ;
        RECT 1136.3400 815.9200 1139.3400 816.4000 ;
        RECT 1093.1000 832.2400 1094.1000 832.7200 ;
        RECT 1093.1000 837.6800 1094.1000 838.1600 ;
        RECT 1093.1000 815.9200 1094.1000 816.4000 ;
        RECT 1093.1000 821.3600 1094.1000 821.8400 ;
        RECT 1093.1000 826.8000 1094.1000 827.2800 ;
        RECT 1048.1000 859.4400 1049.1000 859.9200 ;
        RECT 1048.1000 864.8800 1049.1000 865.3600 ;
        RECT 1048.1000 870.3200 1049.1000 870.8000 ;
        RECT 1048.1000 843.1200 1049.1000 843.6000 ;
        RECT 1048.1000 848.5600 1049.1000 849.0400 ;
        RECT 1048.1000 854.0000 1049.1000 854.4800 ;
        RECT 1048.1000 832.2400 1049.1000 832.7200 ;
        RECT 1048.1000 837.6800 1049.1000 838.1600 ;
        RECT 1048.1000 815.9200 1049.1000 816.4000 ;
        RECT 1048.1000 821.3600 1049.1000 821.8400 ;
        RECT 1048.1000 826.8000 1049.1000 827.2800 ;
        RECT 1136.3400 799.6000 1139.3400 800.0800 ;
        RECT 1136.3400 805.0400 1139.3400 805.5200 ;
        RECT 1136.3400 810.4800 1139.3400 810.9600 ;
        RECT 1136.3400 794.1600 1139.3400 794.6400 ;
        RECT 1136.3400 783.2800 1139.3400 783.7600 ;
        RECT 1136.3400 788.7200 1139.3400 789.2000 ;
        RECT 1093.1000 799.6000 1094.1000 800.0800 ;
        RECT 1093.1000 805.0400 1094.1000 805.5200 ;
        RECT 1093.1000 810.4800 1094.1000 810.9600 ;
        RECT 1093.1000 783.2800 1094.1000 783.7600 ;
        RECT 1093.1000 788.7200 1094.1000 789.2000 ;
        RECT 1093.1000 794.1600 1094.1000 794.6400 ;
        RECT 1136.3400 772.4000 1139.3400 772.8800 ;
        RECT 1136.3400 777.8400 1139.3400 778.3200 ;
        RECT 1093.1000 772.4000 1094.1000 772.8800 ;
        RECT 1093.1000 777.8400 1094.1000 778.3200 ;
        RECT 1048.1000 799.6000 1049.1000 800.0800 ;
        RECT 1048.1000 805.0400 1049.1000 805.5200 ;
        RECT 1048.1000 810.4800 1049.1000 810.9600 ;
        RECT 1048.1000 783.2800 1049.1000 783.7600 ;
        RECT 1048.1000 788.7200 1049.1000 789.2000 ;
        RECT 1048.1000 794.1600 1049.1000 794.6400 ;
        RECT 1048.1000 772.4000 1049.1000 772.8800 ;
        RECT 1048.1000 777.8400 1049.1000 778.3200 ;
        RECT 1003.1000 859.4400 1004.1000 859.9200 ;
        RECT 1003.1000 864.8800 1004.1000 865.3600 ;
        RECT 1003.1000 870.3200 1004.1000 870.8000 ;
        RECT 1003.1000 843.1200 1004.1000 843.6000 ;
        RECT 1003.1000 848.5600 1004.1000 849.0400 ;
        RECT 1003.1000 854.0000 1004.1000 854.4800 ;
        RECT 1003.1000 832.2400 1004.1000 832.7200 ;
        RECT 1003.1000 837.6800 1004.1000 838.1600 ;
        RECT 1003.1000 815.9200 1004.1000 816.4000 ;
        RECT 1003.1000 821.3600 1004.1000 821.8400 ;
        RECT 1003.1000 826.8000 1004.1000 827.2800 ;
        RECT 958.1000 859.4400 959.1000 859.9200 ;
        RECT 958.1000 864.8800 959.1000 865.3600 ;
        RECT 958.1000 870.3200 959.1000 870.8000 ;
        RECT 958.1000 843.1200 959.1000 843.6000 ;
        RECT 958.1000 848.5600 959.1000 849.0400 ;
        RECT 958.1000 854.0000 959.1000 854.4800 ;
        RECT 902.3400 870.3200 905.3400 870.8000 ;
        RECT 913.1000 870.3200 914.1000 870.8000 ;
        RECT 902.3400 859.4400 905.3400 859.9200 ;
        RECT 913.1000 859.4400 914.1000 859.9200 ;
        RECT 902.3400 864.8800 905.3400 865.3600 ;
        RECT 913.1000 864.8800 914.1000 865.3600 ;
        RECT 902.3400 854.0000 905.3400 854.4800 ;
        RECT 913.1000 854.0000 914.1000 854.4800 ;
        RECT 913.1000 848.5600 914.1000 849.0400 ;
        RECT 913.1000 843.1200 914.1000 843.6000 ;
        RECT 902.3400 848.5600 905.3400 849.0400 ;
        RECT 902.3400 843.1200 905.3400 843.6000 ;
        RECT 958.1000 832.2400 959.1000 832.7200 ;
        RECT 958.1000 837.6800 959.1000 838.1600 ;
        RECT 958.1000 815.9200 959.1000 816.4000 ;
        RECT 958.1000 821.3600 959.1000 821.8400 ;
        RECT 958.1000 826.8000 959.1000 827.2800 ;
        RECT 902.3400 837.6800 905.3400 838.1600 ;
        RECT 913.1000 837.6800 914.1000 838.1600 ;
        RECT 902.3400 832.2400 905.3400 832.7200 ;
        RECT 913.1000 832.2400 914.1000 832.7200 ;
        RECT 913.1000 826.8000 914.1000 827.2800 ;
        RECT 913.1000 821.3600 914.1000 821.8400 ;
        RECT 902.3400 826.8000 905.3400 827.2800 ;
        RECT 902.3400 821.3600 905.3400 821.8400 ;
        RECT 902.3400 815.9200 905.3400 816.4000 ;
        RECT 913.1000 815.9200 914.1000 816.4000 ;
        RECT 1003.1000 799.6000 1004.1000 800.0800 ;
        RECT 1003.1000 805.0400 1004.1000 805.5200 ;
        RECT 1003.1000 810.4800 1004.1000 810.9600 ;
        RECT 1003.1000 783.2800 1004.1000 783.7600 ;
        RECT 1003.1000 788.7200 1004.1000 789.2000 ;
        RECT 1003.1000 794.1600 1004.1000 794.6400 ;
        RECT 1003.1000 772.4000 1004.1000 772.8800 ;
        RECT 1003.1000 777.8400 1004.1000 778.3200 ;
        RECT 958.1000 799.6000 959.1000 800.0800 ;
        RECT 958.1000 805.0400 959.1000 805.5200 ;
        RECT 958.1000 810.4800 959.1000 810.9600 ;
        RECT 958.1000 783.2800 959.1000 783.7600 ;
        RECT 958.1000 788.7200 959.1000 789.2000 ;
        RECT 958.1000 794.1600 959.1000 794.6400 ;
        RECT 902.3400 810.4800 905.3400 810.9600 ;
        RECT 913.1000 810.4800 914.1000 810.9600 ;
        RECT 902.3400 799.6000 905.3400 800.0800 ;
        RECT 913.1000 799.6000 914.1000 800.0800 ;
        RECT 902.3400 805.0400 905.3400 805.5200 ;
        RECT 913.1000 805.0400 914.1000 805.5200 ;
        RECT 902.3400 794.1600 905.3400 794.6400 ;
        RECT 913.1000 794.1600 914.1000 794.6400 ;
        RECT 913.1000 788.7200 914.1000 789.2000 ;
        RECT 913.1000 783.2800 914.1000 783.7600 ;
        RECT 902.3400 788.7200 905.3400 789.2000 ;
        RECT 902.3400 783.2800 905.3400 783.7600 ;
        RECT 958.1000 772.4000 959.1000 772.8800 ;
        RECT 958.1000 777.8400 959.1000 778.3200 ;
        RECT 902.3400 777.8400 905.3400 778.3200 ;
        RECT 913.1000 777.8400 914.1000 778.3200 ;
        RECT 902.3400 772.4000 905.3400 772.8800 ;
        RECT 913.1000 772.4000 914.1000 772.8800 ;
        RECT 902.3400 977.3100 1139.3400 980.3100 ;
        RECT 902.3400 764.2100 1139.3400 767.2100 ;
    END
# end of P/G pin shape extracted from block 'RegFile'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1153.4600 2830.6100 1155.4600 2857.5400 ;
        RECT 1356.5600 2830.6100 1358.5600 2857.5400 ;
      LAYER met3 ;
        RECT 1356.5600 2847.3200 1358.5600 2847.8000 ;
        RECT 1153.4600 2847.3200 1155.4600 2847.8000 ;
        RECT 1356.5600 2841.8800 1358.5600 2842.3600 ;
        RECT 1356.5600 2836.4400 1358.5600 2836.9200 ;
        RECT 1153.4600 2841.8800 1155.4600 2842.3600 ;
        RECT 1153.4600 2836.4400 1155.4600 2836.9200 ;
        RECT 1153.4600 2855.5400 1358.5600 2857.5400 ;
        RECT 1153.4600 2830.6100 1358.5600 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 534.5700 1345.8200 750.6700 ;
        RECT 1299.2200 534.5700 1300.8200 750.6700 ;
        RECT 1254.2200 534.5700 1255.8200 750.6700 ;
        RECT 1209.2200 534.5700 1210.8200 750.6700 ;
        RECT 1164.2200 534.5700 1165.8200 750.6700 ;
        RECT 1356.5600 534.5700 1359.5600 750.6700 ;
        RECT 1152.4600 534.5700 1155.4600 750.6700 ;
      LAYER met3 ;
        RECT 1356.5600 727.7200 1359.5600 728.2000 ;
        RECT 1356.5600 733.1600 1359.5600 733.6400 ;
        RECT 1344.2200 727.7200 1345.8200 728.2000 ;
        RECT 1344.2200 733.1600 1345.8200 733.6400 ;
        RECT 1356.5600 738.6000 1359.5600 739.0800 ;
        RECT 1344.2200 738.6000 1345.8200 739.0800 ;
        RECT 1356.5600 716.8400 1359.5600 717.3200 ;
        RECT 1356.5600 722.2800 1359.5600 722.7600 ;
        RECT 1344.2200 716.8400 1345.8200 717.3200 ;
        RECT 1344.2200 722.2800 1345.8200 722.7600 ;
        RECT 1356.5600 700.5200 1359.5600 701.0000 ;
        RECT 1356.5600 705.9600 1359.5600 706.4400 ;
        RECT 1344.2200 700.5200 1345.8200 701.0000 ;
        RECT 1344.2200 705.9600 1345.8200 706.4400 ;
        RECT 1356.5600 711.4000 1359.5600 711.8800 ;
        RECT 1344.2200 711.4000 1345.8200 711.8800 ;
        RECT 1299.2200 727.7200 1300.8200 728.2000 ;
        RECT 1299.2200 733.1600 1300.8200 733.6400 ;
        RECT 1299.2200 738.6000 1300.8200 739.0800 ;
        RECT 1299.2200 716.8400 1300.8200 717.3200 ;
        RECT 1299.2200 722.2800 1300.8200 722.7600 ;
        RECT 1299.2200 700.5200 1300.8200 701.0000 ;
        RECT 1299.2200 705.9600 1300.8200 706.4400 ;
        RECT 1299.2200 711.4000 1300.8200 711.8800 ;
        RECT 1356.5600 684.2000 1359.5600 684.6800 ;
        RECT 1356.5600 689.6400 1359.5600 690.1200 ;
        RECT 1356.5600 695.0800 1359.5600 695.5600 ;
        RECT 1344.2200 684.2000 1345.8200 684.6800 ;
        RECT 1344.2200 689.6400 1345.8200 690.1200 ;
        RECT 1344.2200 695.0800 1345.8200 695.5600 ;
        RECT 1356.5600 673.3200 1359.5600 673.8000 ;
        RECT 1356.5600 678.7600 1359.5600 679.2400 ;
        RECT 1344.2200 673.3200 1345.8200 673.8000 ;
        RECT 1344.2200 678.7600 1345.8200 679.2400 ;
        RECT 1356.5600 657.0000 1359.5600 657.4800 ;
        RECT 1356.5600 662.4400 1359.5600 662.9200 ;
        RECT 1356.5600 667.8800 1359.5600 668.3600 ;
        RECT 1344.2200 657.0000 1345.8200 657.4800 ;
        RECT 1344.2200 662.4400 1345.8200 662.9200 ;
        RECT 1344.2200 667.8800 1345.8200 668.3600 ;
        RECT 1356.5600 646.1200 1359.5600 646.6000 ;
        RECT 1356.5600 651.5600 1359.5600 652.0400 ;
        RECT 1344.2200 646.1200 1345.8200 646.6000 ;
        RECT 1344.2200 651.5600 1345.8200 652.0400 ;
        RECT 1299.2200 684.2000 1300.8200 684.6800 ;
        RECT 1299.2200 689.6400 1300.8200 690.1200 ;
        RECT 1299.2200 695.0800 1300.8200 695.5600 ;
        RECT 1299.2200 673.3200 1300.8200 673.8000 ;
        RECT 1299.2200 678.7600 1300.8200 679.2400 ;
        RECT 1299.2200 657.0000 1300.8200 657.4800 ;
        RECT 1299.2200 662.4400 1300.8200 662.9200 ;
        RECT 1299.2200 667.8800 1300.8200 668.3600 ;
        RECT 1299.2200 646.1200 1300.8200 646.6000 ;
        RECT 1299.2200 651.5600 1300.8200 652.0400 ;
        RECT 1254.2200 727.7200 1255.8200 728.2000 ;
        RECT 1254.2200 733.1600 1255.8200 733.6400 ;
        RECT 1254.2200 738.6000 1255.8200 739.0800 ;
        RECT 1209.2200 727.7200 1210.8200 728.2000 ;
        RECT 1209.2200 733.1600 1210.8200 733.6400 ;
        RECT 1209.2200 738.6000 1210.8200 739.0800 ;
        RECT 1254.2200 716.8400 1255.8200 717.3200 ;
        RECT 1254.2200 722.2800 1255.8200 722.7600 ;
        RECT 1254.2200 700.5200 1255.8200 701.0000 ;
        RECT 1254.2200 705.9600 1255.8200 706.4400 ;
        RECT 1254.2200 711.4000 1255.8200 711.8800 ;
        RECT 1209.2200 716.8400 1210.8200 717.3200 ;
        RECT 1209.2200 722.2800 1210.8200 722.7600 ;
        RECT 1209.2200 700.5200 1210.8200 701.0000 ;
        RECT 1209.2200 705.9600 1210.8200 706.4400 ;
        RECT 1209.2200 711.4000 1210.8200 711.8800 ;
        RECT 1164.2200 727.7200 1165.8200 728.2000 ;
        RECT 1164.2200 733.1600 1165.8200 733.6400 ;
        RECT 1152.4600 733.1600 1155.4600 733.6400 ;
        RECT 1152.4600 727.7200 1155.4600 728.2000 ;
        RECT 1152.4600 738.6000 1155.4600 739.0800 ;
        RECT 1164.2200 738.6000 1165.8200 739.0800 ;
        RECT 1164.2200 716.8400 1165.8200 717.3200 ;
        RECT 1164.2200 722.2800 1165.8200 722.7600 ;
        RECT 1152.4600 722.2800 1155.4600 722.7600 ;
        RECT 1152.4600 716.8400 1155.4600 717.3200 ;
        RECT 1164.2200 700.5200 1165.8200 701.0000 ;
        RECT 1164.2200 705.9600 1165.8200 706.4400 ;
        RECT 1152.4600 705.9600 1155.4600 706.4400 ;
        RECT 1152.4600 700.5200 1155.4600 701.0000 ;
        RECT 1152.4600 711.4000 1155.4600 711.8800 ;
        RECT 1164.2200 711.4000 1165.8200 711.8800 ;
        RECT 1254.2200 684.2000 1255.8200 684.6800 ;
        RECT 1254.2200 689.6400 1255.8200 690.1200 ;
        RECT 1254.2200 695.0800 1255.8200 695.5600 ;
        RECT 1254.2200 673.3200 1255.8200 673.8000 ;
        RECT 1254.2200 678.7600 1255.8200 679.2400 ;
        RECT 1209.2200 684.2000 1210.8200 684.6800 ;
        RECT 1209.2200 689.6400 1210.8200 690.1200 ;
        RECT 1209.2200 695.0800 1210.8200 695.5600 ;
        RECT 1209.2200 673.3200 1210.8200 673.8000 ;
        RECT 1209.2200 678.7600 1210.8200 679.2400 ;
        RECT 1254.2200 657.0000 1255.8200 657.4800 ;
        RECT 1254.2200 662.4400 1255.8200 662.9200 ;
        RECT 1254.2200 667.8800 1255.8200 668.3600 ;
        RECT 1254.2200 646.1200 1255.8200 646.6000 ;
        RECT 1254.2200 651.5600 1255.8200 652.0400 ;
        RECT 1209.2200 657.0000 1210.8200 657.4800 ;
        RECT 1209.2200 662.4400 1210.8200 662.9200 ;
        RECT 1209.2200 667.8800 1210.8200 668.3600 ;
        RECT 1209.2200 646.1200 1210.8200 646.6000 ;
        RECT 1209.2200 651.5600 1210.8200 652.0400 ;
        RECT 1164.2200 684.2000 1165.8200 684.6800 ;
        RECT 1164.2200 689.6400 1165.8200 690.1200 ;
        RECT 1164.2200 695.0800 1165.8200 695.5600 ;
        RECT 1152.4600 684.2000 1155.4600 684.6800 ;
        RECT 1152.4600 689.6400 1155.4600 690.1200 ;
        RECT 1152.4600 695.0800 1155.4600 695.5600 ;
        RECT 1164.2200 673.3200 1165.8200 673.8000 ;
        RECT 1164.2200 678.7600 1165.8200 679.2400 ;
        RECT 1152.4600 673.3200 1155.4600 673.8000 ;
        RECT 1152.4600 678.7600 1155.4600 679.2400 ;
        RECT 1164.2200 657.0000 1165.8200 657.4800 ;
        RECT 1164.2200 662.4400 1165.8200 662.9200 ;
        RECT 1164.2200 667.8800 1165.8200 668.3600 ;
        RECT 1152.4600 657.0000 1155.4600 657.4800 ;
        RECT 1152.4600 662.4400 1155.4600 662.9200 ;
        RECT 1152.4600 667.8800 1155.4600 668.3600 ;
        RECT 1164.2200 646.1200 1165.8200 646.6000 ;
        RECT 1164.2200 651.5600 1165.8200 652.0400 ;
        RECT 1152.4600 646.1200 1155.4600 646.6000 ;
        RECT 1152.4600 651.5600 1155.4600 652.0400 ;
        RECT 1356.5600 629.8000 1359.5600 630.2800 ;
        RECT 1356.5600 635.2400 1359.5600 635.7200 ;
        RECT 1356.5600 640.6800 1359.5600 641.1600 ;
        RECT 1344.2200 629.8000 1345.8200 630.2800 ;
        RECT 1344.2200 635.2400 1345.8200 635.7200 ;
        RECT 1344.2200 640.6800 1345.8200 641.1600 ;
        RECT 1356.5600 618.9200 1359.5600 619.4000 ;
        RECT 1356.5600 624.3600 1359.5600 624.8400 ;
        RECT 1344.2200 618.9200 1345.8200 619.4000 ;
        RECT 1344.2200 624.3600 1345.8200 624.8400 ;
        RECT 1356.5600 602.6000 1359.5600 603.0800 ;
        RECT 1356.5600 608.0400 1359.5600 608.5200 ;
        RECT 1356.5600 613.4800 1359.5600 613.9600 ;
        RECT 1344.2200 602.6000 1345.8200 603.0800 ;
        RECT 1344.2200 608.0400 1345.8200 608.5200 ;
        RECT 1344.2200 613.4800 1345.8200 613.9600 ;
        RECT 1356.5600 591.7200 1359.5600 592.2000 ;
        RECT 1356.5600 597.1600 1359.5600 597.6400 ;
        RECT 1344.2200 591.7200 1345.8200 592.2000 ;
        RECT 1344.2200 597.1600 1345.8200 597.6400 ;
        RECT 1299.2200 629.8000 1300.8200 630.2800 ;
        RECT 1299.2200 635.2400 1300.8200 635.7200 ;
        RECT 1299.2200 640.6800 1300.8200 641.1600 ;
        RECT 1299.2200 618.9200 1300.8200 619.4000 ;
        RECT 1299.2200 624.3600 1300.8200 624.8400 ;
        RECT 1299.2200 602.6000 1300.8200 603.0800 ;
        RECT 1299.2200 608.0400 1300.8200 608.5200 ;
        RECT 1299.2200 613.4800 1300.8200 613.9600 ;
        RECT 1299.2200 591.7200 1300.8200 592.2000 ;
        RECT 1299.2200 597.1600 1300.8200 597.6400 ;
        RECT 1356.5600 575.4000 1359.5600 575.8800 ;
        RECT 1356.5600 580.8400 1359.5600 581.3200 ;
        RECT 1356.5600 586.2800 1359.5600 586.7600 ;
        RECT 1344.2200 575.4000 1345.8200 575.8800 ;
        RECT 1344.2200 580.8400 1345.8200 581.3200 ;
        RECT 1344.2200 586.2800 1345.8200 586.7600 ;
        RECT 1356.5600 564.5200 1359.5600 565.0000 ;
        RECT 1356.5600 569.9600 1359.5600 570.4400 ;
        RECT 1344.2200 564.5200 1345.8200 565.0000 ;
        RECT 1344.2200 569.9600 1345.8200 570.4400 ;
        RECT 1356.5600 548.2000 1359.5600 548.6800 ;
        RECT 1356.5600 553.6400 1359.5600 554.1200 ;
        RECT 1356.5600 559.0800 1359.5600 559.5600 ;
        RECT 1344.2200 548.2000 1345.8200 548.6800 ;
        RECT 1344.2200 553.6400 1345.8200 554.1200 ;
        RECT 1344.2200 559.0800 1345.8200 559.5600 ;
        RECT 1356.5600 542.7600 1359.5600 543.2400 ;
        RECT 1344.2200 542.7600 1345.8200 543.2400 ;
        RECT 1299.2200 575.4000 1300.8200 575.8800 ;
        RECT 1299.2200 580.8400 1300.8200 581.3200 ;
        RECT 1299.2200 586.2800 1300.8200 586.7600 ;
        RECT 1299.2200 564.5200 1300.8200 565.0000 ;
        RECT 1299.2200 569.9600 1300.8200 570.4400 ;
        RECT 1299.2200 548.2000 1300.8200 548.6800 ;
        RECT 1299.2200 553.6400 1300.8200 554.1200 ;
        RECT 1299.2200 559.0800 1300.8200 559.5600 ;
        RECT 1299.2200 542.7600 1300.8200 543.2400 ;
        RECT 1254.2200 629.8000 1255.8200 630.2800 ;
        RECT 1254.2200 635.2400 1255.8200 635.7200 ;
        RECT 1254.2200 640.6800 1255.8200 641.1600 ;
        RECT 1254.2200 618.9200 1255.8200 619.4000 ;
        RECT 1254.2200 624.3600 1255.8200 624.8400 ;
        RECT 1209.2200 629.8000 1210.8200 630.2800 ;
        RECT 1209.2200 635.2400 1210.8200 635.7200 ;
        RECT 1209.2200 640.6800 1210.8200 641.1600 ;
        RECT 1209.2200 618.9200 1210.8200 619.4000 ;
        RECT 1209.2200 624.3600 1210.8200 624.8400 ;
        RECT 1254.2200 602.6000 1255.8200 603.0800 ;
        RECT 1254.2200 608.0400 1255.8200 608.5200 ;
        RECT 1254.2200 613.4800 1255.8200 613.9600 ;
        RECT 1254.2200 591.7200 1255.8200 592.2000 ;
        RECT 1254.2200 597.1600 1255.8200 597.6400 ;
        RECT 1209.2200 602.6000 1210.8200 603.0800 ;
        RECT 1209.2200 608.0400 1210.8200 608.5200 ;
        RECT 1209.2200 613.4800 1210.8200 613.9600 ;
        RECT 1209.2200 591.7200 1210.8200 592.2000 ;
        RECT 1209.2200 597.1600 1210.8200 597.6400 ;
        RECT 1164.2200 629.8000 1165.8200 630.2800 ;
        RECT 1164.2200 635.2400 1165.8200 635.7200 ;
        RECT 1164.2200 640.6800 1165.8200 641.1600 ;
        RECT 1152.4600 629.8000 1155.4600 630.2800 ;
        RECT 1152.4600 635.2400 1155.4600 635.7200 ;
        RECT 1152.4600 640.6800 1155.4600 641.1600 ;
        RECT 1164.2200 618.9200 1165.8200 619.4000 ;
        RECT 1164.2200 624.3600 1165.8200 624.8400 ;
        RECT 1152.4600 618.9200 1155.4600 619.4000 ;
        RECT 1152.4600 624.3600 1155.4600 624.8400 ;
        RECT 1164.2200 602.6000 1165.8200 603.0800 ;
        RECT 1164.2200 608.0400 1165.8200 608.5200 ;
        RECT 1164.2200 613.4800 1165.8200 613.9600 ;
        RECT 1152.4600 602.6000 1155.4600 603.0800 ;
        RECT 1152.4600 608.0400 1155.4600 608.5200 ;
        RECT 1152.4600 613.4800 1155.4600 613.9600 ;
        RECT 1164.2200 591.7200 1165.8200 592.2000 ;
        RECT 1164.2200 597.1600 1165.8200 597.6400 ;
        RECT 1152.4600 591.7200 1155.4600 592.2000 ;
        RECT 1152.4600 597.1600 1155.4600 597.6400 ;
        RECT 1254.2200 575.4000 1255.8200 575.8800 ;
        RECT 1254.2200 580.8400 1255.8200 581.3200 ;
        RECT 1254.2200 586.2800 1255.8200 586.7600 ;
        RECT 1254.2200 564.5200 1255.8200 565.0000 ;
        RECT 1254.2200 569.9600 1255.8200 570.4400 ;
        RECT 1209.2200 575.4000 1210.8200 575.8800 ;
        RECT 1209.2200 580.8400 1210.8200 581.3200 ;
        RECT 1209.2200 586.2800 1210.8200 586.7600 ;
        RECT 1209.2200 564.5200 1210.8200 565.0000 ;
        RECT 1209.2200 569.9600 1210.8200 570.4400 ;
        RECT 1254.2200 548.2000 1255.8200 548.6800 ;
        RECT 1254.2200 553.6400 1255.8200 554.1200 ;
        RECT 1254.2200 559.0800 1255.8200 559.5600 ;
        RECT 1254.2200 542.7600 1255.8200 543.2400 ;
        RECT 1209.2200 548.2000 1210.8200 548.6800 ;
        RECT 1209.2200 553.6400 1210.8200 554.1200 ;
        RECT 1209.2200 559.0800 1210.8200 559.5600 ;
        RECT 1209.2200 542.7600 1210.8200 543.2400 ;
        RECT 1164.2200 575.4000 1165.8200 575.8800 ;
        RECT 1164.2200 580.8400 1165.8200 581.3200 ;
        RECT 1164.2200 586.2800 1165.8200 586.7600 ;
        RECT 1152.4600 575.4000 1155.4600 575.8800 ;
        RECT 1152.4600 580.8400 1155.4600 581.3200 ;
        RECT 1152.4600 586.2800 1155.4600 586.7600 ;
        RECT 1164.2200 564.5200 1165.8200 565.0000 ;
        RECT 1164.2200 569.9600 1165.8200 570.4400 ;
        RECT 1152.4600 564.5200 1155.4600 565.0000 ;
        RECT 1152.4600 569.9600 1155.4600 570.4400 ;
        RECT 1164.2200 548.2000 1165.8200 548.6800 ;
        RECT 1164.2200 553.6400 1165.8200 554.1200 ;
        RECT 1164.2200 559.0800 1165.8200 559.5600 ;
        RECT 1152.4600 548.2000 1155.4600 548.6800 ;
        RECT 1152.4600 553.6400 1155.4600 554.1200 ;
        RECT 1152.4600 559.0800 1155.4600 559.5600 ;
        RECT 1152.4600 542.7600 1155.4600 543.2400 ;
        RECT 1164.2200 542.7600 1165.8200 543.2400 ;
        RECT 1152.4600 747.6700 1359.5600 750.6700 ;
        RECT 1152.4600 534.5700 1359.5600 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 304.9300 1345.8200 521.0300 ;
        RECT 1299.2200 304.9300 1300.8200 521.0300 ;
        RECT 1254.2200 304.9300 1255.8200 521.0300 ;
        RECT 1209.2200 304.9300 1210.8200 521.0300 ;
        RECT 1164.2200 304.9300 1165.8200 521.0300 ;
        RECT 1356.5600 304.9300 1359.5600 521.0300 ;
        RECT 1152.4600 304.9300 1155.4600 521.0300 ;
      LAYER met3 ;
        RECT 1356.5600 498.0800 1359.5600 498.5600 ;
        RECT 1356.5600 503.5200 1359.5600 504.0000 ;
        RECT 1344.2200 498.0800 1345.8200 498.5600 ;
        RECT 1344.2200 503.5200 1345.8200 504.0000 ;
        RECT 1356.5600 508.9600 1359.5600 509.4400 ;
        RECT 1344.2200 508.9600 1345.8200 509.4400 ;
        RECT 1356.5600 487.2000 1359.5600 487.6800 ;
        RECT 1356.5600 492.6400 1359.5600 493.1200 ;
        RECT 1344.2200 487.2000 1345.8200 487.6800 ;
        RECT 1344.2200 492.6400 1345.8200 493.1200 ;
        RECT 1356.5600 470.8800 1359.5600 471.3600 ;
        RECT 1356.5600 476.3200 1359.5600 476.8000 ;
        RECT 1344.2200 470.8800 1345.8200 471.3600 ;
        RECT 1344.2200 476.3200 1345.8200 476.8000 ;
        RECT 1356.5600 481.7600 1359.5600 482.2400 ;
        RECT 1344.2200 481.7600 1345.8200 482.2400 ;
        RECT 1299.2200 498.0800 1300.8200 498.5600 ;
        RECT 1299.2200 503.5200 1300.8200 504.0000 ;
        RECT 1299.2200 508.9600 1300.8200 509.4400 ;
        RECT 1299.2200 487.2000 1300.8200 487.6800 ;
        RECT 1299.2200 492.6400 1300.8200 493.1200 ;
        RECT 1299.2200 470.8800 1300.8200 471.3600 ;
        RECT 1299.2200 476.3200 1300.8200 476.8000 ;
        RECT 1299.2200 481.7600 1300.8200 482.2400 ;
        RECT 1356.5600 454.5600 1359.5600 455.0400 ;
        RECT 1356.5600 460.0000 1359.5600 460.4800 ;
        RECT 1356.5600 465.4400 1359.5600 465.9200 ;
        RECT 1344.2200 454.5600 1345.8200 455.0400 ;
        RECT 1344.2200 460.0000 1345.8200 460.4800 ;
        RECT 1344.2200 465.4400 1345.8200 465.9200 ;
        RECT 1356.5600 443.6800 1359.5600 444.1600 ;
        RECT 1356.5600 449.1200 1359.5600 449.6000 ;
        RECT 1344.2200 443.6800 1345.8200 444.1600 ;
        RECT 1344.2200 449.1200 1345.8200 449.6000 ;
        RECT 1356.5600 427.3600 1359.5600 427.8400 ;
        RECT 1356.5600 432.8000 1359.5600 433.2800 ;
        RECT 1356.5600 438.2400 1359.5600 438.7200 ;
        RECT 1344.2200 427.3600 1345.8200 427.8400 ;
        RECT 1344.2200 432.8000 1345.8200 433.2800 ;
        RECT 1344.2200 438.2400 1345.8200 438.7200 ;
        RECT 1356.5600 416.4800 1359.5600 416.9600 ;
        RECT 1356.5600 421.9200 1359.5600 422.4000 ;
        RECT 1344.2200 416.4800 1345.8200 416.9600 ;
        RECT 1344.2200 421.9200 1345.8200 422.4000 ;
        RECT 1299.2200 454.5600 1300.8200 455.0400 ;
        RECT 1299.2200 460.0000 1300.8200 460.4800 ;
        RECT 1299.2200 465.4400 1300.8200 465.9200 ;
        RECT 1299.2200 443.6800 1300.8200 444.1600 ;
        RECT 1299.2200 449.1200 1300.8200 449.6000 ;
        RECT 1299.2200 427.3600 1300.8200 427.8400 ;
        RECT 1299.2200 432.8000 1300.8200 433.2800 ;
        RECT 1299.2200 438.2400 1300.8200 438.7200 ;
        RECT 1299.2200 416.4800 1300.8200 416.9600 ;
        RECT 1299.2200 421.9200 1300.8200 422.4000 ;
        RECT 1254.2200 498.0800 1255.8200 498.5600 ;
        RECT 1254.2200 503.5200 1255.8200 504.0000 ;
        RECT 1254.2200 508.9600 1255.8200 509.4400 ;
        RECT 1209.2200 498.0800 1210.8200 498.5600 ;
        RECT 1209.2200 503.5200 1210.8200 504.0000 ;
        RECT 1209.2200 508.9600 1210.8200 509.4400 ;
        RECT 1254.2200 487.2000 1255.8200 487.6800 ;
        RECT 1254.2200 492.6400 1255.8200 493.1200 ;
        RECT 1254.2200 470.8800 1255.8200 471.3600 ;
        RECT 1254.2200 476.3200 1255.8200 476.8000 ;
        RECT 1254.2200 481.7600 1255.8200 482.2400 ;
        RECT 1209.2200 487.2000 1210.8200 487.6800 ;
        RECT 1209.2200 492.6400 1210.8200 493.1200 ;
        RECT 1209.2200 470.8800 1210.8200 471.3600 ;
        RECT 1209.2200 476.3200 1210.8200 476.8000 ;
        RECT 1209.2200 481.7600 1210.8200 482.2400 ;
        RECT 1164.2200 498.0800 1165.8200 498.5600 ;
        RECT 1164.2200 503.5200 1165.8200 504.0000 ;
        RECT 1152.4600 503.5200 1155.4600 504.0000 ;
        RECT 1152.4600 498.0800 1155.4600 498.5600 ;
        RECT 1152.4600 508.9600 1155.4600 509.4400 ;
        RECT 1164.2200 508.9600 1165.8200 509.4400 ;
        RECT 1164.2200 487.2000 1165.8200 487.6800 ;
        RECT 1164.2200 492.6400 1165.8200 493.1200 ;
        RECT 1152.4600 492.6400 1155.4600 493.1200 ;
        RECT 1152.4600 487.2000 1155.4600 487.6800 ;
        RECT 1164.2200 470.8800 1165.8200 471.3600 ;
        RECT 1164.2200 476.3200 1165.8200 476.8000 ;
        RECT 1152.4600 476.3200 1155.4600 476.8000 ;
        RECT 1152.4600 470.8800 1155.4600 471.3600 ;
        RECT 1152.4600 481.7600 1155.4600 482.2400 ;
        RECT 1164.2200 481.7600 1165.8200 482.2400 ;
        RECT 1254.2200 454.5600 1255.8200 455.0400 ;
        RECT 1254.2200 460.0000 1255.8200 460.4800 ;
        RECT 1254.2200 465.4400 1255.8200 465.9200 ;
        RECT 1254.2200 443.6800 1255.8200 444.1600 ;
        RECT 1254.2200 449.1200 1255.8200 449.6000 ;
        RECT 1209.2200 454.5600 1210.8200 455.0400 ;
        RECT 1209.2200 460.0000 1210.8200 460.4800 ;
        RECT 1209.2200 465.4400 1210.8200 465.9200 ;
        RECT 1209.2200 443.6800 1210.8200 444.1600 ;
        RECT 1209.2200 449.1200 1210.8200 449.6000 ;
        RECT 1254.2200 427.3600 1255.8200 427.8400 ;
        RECT 1254.2200 432.8000 1255.8200 433.2800 ;
        RECT 1254.2200 438.2400 1255.8200 438.7200 ;
        RECT 1254.2200 416.4800 1255.8200 416.9600 ;
        RECT 1254.2200 421.9200 1255.8200 422.4000 ;
        RECT 1209.2200 427.3600 1210.8200 427.8400 ;
        RECT 1209.2200 432.8000 1210.8200 433.2800 ;
        RECT 1209.2200 438.2400 1210.8200 438.7200 ;
        RECT 1209.2200 416.4800 1210.8200 416.9600 ;
        RECT 1209.2200 421.9200 1210.8200 422.4000 ;
        RECT 1164.2200 454.5600 1165.8200 455.0400 ;
        RECT 1164.2200 460.0000 1165.8200 460.4800 ;
        RECT 1164.2200 465.4400 1165.8200 465.9200 ;
        RECT 1152.4600 454.5600 1155.4600 455.0400 ;
        RECT 1152.4600 460.0000 1155.4600 460.4800 ;
        RECT 1152.4600 465.4400 1155.4600 465.9200 ;
        RECT 1164.2200 443.6800 1165.8200 444.1600 ;
        RECT 1164.2200 449.1200 1165.8200 449.6000 ;
        RECT 1152.4600 443.6800 1155.4600 444.1600 ;
        RECT 1152.4600 449.1200 1155.4600 449.6000 ;
        RECT 1164.2200 427.3600 1165.8200 427.8400 ;
        RECT 1164.2200 432.8000 1165.8200 433.2800 ;
        RECT 1164.2200 438.2400 1165.8200 438.7200 ;
        RECT 1152.4600 427.3600 1155.4600 427.8400 ;
        RECT 1152.4600 432.8000 1155.4600 433.2800 ;
        RECT 1152.4600 438.2400 1155.4600 438.7200 ;
        RECT 1164.2200 416.4800 1165.8200 416.9600 ;
        RECT 1164.2200 421.9200 1165.8200 422.4000 ;
        RECT 1152.4600 416.4800 1155.4600 416.9600 ;
        RECT 1152.4600 421.9200 1155.4600 422.4000 ;
        RECT 1356.5600 400.1600 1359.5600 400.6400 ;
        RECT 1356.5600 405.6000 1359.5600 406.0800 ;
        RECT 1356.5600 411.0400 1359.5600 411.5200 ;
        RECT 1344.2200 400.1600 1345.8200 400.6400 ;
        RECT 1344.2200 405.6000 1345.8200 406.0800 ;
        RECT 1344.2200 411.0400 1345.8200 411.5200 ;
        RECT 1356.5600 389.2800 1359.5600 389.7600 ;
        RECT 1356.5600 394.7200 1359.5600 395.2000 ;
        RECT 1344.2200 389.2800 1345.8200 389.7600 ;
        RECT 1344.2200 394.7200 1345.8200 395.2000 ;
        RECT 1356.5600 372.9600 1359.5600 373.4400 ;
        RECT 1356.5600 378.4000 1359.5600 378.8800 ;
        RECT 1356.5600 383.8400 1359.5600 384.3200 ;
        RECT 1344.2200 372.9600 1345.8200 373.4400 ;
        RECT 1344.2200 378.4000 1345.8200 378.8800 ;
        RECT 1344.2200 383.8400 1345.8200 384.3200 ;
        RECT 1356.5600 362.0800 1359.5600 362.5600 ;
        RECT 1356.5600 367.5200 1359.5600 368.0000 ;
        RECT 1344.2200 362.0800 1345.8200 362.5600 ;
        RECT 1344.2200 367.5200 1345.8200 368.0000 ;
        RECT 1299.2200 400.1600 1300.8200 400.6400 ;
        RECT 1299.2200 405.6000 1300.8200 406.0800 ;
        RECT 1299.2200 411.0400 1300.8200 411.5200 ;
        RECT 1299.2200 389.2800 1300.8200 389.7600 ;
        RECT 1299.2200 394.7200 1300.8200 395.2000 ;
        RECT 1299.2200 372.9600 1300.8200 373.4400 ;
        RECT 1299.2200 378.4000 1300.8200 378.8800 ;
        RECT 1299.2200 383.8400 1300.8200 384.3200 ;
        RECT 1299.2200 362.0800 1300.8200 362.5600 ;
        RECT 1299.2200 367.5200 1300.8200 368.0000 ;
        RECT 1356.5600 345.7600 1359.5600 346.2400 ;
        RECT 1356.5600 351.2000 1359.5600 351.6800 ;
        RECT 1356.5600 356.6400 1359.5600 357.1200 ;
        RECT 1344.2200 345.7600 1345.8200 346.2400 ;
        RECT 1344.2200 351.2000 1345.8200 351.6800 ;
        RECT 1344.2200 356.6400 1345.8200 357.1200 ;
        RECT 1356.5600 334.8800 1359.5600 335.3600 ;
        RECT 1356.5600 340.3200 1359.5600 340.8000 ;
        RECT 1344.2200 334.8800 1345.8200 335.3600 ;
        RECT 1344.2200 340.3200 1345.8200 340.8000 ;
        RECT 1356.5600 318.5600 1359.5600 319.0400 ;
        RECT 1356.5600 324.0000 1359.5600 324.4800 ;
        RECT 1356.5600 329.4400 1359.5600 329.9200 ;
        RECT 1344.2200 318.5600 1345.8200 319.0400 ;
        RECT 1344.2200 324.0000 1345.8200 324.4800 ;
        RECT 1344.2200 329.4400 1345.8200 329.9200 ;
        RECT 1356.5600 313.1200 1359.5600 313.6000 ;
        RECT 1344.2200 313.1200 1345.8200 313.6000 ;
        RECT 1299.2200 345.7600 1300.8200 346.2400 ;
        RECT 1299.2200 351.2000 1300.8200 351.6800 ;
        RECT 1299.2200 356.6400 1300.8200 357.1200 ;
        RECT 1299.2200 334.8800 1300.8200 335.3600 ;
        RECT 1299.2200 340.3200 1300.8200 340.8000 ;
        RECT 1299.2200 318.5600 1300.8200 319.0400 ;
        RECT 1299.2200 324.0000 1300.8200 324.4800 ;
        RECT 1299.2200 329.4400 1300.8200 329.9200 ;
        RECT 1299.2200 313.1200 1300.8200 313.6000 ;
        RECT 1254.2200 400.1600 1255.8200 400.6400 ;
        RECT 1254.2200 405.6000 1255.8200 406.0800 ;
        RECT 1254.2200 411.0400 1255.8200 411.5200 ;
        RECT 1254.2200 389.2800 1255.8200 389.7600 ;
        RECT 1254.2200 394.7200 1255.8200 395.2000 ;
        RECT 1209.2200 400.1600 1210.8200 400.6400 ;
        RECT 1209.2200 405.6000 1210.8200 406.0800 ;
        RECT 1209.2200 411.0400 1210.8200 411.5200 ;
        RECT 1209.2200 389.2800 1210.8200 389.7600 ;
        RECT 1209.2200 394.7200 1210.8200 395.2000 ;
        RECT 1254.2200 372.9600 1255.8200 373.4400 ;
        RECT 1254.2200 378.4000 1255.8200 378.8800 ;
        RECT 1254.2200 383.8400 1255.8200 384.3200 ;
        RECT 1254.2200 362.0800 1255.8200 362.5600 ;
        RECT 1254.2200 367.5200 1255.8200 368.0000 ;
        RECT 1209.2200 372.9600 1210.8200 373.4400 ;
        RECT 1209.2200 378.4000 1210.8200 378.8800 ;
        RECT 1209.2200 383.8400 1210.8200 384.3200 ;
        RECT 1209.2200 362.0800 1210.8200 362.5600 ;
        RECT 1209.2200 367.5200 1210.8200 368.0000 ;
        RECT 1164.2200 400.1600 1165.8200 400.6400 ;
        RECT 1164.2200 405.6000 1165.8200 406.0800 ;
        RECT 1164.2200 411.0400 1165.8200 411.5200 ;
        RECT 1152.4600 400.1600 1155.4600 400.6400 ;
        RECT 1152.4600 405.6000 1155.4600 406.0800 ;
        RECT 1152.4600 411.0400 1155.4600 411.5200 ;
        RECT 1164.2200 389.2800 1165.8200 389.7600 ;
        RECT 1164.2200 394.7200 1165.8200 395.2000 ;
        RECT 1152.4600 389.2800 1155.4600 389.7600 ;
        RECT 1152.4600 394.7200 1155.4600 395.2000 ;
        RECT 1164.2200 372.9600 1165.8200 373.4400 ;
        RECT 1164.2200 378.4000 1165.8200 378.8800 ;
        RECT 1164.2200 383.8400 1165.8200 384.3200 ;
        RECT 1152.4600 372.9600 1155.4600 373.4400 ;
        RECT 1152.4600 378.4000 1155.4600 378.8800 ;
        RECT 1152.4600 383.8400 1155.4600 384.3200 ;
        RECT 1164.2200 362.0800 1165.8200 362.5600 ;
        RECT 1164.2200 367.5200 1165.8200 368.0000 ;
        RECT 1152.4600 362.0800 1155.4600 362.5600 ;
        RECT 1152.4600 367.5200 1155.4600 368.0000 ;
        RECT 1254.2200 345.7600 1255.8200 346.2400 ;
        RECT 1254.2200 351.2000 1255.8200 351.6800 ;
        RECT 1254.2200 356.6400 1255.8200 357.1200 ;
        RECT 1254.2200 334.8800 1255.8200 335.3600 ;
        RECT 1254.2200 340.3200 1255.8200 340.8000 ;
        RECT 1209.2200 345.7600 1210.8200 346.2400 ;
        RECT 1209.2200 351.2000 1210.8200 351.6800 ;
        RECT 1209.2200 356.6400 1210.8200 357.1200 ;
        RECT 1209.2200 334.8800 1210.8200 335.3600 ;
        RECT 1209.2200 340.3200 1210.8200 340.8000 ;
        RECT 1254.2200 318.5600 1255.8200 319.0400 ;
        RECT 1254.2200 324.0000 1255.8200 324.4800 ;
        RECT 1254.2200 329.4400 1255.8200 329.9200 ;
        RECT 1254.2200 313.1200 1255.8200 313.6000 ;
        RECT 1209.2200 318.5600 1210.8200 319.0400 ;
        RECT 1209.2200 324.0000 1210.8200 324.4800 ;
        RECT 1209.2200 329.4400 1210.8200 329.9200 ;
        RECT 1209.2200 313.1200 1210.8200 313.6000 ;
        RECT 1164.2200 345.7600 1165.8200 346.2400 ;
        RECT 1164.2200 351.2000 1165.8200 351.6800 ;
        RECT 1164.2200 356.6400 1165.8200 357.1200 ;
        RECT 1152.4600 345.7600 1155.4600 346.2400 ;
        RECT 1152.4600 351.2000 1155.4600 351.6800 ;
        RECT 1152.4600 356.6400 1155.4600 357.1200 ;
        RECT 1164.2200 334.8800 1165.8200 335.3600 ;
        RECT 1164.2200 340.3200 1165.8200 340.8000 ;
        RECT 1152.4600 334.8800 1155.4600 335.3600 ;
        RECT 1152.4600 340.3200 1155.4600 340.8000 ;
        RECT 1164.2200 318.5600 1165.8200 319.0400 ;
        RECT 1164.2200 324.0000 1165.8200 324.4800 ;
        RECT 1164.2200 329.4400 1165.8200 329.9200 ;
        RECT 1152.4600 318.5600 1155.4600 319.0400 ;
        RECT 1152.4600 324.0000 1155.4600 324.4800 ;
        RECT 1152.4600 329.4400 1155.4600 329.9200 ;
        RECT 1152.4600 313.1200 1155.4600 313.6000 ;
        RECT 1164.2200 313.1200 1165.8200 313.6000 ;
        RECT 1152.4600 518.0300 1359.5600 521.0300 ;
        RECT 1152.4600 304.9300 1359.5600 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 75.2900 1345.8200 291.3900 ;
        RECT 1299.2200 75.2900 1300.8200 291.3900 ;
        RECT 1254.2200 75.2900 1255.8200 291.3900 ;
        RECT 1209.2200 75.2900 1210.8200 291.3900 ;
        RECT 1164.2200 75.2900 1165.8200 291.3900 ;
        RECT 1356.5600 75.2900 1359.5600 291.3900 ;
        RECT 1152.4600 75.2900 1155.4600 291.3900 ;
      LAYER met3 ;
        RECT 1356.5600 268.4400 1359.5600 268.9200 ;
        RECT 1356.5600 273.8800 1359.5600 274.3600 ;
        RECT 1344.2200 268.4400 1345.8200 268.9200 ;
        RECT 1344.2200 273.8800 1345.8200 274.3600 ;
        RECT 1356.5600 279.3200 1359.5600 279.8000 ;
        RECT 1344.2200 279.3200 1345.8200 279.8000 ;
        RECT 1356.5600 257.5600 1359.5600 258.0400 ;
        RECT 1356.5600 263.0000 1359.5600 263.4800 ;
        RECT 1344.2200 257.5600 1345.8200 258.0400 ;
        RECT 1344.2200 263.0000 1345.8200 263.4800 ;
        RECT 1356.5600 241.2400 1359.5600 241.7200 ;
        RECT 1356.5600 246.6800 1359.5600 247.1600 ;
        RECT 1344.2200 241.2400 1345.8200 241.7200 ;
        RECT 1344.2200 246.6800 1345.8200 247.1600 ;
        RECT 1356.5600 252.1200 1359.5600 252.6000 ;
        RECT 1344.2200 252.1200 1345.8200 252.6000 ;
        RECT 1299.2200 268.4400 1300.8200 268.9200 ;
        RECT 1299.2200 273.8800 1300.8200 274.3600 ;
        RECT 1299.2200 279.3200 1300.8200 279.8000 ;
        RECT 1299.2200 257.5600 1300.8200 258.0400 ;
        RECT 1299.2200 263.0000 1300.8200 263.4800 ;
        RECT 1299.2200 241.2400 1300.8200 241.7200 ;
        RECT 1299.2200 246.6800 1300.8200 247.1600 ;
        RECT 1299.2200 252.1200 1300.8200 252.6000 ;
        RECT 1356.5600 224.9200 1359.5600 225.4000 ;
        RECT 1356.5600 230.3600 1359.5600 230.8400 ;
        RECT 1356.5600 235.8000 1359.5600 236.2800 ;
        RECT 1344.2200 224.9200 1345.8200 225.4000 ;
        RECT 1344.2200 230.3600 1345.8200 230.8400 ;
        RECT 1344.2200 235.8000 1345.8200 236.2800 ;
        RECT 1356.5600 214.0400 1359.5600 214.5200 ;
        RECT 1356.5600 219.4800 1359.5600 219.9600 ;
        RECT 1344.2200 214.0400 1345.8200 214.5200 ;
        RECT 1344.2200 219.4800 1345.8200 219.9600 ;
        RECT 1356.5600 197.7200 1359.5600 198.2000 ;
        RECT 1356.5600 203.1600 1359.5600 203.6400 ;
        RECT 1356.5600 208.6000 1359.5600 209.0800 ;
        RECT 1344.2200 197.7200 1345.8200 198.2000 ;
        RECT 1344.2200 203.1600 1345.8200 203.6400 ;
        RECT 1344.2200 208.6000 1345.8200 209.0800 ;
        RECT 1356.5600 186.8400 1359.5600 187.3200 ;
        RECT 1356.5600 192.2800 1359.5600 192.7600 ;
        RECT 1344.2200 186.8400 1345.8200 187.3200 ;
        RECT 1344.2200 192.2800 1345.8200 192.7600 ;
        RECT 1299.2200 224.9200 1300.8200 225.4000 ;
        RECT 1299.2200 230.3600 1300.8200 230.8400 ;
        RECT 1299.2200 235.8000 1300.8200 236.2800 ;
        RECT 1299.2200 214.0400 1300.8200 214.5200 ;
        RECT 1299.2200 219.4800 1300.8200 219.9600 ;
        RECT 1299.2200 197.7200 1300.8200 198.2000 ;
        RECT 1299.2200 203.1600 1300.8200 203.6400 ;
        RECT 1299.2200 208.6000 1300.8200 209.0800 ;
        RECT 1299.2200 186.8400 1300.8200 187.3200 ;
        RECT 1299.2200 192.2800 1300.8200 192.7600 ;
        RECT 1254.2200 268.4400 1255.8200 268.9200 ;
        RECT 1254.2200 273.8800 1255.8200 274.3600 ;
        RECT 1254.2200 279.3200 1255.8200 279.8000 ;
        RECT 1209.2200 268.4400 1210.8200 268.9200 ;
        RECT 1209.2200 273.8800 1210.8200 274.3600 ;
        RECT 1209.2200 279.3200 1210.8200 279.8000 ;
        RECT 1254.2200 257.5600 1255.8200 258.0400 ;
        RECT 1254.2200 263.0000 1255.8200 263.4800 ;
        RECT 1254.2200 241.2400 1255.8200 241.7200 ;
        RECT 1254.2200 246.6800 1255.8200 247.1600 ;
        RECT 1254.2200 252.1200 1255.8200 252.6000 ;
        RECT 1209.2200 257.5600 1210.8200 258.0400 ;
        RECT 1209.2200 263.0000 1210.8200 263.4800 ;
        RECT 1209.2200 241.2400 1210.8200 241.7200 ;
        RECT 1209.2200 246.6800 1210.8200 247.1600 ;
        RECT 1209.2200 252.1200 1210.8200 252.6000 ;
        RECT 1164.2200 268.4400 1165.8200 268.9200 ;
        RECT 1164.2200 273.8800 1165.8200 274.3600 ;
        RECT 1152.4600 273.8800 1155.4600 274.3600 ;
        RECT 1152.4600 268.4400 1155.4600 268.9200 ;
        RECT 1152.4600 279.3200 1155.4600 279.8000 ;
        RECT 1164.2200 279.3200 1165.8200 279.8000 ;
        RECT 1164.2200 257.5600 1165.8200 258.0400 ;
        RECT 1164.2200 263.0000 1165.8200 263.4800 ;
        RECT 1152.4600 263.0000 1155.4600 263.4800 ;
        RECT 1152.4600 257.5600 1155.4600 258.0400 ;
        RECT 1164.2200 241.2400 1165.8200 241.7200 ;
        RECT 1164.2200 246.6800 1165.8200 247.1600 ;
        RECT 1152.4600 246.6800 1155.4600 247.1600 ;
        RECT 1152.4600 241.2400 1155.4600 241.7200 ;
        RECT 1152.4600 252.1200 1155.4600 252.6000 ;
        RECT 1164.2200 252.1200 1165.8200 252.6000 ;
        RECT 1254.2200 224.9200 1255.8200 225.4000 ;
        RECT 1254.2200 230.3600 1255.8200 230.8400 ;
        RECT 1254.2200 235.8000 1255.8200 236.2800 ;
        RECT 1254.2200 214.0400 1255.8200 214.5200 ;
        RECT 1254.2200 219.4800 1255.8200 219.9600 ;
        RECT 1209.2200 224.9200 1210.8200 225.4000 ;
        RECT 1209.2200 230.3600 1210.8200 230.8400 ;
        RECT 1209.2200 235.8000 1210.8200 236.2800 ;
        RECT 1209.2200 214.0400 1210.8200 214.5200 ;
        RECT 1209.2200 219.4800 1210.8200 219.9600 ;
        RECT 1254.2200 197.7200 1255.8200 198.2000 ;
        RECT 1254.2200 203.1600 1255.8200 203.6400 ;
        RECT 1254.2200 208.6000 1255.8200 209.0800 ;
        RECT 1254.2200 186.8400 1255.8200 187.3200 ;
        RECT 1254.2200 192.2800 1255.8200 192.7600 ;
        RECT 1209.2200 197.7200 1210.8200 198.2000 ;
        RECT 1209.2200 203.1600 1210.8200 203.6400 ;
        RECT 1209.2200 208.6000 1210.8200 209.0800 ;
        RECT 1209.2200 186.8400 1210.8200 187.3200 ;
        RECT 1209.2200 192.2800 1210.8200 192.7600 ;
        RECT 1164.2200 224.9200 1165.8200 225.4000 ;
        RECT 1164.2200 230.3600 1165.8200 230.8400 ;
        RECT 1164.2200 235.8000 1165.8200 236.2800 ;
        RECT 1152.4600 224.9200 1155.4600 225.4000 ;
        RECT 1152.4600 230.3600 1155.4600 230.8400 ;
        RECT 1152.4600 235.8000 1155.4600 236.2800 ;
        RECT 1164.2200 214.0400 1165.8200 214.5200 ;
        RECT 1164.2200 219.4800 1165.8200 219.9600 ;
        RECT 1152.4600 214.0400 1155.4600 214.5200 ;
        RECT 1152.4600 219.4800 1155.4600 219.9600 ;
        RECT 1164.2200 197.7200 1165.8200 198.2000 ;
        RECT 1164.2200 203.1600 1165.8200 203.6400 ;
        RECT 1164.2200 208.6000 1165.8200 209.0800 ;
        RECT 1152.4600 197.7200 1155.4600 198.2000 ;
        RECT 1152.4600 203.1600 1155.4600 203.6400 ;
        RECT 1152.4600 208.6000 1155.4600 209.0800 ;
        RECT 1164.2200 186.8400 1165.8200 187.3200 ;
        RECT 1164.2200 192.2800 1165.8200 192.7600 ;
        RECT 1152.4600 186.8400 1155.4600 187.3200 ;
        RECT 1152.4600 192.2800 1155.4600 192.7600 ;
        RECT 1356.5600 170.5200 1359.5600 171.0000 ;
        RECT 1356.5600 175.9600 1359.5600 176.4400 ;
        RECT 1356.5600 181.4000 1359.5600 181.8800 ;
        RECT 1344.2200 170.5200 1345.8200 171.0000 ;
        RECT 1344.2200 175.9600 1345.8200 176.4400 ;
        RECT 1344.2200 181.4000 1345.8200 181.8800 ;
        RECT 1356.5600 159.6400 1359.5600 160.1200 ;
        RECT 1356.5600 165.0800 1359.5600 165.5600 ;
        RECT 1344.2200 159.6400 1345.8200 160.1200 ;
        RECT 1344.2200 165.0800 1345.8200 165.5600 ;
        RECT 1356.5600 143.3200 1359.5600 143.8000 ;
        RECT 1356.5600 148.7600 1359.5600 149.2400 ;
        RECT 1356.5600 154.2000 1359.5600 154.6800 ;
        RECT 1344.2200 143.3200 1345.8200 143.8000 ;
        RECT 1344.2200 148.7600 1345.8200 149.2400 ;
        RECT 1344.2200 154.2000 1345.8200 154.6800 ;
        RECT 1356.5600 132.4400 1359.5600 132.9200 ;
        RECT 1356.5600 137.8800 1359.5600 138.3600 ;
        RECT 1344.2200 132.4400 1345.8200 132.9200 ;
        RECT 1344.2200 137.8800 1345.8200 138.3600 ;
        RECT 1299.2200 170.5200 1300.8200 171.0000 ;
        RECT 1299.2200 175.9600 1300.8200 176.4400 ;
        RECT 1299.2200 181.4000 1300.8200 181.8800 ;
        RECT 1299.2200 159.6400 1300.8200 160.1200 ;
        RECT 1299.2200 165.0800 1300.8200 165.5600 ;
        RECT 1299.2200 143.3200 1300.8200 143.8000 ;
        RECT 1299.2200 148.7600 1300.8200 149.2400 ;
        RECT 1299.2200 154.2000 1300.8200 154.6800 ;
        RECT 1299.2200 132.4400 1300.8200 132.9200 ;
        RECT 1299.2200 137.8800 1300.8200 138.3600 ;
        RECT 1356.5600 116.1200 1359.5600 116.6000 ;
        RECT 1356.5600 121.5600 1359.5600 122.0400 ;
        RECT 1356.5600 127.0000 1359.5600 127.4800 ;
        RECT 1344.2200 116.1200 1345.8200 116.6000 ;
        RECT 1344.2200 121.5600 1345.8200 122.0400 ;
        RECT 1344.2200 127.0000 1345.8200 127.4800 ;
        RECT 1356.5600 105.2400 1359.5600 105.7200 ;
        RECT 1356.5600 110.6800 1359.5600 111.1600 ;
        RECT 1344.2200 105.2400 1345.8200 105.7200 ;
        RECT 1344.2200 110.6800 1345.8200 111.1600 ;
        RECT 1356.5600 88.9200 1359.5600 89.4000 ;
        RECT 1356.5600 94.3600 1359.5600 94.8400 ;
        RECT 1356.5600 99.8000 1359.5600 100.2800 ;
        RECT 1344.2200 88.9200 1345.8200 89.4000 ;
        RECT 1344.2200 94.3600 1345.8200 94.8400 ;
        RECT 1344.2200 99.8000 1345.8200 100.2800 ;
        RECT 1356.5600 83.4800 1359.5600 83.9600 ;
        RECT 1344.2200 83.4800 1345.8200 83.9600 ;
        RECT 1299.2200 116.1200 1300.8200 116.6000 ;
        RECT 1299.2200 121.5600 1300.8200 122.0400 ;
        RECT 1299.2200 127.0000 1300.8200 127.4800 ;
        RECT 1299.2200 105.2400 1300.8200 105.7200 ;
        RECT 1299.2200 110.6800 1300.8200 111.1600 ;
        RECT 1299.2200 88.9200 1300.8200 89.4000 ;
        RECT 1299.2200 94.3600 1300.8200 94.8400 ;
        RECT 1299.2200 99.8000 1300.8200 100.2800 ;
        RECT 1299.2200 83.4800 1300.8200 83.9600 ;
        RECT 1254.2200 170.5200 1255.8200 171.0000 ;
        RECT 1254.2200 175.9600 1255.8200 176.4400 ;
        RECT 1254.2200 181.4000 1255.8200 181.8800 ;
        RECT 1254.2200 159.6400 1255.8200 160.1200 ;
        RECT 1254.2200 165.0800 1255.8200 165.5600 ;
        RECT 1209.2200 170.5200 1210.8200 171.0000 ;
        RECT 1209.2200 175.9600 1210.8200 176.4400 ;
        RECT 1209.2200 181.4000 1210.8200 181.8800 ;
        RECT 1209.2200 159.6400 1210.8200 160.1200 ;
        RECT 1209.2200 165.0800 1210.8200 165.5600 ;
        RECT 1254.2200 143.3200 1255.8200 143.8000 ;
        RECT 1254.2200 148.7600 1255.8200 149.2400 ;
        RECT 1254.2200 154.2000 1255.8200 154.6800 ;
        RECT 1254.2200 132.4400 1255.8200 132.9200 ;
        RECT 1254.2200 137.8800 1255.8200 138.3600 ;
        RECT 1209.2200 143.3200 1210.8200 143.8000 ;
        RECT 1209.2200 148.7600 1210.8200 149.2400 ;
        RECT 1209.2200 154.2000 1210.8200 154.6800 ;
        RECT 1209.2200 132.4400 1210.8200 132.9200 ;
        RECT 1209.2200 137.8800 1210.8200 138.3600 ;
        RECT 1164.2200 170.5200 1165.8200 171.0000 ;
        RECT 1164.2200 175.9600 1165.8200 176.4400 ;
        RECT 1164.2200 181.4000 1165.8200 181.8800 ;
        RECT 1152.4600 170.5200 1155.4600 171.0000 ;
        RECT 1152.4600 175.9600 1155.4600 176.4400 ;
        RECT 1152.4600 181.4000 1155.4600 181.8800 ;
        RECT 1164.2200 159.6400 1165.8200 160.1200 ;
        RECT 1164.2200 165.0800 1165.8200 165.5600 ;
        RECT 1152.4600 159.6400 1155.4600 160.1200 ;
        RECT 1152.4600 165.0800 1155.4600 165.5600 ;
        RECT 1164.2200 143.3200 1165.8200 143.8000 ;
        RECT 1164.2200 148.7600 1165.8200 149.2400 ;
        RECT 1164.2200 154.2000 1165.8200 154.6800 ;
        RECT 1152.4600 143.3200 1155.4600 143.8000 ;
        RECT 1152.4600 148.7600 1155.4600 149.2400 ;
        RECT 1152.4600 154.2000 1155.4600 154.6800 ;
        RECT 1164.2200 132.4400 1165.8200 132.9200 ;
        RECT 1164.2200 137.8800 1165.8200 138.3600 ;
        RECT 1152.4600 132.4400 1155.4600 132.9200 ;
        RECT 1152.4600 137.8800 1155.4600 138.3600 ;
        RECT 1254.2200 116.1200 1255.8200 116.6000 ;
        RECT 1254.2200 121.5600 1255.8200 122.0400 ;
        RECT 1254.2200 127.0000 1255.8200 127.4800 ;
        RECT 1254.2200 105.2400 1255.8200 105.7200 ;
        RECT 1254.2200 110.6800 1255.8200 111.1600 ;
        RECT 1209.2200 116.1200 1210.8200 116.6000 ;
        RECT 1209.2200 121.5600 1210.8200 122.0400 ;
        RECT 1209.2200 127.0000 1210.8200 127.4800 ;
        RECT 1209.2200 105.2400 1210.8200 105.7200 ;
        RECT 1209.2200 110.6800 1210.8200 111.1600 ;
        RECT 1254.2200 88.9200 1255.8200 89.4000 ;
        RECT 1254.2200 94.3600 1255.8200 94.8400 ;
        RECT 1254.2200 99.8000 1255.8200 100.2800 ;
        RECT 1254.2200 83.4800 1255.8200 83.9600 ;
        RECT 1209.2200 88.9200 1210.8200 89.4000 ;
        RECT 1209.2200 94.3600 1210.8200 94.8400 ;
        RECT 1209.2200 99.8000 1210.8200 100.2800 ;
        RECT 1209.2200 83.4800 1210.8200 83.9600 ;
        RECT 1164.2200 116.1200 1165.8200 116.6000 ;
        RECT 1164.2200 121.5600 1165.8200 122.0400 ;
        RECT 1164.2200 127.0000 1165.8200 127.4800 ;
        RECT 1152.4600 116.1200 1155.4600 116.6000 ;
        RECT 1152.4600 121.5600 1155.4600 122.0400 ;
        RECT 1152.4600 127.0000 1155.4600 127.4800 ;
        RECT 1164.2200 105.2400 1165.8200 105.7200 ;
        RECT 1164.2200 110.6800 1165.8200 111.1600 ;
        RECT 1152.4600 105.2400 1155.4600 105.7200 ;
        RECT 1152.4600 110.6800 1155.4600 111.1600 ;
        RECT 1164.2200 88.9200 1165.8200 89.4000 ;
        RECT 1164.2200 94.3600 1165.8200 94.8400 ;
        RECT 1164.2200 99.8000 1165.8200 100.2800 ;
        RECT 1152.4600 88.9200 1155.4600 89.4000 ;
        RECT 1152.4600 94.3600 1155.4600 94.8400 ;
        RECT 1152.4600 99.8000 1155.4600 100.2800 ;
        RECT 1152.4600 83.4800 1155.4600 83.9600 ;
        RECT 1164.2200 83.4800 1165.8200 83.9600 ;
        RECT 1152.4600 288.3900 1359.5600 291.3900 ;
        RECT 1152.4600 75.2900 1359.5600 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1153.4600 34.6700 1155.4600 61.6000 ;
        RECT 1356.5600 34.6700 1358.5600 61.6000 ;
      LAYER met3 ;
        RECT 1356.5600 51.3800 1358.5600 51.8600 ;
        RECT 1153.4600 51.3800 1155.4600 51.8600 ;
        RECT 1356.5600 45.9400 1358.5600 46.4200 ;
        RECT 1356.5600 40.5000 1358.5600 40.9800 ;
        RECT 1153.4600 45.9400 1155.4600 46.4200 ;
        RECT 1153.4600 40.5000 1155.4600 40.9800 ;
        RECT 1153.4600 59.6000 1358.5600 61.6000 ;
        RECT 1153.4600 34.6700 1358.5600 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 2601.3300 1345.8200 2817.4300 ;
        RECT 1299.2200 2601.3300 1300.8200 2817.4300 ;
        RECT 1254.2200 2601.3300 1255.8200 2817.4300 ;
        RECT 1209.2200 2601.3300 1210.8200 2817.4300 ;
        RECT 1164.2200 2601.3300 1165.8200 2817.4300 ;
        RECT 1356.5600 2601.3300 1359.5600 2817.4300 ;
        RECT 1152.4600 2601.3300 1155.4600 2817.4300 ;
      LAYER met3 ;
        RECT 1356.5600 2794.4800 1359.5600 2794.9600 ;
        RECT 1356.5600 2799.9200 1359.5600 2800.4000 ;
        RECT 1344.2200 2794.4800 1345.8200 2794.9600 ;
        RECT 1344.2200 2799.9200 1345.8200 2800.4000 ;
        RECT 1356.5600 2805.3600 1359.5600 2805.8400 ;
        RECT 1344.2200 2805.3600 1345.8200 2805.8400 ;
        RECT 1356.5600 2783.6000 1359.5600 2784.0800 ;
        RECT 1356.5600 2789.0400 1359.5600 2789.5200 ;
        RECT 1344.2200 2783.6000 1345.8200 2784.0800 ;
        RECT 1344.2200 2789.0400 1345.8200 2789.5200 ;
        RECT 1356.5600 2767.2800 1359.5600 2767.7600 ;
        RECT 1356.5600 2772.7200 1359.5600 2773.2000 ;
        RECT 1344.2200 2767.2800 1345.8200 2767.7600 ;
        RECT 1344.2200 2772.7200 1345.8200 2773.2000 ;
        RECT 1356.5600 2778.1600 1359.5600 2778.6400 ;
        RECT 1344.2200 2778.1600 1345.8200 2778.6400 ;
        RECT 1299.2200 2794.4800 1300.8200 2794.9600 ;
        RECT 1299.2200 2799.9200 1300.8200 2800.4000 ;
        RECT 1299.2200 2805.3600 1300.8200 2805.8400 ;
        RECT 1299.2200 2783.6000 1300.8200 2784.0800 ;
        RECT 1299.2200 2789.0400 1300.8200 2789.5200 ;
        RECT 1299.2200 2767.2800 1300.8200 2767.7600 ;
        RECT 1299.2200 2772.7200 1300.8200 2773.2000 ;
        RECT 1299.2200 2778.1600 1300.8200 2778.6400 ;
        RECT 1356.5600 2750.9600 1359.5600 2751.4400 ;
        RECT 1356.5600 2756.4000 1359.5600 2756.8800 ;
        RECT 1356.5600 2761.8400 1359.5600 2762.3200 ;
        RECT 1344.2200 2750.9600 1345.8200 2751.4400 ;
        RECT 1344.2200 2756.4000 1345.8200 2756.8800 ;
        RECT 1344.2200 2761.8400 1345.8200 2762.3200 ;
        RECT 1356.5600 2740.0800 1359.5600 2740.5600 ;
        RECT 1356.5600 2745.5200 1359.5600 2746.0000 ;
        RECT 1344.2200 2740.0800 1345.8200 2740.5600 ;
        RECT 1344.2200 2745.5200 1345.8200 2746.0000 ;
        RECT 1356.5600 2723.7600 1359.5600 2724.2400 ;
        RECT 1356.5600 2729.2000 1359.5600 2729.6800 ;
        RECT 1356.5600 2734.6400 1359.5600 2735.1200 ;
        RECT 1344.2200 2723.7600 1345.8200 2724.2400 ;
        RECT 1344.2200 2729.2000 1345.8200 2729.6800 ;
        RECT 1344.2200 2734.6400 1345.8200 2735.1200 ;
        RECT 1356.5600 2712.8800 1359.5600 2713.3600 ;
        RECT 1356.5600 2718.3200 1359.5600 2718.8000 ;
        RECT 1344.2200 2712.8800 1345.8200 2713.3600 ;
        RECT 1344.2200 2718.3200 1345.8200 2718.8000 ;
        RECT 1299.2200 2750.9600 1300.8200 2751.4400 ;
        RECT 1299.2200 2756.4000 1300.8200 2756.8800 ;
        RECT 1299.2200 2761.8400 1300.8200 2762.3200 ;
        RECT 1299.2200 2740.0800 1300.8200 2740.5600 ;
        RECT 1299.2200 2745.5200 1300.8200 2746.0000 ;
        RECT 1299.2200 2723.7600 1300.8200 2724.2400 ;
        RECT 1299.2200 2729.2000 1300.8200 2729.6800 ;
        RECT 1299.2200 2734.6400 1300.8200 2735.1200 ;
        RECT 1299.2200 2712.8800 1300.8200 2713.3600 ;
        RECT 1299.2200 2718.3200 1300.8200 2718.8000 ;
        RECT 1254.2200 2794.4800 1255.8200 2794.9600 ;
        RECT 1254.2200 2799.9200 1255.8200 2800.4000 ;
        RECT 1254.2200 2805.3600 1255.8200 2805.8400 ;
        RECT 1209.2200 2794.4800 1210.8200 2794.9600 ;
        RECT 1209.2200 2799.9200 1210.8200 2800.4000 ;
        RECT 1209.2200 2805.3600 1210.8200 2805.8400 ;
        RECT 1254.2200 2783.6000 1255.8200 2784.0800 ;
        RECT 1254.2200 2789.0400 1255.8200 2789.5200 ;
        RECT 1254.2200 2767.2800 1255.8200 2767.7600 ;
        RECT 1254.2200 2772.7200 1255.8200 2773.2000 ;
        RECT 1254.2200 2778.1600 1255.8200 2778.6400 ;
        RECT 1209.2200 2783.6000 1210.8200 2784.0800 ;
        RECT 1209.2200 2789.0400 1210.8200 2789.5200 ;
        RECT 1209.2200 2767.2800 1210.8200 2767.7600 ;
        RECT 1209.2200 2772.7200 1210.8200 2773.2000 ;
        RECT 1209.2200 2778.1600 1210.8200 2778.6400 ;
        RECT 1164.2200 2794.4800 1165.8200 2794.9600 ;
        RECT 1164.2200 2799.9200 1165.8200 2800.4000 ;
        RECT 1152.4600 2799.9200 1155.4600 2800.4000 ;
        RECT 1152.4600 2794.4800 1155.4600 2794.9600 ;
        RECT 1152.4600 2805.3600 1155.4600 2805.8400 ;
        RECT 1164.2200 2805.3600 1165.8200 2805.8400 ;
        RECT 1164.2200 2783.6000 1165.8200 2784.0800 ;
        RECT 1164.2200 2789.0400 1165.8200 2789.5200 ;
        RECT 1152.4600 2789.0400 1155.4600 2789.5200 ;
        RECT 1152.4600 2783.6000 1155.4600 2784.0800 ;
        RECT 1164.2200 2767.2800 1165.8200 2767.7600 ;
        RECT 1164.2200 2772.7200 1165.8200 2773.2000 ;
        RECT 1152.4600 2772.7200 1155.4600 2773.2000 ;
        RECT 1152.4600 2767.2800 1155.4600 2767.7600 ;
        RECT 1152.4600 2778.1600 1155.4600 2778.6400 ;
        RECT 1164.2200 2778.1600 1165.8200 2778.6400 ;
        RECT 1254.2200 2750.9600 1255.8200 2751.4400 ;
        RECT 1254.2200 2756.4000 1255.8200 2756.8800 ;
        RECT 1254.2200 2761.8400 1255.8200 2762.3200 ;
        RECT 1254.2200 2740.0800 1255.8200 2740.5600 ;
        RECT 1254.2200 2745.5200 1255.8200 2746.0000 ;
        RECT 1209.2200 2750.9600 1210.8200 2751.4400 ;
        RECT 1209.2200 2756.4000 1210.8200 2756.8800 ;
        RECT 1209.2200 2761.8400 1210.8200 2762.3200 ;
        RECT 1209.2200 2740.0800 1210.8200 2740.5600 ;
        RECT 1209.2200 2745.5200 1210.8200 2746.0000 ;
        RECT 1254.2200 2723.7600 1255.8200 2724.2400 ;
        RECT 1254.2200 2729.2000 1255.8200 2729.6800 ;
        RECT 1254.2200 2734.6400 1255.8200 2735.1200 ;
        RECT 1254.2200 2712.8800 1255.8200 2713.3600 ;
        RECT 1254.2200 2718.3200 1255.8200 2718.8000 ;
        RECT 1209.2200 2723.7600 1210.8200 2724.2400 ;
        RECT 1209.2200 2729.2000 1210.8200 2729.6800 ;
        RECT 1209.2200 2734.6400 1210.8200 2735.1200 ;
        RECT 1209.2200 2712.8800 1210.8200 2713.3600 ;
        RECT 1209.2200 2718.3200 1210.8200 2718.8000 ;
        RECT 1164.2200 2750.9600 1165.8200 2751.4400 ;
        RECT 1164.2200 2756.4000 1165.8200 2756.8800 ;
        RECT 1164.2200 2761.8400 1165.8200 2762.3200 ;
        RECT 1152.4600 2750.9600 1155.4600 2751.4400 ;
        RECT 1152.4600 2756.4000 1155.4600 2756.8800 ;
        RECT 1152.4600 2761.8400 1155.4600 2762.3200 ;
        RECT 1164.2200 2740.0800 1165.8200 2740.5600 ;
        RECT 1164.2200 2745.5200 1165.8200 2746.0000 ;
        RECT 1152.4600 2740.0800 1155.4600 2740.5600 ;
        RECT 1152.4600 2745.5200 1155.4600 2746.0000 ;
        RECT 1164.2200 2723.7600 1165.8200 2724.2400 ;
        RECT 1164.2200 2729.2000 1165.8200 2729.6800 ;
        RECT 1164.2200 2734.6400 1165.8200 2735.1200 ;
        RECT 1152.4600 2723.7600 1155.4600 2724.2400 ;
        RECT 1152.4600 2729.2000 1155.4600 2729.6800 ;
        RECT 1152.4600 2734.6400 1155.4600 2735.1200 ;
        RECT 1164.2200 2712.8800 1165.8200 2713.3600 ;
        RECT 1164.2200 2718.3200 1165.8200 2718.8000 ;
        RECT 1152.4600 2712.8800 1155.4600 2713.3600 ;
        RECT 1152.4600 2718.3200 1155.4600 2718.8000 ;
        RECT 1356.5600 2696.5600 1359.5600 2697.0400 ;
        RECT 1356.5600 2702.0000 1359.5600 2702.4800 ;
        RECT 1356.5600 2707.4400 1359.5600 2707.9200 ;
        RECT 1344.2200 2696.5600 1345.8200 2697.0400 ;
        RECT 1344.2200 2702.0000 1345.8200 2702.4800 ;
        RECT 1344.2200 2707.4400 1345.8200 2707.9200 ;
        RECT 1356.5600 2685.6800 1359.5600 2686.1600 ;
        RECT 1356.5600 2691.1200 1359.5600 2691.6000 ;
        RECT 1344.2200 2685.6800 1345.8200 2686.1600 ;
        RECT 1344.2200 2691.1200 1345.8200 2691.6000 ;
        RECT 1356.5600 2669.3600 1359.5600 2669.8400 ;
        RECT 1356.5600 2674.8000 1359.5600 2675.2800 ;
        RECT 1356.5600 2680.2400 1359.5600 2680.7200 ;
        RECT 1344.2200 2669.3600 1345.8200 2669.8400 ;
        RECT 1344.2200 2674.8000 1345.8200 2675.2800 ;
        RECT 1344.2200 2680.2400 1345.8200 2680.7200 ;
        RECT 1356.5600 2658.4800 1359.5600 2658.9600 ;
        RECT 1356.5600 2663.9200 1359.5600 2664.4000 ;
        RECT 1344.2200 2658.4800 1345.8200 2658.9600 ;
        RECT 1344.2200 2663.9200 1345.8200 2664.4000 ;
        RECT 1299.2200 2696.5600 1300.8200 2697.0400 ;
        RECT 1299.2200 2702.0000 1300.8200 2702.4800 ;
        RECT 1299.2200 2707.4400 1300.8200 2707.9200 ;
        RECT 1299.2200 2685.6800 1300.8200 2686.1600 ;
        RECT 1299.2200 2691.1200 1300.8200 2691.6000 ;
        RECT 1299.2200 2669.3600 1300.8200 2669.8400 ;
        RECT 1299.2200 2674.8000 1300.8200 2675.2800 ;
        RECT 1299.2200 2680.2400 1300.8200 2680.7200 ;
        RECT 1299.2200 2658.4800 1300.8200 2658.9600 ;
        RECT 1299.2200 2663.9200 1300.8200 2664.4000 ;
        RECT 1356.5600 2642.1600 1359.5600 2642.6400 ;
        RECT 1356.5600 2647.6000 1359.5600 2648.0800 ;
        RECT 1356.5600 2653.0400 1359.5600 2653.5200 ;
        RECT 1344.2200 2642.1600 1345.8200 2642.6400 ;
        RECT 1344.2200 2647.6000 1345.8200 2648.0800 ;
        RECT 1344.2200 2653.0400 1345.8200 2653.5200 ;
        RECT 1356.5600 2631.2800 1359.5600 2631.7600 ;
        RECT 1356.5600 2636.7200 1359.5600 2637.2000 ;
        RECT 1344.2200 2631.2800 1345.8200 2631.7600 ;
        RECT 1344.2200 2636.7200 1345.8200 2637.2000 ;
        RECT 1356.5600 2614.9600 1359.5600 2615.4400 ;
        RECT 1356.5600 2620.4000 1359.5600 2620.8800 ;
        RECT 1356.5600 2625.8400 1359.5600 2626.3200 ;
        RECT 1344.2200 2614.9600 1345.8200 2615.4400 ;
        RECT 1344.2200 2620.4000 1345.8200 2620.8800 ;
        RECT 1344.2200 2625.8400 1345.8200 2626.3200 ;
        RECT 1356.5600 2609.5200 1359.5600 2610.0000 ;
        RECT 1344.2200 2609.5200 1345.8200 2610.0000 ;
        RECT 1299.2200 2642.1600 1300.8200 2642.6400 ;
        RECT 1299.2200 2647.6000 1300.8200 2648.0800 ;
        RECT 1299.2200 2653.0400 1300.8200 2653.5200 ;
        RECT 1299.2200 2631.2800 1300.8200 2631.7600 ;
        RECT 1299.2200 2636.7200 1300.8200 2637.2000 ;
        RECT 1299.2200 2614.9600 1300.8200 2615.4400 ;
        RECT 1299.2200 2620.4000 1300.8200 2620.8800 ;
        RECT 1299.2200 2625.8400 1300.8200 2626.3200 ;
        RECT 1299.2200 2609.5200 1300.8200 2610.0000 ;
        RECT 1254.2200 2696.5600 1255.8200 2697.0400 ;
        RECT 1254.2200 2702.0000 1255.8200 2702.4800 ;
        RECT 1254.2200 2707.4400 1255.8200 2707.9200 ;
        RECT 1254.2200 2685.6800 1255.8200 2686.1600 ;
        RECT 1254.2200 2691.1200 1255.8200 2691.6000 ;
        RECT 1209.2200 2696.5600 1210.8200 2697.0400 ;
        RECT 1209.2200 2702.0000 1210.8200 2702.4800 ;
        RECT 1209.2200 2707.4400 1210.8200 2707.9200 ;
        RECT 1209.2200 2685.6800 1210.8200 2686.1600 ;
        RECT 1209.2200 2691.1200 1210.8200 2691.6000 ;
        RECT 1254.2200 2669.3600 1255.8200 2669.8400 ;
        RECT 1254.2200 2674.8000 1255.8200 2675.2800 ;
        RECT 1254.2200 2680.2400 1255.8200 2680.7200 ;
        RECT 1254.2200 2658.4800 1255.8200 2658.9600 ;
        RECT 1254.2200 2663.9200 1255.8200 2664.4000 ;
        RECT 1209.2200 2669.3600 1210.8200 2669.8400 ;
        RECT 1209.2200 2674.8000 1210.8200 2675.2800 ;
        RECT 1209.2200 2680.2400 1210.8200 2680.7200 ;
        RECT 1209.2200 2658.4800 1210.8200 2658.9600 ;
        RECT 1209.2200 2663.9200 1210.8200 2664.4000 ;
        RECT 1164.2200 2696.5600 1165.8200 2697.0400 ;
        RECT 1164.2200 2702.0000 1165.8200 2702.4800 ;
        RECT 1164.2200 2707.4400 1165.8200 2707.9200 ;
        RECT 1152.4600 2696.5600 1155.4600 2697.0400 ;
        RECT 1152.4600 2702.0000 1155.4600 2702.4800 ;
        RECT 1152.4600 2707.4400 1155.4600 2707.9200 ;
        RECT 1164.2200 2685.6800 1165.8200 2686.1600 ;
        RECT 1164.2200 2691.1200 1165.8200 2691.6000 ;
        RECT 1152.4600 2685.6800 1155.4600 2686.1600 ;
        RECT 1152.4600 2691.1200 1155.4600 2691.6000 ;
        RECT 1164.2200 2669.3600 1165.8200 2669.8400 ;
        RECT 1164.2200 2674.8000 1165.8200 2675.2800 ;
        RECT 1164.2200 2680.2400 1165.8200 2680.7200 ;
        RECT 1152.4600 2669.3600 1155.4600 2669.8400 ;
        RECT 1152.4600 2674.8000 1155.4600 2675.2800 ;
        RECT 1152.4600 2680.2400 1155.4600 2680.7200 ;
        RECT 1164.2200 2658.4800 1165.8200 2658.9600 ;
        RECT 1164.2200 2663.9200 1165.8200 2664.4000 ;
        RECT 1152.4600 2658.4800 1155.4600 2658.9600 ;
        RECT 1152.4600 2663.9200 1155.4600 2664.4000 ;
        RECT 1254.2200 2642.1600 1255.8200 2642.6400 ;
        RECT 1254.2200 2647.6000 1255.8200 2648.0800 ;
        RECT 1254.2200 2653.0400 1255.8200 2653.5200 ;
        RECT 1254.2200 2631.2800 1255.8200 2631.7600 ;
        RECT 1254.2200 2636.7200 1255.8200 2637.2000 ;
        RECT 1209.2200 2642.1600 1210.8200 2642.6400 ;
        RECT 1209.2200 2647.6000 1210.8200 2648.0800 ;
        RECT 1209.2200 2653.0400 1210.8200 2653.5200 ;
        RECT 1209.2200 2631.2800 1210.8200 2631.7600 ;
        RECT 1209.2200 2636.7200 1210.8200 2637.2000 ;
        RECT 1254.2200 2614.9600 1255.8200 2615.4400 ;
        RECT 1254.2200 2620.4000 1255.8200 2620.8800 ;
        RECT 1254.2200 2625.8400 1255.8200 2626.3200 ;
        RECT 1254.2200 2609.5200 1255.8200 2610.0000 ;
        RECT 1209.2200 2614.9600 1210.8200 2615.4400 ;
        RECT 1209.2200 2620.4000 1210.8200 2620.8800 ;
        RECT 1209.2200 2625.8400 1210.8200 2626.3200 ;
        RECT 1209.2200 2609.5200 1210.8200 2610.0000 ;
        RECT 1164.2200 2642.1600 1165.8200 2642.6400 ;
        RECT 1164.2200 2647.6000 1165.8200 2648.0800 ;
        RECT 1164.2200 2653.0400 1165.8200 2653.5200 ;
        RECT 1152.4600 2642.1600 1155.4600 2642.6400 ;
        RECT 1152.4600 2647.6000 1155.4600 2648.0800 ;
        RECT 1152.4600 2653.0400 1155.4600 2653.5200 ;
        RECT 1164.2200 2631.2800 1165.8200 2631.7600 ;
        RECT 1164.2200 2636.7200 1165.8200 2637.2000 ;
        RECT 1152.4600 2631.2800 1155.4600 2631.7600 ;
        RECT 1152.4600 2636.7200 1155.4600 2637.2000 ;
        RECT 1164.2200 2614.9600 1165.8200 2615.4400 ;
        RECT 1164.2200 2620.4000 1165.8200 2620.8800 ;
        RECT 1164.2200 2625.8400 1165.8200 2626.3200 ;
        RECT 1152.4600 2614.9600 1155.4600 2615.4400 ;
        RECT 1152.4600 2620.4000 1155.4600 2620.8800 ;
        RECT 1152.4600 2625.8400 1155.4600 2626.3200 ;
        RECT 1152.4600 2609.5200 1155.4600 2610.0000 ;
        RECT 1164.2200 2609.5200 1165.8200 2610.0000 ;
        RECT 1152.4600 2814.4300 1359.5600 2817.4300 ;
        RECT 1152.4600 2601.3300 1359.5600 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 2371.6900 1345.8200 2587.7900 ;
        RECT 1299.2200 2371.6900 1300.8200 2587.7900 ;
        RECT 1254.2200 2371.6900 1255.8200 2587.7900 ;
        RECT 1209.2200 2371.6900 1210.8200 2587.7900 ;
        RECT 1164.2200 2371.6900 1165.8200 2587.7900 ;
        RECT 1356.5600 2371.6900 1359.5600 2587.7900 ;
        RECT 1152.4600 2371.6900 1155.4600 2587.7900 ;
      LAYER met3 ;
        RECT 1356.5600 2564.8400 1359.5600 2565.3200 ;
        RECT 1356.5600 2570.2800 1359.5600 2570.7600 ;
        RECT 1344.2200 2564.8400 1345.8200 2565.3200 ;
        RECT 1344.2200 2570.2800 1345.8200 2570.7600 ;
        RECT 1356.5600 2575.7200 1359.5600 2576.2000 ;
        RECT 1344.2200 2575.7200 1345.8200 2576.2000 ;
        RECT 1356.5600 2553.9600 1359.5600 2554.4400 ;
        RECT 1356.5600 2559.4000 1359.5600 2559.8800 ;
        RECT 1344.2200 2553.9600 1345.8200 2554.4400 ;
        RECT 1344.2200 2559.4000 1345.8200 2559.8800 ;
        RECT 1356.5600 2537.6400 1359.5600 2538.1200 ;
        RECT 1356.5600 2543.0800 1359.5600 2543.5600 ;
        RECT 1344.2200 2537.6400 1345.8200 2538.1200 ;
        RECT 1344.2200 2543.0800 1345.8200 2543.5600 ;
        RECT 1356.5600 2548.5200 1359.5600 2549.0000 ;
        RECT 1344.2200 2548.5200 1345.8200 2549.0000 ;
        RECT 1299.2200 2564.8400 1300.8200 2565.3200 ;
        RECT 1299.2200 2570.2800 1300.8200 2570.7600 ;
        RECT 1299.2200 2575.7200 1300.8200 2576.2000 ;
        RECT 1299.2200 2553.9600 1300.8200 2554.4400 ;
        RECT 1299.2200 2559.4000 1300.8200 2559.8800 ;
        RECT 1299.2200 2537.6400 1300.8200 2538.1200 ;
        RECT 1299.2200 2543.0800 1300.8200 2543.5600 ;
        RECT 1299.2200 2548.5200 1300.8200 2549.0000 ;
        RECT 1356.5600 2521.3200 1359.5600 2521.8000 ;
        RECT 1356.5600 2526.7600 1359.5600 2527.2400 ;
        RECT 1356.5600 2532.2000 1359.5600 2532.6800 ;
        RECT 1344.2200 2521.3200 1345.8200 2521.8000 ;
        RECT 1344.2200 2526.7600 1345.8200 2527.2400 ;
        RECT 1344.2200 2532.2000 1345.8200 2532.6800 ;
        RECT 1356.5600 2510.4400 1359.5600 2510.9200 ;
        RECT 1356.5600 2515.8800 1359.5600 2516.3600 ;
        RECT 1344.2200 2510.4400 1345.8200 2510.9200 ;
        RECT 1344.2200 2515.8800 1345.8200 2516.3600 ;
        RECT 1356.5600 2494.1200 1359.5600 2494.6000 ;
        RECT 1356.5600 2499.5600 1359.5600 2500.0400 ;
        RECT 1356.5600 2505.0000 1359.5600 2505.4800 ;
        RECT 1344.2200 2494.1200 1345.8200 2494.6000 ;
        RECT 1344.2200 2499.5600 1345.8200 2500.0400 ;
        RECT 1344.2200 2505.0000 1345.8200 2505.4800 ;
        RECT 1356.5600 2483.2400 1359.5600 2483.7200 ;
        RECT 1356.5600 2488.6800 1359.5600 2489.1600 ;
        RECT 1344.2200 2483.2400 1345.8200 2483.7200 ;
        RECT 1344.2200 2488.6800 1345.8200 2489.1600 ;
        RECT 1299.2200 2521.3200 1300.8200 2521.8000 ;
        RECT 1299.2200 2526.7600 1300.8200 2527.2400 ;
        RECT 1299.2200 2532.2000 1300.8200 2532.6800 ;
        RECT 1299.2200 2510.4400 1300.8200 2510.9200 ;
        RECT 1299.2200 2515.8800 1300.8200 2516.3600 ;
        RECT 1299.2200 2494.1200 1300.8200 2494.6000 ;
        RECT 1299.2200 2499.5600 1300.8200 2500.0400 ;
        RECT 1299.2200 2505.0000 1300.8200 2505.4800 ;
        RECT 1299.2200 2483.2400 1300.8200 2483.7200 ;
        RECT 1299.2200 2488.6800 1300.8200 2489.1600 ;
        RECT 1254.2200 2564.8400 1255.8200 2565.3200 ;
        RECT 1254.2200 2570.2800 1255.8200 2570.7600 ;
        RECT 1254.2200 2575.7200 1255.8200 2576.2000 ;
        RECT 1209.2200 2564.8400 1210.8200 2565.3200 ;
        RECT 1209.2200 2570.2800 1210.8200 2570.7600 ;
        RECT 1209.2200 2575.7200 1210.8200 2576.2000 ;
        RECT 1254.2200 2553.9600 1255.8200 2554.4400 ;
        RECT 1254.2200 2559.4000 1255.8200 2559.8800 ;
        RECT 1254.2200 2537.6400 1255.8200 2538.1200 ;
        RECT 1254.2200 2543.0800 1255.8200 2543.5600 ;
        RECT 1254.2200 2548.5200 1255.8200 2549.0000 ;
        RECT 1209.2200 2553.9600 1210.8200 2554.4400 ;
        RECT 1209.2200 2559.4000 1210.8200 2559.8800 ;
        RECT 1209.2200 2537.6400 1210.8200 2538.1200 ;
        RECT 1209.2200 2543.0800 1210.8200 2543.5600 ;
        RECT 1209.2200 2548.5200 1210.8200 2549.0000 ;
        RECT 1164.2200 2564.8400 1165.8200 2565.3200 ;
        RECT 1164.2200 2570.2800 1165.8200 2570.7600 ;
        RECT 1152.4600 2570.2800 1155.4600 2570.7600 ;
        RECT 1152.4600 2564.8400 1155.4600 2565.3200 ;
        RECT 1152.4600 2575.7200 1155.4600 2576.2000 ;
        RECT 1164.2200 2575.7200 1165.8200 2576.2000 ;
        RECT 1164.2200 2553.9600 1165.8200 2554.4400 ;
        RECT 1164.2200 2559.4000 1165.8200 2559.8800 ;
        RECT 1152.4600 2559.4000 1155.4600 2559.8800 ;
        RECT 1152.4600 2553.9600 1155.4600 2554.4400 ;
        RECT 1164.2200 2537.6400 1165.8200 2538.1200 ;
        RECT 1164.2200 2543.0800 1165.8200 2543.5600 ;
        RECT 1152.4600 2543.0800 1155.4600 2543.5600 ;
        RECT 1152.4600 2537.6400 1155.4600 2538.1200 ;
        RECT 1152.4600 2548.5200 1155.4600 2549.0000 ;
        RECT 1164.2200 2548.5200 1165.8200 2549.0000 ;
        RECT 1254.2200 2521.3200 1255.8200 2521.8000 ;
        RECT 1254.2200 2526.7600 1255.8200 2527.2400 ;
        RECT 1254.2200 2532.2000 1255.8200 2532.6800 ;
        RECT 1254.2200 2510.4400 1255.8200 2510.9200 ;
        RECT 1254.2200 2515.8800 1255.8200 2516.3600 ;
        RECT 1209.2200 2521.3200 1210.8200 2521.8000 ;
        RECT 1209.2200 2526.7600 1210.8200 2527.2400 ;
        RECT 1209.2200 2532.2000 1210.8200 2532.6800 ;
        RECT 1209.2200 2510.4400 1210.8200 2510.9200 ;
        RECT 1209.2200 2515.8800 1210.8200 2516.3600 ;
        RECT 1254.2200 2494.1200 1255.8200 2494.6000 ;
        RECT 1254.2200 2499.5600 1255.8200 2500.0400 ;
        RECT 1254.2200 2505.0000 1255.8200 2505.4800 ;
        RECT 1254.2200 2483.2400 1255.8200 2483.7200 ;
        RECT 1254.2200 2488.6800 1255.8200 2489.1600 ;
        RECT 1209.2200 2494.1200 1210.8200 2494.6000 ;
        RECT 1209.2200 2499.5600 1210.8200 2500.0400 ;
        RECT 1209.2200 2505.0000 1210.8200 2505.4800 ;
        RECT 1209.2200 2483.2400 1210.8200 2483.7200 ;
        RECT 1209.2200 2488.6800 1210.8200 2489.1600 ;
        RECT 1164.2200 2521.3200 1165.8200 2521.8000 ;
        RECT 1164.2200 2526.7600 1165.8200 2527.2400 ;
        RECT 1164.2200 2532.2000 1165.8200 2532.6800 ;
        RECT 1152.4600 2521.3200 1155.4600 2521.8000 ;
        RECT 1152.4600 2526.7600 1155.4600 2527.2400 ;
        RECT 1152.4600 2532.2000 1155.4600 2532.6800 ;
        RECT 1164.2200 2510.4400 1165.8200 2510.9200 ;
        RECT 1164.2200 2515.8800 1165.8200 2516.3600 ;
        RECT 1152.4600 2510.4400 1155.4600 2510.9200 ;
        RECT 1152.4600 2515.8800 1155.4600 2516.3600 ;
        RECT 1164.2200 2494.1200 1165.8200 2494.6000 ;
        RECT 1164.2200 2499.5600 1165.8200 2500.0400 ;
        RECT 1164.2200 2505.0000 1165.8200 2505.4800 ;
        RECT 1152.4600 2494.1200 1155.4600 2494.6000 ;
        RECT 1152.4600 2499.5600 1155.4600 2500.0400 ;
        RECT 1152.4600 2505.0000 1155.4600 2505.4800 ;
        RECT 1164.2200 2483.2400 1165.8200 2483.7200 ;
        RECT 1164.2200 2488.6800 1165.8200 2489.1600 ;
        RECT 1152.4600 2483.2400 1155.4600 2483.7200 ;
        RECT 1152.4600 2488.6800 1155.4600 2489.1600 ;
        RECT 1356.5600 2466.9200 1359.5600 2467.4000 ;
        RECT 1356.5600 2472.3600 1359.5600 2472.8400 ;
        RECT 1356.5600 2477.8000 1359.5600 2478.2800 ;
        RECT 1344.2200 2466.9200 1345.8200 2467.4000 ;
        RECT 1344.2200 2472.3600 1345.8200 2472.8400 ;
        RECT 1344.2200 2477.8000 1345.8200 2478.2800 ;
        RECT 1356.5600 2456.0400 1359.5600 2456.5200 ;
        RECT 1356.5600 2461.4800 1359.5600 2461.9600 ;
        RECT 1344.2200 2456.0400 1345.8200 2456.5200 ;
        RECT 1344.2200 2461.4800 1345.8200 2461.9600 ;
        RECT 1356.5600 2439.7200 1359.5600 2440.2000 ;
        RECT 1356.5600 2445.1600 1359.5600 2445.6400 ;
        RECT 1356.5600 2450.6000 1359.5600 2451.0800 ;
        RECT 1344.2200 2439.7200 1345.8200 2440.2000 ;
        RECT 1344.2200 2445.1600 1345.8200 2445.6400 ;
        RECT 1344.2200 2450.6000 1345.8200 2451.0800 ;
        RECT 1356.5600 2428.8400 1359.5600 2429.3200 ;
        RECT 1356.5600 2434.2800 1359.5600 2434.7600 ;
        RECT 1344.2200 2428.8400 1345.8200 2429.3200 ;
        RECT 1344.2200 2434.2800 1345.8200 2434.7600 ;
        RECT 1299.2200 2466.9200 1300.8200 2467.4000 ;
        RECT 1299.2200 2472.3600 1300.8200 2472.8400 ;
        RECT 1299.2200 2477.8000 1300.8200 2478.2800 ;
        RECT 1299.2200 2456.0400 1300.8200 2456.5200 ;
        RECT 1299.2200 2461.4800 1300.8200 2461.9600 ;
        RECT 1299.2200 2439.7200 1300.8200 2440.2000 ;
        RECT 1299.2200 2445.1600 1300.8200 2445.6400 ;
        RECT 1299.2200 2450.6000 1300.8200 2451.0800 ;
        RECT 1299.2200 2428.8400 1300.8200 2429.3200 ;
        RECT 1299.2200 2434.2800 1300.8200 2434.7600 ;
        RECT 1356.5600 2412.5200 1359.5600 2413.0000 ;
        RECT 1356.5600 2417.9600 1359.5600 2418.4400 ;
        RECT 1356.5600 2423.4000 1359.5600 2423.8800 ;
        RECT 1344.2200 2412.5200 1345.8200 2413.0000 ;
        RECT 1344.2200 2417.9600 1345.8200 2418.4400 ;
        RECT 1344.2200 2423.4000 1345.8200 2423.8800 ;
        RECT 1356.5600 2401.6400 1359.5600 2402.1200 ;
        RECT 1356.5600 2407.0800 1359.5600 2407.5600 ;
        RECT 1344.2200 2401.6400 1345.8200 2402.1200 ;
        RECT 1344.2200 2407.0800 1345.8200 2407.5600 ;
        RECT 1356.5600 2385.3200 1359.5600 2385.8000 ;
        RECT 1356.5600 2390.7600 1359.5600 2391.2400 ;
        RECT 1356.5600 2396.2000 1359.5600 2396.6800 ;
        RECT 1344.2200 2385.3200 1345.8200 2385.8000 ;
        RECT 1344.2200 2390.7600 1345.8200 2391.2400 ;
        RECT 1344.2200 2396.2000 1345.8200 2396.6800 ;
        RECT 1356.5600 2379.8800 1359.5600 2380.3600 ;
        RECT 1344.2200 2379.8800 1345.8200 2380.3600 ;
        RECT 1299.2200 2412.5200 1300.8200 2413.0000 ;
        RECT 1299.2200 2417.9600 1300.8200 2418.4400 ;
        RECT 1299.2200 2423.4000 1300.8200 2423.8800 ;
        RECT 1299.2200 2401.6400 1300.8200 2402.1200 ;
        RECT 1299.2200 2407.0800 1300.8200 2407.5600 ;
        RECT 1299.2200 2385.3200 1300.8200 2385.8000 ;
        RECT 1299.2200 2390.7600 1300.8200 2391.2400 ;
        RECT 1299.2200 2396.2000 1300.8200 2396.6800 ;
        RECT 1299.2200 2379.8800 1300.8200 2380.3600 ;
        RECT 1254.2200 2466.9200 1255.8200 2467.4000 ;
        RECT 1254.2200 2472.3600 1255.8200 2472.8400 ;
        RECT 1254.2200 2477.8000 1255.8200 2478.2800 ;
        RECT 1254.2200 2456.0400 1255.8200 2456.5200 ;
        RECT 1254.2200 2461.4800 1255.8200 2461.9600 ;
        RECT 1209.2200 2466.9200 1210.8200 2467.4000 ;
        RECT 1209.2200 2472.3600 1210.8200 2472.8400 ;
        RECT 1209.2200 2477.8000 1210.8200 2478.2800 ;
        RECT 1209.2200 2456.0400 1210.8200 2456.5200 ;
        RECT 1209.2200 2461.4800 1210.8200 2461.9600 ;
        RECT 1254.2200 2439.7200 1255.8200 2440.2000 ;
        RECT 1254.2200 2445.1600 1255.8200 2445.6400 ;
        RECT 1254.2200 2450.6000 1255.8200 2451.0800 ;
        RECT 1254.2200 2428.8400 1255.8200 2429.3200 ;
        RECT 1254.2200 2434.2800 1255.8200 2434.7600 ;
        RECT 1209.2200 2439.7200 1210.8200 2440.2000 ;
        RECT 1209.2200 2445.1600 1210.8200 2445.6400 ;
        RECT 1209.2200 2450.6000 1210.8200 2451.0800 ;
        RECT 1209.2200 2428.8400 1210.8200 2429.3200 ;
        RECT 1209.2200 2434.2800 1210.8200 2434.7600 ;
        RECT 1164.2200 2466.9200 1165.8200 2467.4000 ;
        RECT 1164.2200 2472.3600 1165.8200 2472.8400 ;
        RECT 1164.2200 2477.8000 1165.8200 2478.2800 ;
        RECT 1152.4600 2466.9200 1155.4600 2467.4000 ;
        RECT 1152.4600 2472.3600 1155.4600 2472.8400 ;
        RECT 1152.4600 2477.8000 1155.4600 2478.2800 ;
        RECT 1164.2200 2456.0400 1165.8200 2456.5200 ;
        RECT 1164.2200 2461.4800 1165.8200 2461.9600 ;
        RECT 1152.4600 2456.0400 1155.4600 2456.5200 ;
        RECT 1152.4600 2461.4800 1155.4600 2461.9600 ;
        RECT 1164.2200 2439.7200 1165.8200 2440.2000 ;
        RECT 1164.2200 2445.1600 1165.8200 2445.6400 ;
        RECT 1164.2200 2450.6000 1165.8200 2451.0800 ;
        RECT 1152.4600 2439.7200 1155.4600 2440.2000 ;
        RECT 1152.4600 2445.1600 1155.4600 2445.6400 ;
        RECT 1152.4600 2450.6000 1155.4600 2451.0800 ;
        RECT 1164.2200 2428.8400 1165.8200 2429.3200 ;
        RECT 1164.2200 2434.2800 1165.8200 2434.7600 ;
        RECT 1152.4600 2428.8400 1155.4600 2429.3200 ;
        RECT 1152.4600 2434.2800 1155.4600 2434.7600 ;
        RECT 1254.2200 2412.5200 1255.8200 2413.0000 ;
        RECT 1254.2200 2417.9600 1255.8200 2418.4400 ;
        RECT 1254.2200 2423.4000 1255.8200 2423.8800 ;
        RECT 1254.2200 2401.6400 1255.8200 2402.1200 ;
        RECT 1254.2200 2407.0800 1255.8200 2407.5600 ;
        RECT 1209.2200 2412.5200 1210.8200 2413.0000 ;
        RECT 1209.2200 2417.9600 1210.8200 2418.4400 ;
        RECT 1209.2200 2423.4000 1210.8200 2423.8800 ;
        RECT 1209.2200 2401.6400 1210.8200 2402.1200 ;
        RECT 1209.2200 2407.0800 1210.8200 2407.5600 ;
        RECT 1254.2200 2385.3200 1255.8200 2385.8000 ;
        RECT 1254.2200 2390.7600 1255.8200 2391.2400 ;
        RECT 1254.2200 2396.2000 1255.8200 2396.6800 ;
        RECT 1254.2200 2379.8800 1255.8200 2380.3600 ;
        RECT 1209.2200 2385.3200 1210.8200 2385.8000 ;
        RECT 1209.2200 2390.7600 1210.8200 2391.2400 ;
        RECT 1209.2200 2396.2000 1210.8200 2396.6800 ;
        RECT 1209.2200 2379.8800 1210.8200 2380.3600 ;
        RECT 1164.2200 2412.5200 1165.8200 2413.0000 ;
        RECT 1164.2200 2417.9600 1165.8200 2418.4400 ;
        RECT 1164.2200 2423.4000 1165.8200 2423.8800 ;
        RECT 1152.4600 2412.5200 1155.4600 2413.0000 ;
        RECT 1152.4600 2417.9600 1155.4600 2418.4400 ;
        RECT 1152.4600 2423.4000 1155.4600 2423.8800 ;
        RECT 1164.2200 2401.6400 1165.8200 2402.1200 ;
        RECT 1164.2200 2407.0800 1165.8200 2407.5600 ;
        RECT 1152.4600 2401.6400 1155.4600 2402.1200 ;
        RECT 1152.4600 2407.0800 1155.4600 2407.5600 ;
        RECT 1164.2200 2385.3200 1165.8200 2385.8000 ;
        RECT 1164.2200 2390.7600 1165.8200 2391.2400 ;
        RECT 1164.2200 2396.2000 1165.8200 2396.6800 ;
        RECT 1152.4600 2385.3200 1155.4600 2385.8000 ;
        RECT 1152.4600 2390.7600 1155.4600 2391.2400 ;
        RECT 1152.4600 2396.2000 1155.4600 2396.6800 ;
        RECT 1152.4600 2379.8800 1155.4600 2380.3600 ;
        RECT 1164.2200 2379.8800 1165.8200 2380.3600 ;
        RECT 1152.4600 2584.7900 1359.5600 2587.7900 ;
        RECT 1152.4600 2371.6900 1359.5600 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 2142.0500 1345.8200 2358.1500 ;
        RECT 1299.2200 2142.0500 1300.8200 2358.1500 ;
        RECT 1254.2200 2142.0500 1255.8200 2358.1500 ;
        RECT 1209.2200 2142.0500 1210.8200 2358.1500 ;
        RECT 1164.2200 2142.0500 1165.8200 2358.1500 ;
        RECT 1356.5600 2142.0500 1359.5600 2358.1500 ;
        RECT 1152.4600 2142.0500 1155.4600 2358.1500 ;
      LAYER met3 ;
        RECT 1356.5600 2335.2000 1359.5600 2335.6800 ;
        RECT 1356.5600 2340.6400 1359.5600 2341.1200 ;
        RECT 1344.2200 2335.2000 1345.8200 2335.6800 ;
        RECT 1344.2200 2340.6400 1345.8200 2341.1200 ;
        RECT 1356.5600 2346.0800 1359.5600 2346.5600 ;
        RECT 1344.2200 2346.0800 1345.8200 2346.5600 ;
        RECT 1356.5600 2324.3200 1359.5600 2324.8000 ;
        RECT 1356.5600 2329.7600 1359.5600 2330.2400 ;
        RECT 1344.2200 2324.3200 1345.8200 2324.8000 ;
        RECT 1344.2200 2329.7600 1345.8200 2330.2400 ;
        RECT 1356.5600 2308.0000 1359.5600 2308.4800 ;
        RECT 1356.5600 2313.4400 1359.5600 2313.9200 ;
        RECT 1344.2200 2308.0000 1345.8200 2308.4800 ;
        RECT 1344.2200 2313.4400 1345.8200 2313.9200 ;
        RECT 1356.5600 2318.8800 1359.5600 2319.3600 ;
        RECT 1344.2200 2318.8800 1345.8200 2319.3600 ;
        RECT 1299.2200 2335.2000 1300.8200 2335.6800 ;
        RECT 1299.2200 2340.6400 1300.8200 2341.1200 ;
        RECT 1299.2200 2346.0800 1300.8200 2346.5600 ;
        RECT 1299.2200 2324.3200 1300.8200 2324.8000 ;
        RECT 1299.2200 2329.7600 1300.8200 2330.2400 ;
        RECT 1299.2200 2308.0000 1300.8200 2308.4800 ;
        RECT 1299.2200 2313.4400 1300.8200 2313.9200 ;
        RECT 1299.2200 2318.8800 1300.8200 2319.3600 ;
        RECT 1356.5600 2291.6800 1359.5600 2292.1600 ;
        RECT 1356.5600 2297.1200 1359.5600 2297.6000 ;
        RECT 1356.5600 2302.5600 1359.5600 2303.0400 ;
        RECT 1344.2200 2291.6800 1345.8200 2292.1600 ;
        RECT 1344.2200 2297.1200 1345.8200 2297.6000 ;
        RECT 1344.2200 2302.5600 1345.8200 2303.0400 ;
        RECT 1356.5600 2280.8000 1359.5600 2281.2800 ;
        RECT 1356.5600 2286.2400 1359.5600 2286.7200 ;
        RECT 1344.2200 2280.8000 1345.8200 2281.2800 ;
        RECT 1344.2200 2286.2400 1345.8200 2286.7200 ;
        RECT 1356.5600 2264.4800 1359.5600 2264.9600 ;
        RECT 1356.5600 2269.9200 1359.5600 2270.4000 ;
        RECT 1356.5600 2275.3600 1359.5600 2275.8400 ;
        RECT 1344.2200 2264.4800 1345.8200 2264.9600 ;
        RECT 1344.2200 2269.9200 1345.8200 2270.4000 ;
        RECT 1344.2200 2275.3600 1345.8200 2275.8400 ;
        RECT 1356.5600 2253.6000 1359.5600 2254.0800 ;
        RECT 1356.5600 2259.0400 1359.5600 2259.5200 ;
        RECT 1344.2200 2253.6000 1345.8200 2254.0800 ;
        RECT 1344.2200 2259.0400 1345.8200 2259.5200 ;
        RECT 1299.2200 2291.6800 1300.8200 2292.1600 ;
        RECT 1299.2200 2297.1200 1300.8200 2297.6000 ;
        RECT 1299.2200 2302.5600 1300.8200 2303.0400 ;
        RECT 1299.2200 2280.8000 1300.8200 2281.2800 ;
        RECT 1299.2200 2286.2400 1300.8200 2286.7200 ;
        RECT 1299.2200 2264.4800 1300.8200 2264.9600 ;
        RECT 1299.2200 2269.9200 1300.8200 2270.4000 ;
        RECT 1299.2200 2275.3600 1300.8200 2275.8400 ;
        RECT 1299.2200 2253.6000 1300.8200 2254.0800 ;
        RECT 1299.2200 2259.0400 1300.8200 2259.5200 ;
        RECT 1254.2200 2335.2000 1255.8200 2335.6800 ;
        RECT 1254.2200 2340.6400 1255.8200 2341.1200 ;
        RECT 1254.2200 2346.0800 1255.8200 2346.5600 ;
        RECT 1209.2200 2335.2000 1210.8200 2335.6800 ;
        RECT 1209.2200 2340.6400 1210.8200 2341.1200 ;
        RECT 1209.2200 2346.0800 1210.8200 2346.5600 ;
        RECT 1254.2200 2324.3200 1255.8200 2324.8000 ;
        RECT 1254.2200 2329.7600 1255.8200 2330.2400 ;
        RECT 1254.2200 2308.0000 1255.8200 2308.4800 ;
        RECT 1254.2200 2313.4400 1255.8200 2313.9200 ;
        RECT 1254.2200 2318.8800 1255.8200 2319.3600 ;
        RECT 1209.2200 2324.3200 1210.8200 2324.8000 ;
        RECT 1209.2200 2329.7600 1210.8200 2330.2400 ;
        RECT 1209.2200 2308.0000 1210.8200 2308.4800 ;
        RECT 1209.2200 2313.4400 1210.8200 2313.9200 ;
        RECT 1209.2200 2318.8800 1210.8200 2319.3600 ;
        RECT 1164.2200 2335.2000 1165.8200 2335.6800 ;
        RECT 1164.2200 2340.6400 1165.8200 2341.1200 ;
        RECT 1152.4600 2340.6400 1155.4600 2341.1200 ;
        RECT 1152.4600 2335.2000 1155.4600 2335.6800 ;
        RECT 1152.4600 2346.0800 1155.4600 2346.5600 ;
        RECT 1164.2200 2346.0800 1165.8200 2346.5600 ;
        RECT 1164.2200 2324.3200 1165.8200 2324.8000 ;
        RECT 1164.2200 2329.7600 1165.8200 2330.2400 ;
        RECT 1152.4600 2329.7600 1155.4600 2330.2400 ;
        RECT 1152.4600 2324.3200 1155.4600 2324.8000 ;
        RECT 1164.2200 2308.0000 1165.8200 2308.4800 ;
        RECT 1164.2200 2313.4400 1165.8200 2313.9200 ;
        RECT 1152.4600 2313.4400 1155.4600 2313.9200 ;
        RECT 1152.4600 2308.0000 1155.4600 2308.4800 ;
        RECT 1152.4600 2318.8800 1155.4600 2319.3600 ;
        RECT 1164.2200 2318.8800 1165.8200 2319.3600 ;
        RECT 1254.2200 2291.6800 1255.8200 2292.1600 ;
        RECT 1254.2200 2297.1200 1255.8200 2297.6000 ;
        RECT 1254.2200 2302.5600 1255.8200 2303.0400 ;
        RECT 1254.2200 2280.8000 1255.8200 2281.2800 ;
        RECT 1254.2200 2286.2400 1255.8200 2286.7200 ;
        RECT 1209.2200 2291.6800 1210.8200 2292.1600 ;
        RECT 1209.2200 2297.1200 1210.8200 2297.6000 ;
        RECT 1209.2200 2302.5600 1210.8200 2303.0400 ;
        RECT 1209.2200 2280.8000 1210.8200 2281.2800 ;
        RECT 1209.2200 2286.2400 1210.8200 2286.7200 ;
        RECT 1254.2200 2264.4800 1255.8200 2264.9600 ;
        RECT 1254.2200 2269.9200 1255.8200 2270.4000 ;
        RECT 1254.2200 2275.3600 1255.8200 2275.8400 ;
        RECT 1254.2200 2253.6000 1255.8200 2254.0800 ;
        RECT 1254.2200 2259.0400 1255.8200 2259.5200 ;
        RECT 1209.2200 2264.4800 1210.8200 2264.9600 ;
        RECT 1209.2200 2269.9200 1210.8200 2270.4000 ;
        RECT 1209.2200 2275.3600 1210.8200 2275.8400 ;
        RECT 1209.2200 2253.6000 1210.8200 2254.0800 ;
        RECT 1209.2200 2259.0400 1210.8200 2259.5200 ;
        RECT 1164.2200 2291.6800 1165.8200 2292.1600 ;
        RECT 1164.2200 2297.1200 1165.8200 2297.6000 ;
        RECT 1164.2200 2302.5600 1165.8200 2303.0400 ;
        RECT 1152.4600 2291.6800 1155.4600 2292.1600 ;
        RECT 1152.4600 2297.1200 1155.4600 2297.6000 ;
        RECT 1152.4600 2302.5600 1155.4600 2303.0400 ;
        RECT 1164.2200 2280.8000 1165.8200 2281.2800 ;
        RECT 1164.2200 2286.2400 1165.8200 2286.7200 ;
        RECT 1152.4600 2280.8000 1155.4600 2281.2800 ;
        RECT 1152.4600 2286.2400 1155.4600 2286.7200 ;
        RECT 1164.2200 2264.4800 1165.8200 2264.9600 ;
        RECT 1164.2200 2269.9200 1165.8200 2270.4000 ;
        RECT 1164.2200 2275.3600 1165.8200 2275.8400 ;
        RECT 1152.4600 2264.4800 1155.4600 2264.9600 ;
        RECT 1152.4600 2269.9200 1155.4600 2270.4000 ;
        RECT 1152.4600 2275.3600 1155.4600 2275.8400 ;
        RECT 1164.2200 2253.6000 1165.8200 2254.0800 ;
        RECT 1164.2200 2259.0400 1165.8200 2259.5200 ;
        RECT 1152.4600 2253.6000 1155.4600 2254.0800 ;
        RECT 1152.4600 2259.0400 1155.4600 2259.5200 ;
        RECT 1356.5600 2237.2800 1359.5600 2237.7600 ;
        RECT 1356.5600 2242.7200 1359.5600 2243.2000 ;
        RECT 1356.5600 2248.1600 1359.5600 2248.6400 ;
        RECT 1344.2200 2237.2800 1345.8200 2237.7600 ;
        RECT 1344.2200 2242.7200 1345.8200 2243.2000 ;
        RECT 1344.2200 2248.1600 1345.8200 2248.6400 ;
        RECT 1356.5600 2226.4000 1359.5600 2226.8800 ;
        RECT 1356.5600 2231.8400 1359.5600 2232.3200 ;
        RECT 1344.2200 2226.4000 1345.8200 2226.8800 ;
        RECT 1344.2200 2231.8400 1345.8200 2232.3200 ;
        RECT 1356.5600 2210.0800 1359.5600 2210.5600 ;
        RECT 1356.5600 2215.5200 1359.5600 2216.0000 ;
        RECT 1356.5600 2220.9600 1359.5600 2221.4400 ;
        RECT 1344.2200 2210.0800 1345.8200 2210.5600 ;
        RECT 1344.2200 2215.5200 1345.8200 2216.0000 ;
        RECT 1344.2200 2220.9600 1345.8200 2221.4400 ;
        RECT 1356.5600 2199.2000 1359.5600 2199.6800 ;
        RECT 1356.5600 2204.6400 1359.5600 2205.1200 ;
        RECT 1344.2200 2199.2000 1345.8200 2199.6800 ;
        RECT 1344.2200 2204.6400 1345.8200 2205.1200 ;
        RECT 1299.2200 2237.2800 1300.8200 2237.7600 ;
        RECT 1299.2200 2242.7200 1300.8200 2243.2000 ;
        RECT 1299.2200 2248.1600 1300.8200 2248.6400 ;
        RECT 1299.2200 2226.4000 1300.8200 2226.8800 ;
        RECT 1299.2200 2231.8400 1300.8200 2232.3200 ;
        RECT 1299.2200 2210.0800 1300.8200 2210.5600 ;
        RECT 1299.2200 2215.5200 1300.8200 2216.0000 ;
        RECT 1299.2200 2220.9600 1300.8200 2221.4400 ;
        RECT 1299.2200 2199.2000 1300.8200 2199.6800 ;
        RECT 1299.2200 2204.6400 1300.8200 2205.1200 ;
        RECT 1356.5600 2182.8800 1359.5600 2183.3600 ;
        RECT 1356.5600 2188.3200 1359.5600 2188.8000 ;
        RECT 1356.5600 2193.7600 1359.5600 2194.2400 ;
        RECT 1344.2200 2182.8800 1345.8200 2183.3600 ;
        RECT 1344.2200 2188.3200 1345.8200 2188.8000 ;
        RECT 1344.2200 2193.7600 1345.8200 2194.2400 ;
        RECT 1356.5600 2172.0000 1359.5600 2172.4800 ;
        RECT 1356.5600 2177.4400 1359.5600 2177.9200 ;
        RECT 1344.2200 2172.0000 1345.8200 2172.4800 ;
        RECT 1344.2200 2177.4400 1345.8200 2177.9200 ;
        RECT 1356.5600 2155.6800 1359.5600 2156.1600 ;
        RECT 1356.5600 2161.1200 1359.5600 2161.6000 ;
        RECT 1356.5600 2166.5600 1359.5600 2167.0400 ;
        RECT 1344.2200 2155.6800 1345.8200 2156.1600 ;
        RECT 1344.2200 2161.1200 1345.8200 2161.6000 ;
        RECT 1344.2200 2166.5600 1345.8200 2167.0400 ;
        RECT 1356.5600 2150.2400 1359.5600 2150.7200 ;
        RECT 1344.2200 2150.2400 1345.8200 2150.7200 ;
        RECT 1299.2200 2182.8800 1300.8200 2183.3600 ;
        RECT 1299.2200 2188.3200 1300.8200 2188.8000 ;
        RECT 1299.2200 2193.7600 1300.8200 2194.2400 ;
        RECT 1299.2200 2172.0000 1300.8200 2172.4800 ;
        RECT 1299.2200 2177.4400 1300.8200 2177.9200 ;
        RECT 1299.2200 2155.6800 1300.8200 2156.1600 ;
        RECT 1299.2200 2161.1200 1300.8200 2161.6000 ;
        RECT 1299.2200 2166.5600 1300.8200 2167.0400 ;
        RECT 1299.2200 2150.2400 1300.8200 2150.7200 ;
        RECT 1254.2200 2237.2800 1255.8200 2237.7600 ;
        RECT 1254.2200 2242.7200 1255.8200 2243.2000 ;
        RECT 1254.2200 2248.1600 1255.8200 2248.6400 ;
        RECT 1254.2200 2226.4000 1255.8200 2226.8800 ;
        RECT 1254.2200 2231.8400 1255.8200 2232.3200 ;
        RECT 1209.2200 2237.2800 1210.8200 2237.7600 ;
        RECT 1209.2200 2242.7200 1210.8200 2243.2000 ;
        RECT 1209.2200 2248.1600 1210.8200 2248.6400 ;
        RECT 1209.2200 2226.4000 1210.8200 2226.8800 ;
        RECT 1209.2200 2231.8400 1210.8200 2232.3200 ;
        RECT 1254.2200 2210.0800 1255.8200 2210.5600 ;
        RECT 1254.2200 2215.5200 1255.8200 2216.0000 ;
        RECT 1254.2200 2220.9600 1255.8200 2221.4400 ;
        RECT 1254.2200 2199.2000 1255.8200 2199.6800 ;
        RECT 1254.2200 2204.6400 1255.8200 2205.1200 ;
        RECT 1209.2200 2210.0800 1210.8200 2210.5600 ;
        RECT 1209.2200 2215.5200 1210.8200 2216.0000 ;
        RECT 1209.2200 2220.9600 1210.8200 2221.4400 ;
        RECT 1209.2200 2199.2000 1210.8200 2199.6800 ;
        RECT 1209.2200 2204.6400 1210.8200 2205.1200 ;
        RECT 1164.2200 2237.2800 1165.8200 2237.7600 ;
        RECT 1164.2200 2242.7200 1165.8200 2243.2000 ;
        RECT 1164.2200 2248.1600 1165.8200 2248.6400 ;
        RECT 1152.4600 2237.2800 1155.4600 2237.7600 ;
        RECT 1152.4600 2242.7200 1155.4600 2243.2000 ;
        RECT 1152.4600 2248.1600 1155.4600 2248.6400 ;
        RECT 1164.2200 2226.4000 1165.8200 2226.8800 ;
        RECT 1164.2200 2231.8400 1165.8200 2232.3200 ;
        RECT 1152.4600 2226.4000 1155.4600 2226.8800 ;
        RECT 1152.4600 2231.8400 1155.4600 2232.3200 ;
        RECT 1164.2200 2210.0800 1165.8200 2210.5600 ;
        RECT 1164.2200 2215.5200 1165.8200 2216.0000 ;
        RECT 1164.2200 2220.9600 1165.8200 2221.4400 ;
        RECT 1152.4600 2210.0800 1155.4600 2210.5600 ;
        RECT 1152.4600 2215.5200 1155.4600 2216.0000 ;
        RECT 1152.4600 2220.9600 1155.4600 2221.4400 ;
        RECT 1164.2200 2199.2000 1165.8200 2199.6800 ;
        RECT 1164.2200 2204.6400 1165.8200 2205.1200 ;
        RECT 1152.4600 2199.2000 1155.4600 2199.6800 ;
        RECT 1152.4600 2204.6400 1155.4600 2205.1200 ;
        RECT 1254.2200 2182.8800 1255.8200 2183.3600 ;
        RECT 1254.2200 2188.3200 1255.8200 2188.8000 ;
        RECT 1254.2200 2193.7600 1255.8200 2194.2400 ;
        RECT 1254.2200 2172.0000 1255.8200 2172.4800 ;
        RECT 1254.2200 2177.4400 1255.8200 2177.9200 ;
        RECT 1209.2200 2182.8800 1210.8200 2183.3600 ;
        RECT 1209.2200 2188.3200 1210.8200 2188.8000 ;
        RECT 1209.2200 2193.7600 1210.8200 2194.2400 ;
        RECT 1209.2200 2172.0000 1210.8200 2172.4800 ;
        RECT 1209.2200 2177.4400 1210.8200 2177.9200 ;
        RECT 1254.2200 2155.6800 1255.8200 2156.1600 ;
        RECT 1254.2200 2161.1200 1255.8200 2161.6000 ;
        RECT 1254.2200 2166.5600 1255.8200 2167.0400 ;
        RECT 1254.2200 2150.2400 1255.8200 2150.7200 ;
        RECT 1209.2200 2155.6800 1210.8200 2156.1600 ;
        RECT 1209.2200 2161.1200 1210.8200 2161.6000 ;
        RECT 1209.2200 2166.5600 1210.8200 2167.0400 ;
        RECT 1209.2200 2150.2400 1210.8200 2150.7200 ;
        RECT 1164.2200 2182.8800 1165.8200 2183.3600 ;
        RECT 1164.2200 2188.3200 1165.8200 2188.8000 ;
        RECT 1164.2200 2193.7600 1165.8200 2194.2400 ;
        RECT 1152.4600 2182.8800 1155.4600 2183.3600 ;
        RECT 1152.4600 2188.3200 1155.4600 2188.8000 ;
        RECT 1152.4600 2193.7600 1155.4600 2194.2400 ;
        RECT 1164.2200 2172.0000 1165.8200 2172.4800 ;
        RECT 1164.2200 2177.4400 1165.8200 2177.9200 ;
        RECT 1152.4600 2172.0000 1155.4600 2172.4800 ;
        RECT 1152.4600 2177.4400 1155.4600 2177.9200 ;
        RECT 1164.2200 2155.6800 1165.8200 2156.1600 ;
        RECT 1164.2200 2161.1200 1165.8200 2161.6000 ;
        RECT 1164.2200 2166.5600 1165.8200 2167.0400 ;
        RECT 1152.4600 2155.6800 1155.4600 2156.1600 ;
        RECT 1152.4600 2161.1200 1155.4600 2161.6000 ;
        RECT 1152.4600 2166.5600 1155.4600 2167.0400 ;
        RECT 1152.4600 2150.2400 1155.4600 2150.7200 ;
        RECT 1164.2200 2150.2400 1165.8200 2150.7200 ;
        RECT 1152.4600 2355.1500 1359.5600 2358.1500 ;
        RECT 1152.4600 2142.0500 1359.5600 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 1912.4100 1345.8200 2128.5100 ;
        RECT 1299.2200 1912.4100 1300.8200 2128.5100 ;
        RECT 1254.2200 1912.4100 1255.8200 2128.5100 ;
        RECT 1209.2200 1912.4100 1210.8200 2128.5100 ;
        RECT 1164.2200 1912.4100 1165.8200 2128.5100 ;
        RECT 1356.5600 1912.4100 1359.5600 2128.5100 ;
        RECT 1152.4600 1912.4100 1155.4600 2128.5100 ;
      LAYER met3 ;
        RECT 1356.5600 2105.5600 1359.5600 2106.0400 ;
        RECT 1356.5600 2111.0000 1359.5600 2111.4800 ;
        RECT 1344.2200 2105.5600 1345.8200 2106.0400 ;
        RECT 1344.2200 2111.0000 1345.8200 2111.4800 ;
        RECT 1356.5600 2116.4400 1359.5600 2116.9200 ;
        RECT 1344.2200 2116.4400 1345.8200 2116.9200 ;
        RECT 1356.5600 2094.6800 1359.5600 2095.1600 ;
        RECT 1356.5600 2100.1200 1359.5600 2100.6000 ;
        RECT 1344.2200 2094.6800 1345.8200 2095.1600 ;
        RECT 1344.2200 2100.1200 1345.8200 2100.6000 ;
        RECT 1356.5600 2078.3600 1359.5600 2078.8400 ;
        RECT 1356.5600 2083.8000 1359.5600 2084.2800 ;
        RECT 1344.2200 2078.3600 1345.8200 2078.8400 ;
        RECT 1344.2200 2083.8000 1345.8200 2084.2800 ;
        RECT 1356.5600 2089.2400 1359.5600 2089.7200 ;
        RECT 1344.2200 2089.2400 1345.8200 2089.7200 ;
        RECT 1299.2200 2105.5600 1300.8200 2106.0400 ;
        RECT 1299.2200 2111.0000 1300.8200 2111.4800 ;
        RECT 1299.2200 2116.4400 1300.8200 2116.9200 ;
        RECT 1299.2200 2094.6800 1300.8200 2095.1600 ;
        RECT 1299.2200 2100.1200 1300.8200 2100.6000 ;
        RECT 1299.2200 2078.3600 1300.8200 2078.8400 ;
        RECT 1299.2200 2083.8000 1300.8200 2084.2800 ;
        RECT 1299.2200 2089.2400 1300.8200 2089.7200 ;
        RECT 1356.5600 2062.0400 1359.5600 2062.5200 ;
        RECT 1356.5600 2067.4800 1359.5600 2067.9600 ;
        RECT 1356.5600 2072.9200 1359.5600 2073.4000 ;
        RECT 1344.2200 2062.0400 1345.8200 2062.5200 ;
        RECT 1344.2200 2067.4800 1345.8200 2067.9600 ;
        RECT 1344.2200 2072.9200 1345.8200 2073.4000 ;
        RECT 1356.5600 2051.1600 1359.5600 2051.6400 ;
        RECT 1356.5600 2056.6000 1359.5600 2057.0800 ;
        RECT 1344.2200 2051.1600 1345.8200 2051.6400 ;
        RECT 1344.2200 2056.6000 1345.8200 2057.0800 ;
        RECT 1356.5600 2034.8400 1359.5600 2035.3200 ;
        RECT 1356.5600 2040.2800 1359.5600 2040.7600 ;
        RECT 1356.5600 2045.7200 1359.5600 2046.2000 ;
        RECT 1344.2200 2034.8400 1345.8200 2035.3200 ;
        RECT 1344.2200 2040.2800 1345.8200 2040.7600 ;
        RECT 1344.2200 2045.7200 1345.8200 2046.2000 ;
        RECT 1356.5600 2023.9600 1359.5600 2024.4400 ;
        RECT 1356.5600 2029.4000 1359.5600 2029.8800 ;
        RECT 1344.2200 2023.9600 1345.8200 2024.4400 ;
        RECT 1344.2200 2029.4000 1345.8200 2029.8800 ;
        RECT 1299.2200 2062.0400 1300.8200 2062.5200 ;
        RECT 1299.2200 2067.4800 1300.8200 2067.9600 ;
        RECT 1299.2200 2072.9200 1300.8200 2073.4000 ;
        RECT 1299.2200 2051.1600 1300.8200 2051.6400 ;
        RECT 1299.2200 2056.6000 1300.8200 2057.0800 ;
        RECT 1299.2200 2034.8400 1300.8200 2035.3200 ;
        RECT 1299.2200 2040.2800 1300.8200 2040.7600 ;
        RECT 1299.2200 2045.7200 1300.8200 2046.2000 ;
        RECT 1299.2200 2023.9600 1300.8200 2024.4400 ;
        RECT 1299.2200 2029.4000 1300.8200 2029.8800 ;
        RECT 1254.2200 2105.5600 1255.8200 2106.0400 ;
        RECT 1254.2200 2111.0000 1255.8200 2111.4800 ;
        RECT 1254.2200 2116.4400 1255.8200 2116.9200 ;
        RECT 1209.2200 2105.5600 1210.8200 2106.0400 ;
        RECT 1209.2200 2111.0000 1210.8200 2111.4800 ;
        RECT 1209.2200 2116.4400 1210.8200 2116.9200 ;
        RECT 1254.2200 2094.6800 1255.8200 2095.1600 ;
        RECT 1254.2200 2100.1200 1255.8200 2100.6000 ;
        RECT 1254.2200 2078.3600 1255.8200 2078.8400 ;
        RECT 1254.2200 2083.8000 1255.8200 2084.2800 ;
        RECT 1254.2200 2089.2400 1255.8200 2089.7200 ;
        RECT 1209.2200 2094.6800 1210.8200 2095.1600 ;
        RECT 1209.2200 2100.1200 1210.8200 2100.6000 ;
        RECT 1209.2200 2078.3600 1210.8200 2078.8400 ;
        RECT 1209.2200 2083.8000 1210.8200 2084.2800 ;
        RECT 1209.2200 2089.2400 1210.8200 2089.7200 ;
        RECT 1164.2200 2105.5600 1165.8200 2106.0400 ;
        RECT 1164.2200 2111.0000 1165.8200 2111.4800 ;
        RECT 1152.4600 2111.0000 1155.4600 2111.4800 ;
        RECT 1152.4600 2105.5600 1155.4600 2106.0400 ;
        RECT 1152.4600 2116.4400 1155.4600 2116.9200 ;
        RECT 1164.2200 2116.4400 1165.8200 2116.9200 ;
        RECT 1164.2200 2094.6800 1165.8200 2095.1600 ;
        RECT 1164.2200 2100.1200 1165.8200 2100.6000 ;
        RECT 1152.4600 2100.1200 1155.4600 2100.6000 ;
        RECT 1152.4600 2094.6800 1155.4600 2095.1600 ;
        RECT 1164.2200 2078.3600 1165.8200 2078.8400 ;
        RECT 1164.2200 2083.8000 1165.8200 2084.2800 ;
        RECT 1152.4600 2083.8000 1155.4600 2084.2800 ;
        RECT 1152.4600 2078.3600 1155.4600 2078.8400 ;
        RECT 1152.4600 2089.2400 1155.4600 2089.7200 ;
        RECT 1164.2200 2089.2400 1165.8200 2089.7200 ;
        RECT 1254.2200 2062.0400 1255.8200 2062.5200 ;
        RECT 1254.2200 2067.4800 1255.8200 2067.9600 ;
        RECT 1254.2200 2072.9200 1255.8200 2073.4000 ;
        RECT 1254.2200 2051.1600 1255.8200 2051.6400 ;
        RECT 1254.2200 2056.6000 1255.8200 2057.0800 ;
        RECT 1209.2200 2062.0400 1210.8200 2062.5200 ;
        RECT 1209.2200 2067.4800 1210.8200 2067.9600 ;
        RECT 1209.2200 2072.9200 1210.8200 2073.4000 ;
        RECT 1209.2200 2051.1600 1210.8200 2051.6400 ;
        RECT 1209.2200 2056.6000 1210.8200 2057.0800 ;
        RECT 1254.2200 2034.8400 1255.8200 2035.3200 ;
        RECT 1254.2200 2040.2800 1255.8200 2040.7600 ;
        RECT 1254.2200 2045.7200 1255.8200 2046.2000 ;
        RECT 1254.2200 2023.9600 1255.8200 2024.4400 ;
        RECT 1254.2200 2029.4000 1255.8200 2029.8800 ;
        RECT 1209.2200 2034.8400 1210.8200 2035.3200 ;
        RECT 1209.2200 2040.2800 1210.8200 2040.7600 ;
        RECT 1209.2200 2045.7200 1210.8200 2046.2000 ;
        RECT 1209.2200 2023.9600 1210.8200 2024.4400 ;
        RECT 1209.2200 2029.4000 1210.8200 2029.8800 ;
        RECT 1164.2200 2062.0400 1165.8200 2062.5200 ;
        RECT 1164.2200 2067.4800 1165.8200 2067.9600 ;
        RECT 1164.2200 2072.9200 1165.8200 2073.4000 ;
        RECT 1152.4600 2062.0400 1155.4600 2062.5200 ;
        RECT 1152.4600 2067.4800 1155.4600 2067.9600 ;
        RECT 1152.4600 2072.9200 1155.4600 2073.4000 ;
        RECT 1164.2200 2051.1600 1165.8200 2051.6400 ;
        RECT 1164.2200 2056.6000 1165.8200 2057.0800 ;
        RECT 1152.4600 2051.1600 1155.4600 2051.6400 ;
        RECT 1152.4600 2056.6000 1155.4600 2057.0800 ;
        RECT 1164.2200 2034.8400 1165.8200 2035.3200 ;
        RECT 1164.2200 2040.2800 1165.8200 2040.7600 ;
        RECT 1164.2200 2045.7200 1165.8200 2046.2000 ;
        RECT 1152.4600 2034.8400 1155.4600 2035.3200 ;
        RECT 1152.4600 2040.2800 1155.4600 2040.7600 ;
        RECT 1152.4600 2045.7200 1155.4600 2046.2000 ;
        RECT 1164.2200 2023.9600 1165.8200 2024.4400 ;
        RECT 1164.2200 2029.4000 1165.8200 2029.8800 ;
        RECT 1152.4600 2023.9600 1155.4600 2024.4400 ;
        RECT 1152.4600 2029.4000 1155.4600 2029.8800 ;
        RECT 1356.5600 2007.6400 1359.5600 2008.1200 ;
        RECT 1356.5600 2013.0800 1359.5600 2013.5600 ;
        RECT 1356.5600 2018.5200 1359.5600 2019.0000 ;
        RECT 1344.2200 2007.6400 1345.8200 2008.1200 ;
        RECT 1344.2200 2013.0800 1345.8200 2013.5600 ;
        RECT 1344.2200 2018.5200 1345.8200 2019.0000 ;
        RECT 1356.5600 1996.7600 1359.5600 1997.2400 ;
        RECT 1356.5600 2002.2000 1359.5600 2002.6800 ;
        RECT 1344.2200 1996.7600 1345.8200 1997.2400 ;
        RECT 1344.2200 2002.2000 1345.8200 2002.6800 ;
        RECT 1356.5600 1980.4400 1359.5600 1980.9200 ;
        RECT 1356.5600 1985.8800 1359.5600 1986.3600 ;
        RECT 1356.5600 1991.3200 1359.5600 1991.8000 ;
        RECT 1344.2200 1980.4400 1345.8200 1980.9200 ;
        RECT 1344.2200 1985.8800 1345.8200 1986.3600 ;
        RECT 1344.2200 1991.3200 1345.8200 1991.8000 ;
        RECT 1356.5600 1969.5600 1359.5600 1970.0400 ;
        RECT 1356.5600 1975.0000 1359.5600 1975.4800 ;
        RECT 1344.2200 1969.5600 1345.8200 1970.0400 ;
        RECT 1344.2200 1975.0000 1345.8200 1975.4800 ;
        RECT 1299.2200 2007.6400 1300.8200 2008.1200 ;
        RECT 1299.2200 2013.0800 1300.8200 2013.5600 ;
        RECT 1299.2200 2018.5200 1300.8200 2019.0000 ;
        RECT 1299.2200 1996.7600 1300.8200 1997.2400 ;
        RECT 1299.2200 2002.2000 1300.8200 2002.6800 ;
        RECT 1299.2200 1980.4400 1300.8200 1980.9200 ;
        RECT 1299.2200 1985.8800 1300.8200 1986.3600 ;
        RECT 1299.2200 1991.3200 1300.8200 1991.8000 ;
        RECT 1299.2200 1969.5600 1300.8200 1970.0400 ;
        RECT 1299.2200 1975.0000 1300.8200 1975.4800 ;
        RECT 1356.5600 1953.2400 1359.5600 1953.7200 ;
        RECT 1356.5600 1958.6800 1359.5600 1959.1600 ;
        RECT 1356.5600 1964.1200 1359.5600 1964.6000 ;
        RECT 1344.2200 1953.2400 1345.8200 1953.7200 ;
        RECT 1344.2200 1958.6800 1345.8200 1959.1600 ;
        RECT 1344.2200 1964.1200 1345.8200 1964.6000 ;
        RECT 1356.5600 1942.3600 1359.5600 1942.8400 ;
        RECT 1356.5600 1947.8000 1359.5600 1948.2800 ;
        RECT 1344.2200 1942.3600 1345.8200 1942.8400 ;
        RECT 1344.2200 1947.8000 1345.8200 1948.2800 ;
        RECT 1356.5600 1926.0400 1359.5600 1926.5200 ;
        RECT 1356.5600 1931.4800 1359.5600 1931.9600 ;
        RECT 1356.5600 1936.9200 1359.5600 1937.4000 ;
        RECT 1344.2200 1926.0400 1345.8200 1926.5200 ;
        RECT 1344.2200 1931.4800 1345.8200 1931.9600 ;
        RECT 1344.2200 1936.9200 1345.8200 1937.4000 ;
        RECT 1356.5600 1920.6000 1359.5600 1921.0800 ;
        RECT 1344.2200 1920.6000 1345.8200 1921.0800 ;
        RECT 1299.2200 1953.2400 1300.8200 1953.7200 ;
        RECT 1299.2200 1958.6800 1300.8200 1959.1600 ;
        RECT 1299.2200 1964.1200 1300.8200 1964.6000 ;
        RECT 1299.2200 1942.3600 1300.8200 1942.8400 ;
        RECT 1299.2200 1947.8000 1300.8200 1948.2800 ;
        RECT 1299.2200 1926.0400 1300.8200 1926.5200 ;
        RECT 1299.2200 1931.4800 1300.8200 1931.9600 ;
        RECT 1299.2200 1936.9200 1300.8200 1937.4000 ;
        RECT 1299.2200 1920.6000 1300.8200 1921.0800 ;
        RECT 1254.2200 2007.6400 1255.8200 2008.1200 ;
        RECT 1254.2200 2013.0800 1255.8200 2013.5600 ;
        RECT 1254.2200 2018.5200 1255.8200 2019.0000 ;
        RECT 1254.2200 1996.7600 1255.8200 1997.2400 ;
        RECT 1254.2200 2002.2000 1255.8200 2002.6800 ;
        RECT 1209.2200 2007.6400 1210.8200 2008.1200 ;
        RECT 1209.2200 2013.0800 1210.8200 2013.5600 ;
        RECT 1209.2200 2018.5200 1210.8200 2019.0000 ;
        RECT 1209.2200 1996.7600 1210.8200 1997.2400 ;
        RECT 1209.2200 2002.2000 1210.8200 2002.6800 ;
        RECT 1254.2200 1980.4400 1255.8200 1980.9200 ;
        RECT 1254.2200 1985.8800 1255.8200 1986.3600 ;
        RECT 1254.2200 1991.3200 1255.8200 1991.8000 ;
        RECT 1254.2200 1969.5600 1255.8200 1970.0400 ;
        RECT 1254.2200 1975.0000 1255.8200 1975.4800 ;
        RECT 1209.2200 1980.4400 1210.8200 1980.9200 ;
        RECT 1209.2200 1985.8800 1210.8200 1986.3600 ;
        RECT 1209.2200 1991.3200 1210.8200 1991.8000 ;
        RECT 1209.2200 1969.5600 1210.8200 1970.0400 ;
        RECT 1209.2200 1975.0000 1210.8200 1975.4800 ;
        RECT 1164.2200 2007.6400 1165.8200 2008.1200 ;
        RECT 1164.2200 2013.0800 1165.8200 2013.5600 ;
        RECT 1164.2200 2018.5200 1165.8200 2019.0000 ;
        RECT 1152.4600 2007.6400 1155.4600 2008.1200 ;
        RECT 1152.4600 2013.0800 1155.4600 2013.5600 ;
        RECT 1152.4600 2018.5200 1155.4600 2019.0000 ;
        RECT 1164.2200 1996.7600 1165.8200 1997.2400 ;
        RECT 1164.2200 2002.2000 1165.8200 2002.6800 ;
        RECT 1152.4600 1996.7600 1155.4600 1997.2400 ;
        RECT 1152.4600 2002.2000 1155.4600 2002.6800 ;
        RECT 1164.2200 1980.4400 1165.8200 1980.9200 ;
        RECT 1164.2200 1985.8800 1165.8200 1986.3600 ;
        RECT 1164.2200 1991.3200 1165.8200 1991.8000 ;
        RECT 1152.4600 1980.4400 1155.4600 1980.9200 ;
        RECT 1152.4600 1985.8800 1155.4600 1986.3600 ;
        RECT 1152.4600 1991.3200 1155.4600 1991.8000 ;
        RECT 1164.2200 1969.5600 1165.8200 1970.0400 ;
        RECT 1164.2200 1975.0000 1165.8200 1975.4800 ;
        RECT 1152.4600 1969.5600 1155.4600 1970.0400 ;
        RECT 1152.4600 1975.0000 1155.4600 1975.4800 ;
        RECT 1254.2200 1953.2400 1255.8200 1953.7200 ;
        RECT 1254.2200 1958.6800 1255.8200 1959.1600 ;
        RECT 1254.2200 1964.1200 1255.8200 1964.6000 ;
        RECT 1254.2200 1942.3600 1255.8200 1942.8400 ;
        RECT 1254.2200 1947.8000 1255.8200 1948.2800 ;
        RECT 1209.2200 1953.2400 1210.8200 1953.7200 ;
        RECT 1209.2200 1958.6800 1210.8200 1959.1600 ;
        RECT 1209.2200 1964.1200 1210.8200 1964.6000 ;
        RECT 1209.2200 1942.3600 1210.8200 1942.8400 ;
        RECT 1209.2200 1947.8000 1210.8200 1948.2800 ;
        RECT 1254.2200 1926.0400 1255.8200 1926.5200 ;
        RECT 1254.2200 1931.4800 1255.8200 1931.9600 ;
        RECT 1254.2200 1936.9200 1255.8200 1937.4000 ;
        RECT 1254.2200 1920.6000 1255.8200 1921.0800 ;
        RECT 1209.2200 1926.0400 1210.8200 1926.5200 ;
        RECT 1209.2200 1931.4800 1210.8200 1931.9600 ;
        RECT 1209.2200 1936.9200 1210.8200 1937.4000 ;
        RECT 1209.2200 1920.6000 1210.8200 1921.0800 ;
        RECT 1164.2200 1953.2400 1165.8200 1953.7200 ;
        RECT 1164.2200 1958.6800 1165.8200 1959.1600 ;
        RECT 1164.2200 1964.1200 1165.8200 1964.6000 ;
        RECT 1152.4600 1953.2400 1155.4600 1953.7200 ;
        RECT 1152.4600 1958.6800 1155.4600 1959.1600 ;
        RECT 1152.4600 1964.1200 1155.4600 1964.6000 ;
        RECT 1164.2200 1942.3600 1165.8200 1942.8400 ;
        RECT 1164.2200 1947.8000 1165.8200 1948.2800 ;
        RECT 1152.4600 1942.3600 1155.4600 1942.8400 ;
        RECT 1152.4600 1947.8000 1155.4600 1948.2800 ;
        RECT 1164.2200 1926.0400 1165.8200 1926.5200 ;
        RECT 1164.2200 1931.4800 1165.8200 1931.9600 ;
        RECT 1164.2200 1936.9200 1165.8200 1937.4000 ;
        RECT 1152.4600 1926.0400 1155.4600 1926.5200 ;
        RECT 1152.4600 1931.4800 1155.4600 1931.9600 ;
        RECT 1152.4600 1936.9200 1155.4600 1937.4000 ;
        RECT 1152.4600 1920.6000 1155.4600 1921.0800 ;
        RECT 1164.2200 1920.6000 1165.8200 1921.0800 ;
        RECT 1152.4600 2125.5100 1359.5600 2128.5100 ;
        RECT 1152.4600 1912.4100 1359.5600 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 1682.7700 1345.8200 1898.8700 ;
        RECT 1299.2200 1682.7700 1300.8200 1898.8700 ;
        RECT 1254.2200 1682.7700 1255.8200 1898.8700 ;
        RECT 1209.2200 1682.7700 1210.8200 1898.8700 ;
        RECT 1164.2200 1682.7700 1165.8200 1898.8700 ;
        RECT 1356.5600 1682.7700 1359.5600 1898.8700 ;
        RECT 1152.4600 1682.7700 1155.4600 1898.8700 ;
      LAYER met3 ;
        RECT 1356.5600 1875.9200 1359.5600 1876.4000 ;
        RECT 1356.5600 1881.3600 1359.5600 1881.8400 ;
        RECT 1344.2200 1875.9200 1345.8200 1876.4000 ;
        RECT 1344.2200 1881.3600 1345.8200 1881.8400 ;
        RECT 1356.5600 1886.8000 1359.5600 1887.2800 ;
        RECT 1344.2200 1886.8000 1345.8200 1887.2800 ;
        RECT 1356.5600 1865.0400 1359.5600 1865.5200 ;
        RECT 1356.5600 1870.4800 1359.5600 1870.9600 ;
        RECT 1344.2200 1865.0400 1345.8200 1865.5200 ;
        RECT 1344.2200 1870.4800 1345.8200 1870.9600 ;
        RECT 1356.5600 1848.7200 1359.5600 1849.2000 ;
        RECT 1356.5600 1854.1600 1359.5600 1854.6400 ;
        RECT 1344.2200 1848.7200 1345.8200 1849.2000 ;
        RECT 1344.2200 1854.1600 1345.8200 1854.6400 ;
        RECT 1356.5600 1859.6000 1359.5600 1860.0800 ;
        RECT 1344.2200 1859.6000 1345.8200 1860.0800 ;
        RECT 1299.2200 1875.9200 1300.8200 1876.4000 ;
        RECT 1299.2200 1881.3600 1300.8200 1881.8400 ;
        RECT 1299.2200 1886.8000 1300.8200 1887.2800 ;
        RECT 1299.2200 1865.0400 1300.8200 1865.5200 ;
        RECT 1299.2200 1870.4800 1300.8200 1870.9600 ;
        RECT 1299.2200 1848.7200 1300.8200 1849.2000 ;
        RECT 1299.2200 1854.1600 1300.8200 1854.6400 ;
        RECT 1299.2200 1859.6000 1300.8200 1860.0800 ;
        RECT 1356.5600 1832.4000 1359.5600 1832.8800 ;
        RECT 1356.5600 1837.8400 1359.5600 1838.3200 ;
        RECT 1356.5600 1843.2800 1359.5600 1843.7600 ;
        RECT 1344.2200 1832.4000 1345.8200 1832.8800 ;
        RECT 1344.2200 1837.8400 1345.8200 1838.3200 ;
        RECT 1344.2200 1843.2800 1345.8200 1843.7600 ;
        RECT 1356.5600 1821.5200 1359.5600 1822.0000 ;
        RECT 1356.5600 1826.9600 1359.5600 1827.4400 ;
        RECT 1344.2200 1821.5200 1345.8200 1822.0000 ;
        RECT 1344.2200 1826.9600 1345.8200 1827.4400 ;
        RECT 1356.5600 1805.2000 1359.5600 1805.6800 ;
        RECT 1356.5600 1810.6400 1359.5600 1811.1200 ;
        RECT 1356.5600 1816.0800 1359.5600 1816.5600 ;
        RECT 1344.2200 1805.2000 1345.8200 1805.6800 ;
        RECT 1344.2200 1810.6400 1345.8200 1811.1200 ;
        RECT 1344.2200 1816.0800 1345.8200 1816.5600 ;
        RECT 1356.5600 1794.3200 1359.5600 1794.8000 ;
        RECT 1356.5600 1799.7600 1359.5600 1800.2400 ;
        RECT 1344.2200 1794.3200 1345.8200 1794.8000 ;
        RECT 1344.2200 1799.7600 1345.8200 1800.2400 ;
        RECT 1299.2200 1832.4000 1300.8200 1832.8800 ;
        RECT 1299.2200 1837.8400 1300.8200 1838.3200 ;
        RECT 1299.2200 1843.2800 1300.8200 1843.7600 ;
        RECT 1299.2200 1821.5200 1300.8200 1822.0000 ;
        RECT 1299.2200 1826.9600 1300.8200 1827.4400 ;
        RECT 1299.2200 1805.2000 1300.8200 1805.6800 ;
        RECT 1299.2200 1810.6400 1300.8200 1811.1200 ;
        RECT 1299.2200 1816.0800 1300.8200 1816.5600 ;
        RECT 1299.2200 1794.3200 1300.8200 1794.8000 ;
        RECT 1299.2200 1799.7600 1300.8200 1800.2400 ;
        RECT 1254.2200 1875.9200 1255.8200 1876.4000 ;
        RECT 1254.2200 1881.3600 1255.8200 1881.8400 ;
        RECT 1254.2200 1886.8000 1255.8200 1887.2800 ;
        RECT 1209.2200 1875.9200 1210.8200 1876.4000 ;
        RECT 1209.2200 1881.3600 1210.8200 1881.8400 ;
        RECT 1209.2200 1886.8000 1210.8200 1887.2800 ;
        RECT 1254.2200 1865.0400 1255.8200 1865.5200 ;
        RECT 1254.2200 1870.4800 1255.8200 1870.9600 ;
        RECT 1254.2200 1848.7200 1255.8200 1849.2000 ;
        RECT 1254.2200 1854.1600 1255.8200 1854.6400 ;
        RECT 1254.2200 1859.6000 1255.8200 1860.0800 ;
        RECT 1209.2200 1865.0400 1210.8200 1865.5200 ;
        RECT 1209.2200 1870.4800 1210.8200 1870.9600 ;
        RECT 1209.2200 1848.7200 1210.8200 1849.2000 ;
        RECT 1209.2200 1854.1600 1210.8200 1854.6400 ;
        RECT 1209.2200 1859.6000 1210.8200 1860.0800 ;
        RECT 1164.2200 1875.9200 1165.8200 1876.4000 ;
        RECT 1164.2200 1881.3600 1165.8200 1881.8400 ;
        RECT 1152.4600 1881.3600 1155.4600 1881.8400 ;
        RECT 1152.4600 1875.9200 1155.4600 1876.4000 ;
        RECT 1152.4600 1886.8000 1155.4600 1887.2800 ;
        RECT 1164.2200 1886.8000 1165.8200 1887.2800 ;
        RECT 1164.2200 1865.0400 1165.8200 1865.5200 ;
        RECT 1164.2200 1870.4800 1165.8200 1870.9600 ;
        RECT 1152.4600 1870.4800 1155.4600 1870.9600 ;
        RECT 1152.4600 1865.0400 1155.4600 1865.5200 ;
        RECT 1164.2200 1848.7200 1165.8200 1849.2000 ;
        RECT 1164.2200 1854.1600 1165.8200 1854.6400 ;
        RECT 1152.4600 1854.1600 1155.4600 1854.6400 ;
        RECT 1152.4600 1848.7200 1155.4600 1849.2000 ;
        RECT 1152.4600 1859.6000 1155.4600 1860.0800 ;
        RECT 1164.2200 1859.6000 1165.8200 1860.0800 ;
        RECT 1254.2200 1832.4000 1255.8200 1832.8800 ;
        RECT 1254.2200 1837.8400 1255.8200 1838.3200 ;
        RECT 1254.2200 1843.2800 1255.8200 1843.7600 ;
        RECT 1254.2200 1821.5200 1255.8200 1822.0000 ;
        RECT 1254.2200 1826.9600 1255.8200 1827.4400 ;
        RECT 1209.2200 1832.4000 1210.8200 1832.8800 ;
        RECT 1209.2200 1837.8400 1210.8200 1838.3200 ;
        RECT 1209.2200 1843.2800 1210.8200 1843.7600 ;
        RECT 1209.2200 1821.5200 1210.8200 1822.0000 ;
        RECT 1209.2200 1826.9600 1210.8200 1827.4400 ;
        RECT 1254.2200 1805.2000 1255.8200 1805.6800 ;
        RECT 1254.2200 1810.6400 1255.8200 1811.1200 ;
        RECT 1254.2200 1816.0800 1255.8200 1816.5600 ;
        RECT 1254.2200 1794.3200 1255.8200 1794.8000 ;
        RECT 1254.2200 1799.7600 1255.8200 1800.2400 ;
        RECT 1209.2200 1805.2000 1210.8200 1805.6800 ;
        RECT 1209.2200 1810.6400 1210.8200 1811.1200 ;
        RECT 1209.2200 1816.0800 1210.8200 1816.5600 ;
        RECT 1209.2200 1794.3200 1210.8200 1794.8000 ;
        RECT 1209.2200 1799.7600 1210.8200 1800.2400 ;
        RECT 1164.2200 1832.4000 1165.8200 1832.8800 ;
        RECT 1164.2200 1837.8400 1165.8200 1838.3200 ;
        RECT 1164.2200 1843.2800 1165.8200 1843.7600 ;
        RECT 1152.4600 1832.4000 1155.4600 1832.8800 ;
        RECT 1152.4600 1837.8400 1155.4600 1838.3200 ;
        RECT 1152.4600 1843.2800 1155.4600 1843.7600 ;
        RECT 1164.2200 1821.5200 1165.8200 1822.0000 ;
        RECT 1164.2200 1826.9600 1165.8200 1827.4400 ;
        RECT 1152.4600 1821.5200 1155.4600 1822.0000 ;
        RECT 1152.4600 1826.9600 1155.4600 1827.4400 ;
        RECT 1164.2200 1805.2000 1165.8200 1805.6800 ;
        RECT 1164.2200 1810.6400 1165.8200 1811.1200 ;
        RECT 1164.2200 1816.0800 1165.8200 1816.5600 ;
        RECT 1152.4600 1805.2000 1155.4600 1805.6800 ;
        RECT 1152.4600 1810.6400 1155.4600 1811.1200 ;
        RECT 1152.4600 1816.0800 1155.4600 1816.5600 ;
        RECT 1164.2200 1794.3200 1165.8200 1794.8000 ;
        RECT 1164.2200 1799.7600 1165.8200 1800.2400 ;
        RECT 1152.4600 1794.3200 1155.4600 1794.8000 ;
        RECT 1152.4600 1799.7600 1155.4600 1800.2400 ;
        RECT 1356.5600 1778.0000 1359.5600 1778.4800 ;
        RECT 1356.5600 1783.4400 1359.5600 1783.9200 ;
        RECT 1356.5600 1788.8800 1359.5600 1789.3600 ;
        RECT 1344.2200 1778.0000 1345.8200 1778.4800 ;
        RECT 1344.2200 1783.4400 1345.8200 1783.9200 ;
        RECT 1344.2200 1788.8800 1345.8200 1789.3600 ;
        RECT 1356.5600 1767.1200 1359.5600 1767.6000 ;
        RECT 1356.5600 1772.5600 1359.5600 1773.0400 ;
        RECT 1344.2200 1767.1200 1345.8200 1767.6000 ;
        RECT 1344.2200 1772.5600 1345.8200 1773.0400 ;
        RECT 1356.5600 1750.8000 1359.5600 1751.2800 ;
        RECT 1356.5600 1756.2400 1359.5600 1756.7200 ;
        RECT 1356.5600 1761.6800 1359.5600 1762.1600 ;
        RECT 1344.2200 1750.8000 1345.8200 1751.2800 ;
        RECT 1344.2200 1756.2400 1345.8200 1756.7200 ;
        RECT 1344.2200 1761.6800 1345.8200 1762.1600 ;
        RECT 1356.5600 1739.9200 1359.5600 1740.4000 ;
        RECT 1356.5600 1745.3600 1359.5600 1745.8400 ;
        RECT 1344.2200 1739.9200 1345.8200 1740.4000 ;
        RECT 1344.2200 1745.3600 1345.8200 1745.8400 ;
        RECT 1299.2200 1778.0000 1300.8200 1778.4800 ;
        RECT 1299.2200 1783.4400 1300.8200 1783.9200 ;
        RECT 1299.2200 1788.8800 1300.8200 1789.3600 ;
        RECT 1299.2200 1767.1200 1300.8200 1767.6000 ;
        RECT 1299.2200 1772.5600 1300.8200 1773.0400 ;
        RECT 1299.2200 1750.8000 1300.8200 1751.2800 ;
        RECT 1299.2200 1756.2400 1300.8200 1756.7200 ;
        RECT 1299.2200 1761.6800 1300.8200 1762.1600 ;
        RECT 1299.2200 1739.9200 1300.8200 1740.4000 ;
        RECT 1299.2200 1745.3600 1300.8200 1745.8400 ;
        RECT 1356.5600 1723.6000 1359.5600 1724.0800 ;
        RECT 1356.5600 1729.0400 1359.5600 1729.5200 ;
        RECT 1356.5600 1734.4800 1359.5600 1734.9600 ;
        RECT 1344.2200 1723.6000 1345.8200 1724.0800 ;
        RECT 1344.2200 1729.0400 1345.8200 1729.5200 ;
        RECT 1344.2200 1734.4800 1345.8200 1734.9600 ;
        RECT 1356.5600 1712.7200 1359.5600 1713.2000 ;
        RECT 1356.5600 1718.1600 1359.5600 1718.6400 ;
        RECT 1344.2200 1712.7200 1345.8200 1713.2000 ;
        RECT 1344.2200 1718.1600 1345.8200 1718.6400 ;
        RECT 1356.5600 1696.4000 1359.5600 1696.8800 ;
        RECT 1356.5600 1701.8400 1359.5600 1702.3200 ;
        RECT 1356.5600 1707.2800 1359.5600 1707.7600 ;
        RECT 1344.2200 1696.4000 1345.8200 1696.8800 ;
        RECT 1344.2200 1701.8400 1345.8200 1702.3200 ;
        RECT 1344.2200 1707.2800 1345.8200 1707.7600 ;
        RECT 1356.5600 1690.9600 1359.5600 1691.4400 ;
        RECT 1344.2200 1690.9600 1345.8200 1691.4400 ;
        RECT 1299.2200 1723.6000 1300.8200 1724.0800 ;
        RECT 1299.2200 1729.0400 1300.8200 1729.5200 ;
        RECT 1299.2200 1734.4800 1300.8200 1734.9600 ;
        RECT 1299.2200 1712.7200 1300.8200 1713.2000 ;
        RECT 1299.2200 1718.1600 1300.8200 1718.6400 ;
        RECT 1299.2200 1696.4000 1300.8200 1696.8800 ;
        RECT 1299.2200 1701.8400 1300.8200 1702.3200 ;
        RECT 1299.2200 1707.2800 1300.8200 1707.7600 ;
        RECT 1299.2200 1690.9600 1300.8200 1691.4400 ;
        RECT 1254.2200 1778.0000 1255.8200 1778.4800 ;
        RECT 1254.2200 1783.4400 1255.8200 1783.9200 ;
        RECT 1254.2200 1788.8800 1255.8200 1789.3600 ;
        RECT 1254.2200 1767.1200 1255.8200 1767.6000 ;
        RECT 1254.2200 1772.5600 1255.8200 1773.0400 ;
        RECT 1209.2200 1778.0000 1210.8200 1778.4800 ;
        RECT 1209.2200 1783.4400 1210.8200 1783.9200 ;
        RECT 1209.2200 1788.8800 1210.8200 1789.3600 ;
        RECT 1209.2200 1767.1200 1210.8200 1767.6000 ;
        RECT 1209.2200 1772.5600 1210.8200 1773.0400 ;
        RECT 1254.2200 1750.8000 1255.8200 1751.2800 ;
        RECT 1254.2200 1756.2400 1255.8200 1756.7200 ;
        RECT 1254.2200 1761.6800 1255.8200 1762.1600 ;
        RECT 1254.2200 1739.9200 1255.8200 1740.4000 ;
        RECT 1254.2200 1745.3600 1255.8200 1745.8400 ;
        RECT 1209.2200 1750.8000 1210.8200 1751.2800 ;
        RECT 1209.2200 1756.2400 1210.8200 1756.7200 ;
        RECT 1209.2200 1761.6800 1210.8200 1762.1600 ;
        RECT 1209.2200 1739.9200 1210.8200 1740.4000 ;
        RECT 1209.2200 1745.3600 1210.8200 1745.8400 ;
        RECT 1164.2200 1778.0000 1165.8200 1778.4800 ;
        RECT 1164.2200 1783.4400 1165.8200 1783.9200 ;
        RECT 1164.2200 1788.8800 1165.8200 1789.3600 ;
        RECT 1152.4600 1778.0000 1155.4600 1778.4800 ;
        RECT 1152.4600 1783.4400 1155.4600 1783.9200 ;
        RECT 1152.4600 1788.8800 1155.4600 1789.3600 ;
        RECT 1164.2200 1767.1200 1165.8200 1767.6000 ;
        RECT 1164.2200 1772.5600 1165.8200 1773.0400 ;
        RECT 1152.4600 1767.1200 1155.4600 1767.6000 ;
        RECT 1152.4600 1772.5600 1155.4600 1773.0400 ;
        RECT 1164.2200 1750.8000 1165.8200 1751.2800 ;
        RECT 1164.2200 1756.2400 1165.8200 1756.7200 ;
        RECT 1164.2200 1761.6800 1165.8200 1762.1600 ;
        RECT 1152.4600 1750.8000 1155.4600 1751.2800 ;
        RECT 1152.4600 1756.2400 1155.4600 1756.7200 ;
        RECT 1152.4600 1761.6800 1155.4600 1762.1600 ;
        RECT 1164.2200 1739.9200 1165.8200 1740.4000 ;
        RECT 1164.2200 1745.3600 1165.8200 1745.8400 ;
        RECT 1152.4600 1739.9200 1155.4600 1740.4000 ;
        RECT 1152.4600 1745.3600 1155.4600 1745.8400 ;
        RECT 1254.2200 1723.6000 1255.8200 1724.0800 ;
        RECT 1254.2200 1729.0400 1255.8200 1729.5200 ;
        RECT 1254.2200 1734.4800 1255.8200 1734.9600 ;
        RECT 1254.2200 1712.7200 1255.8200 1713.2000 ;
        RECT 1254.2200 1718.1600 1255.8200 1718.6400 ;
        RECT 1209.2200 1723.6000 1210.8200 1724.0800 ;
        RECT 1209.2200 1729.0400 1210.8200 1729.5200 ;
        RECT 1209.2200 1734.4800 1210.8200 1734.9600 ;
        RECT 1209.2200 1712.7200 1210.8200 1713.2000 ;
        RECT 1209.2200 1718.1600 1210.8200 1718.6400 ;
        RECT 1254.2200 1696.4000 1255.8200 1696.8800 ;
        RECT 1254.2200 1701.8400 1255.8200 1702.3200 ;
        RECT 1254.2200 1707.2800 1255.8200 1707.7600 ;
        RECT 1254.2200 1690.9600 1255.8200 1691.4400 ;
        RECT 1209.2200 1696.4000 1210.8200 1696.8800 ;
        RECT 1209.2200 1701.8400 1210.8200 1702.3200 ;
        RECT 1209.2200 1707.2800 1210.8200 1707.7600 ;
        RECT 1209.2200 1690.9600 1210.8200 1691.4400 ;
        RECT 1164.2200 1723.6000 1165.8200 1724.0800 ;
        RECT 1164.2200 1729.0400 1165.8200 1729.5200 ;
        RECT 1164.2200 1734.4800 1165.8200 1734.9600 ;
        RECT 1152.4600 1723.6000 1155.4600 1724.0800 ;
        RECT 1152.4600 1729.0400 1155.4600 1729.5200 ;
        RECT 1152.4600 1734.4800 1155.4600 1734.9600 ;
        RECT 1164.2200 1712.7200 1165.8200 1713.2000 ;
        RECT 1164.2200 1718.1600 1165.8200 1718.6400 ;
        RECT 1152.4600 1712.7200 1155.4600 1713.2000 ;
        RECT 1152.4600 1718.1600 1155.4600 1718.6400 ;
        RECT 1164.2200 1696.4000 1165.8200 1696.8800 ;
        RECT 1164.2200 1701.8400 1165.8200 1702.3200 ;
        RECT 1164.2200 1707.2800 1165.8200 1707.7600 ;
        RECT 1152.4600 1696.4000 1155.4600 1696.8800 ;
        RECT 1152.4600 1701.8400 1155.4600 1702.3200 ;
        RECT 1152.4600 1707.2800 1155.4600 1707.7600 ;
        RECT 1152.4600 1690.9600 1155.4600 1691.4400 ;
        RECT 1164.2200 1690.9600 1165.8200 1691.4400 ;
        RECT 1152.4600 1895.8700 1359.5600 1898.8700 ;
        RECT 1152.4600 1682.7700 1359.5600 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 1453.1300 1345.8200 1669.2300 ;
        RECT 1299.2200 1453.1300 1300.8200 1669.2300 ;
        RECT 1254.2200 1453.1300 1255.8200 1669.2300 ;
        RECT 1209.2200 1453.1300 1210.8200 1669.2300 ;
        RECT 1164.2200 1453.1300 1165.8200 1669.2300 ;
        RECT 1356.5600 1453.1300 1359.5600 1669.2300 ;
        RECT 1152.4600 1453.1300 1155.4600 1669.2300 ;
      LAYER met3 ;
        RECT 1356.5600 1646.2800 1359.5600 1646.7600 ;
        RECT 1356.5600 1651.7200 1359.5600 1652.2000 ;
        RECT 1344.2200 1646.2800 1345.8200 1646.7600 ;
        RECT 1344.2200 1651.7200 1345.8200 1652.2000 ;
        RECT 1356.5600 1657.1600 1359.5600 1657.6400 ;
        RECT 1344.2200 1657.1600 1345.8200 1657.6400 ;
        RECT 1356.5600 1635.4000 1359.5600 1635.8800 ;
        RECT 1356.5600 1640.8400 1359.5600 1641.3200 ;
        RECT 1344.2200 1635.4000 1345.8200 1635.8800 ;
        RECT 1344.2200 1640.8400 1345.8200 1641.3200 ;
        RECT 1356.5600 1619.0800 1359.5600 1619.5600 ;
        RECT 1356.5600 1624.5200 1359.5600 1625.0000 ;
        RECT 1344.2200 1619.0800 1345.8200 1619.5600 ;
        RECT 1344.2200 1624.5200 1345.8200 1625.0000 ;
        RECT 1356.5600 1629.9600 1359.5600 1630.4400 ;
        RECT 1344.2200 1629.9600 1345.8200 1630.4400 ;
        RECT 1299.2200 1646.2800 1300.8200 1646.7600 ;
        RECT 1299.2200 1651.7200 1300.8200 1652.2000 ;
        RECT 1299.2200 1657.1600 1300.8200 1657.6400 ;
        RECT 1299.2200 1635.4000 1300.8200 1635.8800 ;
        RECT 1299.2200 1640.8400 1300.8200 1641.3200 ;
        RECT 1299.2200 1619.0800 1300.8200 1619.5600 ;
        RECT 1299.2200 1624.5200 1300.8200 1625.0000 ;
        RECT 1299.2200 1629.9600 1300.8200 1630.4400 ;
        RECT 1356.5600 1602.7600 1359.5600 1603.2400 ;
        RECT 1356.5600 1608.2000 1359.5600 1608.6800 ;
        RECT 1356.5600 1613.6400 1359.5600 1614.1200 ;
        RECT 1344.2200 1602.7600 1345.8200 1603.2400 ;
        RECT 1344.2200 1608.2000 1345.8200 1608.6800 ;
        RECT 1344.2200 1613.6400 1345.8200 1614.1200 ;
        RECT 1356.5600 1591.8800 1359.5600 1592.3600 ;
        RECT 1356.5600 1597.3200 1359.5600 1597.8000 ;
        RECT 1344.2200 1591.8800 1345.8200 1592.3600 ;
        RECT 1344.2200 1597.3200 1345.8200 1597.8000 ;
        RECT 1356.5600 1575.5600 1359.5600 1576.0400 ;
        RECT 1356.5600 1581.0000 1359.5600 1581.4800 ;
        RECT 1356.5600 1586.4400 1359.5600 1586.9200 ;
        RECT 1344.2200 1575.5600 1345.8200 1576.0400 ;
        RECT 1344.2200 1581.0000 1345.8200 1581.4800 ;
        RECT 1344.2200 1586.4400 1345.8200 1586.9200 ;
        RECT 1356.5600 1564.6800 1359.5600 1565.1600 ;
        RECT 1356.5600 1570.1200 1359.5600 1570.6000 ;
        RECT 1344.2200 1564.6800 1345.8200 1565.1600 ;
        RECT 1344.2200 1570.1200 1345.8200 1570.6000 ;
        RECT 1299.2200 1602.7600 1300.8200 1603.2400 ;
        RECT 1299.2200 1608.2000 1300.8200 1608.6800 ;
        RECT 1299.2200 1613.6400 1300.8200 1614.1200 ;
        RECT 1299.2200 1591.8800 1300.8200 1592.3600 ;
        RECT 1299.2200 1597.3200 1300.8200 1597.8000 ;
        RECT 1299.2200 1575.5600 1300.8200 1576.0400 ;
        RECT 1299.2200 1581.0000 1300.8200 1581.4800 ;
        RECT 1299.2200 1586.4400 1300.8200 1586.9200 ;
        RECT 1299.2200 1564.6800 1300.8200 1565.1600 ;
        RECT 1299.2200 1570.1200 1300.8200 1570.6000 ;
        RECT 1254.2200 1646.2800 1255.8200 1646.7600 ;
        RECT 1254.2200 1651.7200 1255.8200 1652.2000 ;
        RECT 1254.2200 1657.1600 1255.8200 1657.6400 ;
        RECT 1209.2200 1646.2800 1210.8200 1646.7600 ;
        RECT 1209.2200 1651.7200 1210.8200 1652.2000 ;
        RECT 1209.2200 1657.1600 1210.8200 1657.6400 ;
        RECT 1254.2200 1635.4000 1255.8200 1635.8800 ;
        RECT 1254.2200 1640.8400 1255.8200 1641.3200 ;
        RECT 1254.2200 1619.0800 1255.8200 1619.5600 ;
        RECT 1254.2200 1624.5200 1255.8200 1625.0000 ;
        RECT 1254.2200 1629.9600 1255.8200 1630.4400 ;
        RECT 1209.2200 1635.4000 1210.8200 1635.8800 ;
        RECT 1209.2200 1640.8400 1210.8200 1641.3200 ;
        RECT 1209.2200 1619.0800 1210.8200 1619.5600 ;
        RECT 1209.2200 1624.5200 1210.8200 1625.0000 ;
        RECT 1209.2200 1629.9600 1210.8200 1630.4400 ;
        RECT 1164.2200 1646.2800 1165.8200 1646.7600 ;
        RECT 1164.2200 1651.7200 1165.8200 1652.2000 ;
        RECT 1152.4600 1651.7200 1155.4600 1652.2000 ;
        RECT 1152.4600 1646.2800 1155.4600 1646.7600 ;
        RECT 1152.4600 1657.1600 1155.4600 1657.6400 ;
        RECT 1164.2200 1657.1600 1165.8200 1657.6400 ;
        RECT 1164.2200 1635.4000 1165.8200 1635.8800 ;
        RECT 1164.2200 1640.8400 1165.8200 1641.3200 ;
        RECT 1152.4600 1640.8400 1155.4600 1641.3200 ;
        RECT 1152.4600 1635.4000 1155.4600 1635.8800 ;
        RECT 1164.2200 1619.0800 1165.8200 1619.5600 ;
        RECT 1164.2200 1624.5200 1165.8200 1625.0000 ;
        RECT 1152.4600 1624.5200 1155.4600 1625.0000 ;
        RECT 1152.4600 1619.0800 1155.4600 1619.5600 ;
        RECT 1152.4600 1629.9600 1155.4600 1630.4400 ;
        RECT 1164.2200 1629.9600 1165.8200 1630.4400 ;
        RECT 1254.2200 1602.7600 1255.8200 1603.2400 ;
        RECT 1254.2200 1608.2000 1255.8200 1608.6800 ;
        RECT 1254.2200 1613.6400 1255.8200 1614.1200 ;
        RECT 1254.2200 1591.8800 1255.8200 1592.3600 ;
        RECT 1254.2200 1597.3200 1255.8200 1597.8000 ;
        RECT 1209.2200 1602.7600 1210.8200 1603.2400 ;
        RECT 1209.2200 1608.2000 1210.8200 1608.6800 ;
        RECT 1209.2200 1613.6400 1210.8200 1614.1200 ;
        RECT 1209.2200 1591.8800 1210.8200 1592.3600 ;
        RECT 1209.2200 1597.3200 1210.8200 1597.8000 ;
        RECT 1254.2200 1575.5600 1255.8200 1576.0400 ;
        RECT 1254.2200 1581.0000 1255.8200 1581.4800 ;
        RECT 1254.2200 1586.4400 1255.8200 1586.9200 ;
        RECT 1254.2200 1564.6800 1255.8200 1565.1600 ;
        RECT 1254.2200 1570.1200 1255.8200 1570.6000 ;
        RECT 1209.2200 1575.5600 1210.8200 1576.0400 ;
        RECT 1209.2200 1581.0000 1210.8200 1581.4800 ;
        RECT 1209.2200 1586.4400 1210.8200 1586.9200 ;
        RECT 1209.2200 1564.6800 1210.8200 1565.1600 ;
        RECT 1209.2200 1570.1200 1210.8200 1570.6000 ;
        RECT 1164.2200 1602.7600 1165.8200 1603.2400 ;
        RECT 1164.2200 1608.2000 1165.8200 1608.6800 ;
        RECT 1164.2200 1613.6400 1165.8200 1614.1200 ;
        RECT 1152.4600 1602.7600 1155.4600 1603.2400 ;
        RECT 1152.4600 1608.2000 1155.4600 1608.6800 ;
        RECT 1152.4600 1613.6400 1155.4600 1614.1200 ;
        RECT 1164.2200 1591.8800 1165.8200 1592.3600 ;
        RECT 1164.2200 1597.3200 1165.8200 1597.8000 ;
        RECT 1152.4600 1591.8800 1155.4600 1592.3600 ;
        RECT 1152.4600 1597.3200 1155.4600 1597.8000 ;
        RECT 1164.2200 1575.5600 1165.8200 1576.0400 ;
        RECT 1164.2200 1581.0000 1165.8200 1581.4800 ;
        RECT 1164.2200 1586.4400 1165.8200 1586.9200 ;
        RECT 1152.4600 1575.5600 1155.4600 1576.0400 ;
        RECT 1152.4600 1581.0000 1155.4600 1581.4800 ;
        RECT 1152.4600 1586.4400 1155.4600 1586.9200 ;
        RECT 1164.2200 1564.6800 1165.8200 1565.1600 ;
        RECT 1164.2200 1570.1200 1165.8200 1570.6000 ;
        RECT 1152.4600 1564.6800 1155.4600 1565.1600 ;
        RECT 1152.4600 1570.1200 1155.4600 1570.6000 ;
        RECT 1356.5600 1548.3600 1359.5600 1548.8400 ;
        RECT 1356.5600 1553.8000 1359.5600 1554.2800 ;
        RECT 1356.5600 1559.2400 1359.5600 1559.7200 ;
        RECT 1344.2200 1548.3600 1345.8200 1548.8400 ;
        RECT 1344.2200 1553.8000 1345.8200 1554.2800 ;
        RECT 1344.2200 1559.2400 1345.8200 1559.7200 ;
        RECT 1356.5600 1537.4800 1359.5600 1537.9600 ;
        RECT 1356.5600 1542.9200 1359.5600 1543.4000 ;
        RECT 1344.2200 1537.4800 1345.8200 1537.9600 ;
        RECT 1344.2200 1542.9200 1345.8200 1543.4000 ;
        RECT 1356.5600 1521.1600 1359.5600 1521.6400 ;
        RECT 1356.5600 1526.6000 1359.5600 1527.0800 ;
        RECT 1356.5600 1532.0400 1359.5600 1532.5200 ;
        RECT 1344.2200 1521.1600 1345.8200 1521.6400 ;
        RECT 1344.2200 1526.6000 1345.8200 1527.0800 ;
        RECT 1344.2200 1532.0400 1345.8200 1532.5200 ;
        RECT 1356.5600 1510.2800 1359.5600 1510.7600 ;
        RECT 1356.5600 1515.7200 1359.5600 1516.2000 ;
        RECT 1344.2200 1510.2800 1345.8200 1510.7600 ;
        RECT 1344.2200 1515.7200 1345.8200 1516.2000 ;
        RECT 1299.2200 1548.3600 1300.8200 1548.8400 ;
        RECT 1299.2200 1553.8000 1300.8200 1554.2800 ;
        RECT 1299.2200 1559.2400 1300.8200 1559.7200 ;
        RECT 1299.2200 1537.4800 1300.8200 1537.9600 ;
        RECT 1299.2200 1542.9200 1300.8200 1543.4000 ;
        RECT 1299.2200 1521.1600 1300.8200 1521.6400 ;
        RECT 1299.2200 1526.6000 1300.8200 1527.0800 ;
        RECT 1299.2200 1532.0400 1300.8200 1532.5200 ;
        RECT 1299.2200 1510.2800 1300.8200 1510.7600 ;
        RECT 1299.2200 1515.7200 1300.8200 1516.2000 ;
        RECT 1356.5600 1493.9600 1359.5600 1494.4400 ;
        RECT 1356.5600 1499.4000 1359.5600 1499.8800 ;
        RECT 1356.5600 1504.8400 1359.5600 1505.3200 ;
        RECT 1344.2200 1493.9600 1345.8200 1494.4400 ;
        RECT 1344.2200 1499.4000 1345.8200 1499.8800 ;
        RECT 1344.2200 1504.8400 1345.8200 1505.3200 ;
        RECT 1356.5600 1483.0800 1359.5600 1483.5600 ;
        RECT 1356.5600 1488.5200 1359.5600 1489.0000 ;
        RECT 1344.2200 1483.0800 1345.8200 1483.5600 ;
        RECT 1344.2200 1488.5200 1345.8200 1489.0000 ;
        RECT 1356.5600 1466.7600 1359.5600 1467.2400 ;
        RECT 1356.5600 1472.2000 1359.5600 1472.6800 ;
        RECT 1356.5600 1477.6400 1359.5600 1478.1200 ;
        RECT 1344.2200 1466.7600 1345.8200 1467.2400 ;
        RECT 1344.2200 1472.2000 1345.8200 1472.6800 ;
        RECT 1344.2200 1477.6400 1345.8200 1478.1200 ;
        RECT 1356.5600 1461.3200 1359.5600 1461.8000 ;
        RECT 1344.2200 1461.3200 1345.8200 1461.8000 ;
        RECT 1299.2200 1493.9600 1300.8200 1494.4400 ;
        RECT 1299.2200 1499.4000 1300.8200 1499.8800 ;
        RECT 1299.2200 1504.8400 1300.8200 1505.3200 ;
        RECT 1299.2200 1483.0800 1300.8200 1483.5600 ;
        RECT 1299.2200 1488.5200 1300.8200 1489.0000 ;
        RECT 1299.2200 1466.7600 1300.8200 1467.2400 ;
        RECT 1299.2200 1472.2000 1300.8200 1472.6800 ;
        RECT 1299.2200 1477.6400 1300.8200 1478.1200 ;
        RECT 1299.2200 1461.3200 1300.8200 1461.8000 ;
        RECT 1254.2200 1548.3600 1255.8200 1548.8400 ;
        RECT 1254.2200 1553.8000 1255.8200 1554.2800 ;
        RECT 1254.2200 1559.2400 1255.8200 1559.7200 ;
        RECT 1254.2200 1537.4800 1255.8200 1537.9600 ;
        RECT 1254.2200 1542.9200 1255.8200 1543.4000 ;
        RECT 1209.2200 1548.3600 1210.8200 1548.8400 ;
        RECT 1209.2200 1553.8000 1210.8200 1554.2800 ;
        RECT 1209.2200 1559.2400 1210.8200 1559.7200 ;
        RECT 1209.2200 1537.4800 1210.8200 1537.9600 ;
        RECT 1209.2200 1542.9200 1210.8200 1543.4000 ;
        RECT 1254.2200 1521.1600 1255.8200 1521.6400 ;
        RECT 1254.2200 1526.6000 1255.8200 1527.0800 ;
        RECT 1254.2200 1532.0400 1255.8200 1532.5200 ;
        RECT 1254.2200 1510.2800 1255.8200 1510.7600 ;
        RECT 1254.2200 1515.7200 1255.8200 1516.2000 ;
        RECT 1209.2200 1521.1600 1210.8200 1521.6400 ;
        RECT 1209.2200 1526.6000 1210.8200 1527.0800 ;
        RECT 1209.2200 1532.0400 1210.8200 1532.5200 ;
        RECT 1209.2200 1510.2800 1210.8200 1510.7600 ;
        RECT 1209.2200 1515.7200 1210.8200 1516.2000 ;
        RECT 1164.2200 1548.3600 1165.8200 1548.8400 ;
        RECT 1164.2200 1553.8000 1165.8200 1554.2800 ;
        RECT 1164.2200 1559.2400 1165.8200 1559.7200 ;
        RECT 1152.4600 1548.3600 1155.4600 1548.8400 ;
        RECT 1152.4600 1553.8000 1155.4600 1554.2800 ;
        RECT 1152.4600 1559.2400 1155.4600 1559.7200 ;
        RECT 1164.2200 1537.4800 1165.8200 1537.9600 ;
        RECT 1164.2200 1542.9200 1165.8200 1543.4000 ;
        RECT 1152.4600 1537.4800 1155.4600 1537.9600 ;
        RECT 1152.4600 1542.9200 1155.4600 1543.4000 ;
        RECT 1164.2200 1521.1600 1165.8200 1521.6400 ;
        RECT 1164.2200 1526.6000 1165.8200 1527.0800 ;
        RECT 1164.2200 1532.0400 1165.8200 1532.5200 ;
        RECT 1152.4600 1521.1600 1155.4600 1521.6400 ;
        RECT 1152.4600 1526.6000 1155.4600 1527.0800 ;
        RECT 1152.4600 1532.0400 1155.4600 1532.5200 ;
        RECT 1164.2200 1510.2800 1165.8200 1510.7600 ;
        RECT 1164.2200 1515.7200 1165.8200 1516.2000 ;
        RECT 1152.4600 1510.2800 1155.4600 1510.7600 ;
        RECT 1152.4600 1515.7200 1155.4600 1516.2000 ;
        RECT 1254.2200 1493.9600 1255.8200 1494.4400 ;
        RECT 1254.2200 1499.4000 1255.8200 1499.8800 ;
        RECT 1254.2200 1504.8400 1255.8200 1505.3200 ;
        RECT 1254.2200 1483.0800 1255.8200 1483.5600 ;
        RECT 1254.2200 1488.5200 1255.8200 1489.0000 ;
        RECT 1209.2200 1493.9600 1210.8200 1494.4400 ;
        RECT 1209.2200 1499.4000 1210.8200 1499.8800 ;
        RECT 1209.2200 1504.8400 1210.8200 1505.3200 ;
        RECT 1209.2200 1483.0800 1210.8200 1483.5600 ;
        RECT 1209.2200 1488.5200 1210.8200 1489.0000 ;
        RECT 1254.2200 1466.7600 1255.8200 1467.2400 ;
        RECT 1254.2200 1472.2000 1255.8200 1472.6800 ;
        RECT 1254.2200 1477.6400 1255.8200 1478.1200 ;
        RECT 1254.2200 1461.3200 1255.8200 1461.8000 ;
        RECT 1209.2200 1466.7600 1210.8200 1467.2400 ;
        RECT 1209.2200 1472.2000 1210.8200 1472.6800 ;
        RECT 1209.2200 1477.6400 1210.8200 1478.1200 ;
        RECT 1209.2200 1461.3200 1210.8200 1461.8000 ;
        RECT 1164.2200 1493.9600 1165.8200 1494.4400 ;
        RECT 1164.2200 1499.4000 1165.8200 1499.8800 ;
        RECT 1164.2200 1504.8400 1165.8200 1505.3200 ;
        RECT 1152.4600 1493.9600 1155.4600 1494.4400 ;
        RECT 1152.4600 1499.4000 1155.4600 1499.8800 ;
        RECT 1152.4600 1504.8400 1155.4600 1505.3200 ;
        RECT 1164.2200 1483.0800 1165.8200 1483.5600 ;
        RECT 1164.2200 1488.5200 1165.8200 1489.0000 ;
        RECT 1152.4600 1483.0800 1155.4600 1483.5600 ;
        RECT 1152.4600 1488.5200 1155.4600 1489.0000 ;
        RECT 1164.2200 1466.7600 1165.8200 1467.2400 ;
        RECT 1164.2200 1472.2000 1165.8200 1472.6800 ;
        RECT 1164.2200 1477.6400 1165.8200 1478.1200 ;
        RECT 1152.4600 1466.7600 1155.4600 1467.2400 ;
        RECT 1152.4600 1472.2000 1155.4600 1472.6800 ;
        RECT 1152.4600 1477.6400 1155.4600 1478.1200 ;
        RECT 1152.4600 1461.3200 1155.4600 1461.8000 ;
        RECT 1164.2200 1461.3200 1165.8200 1461.8000 ;
        RECT 1152.4600 1666.2300 1359.5600 1669.2300 ;
        RECT 1152.4600 1453.1300 1359.5600 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 1223.4900 1345.8200 1439.5900 ;
        RECT 1299.2200 1223.4900 1300.8200 1439.5900 ;
        RECT 1254.2200 1223.4900 1255.8200 1439.5900 ;
        RECT 1209.2200 1223.4900 1210.8200 1439.5900 ;
        RECT 1164.2200 1223.4900 1165.8200 1439.5900 ;
        RECT 1356.5600 1223.4900 1359.5600 1439.5900 ;
        RECT 1152.4600 1223.4900 1155.4600 1439.5900 ;
      LAYER met3 ;
        RECT 1356.5600 1416.6400 1359.5600 1417.1200 ;
        RECT 1356.5600 1422.0800 1359.5600 1422.5600 ;
        RECT 1344.2200 1416.6400 1345.8200 1417.1200 ;
        RECT 1344.2200 1422.0800 1345.8200 1422.5600 ;
        RECT 1356.5600 1427.5200 1359.5600 1428.0000 ;
        RECT 1344.2200 1427.5200 1345.8200 1428.0000 ;
        RECT 1356.5600 1405.7600 1359.5600 1406.2400 ;
        RECT 1356.5600 1411.2000 1359.5600 1411.6800 ;
        RECT 1344.2200 1405.7600 1345.8200 1406.2400 ;
        RECT 1344.2200 1411.2000 1345.8200 1411.6800 ;
        RECT 1356.5600 1389.4400 1359.5600 1389.9200 ;
        RECT 1356.5600 1394.8800 1359.5600 1395.3600 ;
        RECT 1344.2200 1389.4400 1345.8200 1389.9200 ;
        RECT 1344.2200 1394.8800 1345.8200 1395.3600 ;
        RECT 1356.5600 1400.3200 1359.5600 1400.8000 ;
        RECT 1344.2200 1400.3200 1345.8200 1400.8000 ;
        RECT 1299.2200 1416.6400 1300.8200 1417.1200 ;
        RECT 1299.2200 1422.0800 1300.8200 1422.5600 ;
        RECT 1299.2200 1427.5200 1300.8200 1428.0000 ;
        RECT 1299.2200 1405.7600 1300.8200 1406.2400 ;
        RECT 1299.2200 1411.2000 1300.8200 1411.6800 ;
        RECT 1299.2200 1389.4400 1300.8200 1389.9200 ;
        RECT 1299.2200 1394.8800 1300.8200 1395.3600 ;
        RECT 1299.2200 1400.3200 1300.8200 1400.8000 ;
        RECT 1356.5600 1373.1200 1359.5600 1373.6000 ;
        RECT 1356.5600 1378.5600 1359.5600 1379.0400 ;
        RECT 1356.5600 1384.0000 1359.5600 1384.4800 ;
        RECT 1344.2200 1373.1200 1345.8200 1373.6000 ;
        RECT 1344.2200 1378.5600 1345.8200 1379.0400 ;
        RECT 1344.2200 1384.0000 1345.8200 1384.4800 ;
        RECT 1356.5600 1362.2400 1359.5600 1362.7200 ;
        RECT 1356.5600 1367.6800 1359.5600 1368.1600 ;
        RECT 1344.2200 1362.2400 1345.8200 1362.7200 ;
        RECT 1344.2200 1367.6800 1345.8200 1368.1600 ;
        RECT 1356.5600 1345.9200 1359.5600 1346.4000 ;
        RECT 1356.5600 1351.3600 1359.5600 1351.8400 ;
        RECT 1356.5600 1356.8000 1359.5600 1357.2800 ;
        RECT 1344.2200 1345.9200 1345.8200 1346.4000 ;
        RECT 1344.2200 1351.3600 1345.8200 1351.8400 ;
        RECT 1344.2200 1356.8000 1345.8200 1357.2800 ;
        RECT 1356.5600 1335.0400 1359.5600 1335.5200 ;
        RECT 1356.5600 1340.4800 1359.5600 1340.9600 ;
        RECT 1344.2200 1335.0400 1345.8200 1335.5200 ;
        RECT 1344.2200 1340.4800 1345.8200 1340.9600 ;
        RECT 1299.2200 1373.1200 1300.8200 1373.6000 ;
        RECT 1299.2200 1378.5600 1300.8200 1379.0400 ;
        RECT 1299.2200 1384.0000 1300.8200 1384.4800 ;
        RECT 1299.2200 1362.2400 1300.8200 1362.7200 ;
        RECT 1299.2200 1367.6800 1300.8200 1368.1600 ;
        RECT 1299.2200 1345.9200 1300.8200 1346.4000 ;
        RECT 1299.2200 1351.3600 1300.8200 1351.8400 ;
        RECT 1299.2200 1356.8000 1300.8200 1357.2800 ;
        RECT 1299.2200 1335.0400 1300.8200 1335.5200 ;
        RECT 1299.2200 1340.4800 1300.8200 1340.9600 ;
        RECT 1254.2200 1416.6400 1255.8200 1417.1200 ;
        RECT 1254.2200 1422.0800 1255.8200 1422.5600 ;
        RECT 1254.2200 1427.5200 1255.8200 1428.0000 ;
        RECT 1209.2200 1416.6400 1210.8200 1417.1200 ;
        RECT 1209.2200 1422.0800 1210.8200 1422.5600 ;
        RECT 1209.2200 1427.5200 1210.8200 1428.0000 ;
        RECT 1254.2200 1405.7600 1255.8200 1406.2400 ;
        RECT 1254.2200 1411.2000 1255.8200 1411.6800 ;
        RECT 1254.2200 1389.4400 1255.8200 1389.9200 ;
        RECT 1254.2200 1394.8800 1255.8200 1395.3600 ;
        RECT 1254.2200 1400.3200 1255.8200 1400.8000 ;
        RECT 1209.2200 1405.7600 1210.8200 1406.2400 ;
        RECT 1209.2200 1411.2000 1210.8200 1411.6800 ;
        RECT 1209.2200 1389.4400 1210.8200 1389.9200 ;
        RECT 1209.2200 1394.8800 1210.8200 1395.3600 ;
        RECT 1209.2200 1400.3200 1210.8200 1400.8000 ;
        RECT 1164.2200 1416.6400 1165.8200 1417.1200 ;
        RECT 1164.2200 1422.0800 1165.8200 1422.5600 ;
        RECT 1152.4600 1422.0800 1155.4600 1422.5600 ;
        RECT 1152.4600 1416.6400 1155.4600 1417.1200 ;
        RECT 1152.4600 1427.5200 1155.4600 1428.0000 ;
        RECT 1164.2200 1427.5200 1165.8200 1428.0000 ;
        RECT 1164.2200 1405.7600 1165.8200 1406.2400 ;
        RECT 1164.2200 1411.2000 1165.8200 1411.6800 ;
        RECT 1152.4600 1411.2000 1155.4600 1411.6800 ;
        RECT 1152.4600 1405.7600 1155.4600 1406.2400 ;
        RECT 1164.2200 1389.4400 1165.8200 1389.9200 ;
        RECT 1164.2200 1394.8800 1165.8200 1395.3600 ;
        RECT 1152.4600 1394.8800 1155.4600 1395.3600 ;
        RECT 1152.4600 1389.4400 1155.4600 1389.9200 ;
        RECT 1152.4600 1400.3200 1155.4600 1400.8000 ;
        RECT 1164.2200 1400.3200 1165.8200 1400.8000 ;
        RECT 1254.2200 1373.1200 1255.8200 1373.6000 ;
        RECT 1254.2200 1378.5600 1255.8200 1379.0400 ;
        RECT 1254.2200 1384.0000 1255.8200 1384.4800 ;
        RECT 1254.2200 1362.2400 1255.8200 1362.7200 ;
        RECT 1254.2200 1367.6800 1255.8200 1368.1600 ;
        RECT 1209.2200 1373.1200 1210.8200 1373.6000 ;
        RECT 1209.2200 1378.5600 1210.8200 1379.0400 ;
        RECT 1209.2200 1384.0000 1210.8200 1384.4800 ;
        RECT 1209.2200 1362.2400 1210.8200 1362.7200 ;
        RECT 1209.2200 1367.6800 1210.8200 1368.1600 ;
        RECT 1254.2200 1345.9200 1255.8200 1346.4000 ;
        RECT 1254.2200 1351.3600 1255.8200 1351.8400 ;
        RECT 1254.2200 1356.8000 1255.8200 1357.2800 ;
        RECT 1254.2200 1335.0400 1255.8200 1335.5200 ;
        RECT 1254.2200 1340.4800 1255.8200 1340.9600 ;
        RECT 1209.2200 1345.9200 1210.8200 1346.4000 ;
        RECT 1209.2200 1351.3600 1210.8200 1351.8400 ;
        RECT 1209.2200 1356.8000 1210.8200 1357.2800 ;
        RECT 1209.2200 1335.0400 1210.8200 1335.5200 ;
        RECT 1209.2200 1340.4800 1210.8200 1340.9600 ;
        RECT 1164.2200 1373.1200 1165.8200 1373.6000 ;
        RECT 1164.2200 1378.5600 1165.8200 1379.0400 ;
        RECT 1164.2200 1384.0000 1165.8200 1384.4800 ;
        RECT 1152.4600 1373.1200 1155.4600 1373.6000 ;
        RECT 1152.4600 1378.5600 1155.4600 1379.0400 ;
        RECT 1152.4600 1384.0000 1155.4600 1384.4800 ;
        RECT 1164.2200 1362.2400 1165.8200 1362.7200 ;
        RECT 1164.2200 1367.6800 1165.8200 1368.1600 ;
        RECT 1152.4600 1362.2400 1155.4600 1362.7200 ;
        RECT 1152.4600 1367.6800 1155.4600 1368.1600 ;
        RECT 1164.2200 1345.9200 1165.8200 1346.4000 ;
        RECT 1164.2200 1351.3600 1165.8200 1351.8400 ;
        RECT 1164.2200 1356.8000 1165.8200 1357.2800 ;
        RECT 1152.4600 1345.9200 1155.4600 1346.4000 ;
        RECT 1152.4600 1351.3600 1155.4600 1351.8400 ;
        RECT 1152.4600 1356.8000 1155.4600 1357.2800 ;
        RECT 1164.2200 1335.0400 1165.8200 1335.5200 ;
        RECT 1164.2200 1340.4800 1165.8200 1340.9600 ;
        RECT 1152.4600 1335.0400 1155.4600 1335.5200 ;
        RECT 1152.4600 1340.4800 1155.4600 1340.9600 ;
        RECT 1356.5600 1318.7200 1359.5600 1319.2000 ;
        RECT 1356.5600 1324.1600 1359.5600 1324.6400 ;
        RECT 1356.5600 1329.6000 1359.5600 1330.0800 ;
        RECT 1344.2200 1318.7200 1345.8200 1319.2000 ;
        RECT 1344.2200 1324.1600 1345.8200 1324.6400 ;
        RECT 1344.2200 1329.6000 1345.8200 1330.0800 ;
        RECT 1356.5600 1307.8400 1359.5600 1308.3200 ;
        RECT 1356.5600 1313.2800 1359.5600 1313.7600 ;
        RECT 1344.2200 1307.8400 1345.8200 1308.3200 ;
        RECT 1344.2200 1313.2800 1345.8200 1313.7600 ;
        RECT 1356.5600 1291.5200 1359.5600 1292.0000 ;
        RECT 1356.5600 1296.9600 1359.5600 1297.4400 ;
        RECT 1356.5600 1302.4000 1359.5600 1302.8800 ;
        RECT 1344.2200 1291.5200 1345.8200 1292.0000 ;
        RECT 1344.2200 1296.9600 1345.8200 1297.4400 ;
        RECT 1344.2200 1302.4000 1345.8200 1302.8800 ;
        RECT 1356.5600 1280.6400 1359.5600 1281.1200 ;
        RECT 1356.5600 1286.0800 1359.5600 1286.5600 ;
        RECT 1344.2200 1280.6400 1345.8200 1281.1200 ;
        RECT 1344.2200 1286.0800 1345.8200 1286.5600 ;
        RECT 1299.2200 1318.7200 1300.8200 1319.2000 ;
        RECT 1299.2200 1324.1600 1300.8200 1324.6400 ;
        RECT 1299.2200 1329.6000 1300.8200 1330.0800 ;
        RECT 1299.2200 1307.8400 1300.8200 1308.3200 ;
        RECT 1299.2200 1313.2800 1300.8200 1313.7600 ;
        RECT 1299.2200 1291.5200 1300.8200 1292.0000 ;
        RECT 1299.2200 1296.9600 1300.8200 1297.4400 ;
        RECT 1299.2200 1302.4000 1300.8200 1302.8800 ;
        RECT 1299.2200 1280.6400 1300.8200 1281.1200 ;
        RECT 1299.2200 1286.0800 1300.8200 1286.5600 ;
        RECT 1356.5600 1264.3200 1359.5600 1264.8000 ;
        RECT 1356.5600 1269.7600 1359.5600 1270.2400 ;
        RECT 1356.5600 1275.2000 1359.5600 1275.6800 ;
        RECT 1344.2200 1264.3200 1345.8200 1264.8000 ;
        RECT 1344.2200 1269.7600 1345.8200 1270.2400 ;
        RECT 1344.2200 1275.2000 1345.8200 1275.6800 ;
        RECT 1356.5600 1253.4400 1359.5600 1253.9200 ;
        RECT 1356.5600 1258.8800 1359.5600 1259.3600 ;
        RECT 1344.2200 1253.4400 1345.8200 1253.9200 ;
        RECT 1344.2200 1258.8800 1345.8200 1259.3600 ;
        RECT 1356.5600 1237.1200 1359.5600 1237.6000 ;
        RECT 1356.5600 1242.5600 1359.5600 1243.0400 ;
        RECT 1356.5600 1248.0000 1359.5600 1248.4800 ;
        RECT 1344.2200 1237.1200 1345.8200 1237.6000 ;
        RECT 1344.2200 1242.5600 1345.8200 1243.0400 ;
        RECT 1344.2200 1248.0000 1345.8200 1248.4800 ;
        RECT 1356.5600 1231.6800 1359.5600 1232.1600 ;
        RECT 1344.2200 1231.6800 1345.8200 1232.1600 ;
        RECT 1299.2200 1264.3200 1300.8200 1264.8000 ;
        RECT 1299.2200 1269.7600 1300.8200 1270.2400 ;
        RECT 1299.2200 1275.2000 1300.8200 1275.6800 ;
        RECT 1299.2200 1253.4400 1300.8200 1253.9200 ;
        RECT 1299.2200 1258.8800 1300.8200 1259.3600 ;
        RECT 1299.2200 1237.1200 1300.8200 1237.6000 ;
        RECT 1299.2200 1242.5600 1300.8200 1243.0400 ;
        RECT 1299.2200 1248.0000 1300.8200 1248.4800 ;
        RECT 1299.2200 1231.6800 1300.8200 1232.1600 ;
        RECT 1254.2200 1318.7200 1255.8200 1319.2000 ;
        RECT 1254.2200 1324.1600 1255.8200 1324.6400 ;
        RECT 1254.2200 1329.6000 1255.8200 1330.0800 ;
        RECT 1254.2200 1307.8400 1255.8200 1308.3200 ;
        RECT 1254.2200 1313.2800 1255.8200 1313.7600 ;
        RECT 1209.2200 1318.7200 1210.8200 1319.2000 ;
        RECT 1209.2200 1324.1600 1210.8200 1324.6400 ;
        RECT 1209.2200 1329.6000 1210.8200 1330.0800 ;
        RECT 1209.2200 1307.8400 1210.8200 1308.3200 ;
        RECT 1209.2200 1313.2800 1210.8200 1313.7600 ;
        RECT 1254.2200 1291.5200 1255.8200 1292.0000 ;
        RECT 1254.2200 1296.9600 1255.8200 1297.4400 ;
        RECT 1254.2200 1302.4000 1255.8200 1302.8800 ;
        RECT 1254.2200 1280.6400 1255.8200 1281.1200 ;
        RECT 1254.2200 1286.0800 1255.8200 1286.5600 ;
        RECT 1209.2200 1291.5200 1210.8200 1292.0000 ;
        RECT 1209.2200 1296.9600 1210.8200 1297.4400 ;
        RECT 1209.2200 1302.4000 1210.8200 1302.8800 ;
        RECT 1209.2200 1280.6400 1210.8200 1281.1200 ;
        RECT 1209.2200 1286.0800 1210.8200 1286.5600 ;
        RECT 1164.2200 1318.7200 1165.8200 1319.2000 ;
        RECT 1164.2200 1324.1600 1165.8200 1324.6400 ;
        RECT 1164.2200 1329.6000 1165.8200 1330.0800 ;
        RECT 1152.4600 1318.7200 1155.4600 1319.2000 ;
        RECT 1152.4600 1324.1600 1155.4600 1324.6400 ;
        RECT 1152.4600 1329.6000 1155.4600 1330.0800 ;
        RECT 1164.2200 1307.8400 1165.8200 1308.3200 ;
        RECT 1164.2200 1313.2800 1165.8200 1313.7600 ;
        RECT 1152.4600 1307.8400 1155.4600 1308.3200 ;
        RECT 1152.4600 1313.2800 1155.4600 1313.7600 ;
        RECT 1164.2200 1291.5200 1165.8200 1292.0000 ;
        RECT 1164.2200 1296.9600 1165.8200 1297.4400 ;
        RECT 1164.2200 1302.4000 1165.8200 1302.8800 ;
        RECT 1152.4600 1291.5200 1155.4600 1292.0000 ;
        RECT 1152.4600 1296.9600 1155.4600 1297.4400 ;
        RECT 1152.4600 1302.4000 1155.4600 1302.8800 ;
        RECT 1164.2200 1280.6400 1165.8200 1281.1200 ;
        RECT 1164.2200 1286.0800 1165.8200 1286.5600 ;
        RECT 1152.4600 1280.6400 1155.4600 1281.1200 ;
        RECT 1152.4600 1286.0800 1155.4600 1286.5600 ;
        RECT 1254.2200 1264.3200 1255.8200 1264.8000 ;
        RECT 1254.2200 1269.7600 1255.8200 1270.2400 ;
        RECT 1254.2200 1275.2000 1255.8200 1275.6800 ;
        RECT 1254.2200 1253.4400 1255.8200 1253.9200 ;
        RECT 1254.2200 1258.8800 1255.8200 1259.3600 ;
        RECT 1209.2200 1264.3200 1210.8200 1264.8000 ;
        RECT 1209.2200 1269.7600 1210.8200 1270.2400 ;
        RECT 1209.2200 1275.2000 1210.8200 1275.6800 ;
        RECT 1209.2200 1253.4400 1210.8200 1253.9200 ;
        RECT 1209.2200 1258.8800 1210.8200 1259.3600 ;
        RECT 1254.2200 1237.1200 1255.8200 1237.6000 ;
        RECT 1254.2200 1242.5600 1255.8200 1243.0400 ;
        RECT 1254.2200 1248.0000 1255.8200 1248.4800 ;
        RECT 1254.2200 1231.6800 1255.8200 1232.1600 ;
        RECT 1209.2200 1237.1200 1210.8200 1237.6000 ;
        RECT 1209.2200 1242.5600 1210.8200 1243.0400 ;
        RECT 1209.2200 1248.0000 1210.8200 1248.4800 ;
        RECT 1209.2200 1231.6800 1210.8200 1232.1600 ;
        RECT 1164.2200 1264.3200 1165.8200 1264.8000 ;
        RECT 1164.2200 1269.7600 1165.8200 1270.2400 ;
        RECT 1164.2200 1275.2000 1165.8200 1275.6800 ;
        RECT 1152.4600 1264.3200 1155.4600 1264.8000 ;
        RECT 1152.4600 1269.7600 1155.4600 1270.2400 ;
        RECT 1152.4600 1275.2000 1155.4600 1275.6800 ;
        RECT 1164.2200 1253.4400 1165.8200 1253.9200 ;
        RECT 1164.2200 1258.8800 1165.8200 1259.3600 ;
        RECT 1152.4600 1253.4400 1155.4600 1253.9200 ;
        RECT 1152.4600 1258.8800 1155.4600 1259.3600 ;
        RECT 1164.2200 1237.1200 1165.8200 1237.6000 ;
        RECT 1164.2200 1242.5600 1165.8200 1243.0400 ;
        RECT 1164.2200 1248.0000 1165.8200 1248.4800 ;
        RECT 1152.4600 1237.1200 1155.4600 1237.6000 ;
        RECT 1152.4600 1242.5600 1155.4600 1243.0400 ;
        RECT 1152.4600 1248.0000 1155.4600 1248.4800 ;
        RECT 1152.4600 1231.6800 1155.4600 1232.1600 ;
        RECT 1164.2200 1231.6800 1165.8200 1232.1600 ;
        RECT 1152.4600 1436.5900 1359.5600 1439.5900 ;
        RECT 1152.4600 1223.4900 1359.5600 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 993.8500 1345.8200 1209.9500 ;
        RECT 1299.2200 993.8500 1300.8200 1209.9500 ;
        RECT 1254.2200 993.8500 1255.8200 1209.9500 ;
        RECT 1209.2200 993.8500 1210.8200 1209.9500 ;
        RECT 1164.2200 993.8500 1165.8200 1209.9500 ;
        RECT 1356.5600 993.8500 1359.5600 1209.9500 ;
        RECT 1152.4600 993.8500 1155.4600 1209.9500 ;
      LAYER met3 ;
        RECT 1356.5600 1187.0000 1359.5600 1187.4800 ;
        RECT 1356.5600 1192.4400 1359.5600 1192.9200 ;
        RECT 1344.2200 1187.0000 1345.8200 1187.4800 ;
        RECT 1344.2200 1192.4400 1345.8200 1192.9200 ;
        RECT 1356.5600 1197.8800 1359.5600 1198.3600 ;
        RECT 1344.2200 1197.8800 1345.8200 1198.3600 ;
        RECT 1356.5600 1176.1200 1359.5600 1176.6000 ;
        RECT 1356.5600 1181.5600 1359.5600 1182.0400 ;
        RECT 1344.2200 1176.1200 1345.8200 1176.6000 ;
        RECT 1344.2200 1181.5600 1345.8200 1182.0400 ;
        RECT 1356.5600 1159.8000 1359.5600 1160.2800 ;
        RECT 1356.5600 1165.2400 1359.5600 1165.7200 ;
        RECT 1344.2200 1159.8000 1345.8200 1160.2800 ;
        RECT 1344.2200 1165.2400 1345.8200 1165.7200 ;
        RECT 1356.5600 1170.6800 1359.5600 1171.1600 ;
        RECT 1344.2200 1170.6800 1345.8200 1171.1600 ;
        RECT 1299.2200 1187.0000 1300.8200 1187.4800 ;
        RECT 1299.2200 1192.4400 1300.8200 1192.9200 ;
        RECT 1299.2200 1197.8800 1300.8200 1198.3600 ;
        RECT 1299.2200 1176.1200 1300.8200 1176.6000 ;
        RECT 1299.2200 1181.5600 1300.8200 1182.0400 ;
        RECT 1299.2200 1159.8000 1300.8200 1160.2800 ;
        RECT 1299.2200 1165.2400 1300.8200 1165.7200 ;
        RECT 1299.2200 1170.6800 1300.8200 1171.1600 ;
        RECT 1356.5600 1143.4800 1359.5600 1143.9600 ;
        RECT 1356.5600 1148.9200 1359.5600 1149.4000 ;
        RECT 1356.5600 1154.3600 1359.5600 1154.8400 ;
        RECT 1344.2200 1143.4800 1345.8200 1143.9600 ;
        RECT 1344.2200 1148.9200 1345.8200 1149.4000 ;
        RECT 1344.2200 1154.3600 1345.8200 1154.8400 ;
        RECT 1356.5600 1132.6000 1359.5600 1133.0800 ;
        RECT 1356.5600 1138.0400 1359.5600 1138.5200 ;
        RECT 1344.2200 1132.6000 1345.8200 1133.0800 ;
        RECT 1344.2200 1138.0400 1345.8200 1138.5200 ;
        RECT 1356.5600 1116.2800 1359.5600 1116.7600 ;
        RECT 1356.5600 1121.7200 1359.5600 1122.2000 ;
        RECT 1356.5600 1127.1600 1359.5600 1127.6400 ;
        RECT 1344.2200 1116.2800 1345.8200 1116.7600 ;
        RECT 1344.2200 1121.7200 1345.8200 1122.2000 ;
        RECT 1344.2200 1127.1600 1345.8200 1127.6400 ;
        RECT 1356.5600 1105.4000 1359.5600 1105.8800 ;
        RECT 1356.5600 1110.8400 1359.5600 1111.3200 ;
        RECT 1344.2200 1105.4000 1345.8200 1105.8800 ;
        RECT 1344.2200 1110.8400 1345.8200 1111.3200 ;
        RECT 1299.2200 1143.4800 1300.8200 1143.9600 ;
        RECT 1299.2200 1148.9200 1300.8200 1149.4000 ;
        RECT 1299.2200 1154.3600 1300.8200 1154.8400 ;
        RECT 1299.2200 1132.6000 1300.8200 1133.0800 ;
        RECT 1299.2200 1138.0400 1300.8200 1138.5200 ;
        RECT 1299.2200 1116.2800 1300.8200 1116.7600 ;
        RECT 1299.2200 1121.7200 1300.8200 1122.2000 ;
        RECT 1299.2200 1127.1600 1300.8200 1127.6400 ;
        RECT 1299.2200 1105.4000 1300.8200 1105.8800 ;
        RECT 1299.2200 1110.8400 1300.8200 1111.3200 ;
        RECT 1254.2200 1187.0000 1255.8200 1187.4800 ;
        RECT 1254.2200 1192.4400 1255.8200 1192.9200 ;
        RECT 1254.2200 1197.8800 1255.8200 1198.3600 ;
        RECT 1209.2200 1187.0000 1210.8200 1187.4800 ;
        RECT 1209.2200 1192.4400 1210.8200 1192.9200 ;
        RECT 1209.2200 1197.8800 1210.8200 1198.3600 ;
        RECT 1254.2200 1176.1200 1255.8200 1176.6000 ;
        RECT 1254.2200 1181.5600 1255.8200 1182.0400 ;
        RECT 1254.2200 1159.8000 1255.8200 1160.2800 ;
        RECT 1254.2200 1165.2400 1255.8200 1165.7200 ;
        RECT 1254.2200 1170.6800 1255.8200 1171.1600 ;
        RECT 1209.2200 1176.1200 1210.8200 1176.6000 ;
        RECT 1209.2200 1181.5600 1210.8200 1182.0400 ;
        RECT 1209.2200 1159.8000 1210.8200 1160.2800 ;
        RECT 1209.2200 1165.2400 1210.8200 1165.7200 ;
        RECT 1209.2200 1170.6800 1210.8200 1171.1600 ;
        RECT 1164.2200 1187.0000 1165.8200 1187.4800 ;
        RECT 1164.2200 1192.4400 1165.8200 1192.9200 ;
        RECT 1152.4600 1192.4400 1155.4600 1192.9200 ;
        RECT 1152.4600 1187.0000 1155.4600 1187.4800 ;
        RECT 1152.4600 1197.8800 1155.4600 1198.3600 ;
        RECT 1164.2200 1197.8800 1165.8200 1198.3600 ;
        RECT 1164.2200 1176.1200 1165.8200 1176.6000 ;
        RECT 1164.2200 1181.5600 1165.8200 1182.0400 ;
        RECT 1152.4600 1181.5600 1155.4600 1182.0400 ;
        RECT 1152.4600 1176.1200 1155.4600 1176.6000 ;
        RECT 1164.2200 1159.8000 1165.8200 1160.2800 ;
        RECT 1164.2200 1165.2400 1165.8200 1165.7200 ;
        RECT 1152.4600 1165.2400 1155.4600 1165.7200 ;
        RECT 1152.4600 1159.8000 1155.4600 1160.2800 ;
        RECT 1152.4600 1170.6800 1155.4600 1171.1600 ;
        RECT 1164.2200 1170.6800 1165.8200 1171.1600 ;
        RECT 1254.2200 1143.4800 1255.8200 1143.9600 ;
        RECT 1254.2200 1148.9200 1255.8200 1149.4000 ;
        RECT 1254.2200 1154.3600 1255.8200 1154.8400 ;
        RECT 1254.2200 1132.6000 1255.8200 1133.0800 ;
        RECT 1254.2200 1138.0400 1255.8200 1138.5200 ;
        RECT 1209.2200 1143.4800 1210.8200 1143.9600 ;
        RECT 1209.2200 1148.9200 1210.8200 1149.4000 ;
        RECT 1209.2200 1154.3600 1210.8200 1154.8400 ;
        RECT 1209.2200 1132.6000 1210.8200 1133.0800 ;
        RECT 1209.2200 1138.0400 1210.8200 1138.5200 ;
        RECT 1254.2200 1116.2800 1255.8200 1116.7600 ;
        RECT 1254.2200 1121.7200 1255.8200 1122.2000 ;
        RECT 1254.2200 1127.1600 1255.8200 1127.6400 ;
        RECT 1254.2200 1105.4000 1255.8200 1105.8800 ;
        RECT 1254.2200 1110.8400 1255.8200 1111.3200 ;
        RECT 1209.2200 1116.2800 1210.8200 1116.7600 ;
        RECT 1209.2200 1121.7200 1210.8200 1122.2000 ;
        RECT 1209.2200 1127.1600 1210.8200 1127.6400 ;
        RECT 1209.2200 1105.4000 1210.8200 1105.8800 ;
        RECT 1209.2200 1110.8400 1210.8200 1111.3200 ;
        RECT 1164.2200 1143.4800 1165.8200 1143.9600 ;
        RECT 1164.2200 1148.9200 1165.8200 1149.4000 ;
        RECT 1164.2200 1154.3600 1165.8200 1154.8400 ;
        RECT 1152.4600 1143.4800 1155.4600 1143.9600 ;
        RECT 1152.4600 1148.9200 1155.4600 1149.4000 ;
        RECT 1152.4600 1154.3600 1155.4600 1154.8400 ;
        RECT 1164.2200 1132.6000 1165.8200 1133.0800 ;
        RECT 1164.2200 1138.0400 1165.8200 1138.5200 ;
        RECT 1152.4600 1132.6000 1155.4600 1133.0800 ;
        RECT 1152.4600 1138.0400 1155.4600 1138.5200 ;
        RECT 1164.2200 1116.2800 1165.8200 1116.7600 ;
        RECT 1164.2200 1121.7200 1165.8200 1122.2000 ;
        RECT 1164.2200 1127.1600 1165.8200 1127.6400 ;
        RECT 1152.4600 1116.2800 1155.4600 1116.7600 ;
        RECT 1152.4600 1121.7200 1155.4600 1122.2000 ;
        RECT 1152.4600 1127.1600 1155.4600 1127.6400 ;
        RECT 1164.2200 1105.4000 1165.8200 1105.8800 ;
        RECT 1164.2200 1110.8400 1165.8200 1111.3200 ;
        RECT 1152.4600 1105.4000 1155.4600 1105.8800 ;
        RECT 1152.4600 1110.8400 1155.4600 1111.3200 ;
        RECT 1356.5600 1089.0800 1359.5600 1089.5600 ;
        RECT 1356.5600 1094.5200 1359.5600 1095.0000 ;
        RECT 1356.5600 1099.9600 1359.5600 1100.4400 ;
        RECT 1344.2200 1089.0800 1345.8200 1089.5600 ;
        RECT 1344.2200 1094.5200 1345.8200 1095.0000 ;
        RECT 1344.2200 1099.9600 1345.8200 1100.4400 ;
        RECT 1356.5600 1078.2000 1359.5600 1078.6800 ;
        RECT 1356.5600 1083.6400 1359.5600 1084.1200 ;
        RECT 1344.2200 1078.2000 1345.8200 1078.6800 ;
        RECT 1344.2200 1083.6400 1345.8200 1084.1200 ;
        RECT 1356.5600 1061.8800 1359.5600 1062.3600 ;
        RECT 1356.5600 1067.3200 1359.5600 1067.8000 ;
        RECT 1356.5600 1072.7600 1359.5600 1073.2400 ;
        RECT 1344.2200 1061.8800 1345.8200 1062.3600 ;
        RECT 1344.2200 1067.3200 1345.8200 1067.8000 ;
        RECT 1344.2200 1072.7600 1345.8200 1073.2400 ;
        RECT 1356.5600 1051.0000 1359.5600 1051.4800 ;
        RECT 1356.5600 1056.4400 1359.5600 1056.9200 ;
        RECT 1344.2200 1051.0000 1345.8200 1051.4800 ;
        RECT 1344.2200 1056.4400 1345.8200 1056.9200 ;
        RECT 1299.2200 1089.0800 1300.8200 1089.5600 ;
        RECT 1299.2200 1094.5200 1300.8200 1095.0000 ;
        RECT 1299.2200 1099.9600 1300.8200 1100.4400 ;
        RECT 1299.2200 1078.2000 1300.8200 1078.6800 ;
        RECT 1299.2200 1083.6400 1300.8200 1084.1200 ;
        RECT 1299.2200 1061.8800 1300.8200 1062.3600 ;
        RECT 1299.2200 1067.3200 1300.8200 1067.8000 ;
        RECT 1299.2200 1072.7600 1300.8200 1073.2400 ;
        RECT 1299.2200 1051.0000 1300.8200 1051.4800 ;
        RECT 1299.2200 1056.4400 1300.8200 1056.9200 ;
        RECT 1356.5600 1034.6800 1359.5600 1035.1600 ;
        RECT 1356.5600 1040.1200 1359.5600 1040.6000 ;
        RECT 1356.5600 1045.5600 1359.5600 1046.0400 ;
        RECT 1344.2200 1034.6800 1345.8200 1035.1600 ;
        RECT 1344.2200 1040.1200 1345.8200 1040.6000 ;
        RECT 1344.2200 1045.5600 1345.8200 1046.0400 ;
        RECT 1356.5600 1023.8000 1359.5600 1024.2800 ;
        RECT 1356.5600 1029.2400 1359.5600 1029.7200 ;
        RECT 1344.2200 1023.8000 1345.8200 1024.2800 ;
        RECT 1344.2200 1029.2400 1345.8200 1029.7200 ;
        RECT 1356.5600 1007.4800 1359.5600 1007.9600 ;
        RECT 1356.5600 1012.9200 1359.5600 1013.4000 ;
        RECT 1356.5600 1018.3600 1359.5600 1018.8400 ;
        RECT 1344.2200 1007.4800 1345.8200 1007.9600 ;
        RECT 1344.2200 1012.9200 1345.8200 1013.4000 ;
        RECT 1344.2200 1018.3600 1345.8200 1018.8400 ;
        RECT 1356.5600 1002.0400 1359.5600 1002.5200 ;
        RECT 1344.2200 1002.0400 1345.8200 1002.5200 ;
        RECT 1299.2200 1034.6800 1300.8200 1035.1600 ;
        RECT 1299.2200 1040.1200 1300.8200 1040.6000 ;
        RECT 1299.2200 1045.5600 1300.8200 1046.0400 ;
        RECT 1299.2200 1023.8000 1300.8200 1024.2800 ;
        RECT 1299.2200 1029.2400 1300.8200 1029.7200 ;
        RECT 1299.2200 1007.4800 1300.8200 1007.9600 ;
        RECT 1299.2200 1012.9200 1300.8200 1013.4000 ;
        RECT 1299.2200 1018.3600 1300.8200 1018.8400 ;
        RECT 1299.2200 1002.0400 1300.8200 1002.5200 ;
        RECT 1254.2200 1089.0800 1255.8200 1089.5600 ;
        RECT 1254.2200 1094.5200 1255.8200 1095.0000 ;
        RECT 1254.2200 1099.9600 1255.8200 1100.4400 ;
        RECT 1254.2200 1078.2000 1255.8200 1078.6800 ;
        RECT 1254.2200 1083.6400 1255.8200 1084.1200 ;
        RECT 1209.2200 1089.0800 1210.8200 1089.5600 ;
        RECT 1209.2200 1094.5200 1210.8200 1095.0000 ;
        RECT 1209.2200 1099.9600 1210.8200 1100.4400 ;
        RECT 1209.2200 1078.2000 1210.8200 1078.6800 ;
        RECT 1209.2200 1083.6400 1210.8200 1084.1200 ;
        RECT 1254.2200 1061.8800 1255.8200 1062.3600 ;
        RECT 1254.2200 1067.3200 1255.8200 1067.8000 ;
        RECT 1254.2200 1072.7600 1255.8200 1073.2400 ;
        RECT 1254.2200 1051.0000 1255.8200 1051.4800 ;
        RECT 1254.2200 1056.4400 1255.8200 1056.9200 ;
        RECT 1209.2200 1061.8800 1210.8200 1062.3600 ;
        RECT 1209.2200 1067.3200 1210.8200 1067.8000 ;
        RECT 1209.2200 1072.7600 1210.8200 1073.2400 ;
        RECT 1209.2200 1051.0000 1210.8200 1051.4800 ;
        RECT 1209.2200 1056.4400 1210.8200 1056.9200 ;
        RECT 1164.2200 1089.0800 1165.8200 1089.5600 ;
        RECT 1164.2200 1094.5200 1165.8200 1095.0000 ;
        RECT 1164.2200 1099.9600 1165.8200 1100.4400 ;
        RECT 1152.4600 1089.0800 1155.4600 1089.5600 ;
        RECT 1152.4600 1094.5200 1155.4600 1095.0000 ;
        RECT 1152.4600 1099.9600 1155.4600 1100.4400 ;
        RECT 1164.2200 1078.2000 1165.8200 1078.6800 ;
        RECT 1164.2200 1083.6400 1165.8200 1084.1200 ;
        RECT 1152.4600 1078.2000 1155.4600 1078.6800 ;
        RECT 1152.4600 1083.6400 1155.4600 1084.1200 ;
        RECT 1164.2200 1061.8800 1165.8200 1062.3600 ;
        RECT 1164.2200 1067.3200 1165.8200 1067.8000 ;
        RECT 1164.2200 1072.7600 1165.8200 1073.2400 ;
        RECT 1152.4600 1061.8800 1155.4600 1062.3600 ;
        RECT 1152.4600 1067.3200 1155.4600 1067.8000 ;
        RECT 1152.4600 1072.7600 1155.4600 1073.2400 ;
        RECT 1164.2200 1051.0000 1165.8200 1051.4800 ;
        RECT 1164.2200 1056.4400 1165.8200 1056.9200 ;
        RECT 1152.4600 1051.0000 1155.4600 1051.4800 ;
        RECT 1152.4600 1056.4400 1155.4600 1056.9200 ;
        RECT 1254.2200 1034.6800 1255.8200 1035.1600 ;
        RECT 1254.2200 1040.1200 1255.8200 1040.6000 ;
        RECT 1254.2200 1045.5600 1255.8200 1046.0400 ;
        RECT 1254.2200 1023.8000 1255.8200 1024.2800 ;
        RECT 1254.2200 1029.2400 1255.8200 1029.7200 ;
        RECT 1209.2200 1034.6800 1210.8200 1035.1600 ;
        RECT 1209.2200 1040.1200 1210.8200 1040.6000 ;
        RECT 1209.2200 1045.5600 1210.8200 1046.0400 ;
        RECT 1209.2200 1023.8000 1210.8200 1024.2800 ;
        RECT 1209.2200 1029.2400 1210.8200 1029.7200 ;
        RECT 1254.2200 1007.4800 1255.8200 1007.9600 ;
        RECT 1254.2200 1012.9200 1255.8200 1013.4000 ;
        RECT 1254.2200 1018.3600 1255.8200 1018.8400 ;
        RECT 1254.2200 1002.0400 1255.8200 1002.5200 ;
        RECT 1209.2200 1007.4800 1210.8200 1007.9600 ;
        RECT 1209.2200 1012.9200 1210.8200 1013.4000 ;
        RECT 1209.2200 1018.3600 1210.8200 1018.8400 ;
        RECT 1209.2200 1002.0400 1210.8200 1002.5200 ;
        RECT 1164.2200 1034.6800 1165.8200 1035.1600 ;
        RECT 1164.2200 1040.1200 1165.8200 1040.6000 ;
        RECT 1164.2200 1045.5600 1165.8200 1046.0400 ;
        RECT 1152.4600 1034.6800 1155.4600 1035.1600 ;
        RECT 1152.4600 1040.1200 1155.4600 1040.6000 ;
        RECT 1152.4600 1045.5600 1155.4600 1046.0400 ;
        RECT 1164.2200 1023.8000 1165.8200 1024.2800 ;
        RECT 1164.2200 1029.2400 1165.8200 1029.7200 ;
        RECT 1152.4600 1023.8000 1155.4600 1024.2800 ;
        RECT 1152.4600 1029.2400 1155.4600 1029.7200 ;
        RECT 1164.2200 1007.4800 1165.8200 1007.9600 ;
        RECT 1164.2200 1012.9200 1165.8200 1013.4000 ;
        RECT 1164.2200 1018.3600 1165.8200 1018.8400 ;
        RECT 1152.4600 1007.4800 1155.4600 1007.9600 ;
        RECT 1152.4600 1012.9200 1155.4600 1013.4000 ;
        RECT 1152.4600 1018.3600 1155.4600 1018.8400 ;
        RECT 1152.4600 1002.0400 1155.4600 1002.5200 ;
        RECT 1164.2200 1002.0400 1165.8200 1002.5200 ;
        RECT 1152.4600 1206.9500 1359.5600 1209.9500 ;
        RECT 1152.4600 993.8500 1359.5600 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1344.2200 764.2100 1345.8200 980.3100 ;
        RECT 1299.2200 764.2100 1300.8200 980.3100 ;
        RECT 1254.2200 764.2100 1255.8200 980.3100 ;
        RECT 1209.2200 764.2100 1210.8200 980.3100 ;
        RECT 1164.2200 764.2100 1165.8200 980.3100 ;
        RECT 1356.5600 764.2100 1359.5600 980.3100 ;
        RECT 1152.4600 764.2100 1155.4600 980.3100 ;
      LAYER met3 ;
        RECT 1356.5600 957.3600 1359.5600 957.8400 ;
        RECT 1356.5600 962.8000 1359.5600 963.2800 ;
        RECT 1344.2200 957.3600 1345.8200 957.8400 ;
        RECT 1344.2200 962.8000 1345.8200 963.2800 ;
        RECT 1356.5600 968.2400 1359.5600 968.7200 ;
        RECT 1344.2200 968.2400 1345.8200 968.7200 ;
        RECT 1356.5600 946.4800 1359.5600 946.9600 ;
        RECT 1356.5600 951.9200 1359.5600 952.4000 ;
        RECT 1344.2200 946.4800 1345.8200 946.9600 ;
        RECT 1344.2200 951.9200 1345.8200 952.4000 ;
        RECT 1356.5600 930.1600 1359.5600 930.6400 ;
        RECT 1356.5600 935.6000 1359.5600 936.0800 ;
        RECT 1344.2200 930.1600 1345.8200 930.6400 ;
        RECT 1344.2200 935.6000 1345.8200 936.0800 ;
        RECT 1356.5600 941.0400 1359.5600 941.5200 ;
        RECT 1344.2200 941.0400 1345.8200 941.5200 ;
        RECT 1299.2200 957.3600 1300.8200 957.8400 ;
        RECT 1299.2200 962.8000 1300.8200 963.2800 ;
        RECT 1299.2200 968.2400 1300.8200 968.7200 ;
        RECT 1299.2200 946.4800 1300.8200 946.9600 ;
        RECT 1299.2200 951.9200 1300.8200 952.4000 ;
        RECT 1299.2200 930.1600 1300.8200 930.6400 ;
        RECT 1299.2200 935.6000 1300.8200 936.0800 ;
        RECT 1299.2200 941.0400 1300.8200 941.5200 ;
        RECT 1356.5600 913.8400 1359.5600 914.3200 ;
        RECT 1356.5600 919.2800 1359.5600 919.7600 ;
        RECT 1356.5600 924.7200 1359.5600 925.2000 ;
        RECT 1344.2200 913.8400 1345.8200 914.3200 ;
        RECT 1344.2200 919.2800 1345.8200 919.7600 ;
        RECT 1344.2200 924.7200 1345.8200 925.2000 ;
        RECT 1356.5600 902.9600 1359.5600 903.4400 ;
        RECT 1356.5600 908.4000 1359.5600 908.8800 ;
        RECT 1344.2200 902.9600 1345.8200 903.4400 ;
        RECT 1344.2200 908.4000 1345.8200 908.8800 ;
        RECT 1356.5600 886.6400 1359.5600 887.1200 ;
        RECT 1356.5600 892.0800 1359.5600 892.5600 ;
        RECT 1356.5600 897.5200 1359.5600 898.0000 ;
        RECT 1344.2200 886.6400 1345.8200 887.1200 ;
        RECT 1344.2200 892.0800 1345.8200 892.5600 ;
        RECT 1344.2200 897.5200 1345.8200 898.0000 ;
        RECT 1356.5600 875.7600 1359.5600 876.2400 ;
        RECT 1356.5600 881.2000 1359.5600 881.6800 ;
        RECT 1344.2200 875.7600 1345.8200 876.2400 ;
        RECT 1344.2200 881.2000 1345.8200 881.6800 ;
        RECT 1299.2200 913.8400 1300.8200 914.3200 ;
        RECT 1299.2200 919.2800 1300.8200 919.7600 ;
        RECT 1299.2200 924.7200 1300.8200 925.2000 ;
        RECT 1299.2200 902.9600 1300.8200 903.4400 ;
        RECT 1299.2200 908.4000 1300.8200 908.8800 ;
        RECT 1299.2200 886.6400 1300.8200 887.1200 ;
        RECT 1299.2200 892.0800 1300.8200 892.5600 ;
        RECT 1299.2200 897.5200 1300.8200 898.0000 ;
        RECT 1299.2200 875.7600 1300.8200 876.2400 ;
        RECT 1299.2200 881.2000 1300.8200 881.6800 ;
        RECT 1254.2200 957.3600 1255.8200 957.8400 ;
        RECT 1254.2200 962.8000 1255.8200 963.2800 ;
        RECT 1254.2200 968.2400 1255.8200 968.7200 ;
        RECT 1209.2200 957.3600 1210.8200 957.8400 ;
        RECT 1209.2200 962.8000 1210.8200 963.2800 ;
        RECT 1209.2200 968.2400 1210.8200 968.7200 ;
        RECT 1254.2200 946.4800 1255.8200 946.9600 ;
        RECT 1254.2200 951.9200 1255.8200 952.4000 ;
        RECT 1254.2200 930.1600 1255.8200 930.6400 ;
        RECT 1254.2200 935.6000 1255.8200 936.0800 ;
        RECT 1254.2200 941.0400 1255.8200 941.5200 ;
        RECT 1209.2200 946.4800 1210.8200 946.9600 ;
        RECT 1209.2200 951.9200 1210.8200 952.4000 ;
        RECT 1209.2200 930.1600 1210.8200 930.6400 ;
        RECT 1209.2200 935.6000 1210.8200 936.0800 ;
        RECT 1209.2200 941.0400 1210.8200 941.5200 ;
        RECT 1164.2200 957.3600 1165.8200 957.8400 ;
        RECT 1164.2200 962.8000 1165.8200 963.2800 ;
        RECT 1152.4600 962.8000 1155.4600 963.2800 ;
        RECT 1152.4600 957.3600 1155.4600 957.8400 ;
        RECT 1152.4600 968.2400 1155.4600 968.7200 ;
        RECT 1164.2200 968.2400 1165.8200 968.7200 ;
        RECT 1164.2200 946.4800 1165.8200 946.9600 ;
        RECT 1164.2200 951.9200 1165.8200 952.4000 ;
        RECT 1152.4600 951.9200 1155.4600 952.4000 ;
        RECT 1152.4600 946.4800 1155.4600 946.9600 ;
        RECT 1164.2200 930.1600 1165.8200 930.6400 ;
        RECT 1164.2200 935.6000 1165.8200 936.0800 ;
        RECT 1152.4600 935.6000 1155.4600 936.0800 ;
        RECT 1152.4600 930.1600 1155.4600 930.6400 ;
        RECT 1152.4600 941.0400 1155.4600 941.5200 ;
        RECT 1164.2200 941.0400 1165.8200 941.5200 ;
        RECT 1254.2200 913.8400 1255.8200 914.3200 ;
        RECT 1254.2200 919.2800 1255.8200 919.7600 ;
        RECT 1254.2200 924.7200 1255.8200 925.2000 ;
        RECT 1254.2200 902.9600 1255.8200 903.4400 ;
        RECT 1254.2200 908.4000 1255.8200 908.8800 ;
        RECT 1209.2200 913.8400 1210.8200 914.3200 ;
        RECT 1209.2200 919.2800 1210.8200 919.7600 ;
        RECT 1209.2200 924.7200 1210.8200 925.2000 ;
        RECT 1209.2200 902.9600 1210.8200 903.4400 ;
        RECT 1209.2200 908.4000 1210.8200 908.8800 ;
        RECT 1254.2200 886.6400 1255.8200 887.1200 ;
        RECT 1254.2200 892.0800 1255.8200 892.5600 ;
        RECT 1254.2200 897.5200 1255.8200 898.0000 ;
        RECT 1254.2200 875.7600 1255.8200 876.2400 ;
        RECT 1254.2200 881.2000 1255.8200 881.6800 ;
        RECT 1209.2200 886.6400 1210.8200 887.1200 ;
        RECT 1209.2200 892.0800 1210.8200 892.5600 ;
        RECT 1209.2200 897.5200 1210.8200 898.0000 ;
        RECT 1209.2200 875.7600 1210.8200 876.2400 ;
        RECT 1209.2200 881.2000 1210.8200 881.6800 ;
        RECT 1164.2200 913.8400 1165.8200 914.3200 ;
        RECT 1164.2200 919.2800 1165.8200 919.7600 ;
        RECT 1164.2200 924.7200 1165.8200 925.2000 ;
        RECT 1152.4600 913.8400 1155.4600 914.3200 ;
        RECT 1152.4600 919.2800 1155.4600 919.7600 ;
        RECT 1152.4600 924.7200 1155.4600 925.2000 ;
        RECT 1164.2200 902.9600 1165.8200 903.4400 ;
        RECT 1164.2200 908.4000 1165.8200 908.8800 ;
        RECT 1152.4600 902.9600 1155.4600 903.4400 ;
        RECT 1152.4600 908.4000 1155.4600 908.8800 ;
        RECT 1164.2200 886.6400 1165.8200 887.1200 ;
        RECT 1164.2200 892.0800 1165.8200 892.5600 ;
        RECT 1164.2200 897.5200 1165.8200 898.0000 ;
        RECT 1152.4600 886.6400 1155.4600 887.1200 ;
        RECT 1152.4600 892.0800 1155.4600 892.5600 ;
        RECT 1152.4600 897.5200 1155.4600 898.0000 ;
        RECT 1164.2200 875.7600 1165.8200 876.2400 ;
        RECT 1164.2200 881.2000 1165.8200 881.6800 ;
        RECT 1152.4600 875.7600 1155.4600 876.2400 ;
        RECT 1152.4600 881.2000 1155.4600 881.6800 ;
        RECT 1356.5600 859.4400 1359.5600 859.9200 ;
        RECT 1356.5600 864.8800 1359.5600 865.3600 ;
        RECT 1356.5600 870.3200 1359.5600 870.8000 ;
        RECT 1344.2200 859.4400 1345.8200 859.9200 ;
        RECT 1344.2200 864.8800 1345.8200 865.3600 ;
        RECT 1344.2200 870.3200 1345.8200 870.8000 ;
        RECT 1356.5600 848.5600 1359.5600 849.0400 ;
        RECT 1356.5600 854.0000 1359.5600 854.4800 ;
        RECT 1344.2200 848.5600 1345.8200 849.0400 ;
        RECT 1344.2200 854.0000 1345.8200 854.4800 ;
        RECT 1356.5600 832.2400 1359.5600 832.7200 ;
        RECT 1356.5600 837.6800 1359.5600 838.1600 ;
        RECT 1356.5600 843.1200 1359.5600 843.6000 ;
        RECT 1344.2200 832.2400 1345.8200 832.7200 ;
        RECT 1344.2200 837.6800 1345.8200 838.1600 ;
        RECT 1344.2200 843.1200 1345.8200 843.6000 ;
        RECT 1356.5600 821.3600 1359.5600 821.8400 ;
        RECT 1356.5600 826.8000 1359.5600 827.2800 ;
        RECT 1344.2200 821.3600 1345.8200 821.8400 ;
        RECT 1344.2200 826.8000 1345.8200 827.2800 ;
        RECT 1299.2200 859.4400 1300.8200 859.9200 ;
        RECT 1299.2200 864.8800 1300.8200 865.3600 ;
        RECT 1299.2200 870.3200 1300.8200 870.8000 ;
        RECT 1299.2200 848.5600 1300.8200 849.0400 ;
        RECT 1299.2200 854.0000 1300.8200 854.4800 ;
        RECT 1299.2200 832.2400 1300.8200 832.7200 ;
        RECT 1299.2200 837.6800 1300.8200 838.1600 ;
        RECT 1299.2200 843.1200 1300.8200 843.6000 ;
        RECT 1299.2200 821.3600 1300.8200 821.8400 ;
        RECT 1299.2200 826.8000 1300.8200 827.2800 ;
        RECT 1356.5600 805.0400 1359.5600 805.5200 ;
        RECT 1356.5600 810.4800 1359.5600 810.9600 ;
        RECT 1356.5600 815.9200 1359.5600 816.4000 ;
        RECT 1344.2200 805.0400 1345.8200 805.5200 ;
        RECT 1344.2200 810.4800 1345.8200 810.9600 ;
        RECT 1344.2200 815.9200 1345.8200 816.4000 ;
        RECT 1356.5600 794.1600 1359.5600 794.6400 ;
        RECT 1356.5600 799.6000 1359.5600 800.0800 ;
        RECT 1344.2200 794.1600 1345.8200 794.6400 ;
        RECT 1344.2200 799.6000 1345.8200 800.0800 ;
        RECT 1356.5600 777.8400 1359.5600 778.3200 ;
        RECT 1356.5600 783.2800 1359.5600 783.7600 ;
        RECT 1356.5600 788.7200 1359.5600 789.2000 ;
        RECT 1344.2200 777.8400 1345.8200 778.3200 ;
        RECT 1344.2200 783.2800 1345.8200 783.7600 ;
        RECT 1344.2200 788.7200 1345.8200 789.2000 ;
        RECT 1356.5600 772.4000 1359.5600 772.8800 ;
        RECT 1344.2200 772.4000 1345.8200 772.8800 ;
        RECT 1299.2200 805.0400 1300.8200 805.5200 ;
        RECT 1299.2200 810.4800 1300.8200 810.9600 ;
        RECT 1299.2200 815.9200 1300.8200 816.4000 ;
        RECT 1299.2200 794.1600 1300.8200 794.6400 ;
        RECT 1299.2200 799.6000 1300.8200 800.0800 ;
        RECT 1299.2200 777.8400 1300.8200 778.3200 ;
        RECT 1299.2200 783.2800 1300.8200 783.7600 ;
        RECT 1299.2200 788.7200 1300.8200 789.2000 ;
        RECT 1299.2200 772.4000 1300.8200 772.8800 ;
        RECT 1254.2200 859.4400 1255.8200 859.9200 ;
        RECT 1254.2200 864.8800 1255.8200 865.3600 ;
        RECT 1254.2200 870.3200 1255.8200 870.8000 ;
        RECT 1254.2200 848.5600 1255.8200 849.0400 ;
        RECT 1254.2200 854.0000 1255.8200 854.4800 ;
        RECT 1209.2200 859.4400 1210.8200 859.9200 ;
        RECT 1209.2200 864.8800 1210.8200 865.3600 ;
        RECT 1209.2200 870.3200 1210.8200 870.8000 ;
        RECT 1209.2200 848.5600 1210.8200 849.0400 ;
        RECT 1209.2200 854.0000 1210.8200 854.4800 ;
        RECT 1254.2200 832.2400 1255.8200 832.7200 ;
        RECT 1254.2200 837.6800 1255.8200 838.1600 ;
        RECT 1254.2200 843.1200 1255.8200 843.6000 ;
        RECT 1254.2200 821.3600 1255.8200 821.8400 ;
        RECT 1254.2200 826.8000 1255.8200 827.2800 ;
        RECT 1209.2200 832.2400 1210.8200 832.7200 ;
        RECT 1209.2200 837.6800 1210.8200 838.1600 ;
        RECT 1209.2200 843.1200 1210.8200 843.6000 ;
        RECT 1209.2200 821.3600 1210.8200 821.8400 ;
        RECT 1209.2200 826.8000 1210.8200 827.2800 ;
        RECT 1164.2200 859.4400 1165.8200 859.9200 ;
        RECT 1164.2200 864.8800 1165.8200 865.3600 ;
        RECT 1164.2200 870.3200 1165.8200 870.8000 ;
        RECT 1152.4600 859.4400 1155.4600 859.9200 ;
        RECT 1152.4600 864.8800 1155.4600 865.3600 ;
        RECT 1152.4600 870.3200 1155.4600 870.8000 ;
        RECT 1164.2200 848.5600 1165.8200 849.0400 ;
        RECT 1164.2200 854.0000 1165.8200 854.4800 ;
        RECT 1152.4600 848.5600 1155.4600 849.0400 ;
        RECT 1152.4600 854.0000 1155.4600 854.4800 ;
        RECT 1164.2200 832.2400 1165.8200 832.7200 ;
        RECT 1164.2200 837.6800 1165.8200 838.1600 ;
        RECT 1164.2200 843.1200 1165.8200 843.6000 ;
        RECT 1152.4600 832.2400 1155.4600 832.7200 ;
        RECT 1152.4600 837.6800 1155.4600 838.1600 ;
        RECT 1152.4600 843.1200 1155.4600 843.6000 ;
        RECT 1164.2200 821.3600 1165.8200 821.8400 ;
        RECT 1164.2200 826.8000 1165.8200 827.2800 ;
        RECT 1152.4600 821.3600 1155.4600 821.8400 ;
        RECT 1152.4600 826.8000 1155.4600 827.2800 ;
        RECT 1254.2200 805.0400 1255.8200 805.5200 ;
        RECT 1254.2200 810.4800 1255.8200 810.9600 ;
        RECT 1254.2200 815.9200 1255.8200 816.4000 ;
        RECT 1254.2200 794.1600 1255.8200 794.6400 ;
        RECT 1254.2200 799.6000 1255.8200 800.0800 ;
        RECT 1209.2200 805.0400 1210.8200 805.5200 ;
        RECT 1209.2200 810.4800 1210.8200 810.9600 ;
        RECT 1209.2200 815.9200 1210.8200 816.4000 ;
        RECT 1209.2200 794.1600 1210.8200 794.6400 ;
        RECT 1209.2200 799.6000 1210.8200 800.0800 ;
        RECT 1254.2200 777.8400 1255.8200 778.3200 ;
        RECT 1254.2200 783.2800 1255.8200 783.7600 ;
        RECT 1254.2200 788.7200 1255.8200 789.2000 ;
        RECT 1254.2200 772.4000 1255.8200 772.8800 ;
        RECT 1209.2200 777.8400 1210.8200 778.3200 ;
        RECT 1209.2200 783.2800 1210.8200 783.7600 ;
        RECT 1209.2200 788.7200 1210.8200 789.2000 ;
        RECT 1209.2200 772.4000 1210.8200 772.8800 ;
        RECT 1164.2200 805.0400 1165.8200 805.5200 ;
        RECT 1164.2200 810.4800 1165.8200 810.9600 ;
        RECT 1164.2200 815.9200 1165.8200 816.4000 ;
        RECT 1152.4600 805.0400 1155.4600 805.5200 ;
        RECT 1152.4600 810.4800 1155.4600 810.9600 ;
        RECT 1152.4600 815.9200 1155.4600 816.4000 ;
        RECT 1164.2200 794.1600 1165.8200 794.6400 ;
        RECT 1164.2200 799.6000 1165.8200 800.0800 ;
        RECT 1152.4600 794.1600 1155.4600 794.6400 ;
        RECT 1152.4600 799.6000 1155.4600 800.0800 ;
        RECT 1164.2200 777.8400 1165.8200 778.3200 ;
        RECT 1164.2200 783.2800 1165.8200 783.7600 ;
        RECT 1164.2200 788.7200 1165.8200 789.2000 ;
        RECT 1152.4600 777.8400 1155.4600 778.3200 ;
        RECT 1152.4600 783.2800 1155.4600 783.7600 ;
        RECT 1152.4600 788.7200 1155.4600 789.2000 ;
        RECT 1152.4600 772.4000 1155.4600 772.8800 ;
        RECT 1164.2200 772.4000 1165.8200 772.8800 ;
        RECT 1152.4600 977.3100 1359.5600 980.3100 ;
        RECT 1152.4600 764.2100 1359.5600 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1373.6800 2830.6100 1375.6800 2857.5400 ;
        RECT 1576.7800 2830.6100 1578.7800 2857.5400 ;
      LAYER met3 ;
        RECT 1576.7800 2847.3200 1578.7800 2847.8000 ;
        RECT 1373.6800 2847.3200 1375.6800 2847.8000 ;
        RECT 1576.7800 2841.8800 1578.7800 2842.3600 ;
        RECT 1576.7800 2836.4400 1578.7800 2836.9200 ;
        RECT 1373.6800 2841.8800 1375.6800 2842.3600 ;
        RECT 1373.6800 2836.4400 1375.6800 2836.9200 ;
        RECT 1373.6800 2855.5400 1578.7800 2857.5400 ;
        RECT 1373.6800 2830.6100 1578.7800 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 534.5700 1566.0400 750.6700 ;
        RECT 1519.4400 534.5700 1521.0400 750.6700 ;
        RECT 1474.4400 534.5700 1476.0400 750.6700 ;
        RECT 1429.4400 534.5700 1431.0400 750.6700 ;
        RECT 1384.4400 534.5700 1386.0400 750.6700 ;
        RECT 1576.7800 534.5700 1579.7800 750.6700 ;
        RECT 1372.6800 534.5700 1375.6800 750.6700 ;
      LAYER met3 ;
        RECT 1576.7800 727.7200 1579.7800 728.2000 ;
        RECT 1576.7800 733.1600 1579.7800 733.6400 ;
        RECT 1564.4400 727.7200 1566.0400 728.2000 ;
        RECT 1564.4400 733.1600 1566.0400 733.6400 ;
        RECT 1576.7800 738.6000 1579.7800 739.0800 ;
        RECT 1564.4400 738.6000 1566.0400 739.0800 ;
        RECT 1576.7800 716.8400 1579.7800 717.3200 ;
        RECT 1576.7800 722.2800 1579.7800 722.7600 ;
        RECT 1564.4400 716.8400 1566.0400 717.3200 ;
        RECT 1564.4400 722.2800 1566.0400 722.7600 ;
        RECT 1576.7800 700.5200 1579.7800 701.0000 ;
        RECT 1576.7800 705.9600 1579.7800 706.4400 ;
        RECT 1564.4400 700.5200 1566.0400 701.0000 ;
        RECT 1564.4400 705.9600 1566.0400 706.4400 ;
        RECT 1576.7800 711.4000 1579.7800 711.8800 ;
        RECT 1564.4400 711.4000 1566.0400 711.8800 ;
        RECT 1519.4400 727.7200 1521.0400 728.2000 ;
        RECT 1519.4400 733.1600 1521.0400 733.6400 ;
        RECT 1519.4400 738.6000 1521.0400 739.0800 ;
        RECT 1519.4400 716.8400 1521.0400 717.3200 ;
        RECT 1519.4400 722.2800 1521.0400 722.7600 ;
        RECT 1519.4400 700.5200 1521.0400 701.0000 ;
        RECT 1519.4400 705.9600 1521.0400 706.4400 ;
        RECT 1519.4400 711.4000 1521.0400 711.8800 ;
        RECT 1576.7800 684.2000 1579.7800 684.6800 ;
        RECT 1576.7800 689.6400 1579.7800 690.1200 ;
        RECT 1576.7800 695.0800 1579.7800 695.5600 ;
        RECT 1564.4400 684.2000 1566.0400 684.6800 ;
        RECT 1564.4400 689.6400 1566.0400 690.1200 ;
        RECT 1564.4400 695.0800 1566.0400 695.5600 ;
        RECT 1576.7800 673.3200 1579.7800 673.8000 ;
        RECT 1576.7800 678.7600 1579.7800 679.2400 ;
        RECT 1564.4400 673.3200 1566.0400 673.8000 ;
        RECT 1564.4400 678.7600 1566.0400 679.2400 ;
        RECT 1576.7800 657.0000 1579.7800 657.4800 ;
        RECT 1576.7800 662.4400 1579.7800 662.9200 ;
        RECT 1576.7800 667.8800 1579.7800 668.3600 ;
        RECT 1564.4400 657.0000 1566.0400 657.4800 ;
        RECT 1564.4400 662.4400 1566.0400 662.9200 ;
        RECT 1564.4400 667.8800 1566.0400 668.3600 ;
        RECT 1576.7800 646.1200 1579.7800 646.6000 ;
        RECT 1576.7800 651.5600 1579.7800 652.0400 ;
        RECT 1564.4400 646.1200 1566.0400 646.6000 ;
        RECT 1564.4400 651.5600 1566.0400 652.0400 ;
        RECT 1519.4400 684.2000 1521.0400 684.6800 ;
        RECT 1519.4400 689.6400 1521.0400 690.1200 ;
        RECT 1519.4400 695.0800 1521.0400 695.5600 ;
        RECT 1519.4400 673.3200 1521.0400 673.8000 ;
        RECT 1519.4400 678.7600 1521.0400 679.2400 ;
        RECT 1519.4400 657.0000 1521.0400 657.4800 ;
        RECT 1519.4400 662.4400 1521.0400 662.9200 ;
        RECT 1519.4400 667.8800 1521.0400 668.3600 ;
        RECT 1519.4400 646.1200 1521.0400 646.6000 ;
        RECT 1519.4400 651.5600 1521.0400 652.0400 ;
        RECT 1474.4400 727.7200 1476.0400 728.2000 ;
        RECT 1474.4400 733.1600 1476.0400 733.6400 ;
        RECT 1474.4400 738.6000 1476.0400 739.0800 ;
        RECT 1429.4400 727.7200 1431.0400 728.2000 ;
        RECT 1429.4400 733.1600 1431.0400 733.6400 ;
        RECT 1429.4400 738.6000 1431.0400 739.0800 ;
        RECT 1474.4400 716.8400 1476.0400 717.3200 ;
        RECT 1474.4400 722.2800 1476.0400 722.7600 ;
        RECT 1474.4400 700.5200 1476.0400 701.0000 ;
        RECT 1474.4400 705.9600 1476.0400 706.4400 ;
        RECT 1474.4400 711.4000 1476.0400 711.8800 ;
        RECT 1429.4400 716.8400 1431.0400 717.3200 ;
        RECT 1429.4400 722.2800 1431.0400 722.7600 ;
        RECT 1429.4400 700.5200 1431.0400 701.0000 ;
        RECT 1429.4400 705.9600 1431.0400 706.4400 ;
        RECT 1429.4400 711.4000 1431.0400 711.8800 ;
        RECT 1384.4400 727.7200 1386.0400 728.2000 ;
        RECT 1384.4400 733.1600 1386.0400 733.6400 ;
        RECT 1372.6800 733.1600 1375.6800 733.6400 ;
        RECT 1372.6800 727.7200 1375.6800 728.2000 ;
        RECT 1372.6800 738.6000 1375.6800 739.0800 ;
        RECT 1384.4400 738.6000 1386.0400 739.0800 ;
        RECT 1384.4400 716.8400 1386.0400 717.3200 ;
        RECT 1384.4400 722.2800 1386.0400 722.7600 ;
        RECT 1372.6800 722.2800 1375.6800 722.7600 ;
        RECT 1372.6800 716.8400 1375.6800 717.3200 ;
        RECT 1384.4400 700.5200 1386.0400 701.0000 ;
        RECT 1384.4400 705.9600 1386.0400 706.4400 ;
        RECT 1372.6800 705.9600 1375.6800 706.4400 ;
        RECT 1372.6800 700.5200 1375.6800 701.0000 ;
        RECT 1372.6800 711.4000 1375.6800 711.8800 ;
        RECT 1384.4400 711.4000 1386.0400 711.8800 ;
        RECT 1474.4400 684.2000 1476.0400 684.6800 ;
        RECT 1474.4400 689.6400 1476.0400 690.1200 ;
        RECT 1474.4400 695.0800 1476.0400 695.5600 ;
        RECT 1474.4400 673.3200 1476.0400 673.8000 ;
        RECT 1474.4400 678.7600 1476.0400 679.2400 ;
        RECT 1429.4400 684.2000 1431.0400 684.6800 ;
        RECT 1429.4400 689.6400 1431.0400 690.1200 ;
        RECT 1429.4400 695.0800 1431.0400 695.5600 ;
        RECT 1429.4400 673.3200 1431.0400 673.8000 ;
        RECT 1429.4400 678.7600 1431.0400 679.2400 ;
        RECT 1474.4400 657.0000 1476.0400 657.4800 ;
        RECT 1474.4400 662.4400 1476.0400 662.9200 ;
        RECT 1474.4400 667.8800 1476.0400 668.3600 ;
        RECT 1474.4400 646.1200 1476.0400 646.6000 ;
        RECT 1474.4400 651.5600 1476.0400 652.0400 ;
        RECT 1429.4400 657.0000 1431.0400 657.4800 ;
        RECT 1429.4400 662.4400 1431.0400 662.9200 ;
        RECT 1429.4400 667.8800 1431.0400 668.3600 ;
        RECT 1429.4400 646.1200 1431.0400 646.6000 ;
        RECT 1429.4400 651.5600 1431.0400 652.0400 ;
        RECT 1384.4400 684.2000 1386.0400 684.6800 ;
        RECT 1384.4400 689.6400 1386.0400 690.1200 ;
        RECT 1384.4400 695.0800 1386.0400 695.5600 ;
        RECT 1372.6800 684.2000 1375.6800 684.6800 ;
        RECT 1372.6800 689.6400 1375.6800 690.1200 ;
        RECT 1372.6800 695.0800 1375.6800 695.5600 ;
        RECT 1384.4400 673.3200 1386.0400 673.8000 ;
        RECT 1384.4400 678.7600 1386.0400 679.2400 ;
        RECT 1372.6800 673.3200 1375.6800 673.8000 ;
        RECT 1372.6800 678.7600 1375.6800 679.2400 ;
        RECT 1384.4400 657.0000 1386.0400 657.4800 ;
        RECT 1384.4400 662.4400 1386.0400 662.9200 ;
        RECT 1384.4400 667.8800 1386.0400 668.3600 ;
        RECT 1372.6800 657.0000 1375.6800 657.4800 ;
        RECT 1372.6800 662.4400 1375.6800 662.9200 ;
        RECT 1372.6800 667.8800 1375.6800 668.3600 ;
        RECT 1384.4400 646.1200 1386.0400 646.6000 ;
        RECT 1384.4400 651.5600 1386.0400 652.0400 ;
        RECT 1372.6800 646.1200 1375.6800 646.6000 ;
        RECT 1372.6800 651.5600 1375.6800 652.0400 ;
        RECT 1576.7800 629.8000 1579.7800 630.2800 ;
        RECT 1576.7800 635.2400 1579.7800 635.7200 ;
        RECT 1576.7800 640.6800 1579.7800 641.1600 ;
        RECT 1564.4400 629.8000 1566.0400 630.2800 ;
        RECT 1564.4400 635.2400 1566.0400 635.7200 ;
        RECT 1564.4400 640.6800 1566.0400 641.1600 ;
        RECT 1576.7800 618.9200 1579.7800 619.4000 ;
        RECT 1576.7800 624.3600 1579.7800 624.8400 ;
        RECT 1564.4400 618.9200 1566.0400 619.4000 ;
        RECT 1564.4400 624.3600 1566.0400 624.8400 ;
        RECT 1576.7800 602.6000 1579.7800 603.0800 ;
        RECT 1576.7800 608.0400 1579.7800 608.5200 ;
        RECT 1576.7800 613.4800 1579.7800 613.9600 ;
        RECT 1564.4400 602.6000 1566.0400 603.0800 ;
        RECT 1564.4400 608.0400 1566.0400 608.5200 ;
        RECT 1564.4400 613.4800 1566.0400 613.9600 ;
        RECT 1576.7800 591.7200 1579.7800 592.2000 ;
        RECT 1576.7800 597.1600 1579.7800 597.6400 ;
        RECT 1564.4400 591.7200 1566.0400 592.2000 ;
        RECT 1564.4400 597.1600 1566.0400 597.6400 ;
        RECT 1519.4400 629.8000 1521.0400 630.2800 ;
        RECT 1519.4400 635.2400 1521.0400 635.7200 ;
        RECT 1519.4400 640.6800 1521.0400 641.1600 ;
        RECT 1519.4400 618.9200 1521.0400 619.4000 ;
        RECT 1519.4400 624.3600 1521.0400 624.8400 ;
        RECT 1519.4400 602.6000 1521.0400 603.0800 ;
        RECT 1519.4400 608.0400 1521.0400 608.5200 ;
        RECT 1519.4400 613.4800 1521.0400 613.9600 ;
        RECT 1519.4400 591.7200 1521.0400 592.2000 ;
        RECT 1519.4400 597.1600 1521.0400 597.6400 ;
        RECT 1576.7800 575.4000 1579.7800 575.8800 ;
        RECT 1576.7800 580.8400 1579.7800 581.3200 ;
        RECT 1576.7800 586.2800 1579.7800 586.7600 ;
        RECT 1564.4400 575.4000 1566.0400 575.8800 ;
        RECT 1564.4400 580.8400 1566.0400 581.3200 ;
        RECT 1564.4400 586.2800 1566.0400 586.7600 ;
        RECT 1576.7800 564.5200 1579.7800 565.0000 ;
        RECT 1576.7800 569.9600 1579.7800 570.4400 ;
        RECT 1564.4400 564.5200 1566.0400 565.0000 ;
        RECT 1564.4400 569.9600 1566.0400 570.4400 ;
        RECT 1576.7800 548.2000 1579.7800 548.6800 ;
        RECT 1576.7800 553.6400 1579.7800 554.1200 ;
        RECT 1576.7800 559.0800 1579.7800 559.5600 ;
        RECT 1564.4400 548.2000 1566.0400 548.6800 ;
        RECT 1564.4400 553.6400 1566.0400 554.1200 ;
        RECT 1564.4400 559.0800 1566.0400 559.5600 ;
        RECT 1576.7800 542.7600 1579.7800 543.2400 ;
        RECT 1564.4400 542.7600 1566.0400 543.2400 ;
        RECT 1519.4400 575.4000 1521.0400 575.8800 ;
        RECT 1519.4400 580.8400 1521.0400 581.3200 ;
        RECT 1519.4400 586.2800 1521.0400 586.7600 ;
        RECT 1519.4400 564.5200 1521.0400 565.0000 ;
        RECT 1519.4400 569.9600 1521.0400 570.4400 ;
        RECT 1519.4400 548.2000 1521.0400 548.6800 ;
        RECT 1519.4400 553.6400 1521.0400 554.1200 ;
        RECT 1519.4400 559.0800 1521.0400 559.5600 ;
        RECT 1519.4400 542.7600 1521.0400 543.2400 ;
        RECT 1474.4400 629.8000 1476.0400 630.2800 ;
        RECT 1474.4400 635.2400 1476.0400 635.7200 ;
        RECT 1474.4400 640.6800 1476.0400 641.1600 ;
        RECT 1474.4400 618.9200 1476.0400 619.4000 ;
        RECT 1474.4400 624.3600 1476.0400 624.8400 ;
        RECT 1429.4400 629.8000 1431.0400 630.2800 ;
        RECT 1429.4400 635.2400 1431.0400 635.7200 ;
        RECT 1429.4400 640.6800 1431.0400 641.1600 ;
        RECT 1429.4400 618.9200 1431.0400 619.4000 ;
        RECT 1429.4400 624.3600 1431.0400 624.8400 ;
        RECT 1474.4400 602.6000 1476.0400 603.0800 ;
        RECT 1474.4400 608.0400 1476.0400 608.5200 ;
        RECT 1474.4400 613.4800 1476.0400 613.9600 ;
        RECT 1474.4400 591.7200 1476.0400 592.2000 ;
        RECT 1474.4400 597.1600 1476.0400 597.6400 ;
        RECT 1429.4400 602.6000 1431.0400 603.0800 ;
        RECT 1429.4400 608.0400 1431.0400 608.5200 ;
        RECT 1429.4400 613.4800 1431.0400 613.9600 ;
        RECT 1429.4400 591.7200 1431.0400 592.2000 ;
        RECT 1429.4400 597.1600 1431.0400 597.6400 ;
        RECT 1384.4400 629.8000 1386.0400 630.2800 ;
        RECT 1384.4400 635.2400 1386.0400 635.7200 ;
        RECT 1384.4400 640.6800 1386.0400 641.1600 ;
        RECT 1372.6800 629.8000 1375.6800 630.2800 ;
        RECT 1372.6800 635.2400 1375.6800 635.7200 ;
        RECT 1372.6800 640.6800 1375.6800 641.1600 ;
        RECT 1384.4400 618.9200 1386.0400 619.4000 ;
        RECT 1384.4400 624.3600 1386.0400 624.8400 ;
        RECT 1372.6800 618.9200 1375.6800 619.4000 ;
        RECT 1372.6800 624.3600 1375.6800 624.8400 ;
        RECT 1384.4400 602.6000 1386.0400 603.0800 ;
        RECT 1384.4400 608.0400 1386.0400 608.5200 ;
        RECT 1384.4400 613.4800 1386.0400 613.9600 ;
        RECT 1372.6800 602.6000 1375.6800 603.0800 ;
        RECT 1372.6800 608.0400 1375.6800 608.5200 ;
        RECT 1372.6800 613.4800 1375.6800 613.9600 ;
        RECT 1384.4400 591.7200 1386.0400 592.2000 ;
        RECT 1384.4400 597.1600 1386.0400 597.6400 ;
        RECT 1372.6800 591.7200 1375.6800 592.2000 ;
        RECT 1372.6800 597.1600 1375.6800 597.6400 ;
        RECT 1474.4400 575.4000 1476.0400 575.8800 ;
        RECT 1474.4400 580.8400 1476.0400 581.3200 ;
        RECT 1474.4400 586.2800 1476.0400 586.7600 ;
        RECT 1474.4400 564.5200 1476.0400 565.0000 ;
        RECT 1474.4400 569.9600 1476.0400 570.4400 ;
        RECT 1429.4400 575.4000 1431.0400 575.8800 ;
        RECT 1429.4400 580.8400 1431.0400 581.3200 ;
        RECT 1429.4400 586.2800 1431.0400 586.7600 ;
        RECT 1429.4400 564.5200 1431.0400 565.0000 ;
        RECT 1429.4400 569.9600 1431.0400 570.4400 ;
        RECT 1474.4400 548.2000 1476.0400 548.6800 ;
        RECT 1474.4400 553.6400 1476.0400 554.1200 ;
        RECT 1474.4400 559.0800 1476.0400 559.5600 ;
        RECT 1474.4400 542.7600 1476.0400 543.2400 ;
        RECT 1429.4400 548.2000 1431.0400 548.6800 ;
        RECT 1429.4400 553.6400 1431.0400 554.1200 ;
        RECT 1429.4400 559.0800 1431.0400 559.5600 ;
        RECT 1429.4400 542.7600 1431.0400 543.2400 ;
        RECT 1384.4400 575.4000 1386.0400 575.8800 ;
        RECT 1384.4400 580.8400 1386.0400 581.3200 ;
        RECT 1384.4400 586.2800 1386.0400 586.7600 ;
        RECT 1372.6800 575.4000 1375.6800 575.8800 ;
        RECT 1372.6800 580.8400 1375.6800 581.3200 ;
        RECT 1372.6800 586.2800 1375.6800 586.7600 ;
        RECT 1384.4400 564.5200 1386.0400 565.0000 ;
        RECT 1384.4400 569.9600 1386.0400 570.4400 ;
        RECT 1372.6800 564.5200 1375.6800 565.0000 ;
        RECT 1372.6800 569.9600 1375.6800 570.4400 ;
        RECT 1384.4400 548.2000 1386.0400 548.6800 ;
        RECT 1384.4400 553.6400 1386.0400 554.1200 ;
        RECT 1384.4400 559.0800 1386.0400 559.5600 ;
        RECT 1372.6800 548.2000 1375.6800 548.6800 ;
        RECT 1372.6800 553.6400 1375.6800 554.1200 ;
        RECT 1372.6800 559.0800 1375.6800 559.5600 ;
        RECT 1372.6800 542.7600 1375.6800 543.2400 ;
        RECT 1384.4400 542.7600 1386.0400 543.2400 ;
        RECT 1372.6800 747.6700 1579.7800 750.6700 ;
        RECT 1372.6800 534.5700 1579.7800 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 304.9300 1566.0400 521.0300 ;
        RECT 1519.4400 304.9300 1521.0400 521.0300 ;
        RECT 1474.4400 304.9300 1476.0400 521.0300 ;
        RECT 1429.4400 304.9300 1431.0400 521.0300 ;
        RECT 1384.4400 304.9300 1386.0400 521.0300 ;
        RECT 1576.7800 304.9300 1579.7800 521.0300 ;
        RECT 1372.6800 304.9300 1375.6800 521.0300 ;
      LAYER met3 ;
        RECT 1576.7800 498.0800 1579.7800 498.5600 ;
        RECT 1576.7800 503.5200 1579.7800 504.0000 ;
        RECT 1564.4400 498.0800 1566.0400 498.5600 ;
        RECT 1564.4400 503.5200 1566.0400 504.0000 ;
        RECT 1576.7800 508.9600 1579.7800 509.4400 ;
        RECT 1564.4400 508.9600 1566.0400 509.4400 ;
        RECT 1576.7800 487.2000 1579.7800 487.6800 ;
        RECT 1576.7800 492.6400 1579.7800 493.1200 ;
        RECT 1564.4400 487.2000 1566.0400 487.6800 ;
        RECT 1564.4400 492.6400 1566.0400 493.1200 ;
        RECT 1576.7800 470.8800 1579.7800 471.3600 ;
        RECT 1576.7800 476.3200 1579.7800 476.8000 ;
        RECT 1564.4400 470.8800 1566.0400 471.3600 ;
        RECT 1564.4400 476.3200 1566.0400 476.8000 ;
        RECT 1576.7800 481.7600 1579.7800 482.2400 ;
        RECT 1564.4400 481.7600 1566.0400 482.2400 ;
        RECT 1519.4400 498.0800 1521.0400 498.5600 ;
        RECT 1519.4400 503.5200 1521.0400 504.0000 ;
        RECT 1519.4400 508.9600 1521.0400 509.4400 ;
        RECT 1519.4400 487.2000 1521.0400 487.6800 ;
        RECT 1519.4400 492.6400 1521.0400 493.1200 ;
        RECT 1519.4400 470.8800 1521.0400 471.3600 ;
        RECT 1519.4400 476.3200 1521.0400 476.8000 ;
        RECT 1519.4400 481.7600 1521.0400 482.2400 ;
        RECT 1576.7800 454.5600 1579.7800 455.0400 ;
        RECT 1576.7800 460.0000 1579.7800 460.4800 ;
        RECT 1576.7800 465.4400 1579.7800 465.9200 ;
        RECT 1564.4400 454.5600 1566.0400 455.0400 ;
        RECT 1564.4400 460.0000 1566.0400 460.4800 ;
        RECT 1564.4400 465.4400 1566.0400 465.9200 ;
        RECT 1576.7800 443.6800 1579.7800 444.1600 ;
        RECT 1576.7800 449.1200 1579.7800 449.6000 ;
        RECT 1564.4400 443.6800 1566.0400 444.1600 ;
        RECT 1564.4400 449.1200 1566.0400 449.6000 ;
        RECT 1576.7800 427.3600 1579.7800 427.8400 ;
        RECT 1576.7800 432.8000 1579.7800 433.2800 ;
        RECT 1576.7800 438.2400 1579.7800 438.7200 ;
        RECT 1564.4400 427.3600 1566.0400 427.8400 ;
        RECT 1564.4400 432.8000 1566.0400 433.2800 ;
        RECT 1564.4400 438.2400 1566.0400 438.7200 ;
        RECT 1576.7800 416.4800 1579.7800 416.9600 ;
        RECT 1576.7800 421.9200 1579.7800 422.4000 ;
        RECT 1564.4400 416.4800 1566.0400 416.9600 ;
        RECT 1564.4400 421.9200 1566.0400 422.4000 ;
        RECT 1519.4400 454.5600 1521.0400 455.0400 ;
        RECT 1519.4400 460.0000 1521.0400 460.4800 ;
        RECT 1519.4400 465.4400 1521.0400 465.9200 ;
        RECT 1519.4400 443.6800 1521.0400 444.1600 ;
        RECT 1519.4400 449.1200 1521.0400 449.6000 ;
        RECT 1519.4400 427.3600 1521.0400 427.8400 ;
        RECT 1519.4400 432.8000 1521.0400 433.2800 ;
        RECT 1519.4400 438.2400 1521.0400 438.7200 ;
        RECT 1519.4400 416.4800 1521.0400 416.9600 ;
        RECT 1519.4400 421.9200 1521.0400 422.4000 ;
        RECT 1474.4400 498.0800 1476.0400 498.5600 ;
        RECT 1474.4400 503.5200 1476.0400 504.0000 ;
        RECT 1474.4400 508.9600 1476.0400 509.4400 ;
        RECT 1429.4400 498.0800 1431.0400 498.5600 ;
        RECT 1429.4400 503.5200 1431.0400 504.0000 ;
        RECT 1429.4400 508.9600 1431.0400 509.4400 ;
        RECT 1474.4400 487.2000 1476.0400 487.6800 ;
        RECT 1474.4400 492.6400 1476.0400 493.1200 ;
        RECT 1474.4400 470.8800 1476.0400 471.3600 ;
        RECT 1474.4400 476.3200 1476.0400 476.8000 ;
        RECT 1474.4400 481.7600 1476.0400 482.2400 ;
        RECT 1429.4400 487.2000 1431.0400 487.6800 ;
        RECT 1429.4400 492.6400 1431.0400 493.1200 ;
        RECT 1429.4400 470.8800 1431.0400 471.3600 ;
        RECT 1429.4400 476.3200 1431.0400 476.8000 ;
        RECT 1429.4400 481.7600 1431.0400 482.2400 ;
        RECT 1384.4400 498.0800 1386.0400 498.5600 ;
        RECT 1384.4400 503.5200 1386.0400 504.0000 ;
        RECT 1372.6800 503.5200 1375.6800 504.0000 ;
        RECT 1372.6800 498.0800 1375.6800 498.5600 ;
        RECT 1372.6800 508.9600 1375.6800 509.4400 ;
        RECT 1384.4400 508.9600 1386.0400 509.4400 ;
        RECT 1384.4400 487.2000 1386.0400 487.6800 ;
        RECT 1384.4400 492.6400 1386.0400 493.1200 ;
        RECT 1372.6800 492.6400 1375.6800 493.1200 ;
        RECT 1372.6800 487.2000 1375.6800 487.6800 ;
        RECT 1384.4400 470.8800 1386.0400 471.3600 ;
        RECT 1384.4400 476.3200 1386.0400 476.8000 ;
        RECT 1372.6800 476.3200 1375.6800 476.8000 ;
        RECT 1372.6800 470.8800 1375.6800 471.3600 ;
        RECT 1372.6800 481.7600 1375.6800 482.2400 ;
        RECT 1384.4400 481.7600 1386.0400 482.2400 ;
        RECT 1474.4400 454.5600 1476.0400 455.0400 ;
        RECT 1474.4400 460.0000 1476.0400 460.4800 ;
        RECT 1474.4400 465.4400 1476.0400 465.9200 ;
        RECT 1474.4400 443.6800 1476.0400 444.1600 ;
        RECT 1474.4400 449.1200 1476.0400 449.6000 ;
        RECT 1429.4400 454.5600 1431.0400 455.0400 ;
        RECT 1429.4400 460.0000 1431.0400 460.4800 ;
        RECT 1429.4400 465.4400 1431.0400 465.9200 ;
        RECT 1429.4400 443.6800 1431.0400 444.1600 ;
        RECT 1429.4400 449.1200 1431.0400 449.6000 ;
        RECT 1474.4400 427.3600 1476.0400 427.8400 ;
        RECT 1474.4400 432.8000 1476.0400 433.2800 ;
        RECT 1474.4400 438.2400 1476.0400 438.7200 ;
        RECT 1474.4400 416.4800 1476.0400 416.9600 ;
        RECT 1474.4400 421.9200 1476.0400 422.4000 ;
        RECT 1429.4400 427.3600 1431.0400 427.8400 ;
        RECT 1429.4400 432.8000 1431.0400 433.2800 ;
        RECT 1429.4400 438.2400 1431.0400 438.7200 ;
        RECT 1429.4400 416.4800 1431.0400 416.9600 ;
        RECT 1429.4400 421.9200 1431.0400 422.4000 ;
        RECT 1384.4400 454.5600 1386.0400 455.0400 ;
        RECT 1384.4400 460.0000 1386.0400 460.4800 ;
        RECT 1384.4400 465.4400 1386.0400 465.9200 ;
        RECT 1372.6800 454.5600 1375.6800 455.0400 ;
        RECT 1372.6800 460.0000 1375.6800 460.4800 ;
        RECT 1372.6800 465.4400 1375.6800 465.9200 ;
        RECT 1384.4400 443.6800 1386.0400 444.1600 ;
        RECT 1384.4400 449.1200 1386.0400 449.6000 ;
        RECT 1372.6800 443.6800 1375.6800 444.1600 ;
        RECT 1372.6800 449.1200 1375.6800 449.6000 ;
        RECT 1384.4400 427.3600 1386.0400 427.8400 ;
        RECT 1384.4400 432.8000 1386.0400 433.2800 ;
        RECT 1384.4400 438.2400 1386.0400 438.7200 ;
        RECT 1372.6800 427.3600 1375.6800 427.8400 ;
        RECT 1372.6800 432.8000 1375.6800 433.2800 ;
        RECT 1372.6800 438.2400 1375.6800 438.7200 ;
        RECT 1384.4400 416.4800 1386.0400 416.9600 ;
        RECT 1384.4400 421.9200 1386.0400 422.4000 ;
        RECT 1372.6800 416.4800 1375.6800 416.9600 ;
        RECT 1372.6800 421.9200 1375.6800 422.4000 ;
        RECT 1576.7800 400.1600 1579.7800 400.6400 ;
        RECT 1576.7800 405.6000 1579.7800 406.0800 ;
        RECT 1576.7800 411.0400 1579.7800 411.5200 ;
        RECT 1564.4400 400.1600 1566.0400 400.6400 ;
        RECT 1564.4400 405.6000 1566.0400 406.0800 ;
        RECT 1564.4400 411.0400 1566.0400 411.5200 ;
        RECT 1576.7800 389.2800 1579.7800 389.7600 ;
        RECT 1576.7800 394.7200 1579.7800 395.2000 ;
        RECT 1564.4400 389.2800 1566.0400 389.7600 ;
        RECT 1564.4400 394.7200 1566.0400 395.2000 ;
        RECT 1576.7800 372.9600 1579.7800 373.4400 ;
        RECT 1576.7800 378.4000 1579.7800 378.8800 ;
        RECT 1576.7800 383.8400 1579.7800 384.3200 ;
        RECT 1564.4400 372.9600 1566.0400 373.4400 ;
        RECT 1564.4400 378.4000 1566.0400 378.8800 ;
        RECT 1564.4400 383.8400 1566.0400 384.3200 ;
        RECT 1576.7800 362.0800 1579.7800 362.5600 ;
        RECT 1576.7800 367.5200 1579.7800 368.0000 ;
        RECT 1564.4400 362.0800 1566.0400 362.5600 ;
        RECT 1564.4400 367.5200 1566.0400 368.0000 ;
        RECT 1519.4400 400.1600 1521.0400 400.6400 ;
        RECT 1519.4400 405.6000 1521.0400 406.0800 ;
        RECT 1519.4400 411.0400 1521.0400 411.5200 ;
        RECT 1519.4400 389.2800 1521.0400 389.7600 ;
        RECT 1519.4400 394.7200 1521.0400 395.2000 ;
        RECT 1519.4400 372.9600 1521.0400 373.4400 ;
        RECT 1519.4400 378.4000 1521.0400 378.8800 ;
        RECT 1519.4400 383.8400 1521.0400 384.3200 ;
        RECT 1519.4400 362.0800 1521.0400 362.5600 ;
        RECT 1519.4400 367.5200 1521.0400 368.0000 ;
        RECT 1576.7800 345.7600 1579.7800 346.2400 ;
        RECT 1576.7800 351.2000 1579.7800 351.6800 ;
        RECT 1576.7800 356.6400 1579.7800 357.1200 ;
        RECT 1564.4400 345.7600 1566.0400 346.2400 ;
        RECT 1564.4400 351.2000 1566.0400 351.6800 ;
        RECT 1564.4400 356.6400 1566.0400 357.1200 ;
        RECT 1576.7800 334.8800 1579.7800 335.3600 ;
        RECT 1576.7800 340.3200 1579.7800 340.8000 ;
        RECT 1564.4400 334.8800 1566.0400 335.3600 ;
        RECT 1564.4400 340.3200 1566.0400 340.8000 ;
        RECT 1576.7800 318.5600 1579.7800 319.0400 ;
        RECT 1576.7800 324.0000 1579.7800 324.4800 ;
        RECT 1576.7800 329.4400 1579.7800 329.9200 ;
        RECT 1564.4400 318.5600 1566.0400 319.0400 ;
        RECT 1564.4400 324.0000 1566.0400 324.4800 ;
        RECT 1564.4400 329.4400 1566.0400 329.9200 ;
        RECT 1576.7800 313.1200 1579.7800 313.6000 ;
        RECT 1564.4400 313.1200 1566.0400 313.6000 ;
        RECT 1519.4400 345.7600 1521.0400 346.2400 ;
        RECT 1519.4400 351.2000 1521.0400 351.6800 ;
        RECT 1519.4400 356.6400 1521.0400 357.1200 ;
        RECT 1519.4400 334.8800 1521.0400 335.3600 ;
        RECT 1519.4400 340.3200 1521.0400 340.8000 ;
        RECT 1519.4400 318.5600 1521.0400 319.0400 ;
        RECT 1519.4400 324.0000 1521.0400 324.4800 ;
        RECT 1519.4400 329.4400 1521.0400 329.9200 ;
        RECT 1519.4400 313.1200 1521.0400 313.6000 ;
        RECT 1474.4400 400.1600 1476.0400 400.6400 ;
        RECT 1474.4400 405.6000 1476.0400 406.0800 ;
        RECT 1474.4400 411.0400 1476.0400 411.5200 ;
        RECT 1474.4400 389.2800 1476.0400 389.7600 ;
        RECT 1474.4400 394.7200 1476.0400 395.2000 ;
        RECT 1429.4400 400.1600 1431.0400 400.6400 ;
        RECT 1429.4400 405.6000 1431.0400 406.0800 ;
        RECT 1429.4400 411.0400 1431.0400 411.5200 ;
        RECT 1429.4400 389.2800 1431.0400 389.7600 ;
        RECT 1429.4400 394.7200 1431.0400 395.2000 ;
        RECT 1474.4400 372.9600 1476.0400 373.4400 ;
        RECT 1474.4400 378.4000 1476.0400 378.8800 ;
        RECT 1474.4400 383.8400 1476.0400 384.3200 ;
        RECT 1474.4400 362.0800 1476.0400 362.5600 ;
        RECT 1474.4400 367.5200 1476.0400 368.0000 ;
        RECT 1429.4400 372.9600 1431.0400 373.4400 ;
        RECT 1429.4400 378.4000 1431.0400 378.8800 ;
        RECT 1429.4400 383.8400 1431.0400 384.3200 ;
        RECT 1429.4400 362.0800 1431.0400 362.5600 ;
        RECT 1429.4400 367.5200 1431.0400 368.0000 ;
        RECT 1384.4400 400.1600 1386.0400 400.6400 ;
        RECT 1384.4400 405.6000 1386.0400 406.0800 ;
        RECT 1384.4400 411.0400 1386.0400 411.5200 ;
        RECT 1372.6800 400.1600 1375.6800 400.6400 ;
        RECT 1372.6800 405.6000 1375.6800 406.0800 ;
        RECT 1372.6800 411.0400 1375.6800 411.5200 ;
        RECT 1384.4400 389.2800 1386.0400 389.7600 ;
        RECT 1384.4400 394.7200 1386.0400 395.2000 ;
        RECT 1372.6800 389.2800 1375.6800 389.7600 ;
        RECT 1372.6800 394.7200 1375.6800 395.2000 ;
        RECT 1384.4400 372.9600 1386.0400 373.4400 ;
        RECT 1384.4400 378.4000 1386.0400 378.8800 ;
        RECT 1384.4400 383.8400 1386.0400 384.3200 ;
        RECT 1372.6800 372.9600 1375.6800 373.4400 ;
        RECT 1372.6800 378.4000 1375.6800 378.8800 ;
        RECT 1372.6800 383.8400 1375.6800 384.3200 ;
        RECT 1384.4400 362.0800 1386.0400 362.5600 ;
        RECT 1384.4400 367.5200 1386.0400 368.0000 ;
        RECT 1372.6800 362.0800 1375.6800 362.5600 ;
        RECT 1372.6800 367.5200 1375.6800 368.0000 ;
        RECT 1474.4400 345.7600 1476.0400 346.2400 ;
        RECT 1474.4400 351.2000 1476.0400 351.6800 ;
        RECT 1474.4400 356.6400 1476.0400 357.1200 ;
        RECT 1474.4400 334.8800 1476.0400 335.3600 ;
        RECT 1474.4400 340.3200 1476.0400 340.8000 ;
        RECT 1429.4400 345.7600 1431.0400 346.2400 ;
        RECT 1429.4400 351.2000 1431.0400 351.6800 ;
        RECT 1429.4400 356.6400 1431.0400 357.1200 ;
        RECT 1429.4400 334.8800 1431.0400 335.3600 ;
        RECT 1429.4400 340.3200 1431.0400 340.8000 ;
        RECT 1474.4400 318.5600 1476.0400 319.0400 ;
        RECT 1474.4400 324.0000 1476.0400 324.4800 ;
        RECT 1474.4400 329.4400 1476.0400 329.9200 ;
        RECT 1474.4400 313.1200 1476.0400 313.6000 ;
        RECT 1429.4400 318.5600 1431.0400 319.0400 ;
        RECT 1429.4400 324.0000 1431.0400 324.4800 ;
        RECT 1429.4400 329.4400 1431.0400 329.9200 ;
        RECT 1429.4400 313.1200 1431.0400 313.6000 ;
        RECT 1384.4400 345.7600 1386.0400 346.2400 ;
        RECT 1384.4400 351.2000 1386.0400 351.6800 ;
        RECT 1384.4400 356.6400 1386.0400 357.1200 ;
        RECT 1372.6800 345.7600 1375.6800 346.2400 ;
        RECT 1372.6800 351.2000 1375.6800 351.6800 ;
        RECT 1372.6800 356.6400 1375.6800 357.1200 ;
        RECT 1384.4400 334.8800 1386.0400 335.3600 ;
        RECT 1384.4400 340.3200 1386.0400 340.8000 ;
        RECT 1372.6800 334.8800 1375.6800 335.3600 ;
        RECT 1372.6800 340.3200 1375.6800 340.8000 ;
        RECT 1384.4400 318.5600 1386.0400 319.0400 ;
        RECT 1384.4400 324.0000 1386.0400 324.4800 ;
        RECT 1384.4400 329.4400 1386.0400 329.9200 ;
        RECT 1372.6800 318.5600 1375.6800 319.0400 ;
        RECT 1372.6800 324.0000 1375.6800 324.4800 ;
        RECT 1372.6800 329.4400 1375.6800 329.9200 ;
        RECT 1372.6800 313.1200 1375.6800 313.6000 ;
        RECT 1384.4400 313.1200 1386.0400 313.6000 ;
        RECT 1372.6800 518.0300 1579.7800 521.0300 ;
        RECT 1372.6800 304.9300 1579.7800 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 75.2900 1566.0400 291.3900 ;
        RECT 1519.4400 75.2900 1521.0400 291.3900 ;
        RECT 1474.4400 75.2900 1476.0400 291.3900 ;
        RECT 1429.4400 75.2900 1431.0400 291.3900 ;
        RECT 1384.4400 75.2900 1386.0400 291.3900 ;
        RECT 1576.7800 75.2900 1579.7800 291.3900 ;
        RECT 1372.6800 75.2900 1375.6800 291.3900 ;
      LAYER met3 ;
        RECT 1576.7800 268.4400 1579.7800 268.9200 ;
        RECT 1576.7800 273.8800 1579.7800 274.3600 ;
        RECT 1564.4400 268.4400 1566.0400 268.9200 ;
        RECT 1564.4400 273.8800 1566.0400 274.3600 ;
        RECT 1576.7800 279.3200 1579.7800 279.8000 ;
        RECT 1564.4400 279.3200 1566.0400 279.8000 ;
        RECT 1576.7800 257.5600 1579.7800 258.0400 ;
        RECT 1576.7800 263.0000 1579.7800 263.4800 ;
        RECT 1564.4400 257.5600 1566.0400 258.0400 ;
        RECT 1564.4400 263.0000 1566.0400 263.4800 ;
        RECT 1576.7800 241.2400 1579.7800 241.7200 ;
        RECT 1576.7800 246.6800 1579.7800 247.1600 ;
        RECT 1564.4400 241.2400 1566.0400 241.7200 ;
        RECT 1564.4400 246.6800 1566.0400 247.1600 ;
        RECT 1576.7800 252.1200 1579.7800 252.6000 ;
        RECT 1564.4400 252.1200 1566.0400 252.6000 ;
        RECT 1519.4400 268.4400 1521.0400 268.9200 ;
        RECT 1519.4400 273.8800 1521.0400 274.3600 ;
        RECT 1519.4400 279.3200 1521.0400 279.8000 ;
        RECT 1519.4400 257.5600 1521.0400 258.0400 ;
        RECT 1519.4400 263.0000 1521.0400 263.4800 ;
        RECT 1519.4400 241.2400 1521.0400 241.7200 ;
        RECT 1519.4400 246.6800 1521.0400 247.1600 ;
        RECT 1519.4400 252.1200 1521.0400 252.6000 ;
        RECT 1576.7800 224.9200 1579.7800 225.4000 ;
        RECT 1576.7800 230.3600 1579.7800 230.8400 ;
        RECT 1576.7800 235.8000 1579.7800 236.2800 ;
        RECT 1564.4400 224.9200 1566.0400 225.4000 ;
        RECT 1564.4400 230.3600 1566.0400 230.8400 ;
        RECT 1564.4400 235.8000 1566.0400 236.2800 ;
        RECT 1576.7800 214.0400 1579.7800 214.5200 ;
        RECT 1576.7800 219.4800 1579.7800 219.9600 ;
        RECT 1564.4400 214.0400 1566.0400 214.5200 ;
        RECT 1564.4400 219.4800 1566.0400 219.9600 ;
        RECT 1576.7800 197.7200 1579.7800 198.2000 ;
        RECT 1576.7800 203.1600 1579.7800 203.6400 ;
        RECT 1576.7800 208.6000 1579.7800 209.0800 ;
        RECT 1564.4400 197.7200 1566.0400 198.2000 ;
        RECT 1564.4400 203.1600 1566.0400 203.6400 ;
        RECT 1564.4400 208.6000 1566.0400 209.0800 ;
        RECT 1576.7800 186.8400 1579.7800 187.3200 ;
        RECT 1576.7800 192.2800 1579.7800 192.7600 ;
        RECT 1564.4400 186.8400 1566.0400 187.3200 ;
        RECT 1564.4400 192.2800 1566.0400 192.7600 ;
        RECT 1519.4400 224.9200 1521.0400 225.4000 ;
        RECT 1519.4400 230.3600 1521.0400 230.8400 ;
        RECT 1519.4400 235.8000 1521.0400 236.2800 ;
        RECT 1519.4400 214.0400 1521.0400 214.5200 ;
        RECT 1519.4400 219.4800 1521.0400 219.9600 ;
        RECT 1519.4400 197.7200 1521.0400 198.2000 ;
        RECT 1519.4400 203.1600 1521.0400 203.6400 ;
        RECT 1519.4400 208.6000 1521.0400 209.0800 ;
        RECT 1519.4400 186.8400 1521.0400 187.3200 ;
        RECT 1519.4400 192.2800 1521.0400 192.7600 ;
        RECT 1474.4400 268.4400 1476.0400 268.9200 ;
        RECT 1474.4400 273.8800 1476.0400 274.3600 ;
        RECT 1474.4400 279.3200 1476.0400 279.8000 ;
        RECT 1429.4400 268.4400 1431.0400 268.9200 ;
        RECT 1429.4400 273.8800 1431.0400 274.3600 ;
        RECT 1429.4400 279.3200 1431.0400 279.8000 ;
        RECT 1474.4400 257.5600 1476.0400 258.0400 ;
        RECT 1474.4400 263.0000 1476.0400 263.4800 ;
        RECT 1474.4400 241.2400 1476.0400 241.7200 ;
        RECT 1474.4400 246.6800 1476.0400 247.1600 ;
        RECT 1474.4400 252.1200 1476.0400 252.6000 ;
        RECT 1429.4400 257.5600 1431.0400 258.0400 ;
        RECT 1429.4400 263.0000 1431.0400 263.4800 ;
        RECT 1429.4400 241.2400 1431.0400 241.7200 ;
        RECT 1429.4400 246.6800 1431.0400 247.1600 ;
        RECT 1429.4400 252.1200 1431.0400 252.6000 ;
        RECT 1384.4400 268.4400 1386.0400 268.9200 ;
        RECT 1384.4400 273.8800 1386.0400 274.3600 ;
        RECT 1372.6800 273.8800 1375.6800 274.3600 ;
        RECT 1372.6800 268.4400 1375.6800 268.9200 ;
        RECT 1372.6800 279.3200 1375.6800 279.8000 ;
        RECT 1384.4400 279.3200 1386.0400 279.8000 ;
        RECT 1384.4400 257.5600 1386.0400 258.0400 ;
        RECT 1384.4400 263.0000 1386.0400 263.4800 ;
        RECT 1372.6800 263.0000 1375.6800 263.4800 ;
        RECT 1372.6800 257.5600 1375.6800 258.0400 ;
        RECT 1384.4400 241.2400 1386.0400 241.7200 ;
        RECT 1384.4400 246.6800 1386.0400 247.1600 ;
        RECT 1372.6800 246.6800 1375.6800 247.1600 ;
        RECT 1372.6800 241.2400 1375.6800 241.7200 ;
        RECT 1372.6800 252.1200 1375.6800 252.6000 ;
        RECT 1384.4400 252.1200 1386.0400 252.6000 ;
        RECT 1474.4400 224.9200 1476.0400 225.4000 ;
        RECT 1474.4400 230.3600 1476.0400 230.8400 ;
        RECT 1474.4400 235.8000 1476.0400 236.2800 ;
        RECT 1474.4400 214.0400 1476.0400 214.5200 ;
        RECT 1474.4400 219.4800 1476.0400 219.9600 ;
        RECT 1429.4400 224.9200 1431.0400 225.4000 ;
        RECT 1429.4400 230.3600 1431.0400 230.8400 ;
        RECT 1429.4400 235.8000 1431.0400 236.2800 ;
        RECT 1429.4400 214.0400 1431.0400 214.5200 ;
        RECT 1429.4400 219.4800 1431.0400 219.9600 ;
        RECT 1474.4400 197.7200 1476.0400 198.2000 ;
        RECT 1474.4400 203.1600 1476.0400 203.6400 ;
        RECT 1474.4400 208.6000 1476.0400 209.0800 ;
        RECT 1474.4400 186.8400 1476.0400 187.3200 ;
        RECT 1474.4400 192.2800 1476.0400 192.7600 ;
        RECT 1429.4400 197.7200 1431.0400 198.2000 ;
        RECT 1429.4400 203.1600 1431.0400 203.6400 ;
        RECT 1429.4400 208.6000 1431.0400 209.0800 ;
        RECT 1429.4400 186.8400 1431.0400 187.3200 ;
        RECT 1429.4400 192.2800 1431.0400 192.7600 ;
        RECT 1384.4400 224.9200 1386.0400 225.4000 ;
        RECT 1384.4400 230.3600 1386.0400 230.8400 ;
        RECT 1384.4400 235.8000 1386.0400 236.2800 ;
        RECT 1372.6800 224.9200 1375.6800 225.4000 ;
        RECT 1372.6800 230.3600 1375.6800 230.8400 ;
        RECT 1372.6800 235.8000 1375.6800 236.2800 ;
        RECT 1384.4400 214.0400 1386.0400 214.5200 ;
        RECT 1384.4400 219.4800 1386.0400 219.9600 ;
        RECT 1372.6800 214.0400 1375.6800 214.5200 ;
        RECT 1372.6800 219.4800 1375.6800 219.9600 ;
        RECT 1384.4400 197.7200 1386.0400 198.2000 ;
        RECT 1384.4400 203.1600 1386.0400 203.6400 ;
        RECT 1384.4400 208.6000 1386.0400 209.0800 ;
        RECT 1372.6800 197.7200 1375.6800 198.2000 ;
        RECT 1372.6800 203.1600 1375.6800 203.6400 ;
        RECT 1372.6800 208.6000 1375.6800 209.0800 ;
        RECT 1384.4400 186.8400 1386.0400 187.3200 ;
        RECT 1384.4400 192.2800 1386.0400 192.7600 ;
        RECT 1372.6800 186.8400 1375.6800 187.3200 ;
        RECT 1372.6800 192.2800 1375.6800 192.7600 ;
        RECT 1576.7800 170.5200 1579.7800 171.0000 ;
        RECT 1576.7800 175.9600 1579.7800 176.4400 ;
        RECT 1576.7800 181.4000 1579.7800 181.8800 ;
        RECT 1564.4400 170.5200 1566.0400 171.0000 ;
        RECT 1564.4400 175.9600 1566.0400 176.4400 ;
        RECT 1564.4400 181.4000 1566.0400 181.8800 ;
        RECT 1576.7800 159.6400 1579.7800 160.1200 ;
        RECT 1576.7800 165.0800 1579.7800 165.5600 ;
        RECT 1564.4400 159.6400 1566.0400 160.1200 ;
        RECT 1564.4400 165.0800 1566.0400 165.5600 ;
        RECT 1576.7800 143.3200 1579.7800 143.8000 ;
        RECT 1576.7800 148.7600 1579.7800 149.2400 ;
        RECT 1576.7800 154.2000 1579.7800 154.6800 ;
        RECT 1564.4400 143.3200 1566.0400 143.8000 ;
        RECT 1564.4400 148.7600 1566.0400 149.2400 ;
        RECT 1564.4400 154.2000 1566.0400 154.6800 ;
        RECT 1576.7800 132.4400 1579.7800 132.9200 ;
        RECT 1576.7800 137.8800 1579.7800 138.3600 ;
        RECT 1564.4400 132.4400 1566.0400 132.9200 ;
        RECT 1564.4400 137.8800 1566.0400 138.3600 ;
        RECT 1519.4400 170.5200 1521.0400 171.0000 ;
        RECT 1519.4400 175.9600 1521.0400 176.4400 ;
        RECT 1519.4400 181.4000 1521.0400 181.8800 ;
        RECT 1519.4400 159.6400 1521.0400 160.1200 ;
        RECT 1519.4400 165.0800 1521.0400 165.5600 ;
        RECT 1519.4400 143.3200 1521.0400 143.8000 ;
        RECT 1519.4400 148.7600 1521.0400 149.2400 ;
        RECT 1519.4400 154.2000 1521.0400 154.6800 ;
        RECT 1519.4400 132.4400 1521.0400 132.9200 ;
        RECT 1519.4400 137.8800 1521.0400 138.3600 ;
        RECT 1576.7800 116.1200 1579.7800 116.6000 ;
        RECT 1576.7800 121.5600 1579.7800 122.0400 ;
        RECT 1576.7800 127.0000 1579.7800 127.4800 ;
        RECT 1564.4400 116.1200 1566.0400 116.6000 ;
        RECT 1564.4400 121.5600 1566.0400 122.0400 ;
        RECT 1564.4400 127.0000 1566.0400 127.4800 ;
        RECT 1576.7800 105.2400 1579.7800 105.7200 ;
        RECT 1576.7800 110.6800 1579.7800 111.1600 ;
        RECT 1564.4400 105.2400 1566.0400 105.7200 ;
        RECT 1564.4400 110.6800 1566.0400 111.1600 ;
        RECT 1576.7800 88.9200 1579.7800 89.4000 ;
        RECT 1576.7800 94.3600 1579.7800 94.8400 ;
        RECT 1576.7800 99.8000 1579.7800 100.2800 ;
        RECT 1564.4400 88.9200 1566.0400 89.4000 ;
        RECT 1564.4400 94.3600 1566.0400 94.8400 ;
        RECT 1564.4400 99.8000 1566.0400 100.2800 ;
        RECT 1576.7800 83.4800 1579.7800 83.9600 ;
        RECT 1564.4400 83.4800 1566.0400 83.9600 ;
        RECT 1519.4400 116.1200 1521.0400 116.6000 ;
        RECT 1519.4400 121.5600 1521.0400 122.0400 ;
        RECT 1519.4400 127.0000 1521.0400 127.4800 ;
        RECT 1519.4400 105.2400 1521.0400 105.7200 ;
        RECT 1519.4400 110.6800 1521.0400 111.1600 ;
        RECT 1519.4400 88.9200 1521.0400 89.4000 ;
        RECT 1519.4400 94.3600 1521.0400 94.8400 ;
        RECT 1519.4400 99.8000 1521.0400 100.2800 ;
        RECT 1519.4400 83.4800 1521.0400 83.9600 ;
        RECT 1474.4400 170.5200 1476.0400 171.0000 ;
        RECT 1474.4400 175.9600 1476.0400 176.4400 ;
        RECT 1474.4400 181.4000 1476.0400 181.8800 ;
        RECT 1474.4400 159.6400 1476.0400 160.1200 ;
        RECT 1474.4400 165.0800 1476.0400 165.5600 ;
        RECT 1429.4400 170.5200 1431.0400 171.0000 ;
        RECT 1429.4400 175.9600 1431.0400 176.4400 ;
        RECT 1429.4400 181.4000 1431.0400 181.8800 ;
        RECT 1429.4400 159.6400 1431.0400 160.1200 ;
        RECT 1429.4400 165.0800 1431.0400 165.5600 ;
        RECT 1474.4400 143.3200 1476.0400 143.8000 ;
        RECT 1474.4400 148.7600 1476.0400 149.2400 ;
        RECT 1474.4400 154.2000 1476.0400 154.6800 ;
        RECT 1474.4400 132.4400 1476.0400 132.9200 ;
        RECT 1474.4400 137.8800 1476.0400 138.3600 ;
        RECT 1429.4400 143.3200 1431.0400 143.8000 ;
        RECT 1429.4400 148.7600 1431.0400 149.2400 ;
        RECT 1429.4400 154.2000 1431.0400 154.6800 ;
        RECT 1429.4400 132.4400 1431.0400 132.9200 ;
        RECT 1429.4400 137.8800 1431.0400 138.3600 ;
        RECT 1384.4400 170.5200 1386.0400 171.0000 ;
        RECT 1384.4400 175.9600 1386.0400 176.4400 ;
        RECT 1384.4400 181.4000 1386.0400 181.8800 ;
        RECT 1372.6800 170.5200 1375.6800 171.0000 ;
        RECT 1372.6800 175.9600 1375.6800 176.4400 ;
        RECT 1372.6800 181.4000 1375.6800 181.8800 ;
        RECT 1384.4400 159.6400 1386.0400 160.1200 ;
        RECT 1384.4400 165.0800 1386.0400 165.5600 ;
        RECT 1372.6800 159.6400 1375.6800 160.1200 ;
        RECT 1372.6800 165.0800 1375.6800 165.5600 ;
        RECT 1384.4400 143.3200 1386.0400 143.8000 ;
        RECT 1384.4400 148.7600 1386.0400 149.2400 ;
        RECT 1384.4400 154.2000 1386.0400 154.6800 ;
        RECT 1372.6800 143.3200 1375.6800 143.8000 ;
        RECT 1372.6800 148.7600 1375.6800 149.2400 ;
        RECT 1372.6800 154.2000 1375.6800 154.6800 ;
        RECT 1384.4400 132.4400 1386.0400 132.9200 ;
        RECT 1384.4400 137.8800 1386.0400 138.3600 ;
        RECT 1372.6800 132.4400 1375.6800 132.9200 ;
        RECT 1372.6800 137.8800 1375.6800 138.3600 ;
        RECT 1474.4400 116.1200 1476.0400 116.6000 ;
        RECT 1474.4400 121.5600 1476.0400 122.0400 ;
        RECT 1474.4400 127.0000 1476.0400 127.4800 ;
        RECT 1474.4400 105.2400 1476.0400 105.7200 ;
        RECT 1474.4400 110.6800 1476.0400 111.1600 ;
        RECT 1429.4400 116.1200 1431.0400 116.6000 ;
        RECT 1429.4400 121.5600 1431.0400 122.0400 ;
        RECT 1429.4400 127.0000 1431.0400 127.4800 ;
        RECT 1429.4400 105.2400 1431.0400 105.7200 ;
        RECT 1429.4400 110.6800 1431.0400 111.1600 ;
        RECT 1474.4400 88.9200 1476.0400 89.4000 ;
        RECT 1474.4400 94.3600 1476.0400 94.8400 ;
        RECT 1474.4400 99.8000 1476.0400 100.2800 ;
        RECT 1474.4400 83.4800 1476.0400 83.9600 ;
        RECT 1429.4400 88.9200 1431.0400 89.4000 ;
        RECT 1429.4400 94.3600 1431.0400 94.8400 ;
        RECT 1429.4400 99.8000 1431.0400 100.2800 ;
        RECT 1429.4400 83.4800 1431.0400 83.9600 ;
        RECT 1384.4400 116.1200 1386.0400 116.6000 ;
        RECT 1384.4400 121.5600 1386.0400 122.0400 ;
        RECT 1384.4400 127.0000 1386.0400 127.4800 ;
        RECT 1372.6800 116.1200 1375.6800 116.6000 ;
        RECT 1372.6800 121.5600 1375.6800 122.0400 ;
        RECT 1372.6800 127.0000 1375.6800 127.4800 ;
        RECT 1384.4400 105.2400 1386.0400 105.7200 ;
        RECT 1384.4400 110.6800 1386.0400 111.1600 ;
        RECT 1372.6800 105.2400 1375.6800 105.7200 ;
        RECT 1372.6800 110.6800 1375.6800 111.1600 ;
        RECT 1384.4400 88.9200 1386.0400 89.4000 ;
        RECT 1384.4400 94.3600 1386.0400 94.8400 ;
        RECT 1384.4400 99.8000 1386.0400 100.2800 ;
        RECT 1372.6800 88.9200 1375.6800 89.4000 ;
        RECT 1372.6800 94.3600 1375.6800 94.8400 ;
        RECT 1372.6800 99.8000 1375.6800 100.2800 ;
        RECT 1372.6800 83.4800 1375.6800 83.9600 ;
        RECT 1384.4400 83.4800 1386.0400 83.9600 ;
        RECT 1372.6800 288.3900 1579.7800 291.3900 ;
        RECT 1372.6800 75.2900 1579.7800 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1373.6800 34.6700 1375.6800 61.6000 ;
        RECT 1576.7800 34.6700 1578.7800 61.6000 ;
      LAYER met3 ;
        RECT 1576.7800 51.3800 1578.7800 51.8600 ;
        RECT 1373.6800 51.3800 1375.6800 51.8600 ;
        RECT 1576.7800 45.9400 1578.7800 46.4200 ;
        RECT 1576.7800 40.5000 1578.7800 40.9800 ;
        RECT 1373.6800 45.9400 1375.6800 46.4200 ;
        RECT 1373.6800 40.5000 1375.6800 40.9800 ;
        RECT 1373.6800 59.6000 1578.7800 61.6000 ;
        RECT 1373.6800 34.6700 1578.7800 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 2601.3300 1566.0400 2817.4300 ;
        RECT 1519.4400 2601.3300 1521.0400 2817.4300 ;
        RECT 1474.4400 2601.3300 1476.0400 2817.4300 ;
        RECT 1429.4400 2601.3300 1431.0400 2817.4300 ;
        RECT 1384.4400 2601.3300 1386.0400 2817.4300 ;
        RECT 1576.7800 2601.3300 1579.7800 2817.4300 ;
        RECT 1372.6800 2601.3300 1375.6800 2817.4300 ;
      LAYER met3 ;
        RECT 1576.7800 2794.4800 1579.7800 2794.9600 ;
        RECT 1576.7800 2799.9200 1579.7800 2800.4000 ;
        RECT 1564.4400 2794.4800 1566.0400 2794.9600 ;
        RECT 1564.4400 2799.9200 1566.0400 2800.4000 ;
        RECT 1576.7800 2805.3600 1579.7800 2805.8400 ;
        RECT 1564.4400 2805.3600 1566.0400 2805.8400 ;
        RECT 1576.7800 2783.6000 1579.7800 2784.0800 ;
        RECT 1576.7800 2789.0400 1579.7800 2789.5200 ;
        RECT 1564.4400 2783.6000 1566.0400 2784.0800 ;
        RECT 1564.4400 2789.0400 1566.0400 2789.5200 ;
        RECT 1576.7800 2767.2800 1579.7800 2767.7600 ;
        RECT 1576.7800 2772.7200 1579.7800 2773.2000 ;
        RECT 1564.4400 2767.2800 1566.0400 2767.7600 ;
        RECT 1564.4400 2772.7200 1566.0400 2773.2000 ;
        RECT 1576.7800 2778.1600 1579.7800 2778.6400 ;
        RECT 1564.4400 2778.1600 1566.0400 2778.6400 ;
        RECT 1519.4400 2794.4800 1521.0400 2794.9600 ;
        RECT 1519.4400 2799.9200 1521.0400 2800.4000 ;
        RECT 1519.4400 2805.3600 1521.0400 2805.8400 ;
        RECT 1519.4400 2783.6000 1521.0400 2784.0800 ;
        RECT 1519.4400 2789.0400 1521.0400 2789.5200 ;
        RECT 1519.4400 2767.2800 1521.0400 2767.7600 ;
        RECT 1519.4400 2772.7200 1521.0400 2773.2000 ;
        RECT 1519.4400 2778.1600 1521.0400 2778.6400 ;
        RECT 1576.7800 2750.9600 1579.7800 2751.4400 ;
        RECT 1576.7800 2756.4000 1579.7800 2756.8800 ;
        RECT 1576.7800 2761.8400 1579.7800 2762.3200 ;
        RECT 1564.4400 2750.9600 1566.0400 2751.4400 ;
        RECT 1564.4400 2756.4000 1566.0400 2756.8800 ;
        RECT 1564.4400 2761.8400 1566.0400 2762.3200 ;
        RECT 1576.7800 2740.0800 1579.7800 2740.5600 ;
        RECT 1576.7800 2745.5200 1579.7800 2746.0000 ;
        RECT 1564.4400 2740.0800 1566.0400 2740.5600 ;
        RECT 1564.4400 2745.5200 1566.0400 2746.0000 ;
        RECT 1576.7800 2723.7600 1579.7800 2724.2400 ;
        RECT 1576.7800 2729.2000 1579.7800 2729.6800 ;
        RECT 1576.7800 2734.6400 1579.7800 2735.1200 ;
        RECT 1564.4400 2723.7600 1566.0400 2724.2400 ;
        RECT 1564.4400 2729.2000 1566.0400 2729.6800 ;
        RECT 1564.4400 2734.6400 1566.0400 2735.1200 ;
        RECT 1576.7800 2712.8800 1579.7800 2713.3600 ;
        RECT 1576.7800 2718.3200 1579.7800 2718.8000 ;
        RECT 1564.4400 2712.8800 1566.0400 2713.3600 ;
        RECT 1564.4400 2718.3200 1566.0400 2718.8000 ;
        RECT 1519.4400 2750.9600 1521.0400 2751.4400 ;
        RECT 1519.4400 2756.4000 1521.0400 2756.8800 ;
        RECT 1519.4400 2761.8400 1521.0400 2762.3200 ;
        RECT 1519.4400 2740.0800 1521.0400 2740.5600 ;
        RECT 1519.4400 2745.5200 1521.0400 2746.0000 ;
        RECT 1519.4400 2723.7600 1521.0400 2724.2400 ;
        RECT 1519.4400 2729.2000 1521.0400 2729.6800 ;
        RECT 1519.4400 2734.6400 1521.0400 2735.1200 ;
        RECT 1519.4400 2712.8800 1521.0400 2713.3600 ;
        RECT 1519.4400 2718.3200 1521.0400 2718.8000 ;
        RECT 1474.4400 2794.4800 1476.0400 2794.9600 ;
        RECT 1474.4400 2799.9200 1476.0400 2800.4000 ;
        RECT 1474.4400 2805.3600 1476.0400 2805.8400 ;
        RECT 1429.4400 2794.4800 1431.0400 2794.9600 ;
        RECT 1429.4400 2799.9200 1431.0400 2800.4000 ;
        RECT 1429.4400 2805.3600 1431.0400 2805.8400 ;
        RECT 1474.4400 2783.6000 1476.0400 2784.0800 ;
        RECT 1474.4400 2789.0400 1476.0400 2789.5200 ;
        RECT 1474.4400 2767.2800 1476.0400 2767.7600 ;
        RECT 1474.4400 2772.7200 1476.0400 2773.2000 ;
        RECT 1474.4400 2778.1600 1476.0400 2778.6400 ;
        RECT 1429.4400 2783.6000 1431.0400 2784.0800 ;
        RECT 1429.4400 2789.0400 1431.0400 2789.5200 ;
        RECT 1429.4400 2767.2800 1431.0400 2767.7600 ;
        RECT 1429.4400 2772.7200 1431.0400 2773.2000 ;
        RECT 1429.4400 2778.1600 1431.0400 2778.6400 ;
        RECT 1384.4400 2794.4800 1386.0400 2794.9600 ;
        RECT 1384.4400 2799.9200 1386.0400 2800.4000 ;
        RECT 1372.6800 2799.9200 1375.6800 2800.4000 ;
        RECT 1372.6800 2794.4800 1375.6800 2794.9600 ;
        RECT 1372.6800 2805.3600 1375.6800 2805.8400 ;
        RECT 1384.4400 2805.3600 1386.0400 2805.8400 ;
        RECT 1384.4400 2783.6000 1386.0400 2784.0800 ;
        RECT 1384.4400 2789.0400 1386.0400 2789.5200 ;
        RECT 1372.6800 2789.0400 1375.6800 2789.5200 ;
        RECT 1372.6800 2783.6000 1375.6800 2784.0800 ;
        RECT 1384.4400 2767.2800 1386.0400 2767.7600 ;
        RECT 1384.4400 2772.7200 1386.0400 2773.2000 ;
        RECT 1372.6800 2772.7200 1375.6800 2773.2000 ;
        RECT 1372.6800 2767.2800 1375.6800 2767.7600 ;
        RECT 1372.6800 2778.1600 1375.6800 2778.6400 ;
        RECT 1384.4400 2778.1600 1386.0400 2778.6400 ;
        RECT 1474.4400 2750.9600 1476.0400 2751.4400 ;
        RECT 1474.4400 2756.4000 1476.0400 2756.8800 ;
        RECT 1474.4400 2761.8400 1476.0400 2762.3200 ;
        RECT 1474.4400 2740.0800 1476.0400 2740.5600 ;
        RECT 1474.4400 2745.5200 1476.0400 2746.0000 ;
        RECT 1429.4400 2750.9600 1431.0400 2751.4400 ;
        RECT 1429.4400 2756.4000 1431.0400 2756.8800 ;
        RECT 1429.4400 2761.8400 1431.0400 2762.3200 ;
        RECT 1429.4400 2740.0800 1431.0400 2740.5600 ;
        RECT 1429.4400 2745.5200 1431.0400 2746.0000 ;
        RECT 1474.4400 2723.7600 1476.0400 2724.2400 ;
        RECT 1474.4400 2729.2000 1476.0400 2729.6800 ;
        RECT 1474.4400 2734.6400 1476.0400 2735.1200 ;
        RECT 1474.4400 2712.8800 1476.0400 2713.3600 ;
        RECT 1474.4400 2718.3200 1476.0400 2718.8000 ;
        RECT 1429.4400 2723.7600 1431.0400 2724.2400 ;
        RECT 1429.4400 2729.2000 1431.0400 2729.6800 ;
        RECT 1429.4400 2734.6400 1431.0400 2735.1200 ;
        RECT 1429.4400 2712.8800 1431.0400 2713.3600 ;
        RECT 1429.4400 2718.3200 1431.0400 2718.8000 ;
        RECT 1384.4400 2750.9600 1386.0400 2751.4400 ;
        RECT 1384.4400 2756.4000 1386.0400 2756.8800 ;
        RECT 1384.4400 2761.8400 1386.0400 2762.3200 ;
        RECT 1372.6800 2750.9600 1375.6800 2751.4400 ;
        RECT 1372.6800 2756.4000 1375.6800 2756.8800 ;
        RECT 1372.6800 2761.8400 1375.6800 2762.3200 ;
        RECT 1384.4400 2740.0800 1386.0400 2740.5600 ;
        RECT 1384.4400 2745.5200 1386.0400 2746.0000 ;
        RECT 1372.6800 2740.0800 1375.6800 2740.5600 ;
        RECT 1372.6800 2745.5200 1375.6800 2746.0000 ;
        RECT 1384.4400 2723.7600 1386.0400 2724.2400 ;
        RECT 1384.4400 2729.2000 1386.0400 2729.6800 ;
        RECT 1384.4400 2734.6400 1386.0400 2735.1200 ;
        RECT 1372.6800 2723.7600 1375.6800 2724.2400 ;
        RECT 1372.6800 2729.2000 1375.6800 2729.6800 ;
        RECT 1372.6800 2734.6400 1375.6800 2735.1200 ;
        RECT 1384.4400 2712.8800 1386.0400 2713.3600 ;
        RECT 1384.4400 2718.3200 1386.0400 2718.8000 ;
        RECT 1372.6800 2712.8800 1375.6800 2713.3600 ;
        RECT 1372.6800 2718.3200 1375.6800 2718.8000 ;
        RECT 1576.7800 2696.5600 1579.7800 2697.0400 ;
        RECT 1576.7800 2702.0000 1579.7800 2702.4800 ;
        RECT 1576.7800 2707.4400 1579.7800 2707.9200 ;
        RECT 1564.4400 2696.5600 1566.0400 2697.0400 ;
        RECT 1564.4400 2702.0000 1566.0400 2702.4800 ;
        RECT 1564.4400 2707.4400 1566.0400 2707.9200 ;
        RECT 1576.7800 2685.6800 1579.7800 2686.1600 ;
        RECT 1576.7800 2691.1200 1579.7800 2691.6000 ;
        RECT 1564.4400 2685.6800 1566.0400 2686.1600 ;
        RECT 1564.4400 2691.1200 1566.0400 2691.6000 ;
        RECT 1576.7800 2669.3600 1579.7800 2669.8400 ;
        RECT 1576.7800 2674.8000 1579.7800 2675.2800 ;
        RECT 1576.7800 2680.2400 1579.7800 2680.7200 ;
        RECT 1564.4400 2669.3600 1566.0400 2669.8400 ;
        RECT 1564.4400 2674.8000 1566.0400 2675.2800 ;
        RECT 1564.4400 2680.2400 1566.0400 2680.7200 ;
        RECT 1576.7800 2658.4800 1579.7800 2658.9600 ;
        RECT 1576.7800 2663.9200 1579.7800 2664.4000 ;
        RECT 1564.4400 2658.4800 1566.0400 2658.9600 ;
        RECT 1564.4400 2663.9200 1566.0400 2664.4000 ;
        RECT 1519.4400 2696.5600 1521.0400 2697.0400 ;
        RECT 1519.4400 2702.0000 1521.0400 2702.4800 ;
        RECT 1519.4400 2707.4400 1521.0400 2707.9200 ;
        RECT 1519.4400 2685.6800 1521.0400 2686.1600 ;
        RECT 1519.4400 2691.1200 1521.0400 2691.6000 ;
        RECT 1519.4400 2669.3600 1521.0400 2669.8400 ;
        RECT 1519.4400 2674.8000 1521.0400 2675.2800 ;
        RECT 1519.4400 2680.2400 1521.0400 2680.7200 ;
        RECT 1519.4400 2658.4800 1521.0400 2658.9600 ;
        RECT 1519.4400 2663.9200 1521.0400 2664.4000 ;
        RECT 1576.7800 2642.1600 1579.7800 2642.6400 ;
        RECT 1576.7800 2647.6000 1579.7800 2648.0800 ;
        RECT 1576.7800 2653.0400 1579.7800 2653.5200 ;
        RECT 1564.4400 2642.1600 1566.0400 2642.6400 ;
        RECT 1564.4400 2647.6000 1566.0400 2648.0800 ;
        RECT 1564.4400 2653.0400 1566.0400 2653.5200 ;
        RECT 1576.7800 2631.2800 1579.7800 2631.7600 ;
        RECT 1576.7800 2636.7200 1579.7800 2637.2000 ;
        RECT 1564.4400 2631.2800 1566.0400 2631.7600 ;
        RECT 1564.4400 2636.7200 1566.0400 2637.2000 ;
        RECT 1576.7800 2614.9600 1579.7800 2615.4400 ;
        RECT 1576.7800 2620.4000 1579.7800 2620.8800 ;
        RECT 1576.7800 2625.8400 1579.7800 2626.3200 ;
        RECT 1564.4400 2614.9600 1566.0400 2615.4400 ;
        RECT 1564.4400 2620.4000 1566.0400 2620.8800 ;
        RECT 1564.4400 2625.8400 1566.0400 2626.3200 ;
        RECT 1576.7800 2609.5200 1579.7800 2610.0000 ;
        RECT 1564.4400 2609.5200 1566.0400 2610.0000 ;
        RECT 1519.4400 2642.1600 1521.0400 2642.6400 ;
        RECT 1519.4400 2647.6000 1521.0400 2648.0800 ;
        RECT 1519.4400 2653.0400 1521.0400 2653.5200 ;
        RECT 1519.4400 2631.2800 1521.0400 2631.7600 ;
        RECT 1519.4400 2636.7200 1521.0400 2637.2000 ;
        RECT 1519.4400 2614.9600 1521.0400 2615.4400 ;
        RECT 1519.4400 2620.4000 1521.0400 2620.8800 ;
        RECT 1519.4400 2625.8400 1521.0400 2626.3200 ;
        RECT 1519.4400 2609.5200 1521.0400 2610.0000 ;
        RECT 1474.4400 2696.5600 1476.0400 2697.0400 ;
        RECT 1474.4400 2702.0000 1476.0400 2702.4800 ;
        RECT 1474.4400 2707.4400 1476.0400 2707.9200 ;
        RECT 1474.4400 2685.6800 1476.0400 2686.1600 ;
        RECT 1474.4400 2691.1200 1476.0400 2691.6000 ;
        RECT 1429.4400 2696.5600 1431.0400 2697.0400 ;
        RECT 1429.4400 2702.0000 1431.0400 2702.4800 ;
        RECT 1429.4400 2707.4400 1431.0400 2707.9200 ;
        RECT 1429.4400 2685.6800 1431.0400 2686.1600 ;
        RECT 1429.4400 2691.1200 1431.0400 2691.6000 ;
        RECT 1474.4400 2669.3600 1476.0400 2669.8400 ;
        RECT 1474.4400 2674.8000 1476.0400 2675.2800 ;
        RECT 1474.4400 2680.2400 1476.0400 2680.7200 ;
        RECT 1474.4400 2658.4800 1476.0400 2658.9600 ;
        RECT 1474.4400 2663.9200 1476.0400 2664.4000 ;
        RECT 1429.4400 2669.3600 1431.0400 2669.8400 ;
        RECT 1429.4400 2674.8000 1431.0400 2675.2800 ;
        RECT 1429.4400 2680.2400 1431.0400 2680.7200 ;
        RECT 1429.4400 2658.4800 1431.0400 2658.9600 ;
        RECT 1429.4400 2663.9200 1431.0400 2664.4000 ;
        RECT 1384.4400 2696.5600 1386.0400 2697.0400 ;
        RECT 1384.4400 2702.0000 1386.0400 2702.4800 ;
        RECT 1384.4400 2707.4400 1386.0400 2707.9200 ;
        RECT 1372.6800 2696.5600 1375.6800 2697.0400 ;
        RECT 1372.6800 2702.0000 1375.6800 2702.4800 ;
        RECT 1372.6800 2707.4400 1375.6800 2707.9200 ;
        RECT 1384.4400 2685.6800 1386.0400 2686.1600 ;
        RECT 1384.4400 2691.1200 1386.0400 2691.6000 ;
        RECT 1372.6800 2685.6800 1375.6800 2686.1600 ;
        RECT 1372.6800 2691.1200 1375.6800 2691.6000 ;
        RECT 1384.4400 2669.3600 1386.0400 2669.8400 ;
        RECT 1384.4400 2674.8000 1386.0400 2675.2800 ;
        RECT 1384.4400 2680.2400 1386.0400 2680.7200 ;
        RECT 1372.6800 2669.3600 1375.6800 2669.8400 ;
        RECT 1372.6800 2674.8000 1375.6800 2675.2800 ;
        RECT 1372.6800 2680.2400 1375.6800 2680.7200 ;
        RECT 1384.4400 2658.4800 1386.0400 2658.9600 ;
        RECT 1384.4400 2663.9200 1386.0400 2664.4000 ;
        RECT 1372.6800 2658.4800 1375.6800 2658.9600 ;
        RECT 1372.6800 2663.9200 1375.6800 2664.4000 ;
        RECT 1474.4400 2642.1600 1476.0400 2642.6400 ;
        RECT 1474.4400 2647.6000 1476.0400 2648.0800 ;
        RECT 1474.4400 2653.0400 1476.0400 2653.5200 ;
        RECT 1474.4400 2631.2800 1476.0400 2631.7600 ;
        RECT 1474.4400 2636.7200 1476.0400 2637.2000 ;
        RECT 1429.4400 2642.1600 1431.0400 2642.6400 ;
        RECT 1429.4400 2647.6000 1431.0400 2648.0800 ;
        RECT 1429.4400 2653.0400 1431.0400 2653.5200 ;
        RECT 1429.4400 2631.2800 1431.0400 2631.7600 ;
        RECT 1429.4400 2636.7200 1431.0400 2637.2000 ;
        RECT 1474.4400 2614.9600 1476.0400 2615.4400 ;
        RECT 1474.4400 2620.4000 1476.0400 2620.8800 ;
        RECT 1474.4400 2625.8400 1476.0400 2626.3200 ;
        RECT 1474.4400 2609.5200 1476.0400 2610.0000 ;
        RECT 1429.4400 2614.9600 1431.0400 2615.4400 ;
        RECT 1429.4400 2620.4000 1431.0400 2620.8800 ;
        RECT 1429.4400 2625.8400 1431.0400 2626.3200 ;
        RECT 1429.4400 2609.5200 1431.0400 2610.0000 ;
        RECT 1384.4400 2642.1600 1386.0400 2642.6400 ;
        RECT 1384.4400 2647.6000 1386.0400 2648.0800 ;
        RECT 1384.4400 2653.0400 1386.0400 2653.5200 ;
        RECT 1372.6800 2642.1600 1375.6800 2642.6400 ;
        RECT 1372.6800 2647.6000 1375.6800 2648.0800 ;
        RECT 1372.6800 2653.0400 1375.6800 2653.5200 ;
        RECT 1384.4400 2631.2800 1386.0400 2631.7600 ;
        RECT 1384.4400 2636.7200 1386.0400 2637.2000 ;
        RECT 1372.6800 2631.2800 1375.6800 2631.7600 ;
        RECT 1372.6800 2636.7200 1375.6800 2637.2000 ;
        RECT 1384.4400 2614.9600 1386.0400 2615.4400 ;
        RECT 1384.4400 2620.4000 1386.0400 2620.8800 ;
        RECT 1384.4400 2625.8400 1386.0400 2626.3200 ;
        RECT 1372.6800 2614.9600 1375.6800 2615.4400 ;
        RECT 1372.6800 2620.4000 1375.6800 2620.8800 ;
        RECT 1372.6800 2625.8400 1375.6800 2626.3200 ;
        RECT 1372.6800 2609.5200 1375.6800 2610.0000 ;
        RECT 1384.4400 2609.5200 1386.0400 2610.0000 ;
        RECT 1372.6800 2814.4300 1579.7800 2817.4300 ;
        RECT 1372.6800 2601.3300 1579.7800 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 2371.6900 1566.0400 2587.7900 ;
        RECT 1519.4400 2371.6900 1521.0400 2587.7900 ;
        RECT 1474.4400 2371.6900 1476.0400 2587.7900 ;
        RECT 1429.4400 2371.6900 1431.0400 2587.7900 ;
        RECT 1384.4400 2371.6900 1386.0400 2587.7900 ;
        RECT 1576.7800 2371.6900 1579.7800 2587.7900 ;
        RECT 1372.6800 2371.6900 1375.6800 2587.7900 ;
      LAYER met3 ;
        RECT 1576.7800 2564.8400 1579.7800 2565.3200 ;
        RECT 1576.7800 2570.2800 1579.7800 2570.7600 ;
        RECT 1564.4400 2564.8400 1566.0400 2565.3200 ;
        RECT 1564.4400 2570.2800 1566.0400 2570.7600 ;
        RECT 1576.7800 2575.7200 1579.7800 2576.2000 ;
        RECT 1564.4400 2575.7200 1566.0400 2576.2000 ;
        RECT 1576.7800 2553.9600 1579.7800 2554.4400 ;
        RECT 1576.7800 2559.4000 1579.7800 2559.8800 ;
        RECT 1564.4400 2553.9600 1566.0400 2554.4400 ;
        RECT 1564.4400 2559.4000 1566.0400 2559.8800 ;
        RECT 1576.7800 2537.6400 1579.7800 2538.1200 ;
        RECT 1576.7800 2543.0800 1579.7800 2543.5600 ;
        RECT 1564.4400 2537.6400 1566.0400 2538.1200 ;
        RECT 1564.4400 2543.0800 1566.0400 2543.5600 ;
        RECT 1576.7800 2548.5200 1579.7800 2549.0000 ;
        RECT 1564.4400 2548.5200 1566.0400 2549.0000 ;
        RECT 1519.4400 2564.8400 1521.0400 2565.3200 ;
        RECT 1519.4400 2570.2800 1521.0400 2570.7600 ;
        RECT 1519.4400 2575.7200 1521.0400 2576.2000 ;
        RECT 1519.4400 2553.9600 1521.0400 2554.4400 ;
        RECT 1519.4400 2559.4000 1521.0400 2559.8800 ;
        RECT 1519.4400 2537.6400 1521.0400 2538.1200 ;
        RECT 1519.4400 2543.0800 1521.0400 2543.5600 ;
        RECT 1519.4400 2548.5200 1521.0400 2549.0000 ;
        RECT 1576.7800 2521.3200 1579.7800 2521.8000 ;
        RECT 1576.7800 2526.7600 1579.7800 2527.2400 ;
        RECT 1576.7800 2532.2000 1579.7800 2532.6800 ;
        RECT 1564.4400 2521.3200 1566.0400 2521.8000 ;
        RECT 1564.4400 2526.7600 1566.0400 2527.2400 ;
        RECT 1564.4400 2532.2000 1566.0400 2532.6800 ;
        RECT 1576.7800 2510.4400 1579.7800 2510.9200 ;
        RECT 1576.7800 2515.8800 1579.7800 2516.3600 ;
        RECT 1564.4400 2510.4400 1566.0400 2510.9200 ;
        RECT 1564.4400 2515.8800 1566.0400 2516.3600 ;
        RECT 1576.7800 2494.1200 1579.7800 2494.6000 ;
        RECT 1576.7800 2499.5600 1579.7800 2500.0400 ;
        RECT 1576.7800 2505.0000 1579.7800 2505.4800 ;
        RECT 1564.4400 2494.1200 1566.0400 2494.6000 ;
        RECT 1564.4400 2499.5600 1566.0400 2500.0400 ;
        RECT 1564.4400 2505.0000 1566.0400 2505.4800 ;
        RECT 1576.7800 2483.2400 1579.7800 2483.7200 ;
        RECT 1576.7800 2488.6800 1579.7800 2489.1600 ;
        RECT 1564.4400 2483.2400 1566.0400 2483.7200 ;
        RECT 1564.4400 2488.6800 1566.0400 2489.1600 ;
        RECT 1519.4400 2521.3200 1521.0400 2521.8000 ;
        RECT 1519.4400 2526.7600 1521.0400 2527.2400 ;
        RECT 1519.4400 2532.2000 1521.0400 2532.6800 ;
        RECT 1519.4400 2510.4400 1521.0400 2510.9200 ;
        RECT 1519.4400 2515.8800 1521.0400 2516.3600 ;
        RECT 1519.4400 2494.1200 1521.0400 2494.6000 ;
        RECT 1519.4400 2499.5600 1521.0400 2500.0400 ;
        RECT 1519.4400 2505.0000 1521.0400 2505.4800 ;
        RECT 1519.4400 2483.2400 1521.0400 2483.7200 ;
        RECT 1519.4400 2488.6800 1521.0400 2489.1600 ;
        RECT 1474.4400 2564.8400 1476.0400 2565.3200 ;
        RECT 1474.4400 2570.2800 1476.0400 2570.7600 ;
        RECT 1474.4400 2575.7200 1476.0400 2576.2000 ;
        RECT 1429.4400 2564.8400 1431.0400 2565.3200 ;
        RECT 1429.4400 2570.2800 1431.0400 2570.7600 ;
        RECT 1429.4400 2575.7200 1431.0400 2576.2000 ;
        RECT 1474.4400 2553.9600 1476.0400 2554.4400 ;
        RECT 1474.4400 2559.4000 1476.0400 2559.8800 ;
        RECT 1474.4400 2537.6400 1476.0400 2538.1200 ;
        RECT 1474.4400 2543.0800 1476.0400 2543.5600 ;
        RECT 1474.4400 2548.5200 1476.0400 2549.0000 ;
        RECT 1429.4400 2553.9600 1431.0400 2554.4400 ;
        RECT 1429.4400 2559.4000 1431.0400 2559.8800 ;
        RECT 1429.4400 2537.6400 1431.0400 2538.1200 ;
        RECT 1429.4400 2543.0800 1431.0400 2543.5600 ;
        RECT 1429.4400 2548.5200 1431.0400 2549.0000 ;
        RECT 1384.4400 2564.8400 1386.0400 2565.3200 ;
        RECT 1384.4400 2570.2800 1386.0400 2570.7600 ;
        RECT 1372.6800 2570.2800 1375.6800 2570.7600 ;
        RECT 1372.6800 2564.8400 1375.6800 2565.3200 ;
        RECT 1372.6800 2575.7200 1375.6800 2576.2000 ;
        RECT 1384.4400 2575.7200 1386.0400 2576.2000 ;
        RECT 1384.4400 2553.9600 1386.0400 2554.4400 ;
        RECT 1384.4400 2559.4000 1386.0400 2559.8800 ;
        RECT 1372.6800 2559.4000 1375.6800 2559.8800 ;
        RECT 1372.6800 2553.9600 1375.6800 2554.4400 ;
        RECT 1384.4400 2537.6400 1386.0400 2538.1200 ;
        RECT 1384.4400 2543.0800 1386.0400 2543.5600 ;
        RECT 1372.6800 2543.0800 1375.6800 2543.5600 ;
        RECT 1372.6800 2537.6400 1375.6800 2538.1200 ;
        RECT 1372.6800 2548.5200 1375.6800 2549.0000 ;
        RECT 1384.4400 2548.5200 1386.0400 2549.0000 ;
        RECT 1474.4400 2521.3200 1476.0400 2521.8000 ;
        RECT 1474.4400 2526.7600 1476.0400 2527.2400 ;
        RECT 1474.4400 2532.2000 1476.0400 2532.6800 ;
        RECT 1474.4400 2510.4400 1476.0400 2510.9200 ;
        RECT 1474.4400 2515.8800 1476.0400 2516.3600 ;
        RECT 1429.4400 2521.3200 1431.0400 2521.8000 ;
        RECT 1429.4400 2526.7600 1431.0400 2527.2400 ;
        RECT 1429.4400 2532.2000 1431.0400 2532.6800 ;
        RECT 1429.4400 2510.4400 1431.0400 2510.9200 ;
        RECT 1429.4400 2515.8800 1431.0400 2516.3600 ;
        RECT 1474.4400 2494.1200 1476.0400 2494.6000 ;
        RECT 1474.4400 2499.5600 1476.0400 2500.0400 ;
        RECT 1474.4400 2505.0000 1476.0400 2505.4800 ;
        RECT 1474.4400 2483.2400 1476.0400 2483.7200 ;
        RECT 1474.4400 2488.6800 1476.0400 2489.1600 ;
        RECT 1429.4400 2494.1200 1431.0400 2494.6000 ;
        RECT 1429.4400 2499.5600 1431.0400 2500.0400 ;
        RECT 1429.4400 2505.0000 1431.0400 2505.4800 ;
        RECT 1429.4400 2483.2400 1431.0400 2483.7200 ;
        RECT 1429.4400 2488.6800 1431.0400 2489.1600 ;
        RECT 1384.4400 2521.3200 1386.0400 2521.8000 ;
        RECT 1384.4400 2526.7600 1386.0400 2527.2400 ;
        RECT 1384.4400 2532.2000 1386.0400 2532.6800 ;
        RECT 1372.6800 2521.3200 1375.6800 2521.8000 ;
        RECT 1372.6800 2526.7600 1375.6800 2527.2400 ;
        RECT 1372.6800 2532.2000 1375.6800 2532.6800 ;
        RECT 1384.4400 2510.4400 1386.0400 2510.9200 ;
        RECT 1384.4400 2515.8800 1386.0400 2516.3600 ;
        RECT 1372.6800 2510.4400 1375.6800 2510.9200 ;
        RECT 1372.6800 2515.8800 1375.6800 2516.3600 ;
        RECT 1384.4400 2494.1200 1386.0400 2494.6000 ;
        RECT 1384.4400 2499.5600 1386.0400 2500.0400 ;
        RECT 1384.4400 2505.0000 1386.0400 2505.4800 ;
        RECT 1372.6800 2494.1200 1375.6800 2494.6000 ;
        RECT 1372.6800 2499.5600 1375.6800 2500.0400 ;
        RECT 1372.6800 2505.0000 1375.6800 2505.4800 ;
        RECT 1384.4400 2483.2400 1386.0400 2483.7200 ;
        RECT 1384.4400 2488.6800 1386.0400 2489.1600 ;
        RECT 1372.6800 2483.2400 1375.6800 2483.7200 ;
        RECT 1372.6800 2488.6800 1375.6800 2489.1600 ;
        RECT 1576.7800 2466.9200 1579.7800 2467.4000 ;
        RECT 1576.7800 2472.3600 1579.7800 2472.8400 ;
        RECT 1576.7800 2477.8000 1579.7800 2478.2800 ;
        RECT 1564.4400 2466.9200 1566.0400 2467.4000 ;
        RECT 1564.4400 2472.3600 1566.0400 2472.8400 ;
        RECT 1564.4400 2477.8000 1566.0400 2478.2800 ;
        RECT 1576.7800 2456.0400 1579.7800 2456.5200 ;
        RECT 1576.7800 2461.4800 1579.7800 2461.9600 ;
        RECT 1564.4400 2456.0400 1566.0400 2456.5200 ;
        RECT 1564.4400 2461.4800 1566.0400 2461.9600 ;
        RECT 1576.7800 2439.7200 1579.7800 2440.2000 ;
        RECT 1576.7800 2445.1600 1579.7800 2445.6400 ;
        RECT 1576.7800 2450.6000 1579.7800 2451.0800 ;
        RECT 1564.4400 2439.7200 1566.0400 2440.2000 ;
        RECT 1564.4400 2445.1600 1566.0400 2445.6400 ;
        RECT 1564.4400 2450.6000 1566.0400 2451.0800 ;
        RECT 1576.7800 2428.8400 1579.7800 2429.3200 ;
        RECT 1576.7800 2434.2800 1579.7800 2434.7600 ;
        RECT 1564.4400 2428.8400 1566.0400 2429.3200 ;
        RECT 1564.4400 2434.2800 1566.0400 2434.7600 ;
        RECT 1519.4400 2466.9200 1521.0400 2467.4000 ;
        RECT 1519.4400 2472.3600 1521.0400 2472.8400 ;
        RECT 1519.4400 2477.8000 1521.0400 2478.2800 ;
        RECT 1519.4400 2456.0400 1521.0400 2456.5200 ;
        RECT 1519.4400 2461.4800 1521.0400 2461.9600 ;
        RECT 1519.4400 2439.7200 1521.0400 2440.2000 ;
        RECT 1519.4400 2445.1600 1521.0400 2445.6400 ;
        RECT 1519.4400 2450.6000 1521.0400 2451.0800 ;
        RECT 1519.4400 2428.8400 1521.0400 2429.3200 ;
        RECT 1519.4400 2434.2800 1521.0400 2434.7600 ;
        RECT 1576.7800 2412.5200 1579.7800 2413.0000 ;
        RECT 1576.7800 2417.9600 1579.7800 2418.4400 ;
        RECT 1576.7800 2423.4000 1579.7800 2423.8800 ;
        RECT 1564.4400 2412.5200 1566.0400 2413.0000 ;
        RECT 1564.4400 2417.9600 1566.0400 2418.4400 ;
        RECT 1564.4400 2423.4000 1566.0400 2423.8800 ;
        RECT 1576.7800 2401.6400 1579.7800 2402.1200 ;
        RECT 1576.7800 2407.0800 1579.7800 2407.5600 ;
        RECT 1564.4400 2401.6400 1566.0400 2402.1200 ;
        RECT 1564.4400 2407.0800 1566.0400 2407.5600 ;
        RECT 1576.7800 2385.3200 1579.7800 2385.8000 ;
        RECT 1576.7800 2390.7600 1579.7800 2391.2400 ;
        RECT 1576.7800 2396.2000 1579.7800 2396.6800 ;
        RECT 1564.4400 2385.3200 1566.0400 2385.8000 ;
        RECT 1564.4400 2390.7600 1566.0400 2391.2400 ;
        RECT 1564.4400 2396.2000 1566.0400 2396.6800 ;
        RECT 1576.7800 2379.8800 1579.7800 2380.3600 ;
        RECT 1564.4400 2379.8800 1566.0400 2380.3600 ;
        RECT 1519.4400 2412.5200 1521.0400 2413.0000 ;
        RECT 1519.4400 2417.9600 1521.0400 2418.4400 ;
        RECT 1519.4400 2423.4000 1521.0400 2423.8800 ;
        RECT 1519.4400 2401.6400 1521.0400 2402.1200 ;
        RECT 1519.4400 2407.0800 1521.0400 2407.5600 ;
        RECT 1519.4400 2385.3200 1521.0400 2385.8000 ;
        RECT 1519.4400 2390.7600 1521.0400 2391.2400 ;
        RECT 1519.4400 2396.2000 1521.0400 2396.6800 ;
        RECT 1519.4400 2379.8800 1521.0400 2380.3600 ;
        RECT 1474.4400 2466.9200 1476.0400 2467.4000 ;
        RECT 1474.4400 2472.3600 1476.0400 2472.8400 ;
        RECT 1474.4400 2477.8000 1476.0400 2478.2800 ;
        RECT 1474.4400 2456.0400 1476.0400 2456.5200 ;
        RECT 1474.4400 2461.4800 1476.0400 2461.9600 ;
        RECT 1429.4400 2466.9200 1431.0400 2467.4000 ;
        RECT 1429.4400 2472.3600 1431.0400 2472.8400 ;
        RECT 1429.4400 2477.8000 1431.0400 2478.2800 ;
        RECT 1429.4400 2456.0400 1431.0400 2456.5200 ;
        RECT 1429.4400 2461.4800 1431.0400 2461.9600 ;
        RECT 1474.4400 2439.7200 1476.0400 2440.2000 ;
        RECT 1474.4400 2445.1600 1476.0400 2445.6400 ;
        RECT 1474.4400 2450.6000 1476.0400 2451.0800 ;
        RECT 1474.4400 2428.8400 1476.0400 2429.3200 ;
        RECT 1474.4400 2434.2800 1476.0400 2434.7600 ;
        RECT 1429.4400 2439.7200 1431.0400 2440.2000 ;
        RECT 1429.4400 2445.1600 1431.0400 2445.6400 ;
        RECT 1429.4400 2450.6000 1431.0400 2451.0800 ;
        RECT 1429.4400 2428.8400 1431.0400 2429.3200 ;
        RECT 1429.4400 2434.2800 1431.0400 2434.7600 ;
        RECT 1384.4400 2466.9200 1386.0400 2467.4000 ;
        RECT 1384.4400 2472.3600 1386.0400 2472.8400 ;
        RECT 1384.4400 2477.8000 1386.0400 2478.2800 ;
        RECT 1372.6800 2466.9200 1375.6800 2467.4000 ;
        RECT 1372.6800 2472.3600 1375.6800 2472.8400 ;
        RECT 1372.6800 2477.8000 1375.6800 2478.2800 ;
        RECT 1384.4400 2456.0400 1386.0400 2456.5200 ;
        RECT 1384.4400 2461.4800 1386.0400 2461.9600 ;
        RECT 1372.6800 2456.0400 1375.6800 2456.5200 ;
        RECT 1372.6800 2461.4800 1375.6800 2461.9600 ;
        RECT 1384.4400 2439.7200 1386.0400 2440.2000 ;
        RECT 1384.4400 2445.1600 1386.0400 2445.6400 ;
        RECT 1384.4400 2450.6000 1386.0400 2451.0800 ;
        RECT 1372.6800 2439.7200 1375.6800 2440.2000 ;
        RECT 1372.6800 2445.1600 1375.6800 2445.6400 ;
        RECT 1372.6800 2450.6000 1375.6800 2451.0800 ;
        RECT 1384.4400 2428.8400 1386.0400 2429.3200 ;
        RECT 1384.4400 2434.2800 1386.0400 2434.7600 ;
        RECT 1372.6800 2428.8400 1375.6800 2429.3200 ;
        RECT 1372.6800 2434.2800 1375.6800 2434.7600 ;
        RECT 1474.4400 2412.5200 1476.0400 2413.0000 ;
        RECT 1474.4400 2417.9600 1476.0400 2418.4400 ;
        RECT 1474.4400 2423.4000 1476.0400 2423.8800 ;
        RECT 1474.4400 2401.6400 1476.0400 2402.1200 ;
        RECT 1474.4400 2407.0800 1476.0400 2407.5600 ;
        RECT 1429.4400 2412.5200 1431.0400 2413.0000 ;
        RECT 1429.4400 2417.9600 1431.0400 2418.4400 ;
        RECT 1429.4400 2423.4000 1431.0400 2423.8800 ;
        RECT 1429.4400 2401.6400 1431.0400 2402.1200 ;
        RECT 1429.4400 2407.0800 1431.0400 2407.5600 ;
        RECT 1474.4400 2385.3200 1476.0400 2385.8000 ;
        RECT 1474.4400 2390.7600 1476.0400 2391.2400 ;
        RECT 1474.4400 2396.2000 1476.0400 2396.6800 ;
        RECT 1474.4400 2379.8800 1476.0400 2380.3600 ;
        RECT 1429.4400 2385.3200 1431.0400 2385.8000 ;
        RECT 1429.4400 2390.7600 1431.0400 2391.2400 ;
        RECT 1429.4400 2396.2000 1431.0400 2396.6800 ;
        RECT 1429.4400 2379.8800 1431.0400 2380.3600 ;
        RECT 1384.4400 2412.5200 1386.0400 2413.0000 ;
        RECT 1384.4400 2417.9600 1386.0400 2418.4400 ;
        RECT 1384.4400 2423.4000 1386.0400 2423.8800 ;
        RECT 1372.6800 2412.5200 1375.6800 2413.0000 ;
        RECT 1372.6800 2417.9600 1375.6800 2418.4400 ;
        RECT 1372.6800 2423.4000 1375.6800 2423.8800 ;
        RECT 1384.4400 2401.6400 1386.0400 2402.1200 ;
        RECT 1384.4400 2407.0800 1386.0400 2407.5600 ;
        RECT 1372.6800 2401.6400 1375.6800 2402.1200 ;
        RECT 1372.6800 2407.0800 1375.6800 2407.5600 ;
        RECT 1384.4400 2385.3200 1386.0400 2385.8000 ;
        RECT 1384.4400 2390.7600 1386.0400 2391.2400 ;
        RECT 1384.4400 2396.2000 1386.0400 2396.6800 ;
        RECT 1372.6800 2385.3200 1375.6800 2385.8000 ;
        RECT 1372.6800 2390.7600 1375.6800 2391.2400 ;
        RECT 1372.6800 2396.2000 1375.6800 2396.6800 ;
        RECT 1372.6800 2379.8800 1375.6800 2380.3600 ;
        RECT 1384.4400 2379.8800 1386.0400 2380.3600 ;
        RECT 1372.6800 2584.7900 1579.7800 2587.7900 ;
        RECT 1372.6800 2371.6900 1579.7800 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 2142.0500 1566.0400 2358.1500 ;
        RECT 1519.4400 2142.0500 1521.0400 2358.1500 ;
        RECT 1474.4400 2142.0500 1476.0400 2358.1500 ;
        RECT 1429.4400 2142.0500 1431.0400 2358.1500 ;
        RECT 1384.4400 2142.0500 1386.0400 2358.1500 ;
        RECT 1576.7800 2142.0500 1579.7800 2358.1500 ;
        RECT 1372.6800 2142.0500 1375.6800 2358.1500 ;
      LAYER met3 ;
        RECT 1576.7800 2335.2000 1579.7800 2335.6800 ;
        RECT 1576.7800 2340.6400 1579.7800 2341.1200 ;
        RECT 1564.4400 2335.2000 1566.0400 2335.6800 ;
        RECT 1564.4400 2340.6400 1566.0400 2341.1200 ;
        RECT 1576.7800 2346.0800 1579.7800 2346.5600 ;
        RECT 1564.4400 2346.0800 1566.0400 2346.5600 ;
        RECT 1576.7800 2324.3200 1579.7800 2324.8000 ;
        RECT 1576.7800 2329.7600 1579.7800 2330.2400 ;
        RECT 1564.4400 2324.3200 1566.0400 2324.8000 ;
        RECT 1564.4400 2329.7600 1566.0400 2330.2400 ;
        RECT 1576.7800 2308.0000 1579.7800 2308.4800 ;
        RECT 1576.7800 2313.4400 1579.7800 2313.9200 ;
        RECT 1564.4400 2308.0000 1566.0400 2308.4800 ;
        RECT 1564.4400 2313.4400 1566.0400 2313.9200 ;
        RECT 1576.7800 2318.8800 1579.7800 2319.3600 ;
        RECT 1564.4400 2318.8800 1566.0400 2319.3600 ;
        RECT 1519.4400 2335.2000 1521.0400 2335.6800 ;
        RECT 1519.4400 2340.6400 1521.0400 2341.1200 ;
        RECT 1519.4400 2346.0800 1521.0400 2346.5600 ;
        RECT 1519.4400 2324.3200 1521.0400 2324.8000 ;
        RECT 1519.4400 2329.7600 1521.0400 2330.2400 ;
        RECT 1519.4400 2308.0000 1521.0400 2308.4800 ;
        RECT 1519.4400 2313.4400 1521.0400 2313.9200 ;
        RECT 1519.4400 2318.8800 1521.0400 2319.3600 ;
        RECT 1576.7800 2291.6800 1579.7800 2292.1600 ;
        RECT 1576.7800 2297.1200 1579.7800 2297.6000 ;
        RECT 1576.7800 2302.5600 1579.7800 2303.0400 ;
        RECT 1564.4400 2291.6800 1566.0400 2292.1600 ;
        RECT 1564.4400 2297.1200 1566.0400 2297.6000 ;
        RECT 1564.4400 2302.5600 1566.0400 2303.0400 ;
        RECT 1576.7800 2280.8000 1579.7800 2281.2800 ;
        RECT 1576.7800 2286.2400 1579.7800 2286.7200 ;
        RECT 1564.4400 2280.8000 1566.0400 2281.2800 ;
        RECT 1564.4400 2286.2400 1566.0400 2286.7200 ;
        RECT 1576.7800 2264.4800 1579.7800 2264.9600 ;
        RECT 1576.7800 2269.9200 1579.7800 2270.4000 ;
        RECT 1576.7800 2275.3600 1579.7800 2275.8400 ;
        RECT 1564.4400 2264.4800 1566.0400 2264.9600 ;
        RECT 1564.4400 2269.9200 1566.0400 2270.4000 ;
        RECT 1564.4400 2275.3600 1566.0400 2275.8400 ;
        RECT 1576.7800 2253.6000 1579.7800 2254.0800 ;
        RECT 1576.7800 2259.0400 1579.7800 2259.5200 ;
        RECT 1564.4400 2253.6000 1566.0400 2254.0800 ;
        RECT 1564.4400 2259.0400 1566.0400 2259.5200 ;
        RECT 1519.4400 2291.6800 1521.0400 2292.1600 ;
        RECT 1519.4400 2297.1200 1521.0400 2297.6000 ;
        RECT 1519.4400 2302.5600 1521.0400 2303.0400 ;
        RECT 1519.4400 2280.8000 1521.0400 2281.2800 ;
        RECT 1519.4400 2286.2400 1521.0400 2286.7200 ;
        RECT 1519.4400 2264.4800 1521.0400 2264.9600 ;
        RECT 1519.4400 2269.9200 1521.0400 2270.4000 ;
        RECT 1519.4400 2275.3600 1521.0400 2275.8400 ;
        RECT 1519.4400 2253.6000 1521.0400 2254.0800 ;
        RECT 1519.4400 2259.0400 1521.0400 2259.5200 ;
        RECT 1474.4400 2335.2000 1476.0400 2335.6800 ;
        RECT 1474.4400 2340.6400 1476.0400 2341.1200 ;
        RECT 1474.4400 2346.0800 1476.0400 2346.5600 ;
        RECT 1429.4400 2335.2000 1431.0400 2335.6800 ;
        RECT 1429.4400 2340.6400 1431.0400 2341.1200 ;
        RECT 1429.4400 2346.0800 1431.0400 2346.5600 ;
        RECT 1474.4400 2324.3200 1476.0400 2324.8000 ;
        RECT 1474.4400 2329.7600 1476.0400 2330.2400 ;
        RECT 1474.4400 2308.0000 1476.0400 2308.4800 ;
        RECT 1474.4400 2313.4400 1476.0400 2313.9200 ;
        RECT 1474.4400 2318.8800 1476.0400 2319.3600 ;
        RECT 1429.4400 2324.3200 1431.0400 2324.8000 ;
        RECT 1429.4400 2329.7600 1431.0400 2330.2400 ;
        RECT 1429.4400 2308.0000 1431.0400 2308.4800 ;
        RECT 1429.4400 2313.4400 1431.0400 2313.9200 ;
        RECT 1429.4400 2318.8800 1431.0400 2319.3600 ;
        RECT 1384.4400 2335.2000 1386.0400 2335.6800 ;
        RECT 1384.4400 2340.6400 1386.0400 2341.1200 ;
        RECT 1372.6800 2340.6400 1375.6800 2341.1200 ;
        RECT 1372.6800 2335.2000 1375.6800 2335.6800 ;
        RECT 1372.6800 2346.0800 1375.6800 2346.5600 ;
        RECT 1384.4400 2346.0800 1386.0400 2346.5600 ;
        RECT 1384.4400 2324.3200 1386.0400 2324.8000 ;
        RECT 1384.4400 2329.7600 1386.0400 2330.2400 ;
        RECT 1372.6800 2329.7600 1375.6800 2330.2400 ;
        RECT 1372.6800 2324.3200 1375.6800 2324.8000 ;
        RECT 1384.4400 2308.0000 1386.0400 2308.4800 ;
        RECT 1384.4400 2313.4400 1386.0400 2313.9200 ;
        RECT 1372.6800 2313.4400 1375.6800 2313.9200 ;
        RECT 1372.6800 2308.0000 1375.6800 2308.4800 ;
        RECT 1372.6800 2318.8800 1375.6800 2319.3600 ;
        RECT 1384.4400 2318.8800 1386.0400 2319.3600 ;
        RECT 1474.4400 2291.6800 1476.0400 2292.1600 ;
        RECT 1474.4400 2297.1200 1476.0400 2297.6000 ;
        RECT 1474.4400 2302.5600 1476.0400 2303.0400 ;
        RECT 1474.4400 2280.8000 1476.0400 2281.2800 ;
        RECT 1474.4400 2286.2400 1476.0400 2286.7200 ;
        RECT 1429.4400 2291.6800 1431.0400 2292.1600 ;
        RECT 1429.4400 2297.1200 1431.0400 2297.6000 ;
        RECT 1429.4400 2302.5600 1431.0400 2303.0400 ;
        RECT 1429.4400 2280.8000 1431.0400 2281.2800 ;
        RECT 1429.4400 2286.2400 1431.0400 2286.7200 ;
        RECT 1474.4400 2264.4800 1476.0400 2264.9600 ;
        RECT 1474.4400 2269.9200 1476.0400 2270.4000 ;
        RECT 1474.4400 2275.3600 1476.0400 2275.8400 ;
        RECT 1474.4400 2253.6000 1476.0400 2254.0800 ;
        RECT 1474.4400 2259.0400 1476.0400 2259.5200 ;
        RECT 1429.4400 2264.4800 1431.0400 2264.9600 ;
        RECT 1429.4400 2269.9200 1431.0400 2270.4000 ;
        RECT 1429.4400 2275.3600 1431.0400 2275.8400 ;
        RECT 1429.4400 2253.6000 1431.0400 2254.0800 ;
        RECT 1429.4400 2259.0400 1431.0400 2259.5200 ;
        RECT 1384.4400 2291.6800 1386.0400 2292.1600 ;
        RECT 1384.4400 2297.1200 1386.0400 2297.6000 ;
        RECT 1384.4400 2302.5600 1386.0400 2303.0400 ;
        RECT 1372.6800 2291.6800 1375.6800 2292.1600 ;
        RECT 1372.6800 2297.1200 1375.6800 2297.6000 ;
        RECT 1372.6800 2302.5600 1375.6800 2303.0400 ;
        RECT 1384.4400 2280.8000 1386.0400 2281.2800 ;
        RECT 1384.4400 2286.2400 1386.0400 2286.7200 ;
        RECT 1372.6800 2280.8000 1375.6800 2281.2800 ;
        RECT 1372.6800 2286.2400 1375.6800 2286.7200 ;
        RECT 1384.4400 2264.4800 1386.0400 2264.9600 ;
        RECT 1384.4400 2269.9200 1386.0400 2270.4000 ;
        RECT 1384.4400 2275.3600 1386.0400 2275.8400 ;
        RECT 1372.6800 2264.4800 1375.6800 2264.9600 ;
        RECT 1372.6800 2269.9200 1375.6800 2270.4000 ;
        RECT 1372.6800 2275.3600 1375.6800 2275.8400 ;
        RECT 1384.4400 2253.6000 1386.0400 2254.0800 ;
        RECT 1384.4400 2259.0400 1386.0400 2259.5200 ;
        RECT 1372.6800 2253.6000 1375.6800 2254.0800 ;
        RECT 1372.6800 2259.0400 1375.6800 2259.5200 ;
        RECT 1576.7800 2237.2800 1579.7800 2237.7600 ;
        RECT 1576.7800 2242.7200 1579.7800 2243.2000 ;
        RECT 1576.7800 2248.1600 1579.7800 2248.6400 ;
        RECT 1564.4400 2237.2800 1566.0400 2237.7600 ;
        RECT 1564.4400 2242.7200 1566.0400 2243.2000 ;
        RECT 1564.4400 2248.1600 1566.0400 2248.6400 ;
        RECT 1576.7800 2226.4000 1579.7800 2226.8800 ;
        RECT 1576.7800 2231.8400 1579.7800 2232.3200 ;
        RECT 1564.4400 2226.4000 1566.0400 2226.8800 ;
        RECT 1564.4400 2231.8400 1566.0400 2232.3200 ;
        RECT 1576.7800 2210.0800 1579.7800 2210.5600 ;
        RECT 1576.7800 2215.5200 1579.7800 2216.0000 ;
        RECT 1576.7800 2220.9600 1579.7800 2221.4400 ;
        RECT 1564.4400 2210.0800 1566.0400 2210.5600 ;
        RECT 1564.4400 2215.5200 1566.0400 2216.0000 ;
        RECT 1564.4400 2220.9600 1566.0400 2221.4400 ;
        RECT 1576.7800 2199.2000 1579.7800 2199.6800 ;
        RECT 1576.7800 2204.6400 1579.7800 2205.1200 ;
        RECT 1564.4400 2199.2000 1566.0400 2199.6800 ;
        RECT 1564.4400 2204.6400 1566.0400 2205.1200 ;
        RECT 1519.4400 2237.2800 1521.0400 2237.7600 ;
        RECT 1519.4400 2242.7200 1521.0400 2243.2000 ;
        RECT 1519.4400 2248.1600 1521.0400 2248.6400 ;
        RECT 1519.4400 2226.4000 1521.0400 2226.8800 ;
        RECT 1519.4400 2231.8400 1521.0400 2232.3200 ;
        RECT 1519.4400 2210.0800 1521.0400 2210.5600 ;
        RECT 1519.4400 2215.5200 1521.0400 2216.0000 ;
        RECT 1519.4400 2220.9600 1521.0400 2221.4400 ;
        RECT 1519.4400 2199.2000 1521.0400 2199.6800 ;
        RECT 1519.4400 2204.6400 1521.0400 2205.1200 ;
        RECT 1576.7800 2182.8800 1579.7800 2183.3600 ;
        RECT 1576.7800 2188.3200 1579.7800 2188.8000 ;
        RECT 1576.7800 2193.7600 1579.7800 2194.2400 ;
        RECT 1564.4400 2182.8800 1566.0400 2183.3600 ;
        RECT 1564.4400 2188.3200 1566.0400 2188.8000 ;
        RECT 1564.4400 2193.7600 1566.0400 2194.2400 ;
        RECT 1576.7800 2172.0000 1579.7800 2172.4800 ;
        RECT 1576.7800 2177.4400 1579.7800 2177.9200 ;
        RECT 1564.4400 2172.0000 1566.0400 2172.4800 ;
        RECT 1564.4400 2177.4400 1566.0400 2177.9200 ;
        RECT 1576.7800 2155.6800 1579.7800 2156.1600 ;
        RECT 1576.7800 2161.1200 1579.7800 2161.6000 ;
        RECT 1576.7800 2166.5600 1579.7800 2167.0400 ;
        RECT 1564.4400 2155.6800 1566.0400 2156.1600 ;
        RECT 1564.4400 2161.1200 1566.0400 2161.6000 ;
        RECT 1564.4400 2166.5600 1566.0400 2167.0400 ;
        RECT 1576.7800 2150.2400 1579.7800 2150.7200 ;
        RECT 1564.4400 2150.2400 1566.0400 2150.7200 ;
        RECT 1519.4400 2182.8800 1521.0400 2183.3600 ;
        RECT 1519.4400 2188.3200 1521.0400 2188.8000 ;
        RECT 1519.4400 2193.7600 1521.0400 2194.2400 ;
        RECT 1519.4400 2172.0000 1521.0400 2172.4800 ;
        RECT 1519.4400 2177.4400 1521.0400 2177.9200 ;
        RECT 1519.4400 2155.6800 1521.0400 2156.1600 ;
        RECT 1519.4400 2161.1200 1521.0400 2161.6000 ;
        RECT 1519.4400 2166.5600 1521.0400 2167.0400 ;
        RECT 1519.4400 2150.2400 1521.0400 2150.7200 ;
        RECT 1474.4400 2237.2800 1476.0400 2237.7600 ;
        RECT 1474.4400 2242.7200 1476.0400 2243.2000 ;
        RECT 1474.4400 2248.1600 1476.0400 2248.6400 ;
        RECT 1474.4400 2226.4000 1476.0400 2226.8800 ;
        RECT 1474.4400 2231.8400 1476.0400 2232.3200 ;
        RECT 1429.4400 2237.2800 1431.0400 2237.7600 ;
        RECT 1429.4400 2242.7200 1431.0400 2243.2000 ;
        RECT 1429.4400 2248.1600 1431.0400 2248.6400 ;
        RECT 1429.4400 2226.4000 1431.0400 2226.8800 ;
        RECT 1429.4400 2231.8400 1431.0400 2232.3200 ;
        RECT 1474.4400 2210.0800 1476.0400 2210.5600 ;
        RECT 1474.4400 2215.5200 1476.0400 2216.0000 ;
        RECT 1474.4400 2220.9600 1476.0400 2221.4400 ;
        RECT 1474.4400 2199.2000 1476.0400 2199.6800 ;
        RECT 1474.4400 2204.6400 1476.0400 2205.1200 ;
        RECT 1429.4400 2210.0800 1431.0400 2210.5600 ;
        RECT 1429.4400 2215.5200 1431.0400 2216.0000 ;
        RECT 1429.4400 2220.9600 1431.0400 2221.4400 ;
        RECT 1429.4400 2199.2000 1431.0400 2199.6800 ;
        RECT 1429.4400 2204.6400 1431.0400 2205.1200 ;
        RECT 1384.4400 2237.2800 1386.0400 2237.7600 ;
        RECT 1384.4400 2242.7200 1386.0400 2243.2000 ;
        RECT 1384.4400 2248.1600 1386.0400 2248.6400 ;
        RECT 1372.6800 2237.2800 1375.6800 2237.7600 ;
        RECT 1372.6800 2242.7200 1375.6800 2243.2000 ;
        RECT 1372.6800 2248.1600 1375.6800 2248.6400 ;
        RECT 1384.4400 2226.4000 1386.0400 2226.8800 ;
        RECT 1384.4400 2231.8400 1386.0400 2232.3200 ;
        RECT 1372.6800 2226.4000 1375.6800 2226.8800 ;
        RECT 1372.6800 2231.8400 1375.6800 2232.3200 ;
        RECT 1384.4400 2210.0800 1386.0400 2210.5600 ;
        RECT 1384.4400 2215.5200 1386.0400 2216.0000 ;
        RECT 1384.4400 2220.9600 1386.0400 2221.4400 ;
        RECT 1372.6800 2210.0800 1375.6800 2210.5600 ;
        RECT 1372.6800 2215.5200 1375.6800 2216.0000 ;
        RECT 1372.6800 2220.9600 1375.6800 2221.4400 ;
        RECT 1384.4400 2199.2000 1386.0400 2199.6800 ;
        RECT 1384.4400 2204.6400 1386.0400 2205.1200 ;
        RECT 1372.6800 2199.2000 1375.6800 2199.6800 ;
        RECT 1372.6800 2204.6400 1375.6800 2205.1200 ;
        RECT 1474.4400 2182.8800 1476.0400 2183.3600 ;
        RECT 1474.4400 2188.3200 1476.0400 2188.8000 ;
        RECT 1474.4400 2193.7600 1476.0400 2194.2400 ;
        RECT 1474.4400 2172.0000 1476.0400 2172.4800 ;
        RECT 1474.4400 2177.4400 1476.0400 2177.9200 ;
        RECT 1429.4400 2182.8800 1431.0400 2183.3600 ;
        RECT 1429.4400 2188.3200 1431.0400 2188.8000 ;
        RECT 1429.4400 2193.7600 1431.0400 2194.2400 ;
        RECT 1429.4400 2172.0000 1431.0400 2172.4800 ;
        RECT 1429.4400 2177.4400 1431.0400 2177.9200 ;
        RECT 1474.4400 2155.6800 1476.0400 2156.1600 ;
        RECT 1474.4400 2161.1200 1476.0400 2161.6000 ;
        RECT 1474.4400 2166.5600 1476.0400 2167.0400 ;
        RECT 1474.4400 2150.2400 1476.0400 2150.7200 ;
        RECT 1429.4400 2155.6800 1431.0400 2156.1600 ;
        RECT 1429.4400 2161.1200 1431.0400 2161.6000 ;
        RECT 1429.4400 2166.5600 1431.0400 2167.0400 ;
        RECT 1429.4400 2150.2400 1431.0400 2150.7200 ;
        RECT 1384.4400 2182.8800 1386.0400 2183.3600 ;
        RECT 1384.4400 2188.3200 1386.0400 2188.8000 ;
        RECT 1384.4400 2193.7600 1386.0400 2194.2400 ;
        RECT 1372.6800 2182.8800 1375.6800 2183.3600 ;
        RECT 1372.6800 2188.3200 1375.6800 2188.8000 ;
        RECT 1372.6800 2193.7600 1375.6800 2194.2400 ;
        RECT 1384.4400 2172.0000 1386.0400 2172.4800 ;
        RECT 1384.4400 2177.4400 1386.0400 2177.9200 ;
        RECT 1372.6800 2172.0000 1375.6800 2172.4800 ;
        RECT 1372.6800 2177.4400 1375.6800 2177.9200 ;
        RECT 1384.4400 2155.6800 1386.0400 2156.1600 ;
        RECT 1384.4400 2161.1200 1386.0400 2161.6000 ;
        RECT 1384.4400 2166.5600 1386.0400 2167.0400 ;
        RECT 1372.6800 2155.6800 1375.6800 2156.1600 ;
        RECT 1372.6800 2161.1200 1375.6800 2161.6000 ;
        RECT 1372.6800 2166.5600 1375.6800 2167.0400 ;
        RECT 1372.6800 2150.2400 1375.6800 2150.7200 ;
        RECT 1384.4400 2150.2400 1386.0400 2150.7200 ;
        RECT 1372.6800 2355.1500 1579.7800 2358.1500 ;
        RECT 1372.6800 2142.0500 1579.7800 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 1912.4100 1566.0400 2128.5100 ;
        RECT 1519.4400 1912.4100 1521.0400 2128.5100 ;
        RECT 1474.4400 1912.4100 1476.0400 2128.5100 ;
        RECT 1429.4400 1912.4100 1431.0400 2128.5100 ;
        RECT 1384.4400 1912.4100 1386.0400 2128.5100 ;
        RECT 1576.7800 1912.4100 1579.7800 2128.5100 ;
        RECT 1372.6800 1912.4100 1375.6800 2128.5100 ;
      LAYER met3 ;
        RECT 1576.7800 2105.5600 1579.7800 2106.0400 ;
        RECT 1576.7800 2111.0000 1579.7800 2111.4800 ;
        RECT 1564.4400 2105.5600 1566.0400 2106.0400 ;
        RECT 1564.4400 2111.0000 1566.0400 2111.4800 ;
        RECT 1576.7800 2116.4400 1579.7800 2116.9200 ;
        RECT 1564.4400 2116.4400 1566.0400 2116.9200 ;
        RECT 1576.7800 2094.6800 1579.7800 2095.1600 ;
        RECT 1576.7800 2100.1200 1579.7800 2100.6000 ;
        RECT 1564.4400 2094.6800 1566.0400 2095.1600 ;
        RECT 1564.4400 2100.1200 1566.0400 2100.6000 ;
        RECT 1576.7800 2078.3600 1579.7800 2078.8400 ;
        RECT 1576.7800 2083.8000 1579.7800 2084.2800 ;
        RECT 1564.4400 2078.3600 1566.0400 2078.8400 ;
        RECT 1564.4400 2083.8000 1566.0400 2084.2800 ;
        RECT 1576.7800 2089.2400 1579.7800 2089.7200 ;
        RECT 1564.4400 2089.2400 1566.0400 2089.7200 ;
        RECT 1519.4400 2105.5600 1521.0400 2106.0400 ;
        RECT 1519.4400 2111.0000 1521.0400 2111.4800 ;
        RECT 1519.4400 2116.4400 1521.0400 2116.9200 ;
        RECT 1519.4400 2094.6800 1521.0400 2095.1600 ;
        RECT 1519.4400 2100.1200 1521.0400 2100.6000 ;
        RECT 1519.4400 2078.3600 1521.0400 2078.8400 ;
        RECT 1519.4400 2083.8000 1521.0400 2084.2800 ;
        RECT 1519.4400 2089.2400 1521.0400 2089.7200 ;
        RECT 1576.7800 2062.0400 1579.7800 2062.5200 ;
        RECT 1576.7800 2067.4800 1579.7800 2067.9600 ;
        RECT 1576.7800 2072.9200 1579.7800 2073.4000 ;
        RECT 1564.4400 2062.0400 1566.0400 2062.5200 ;
        RECT 1564.4400 2067.4800 1566.0400 2067.9600 ;
        RECT 1564.4400 2072.9200 1566.0400 2073.4000 ;
        RECT 1576.7800 2051.1600 1579.7800 2051.6400 ;
        RECT 1576.7800 2056.6000 1579.7800 2057.0800 ;
        RECT 1564.4400 2051.1600 1566.0400 2051.6400 ;
        RECT 1564.4400 2056.6000 1566.0400 2057.0800 ;
        RECT 1576.7800 2034.8400 1579.7800 2035.3200 ;
        RECT 1576.7800 2040.2800 1579.7800 2040.7600 ;
        RECT 1576.7800 2045.7200 1579.7800 2046.2000 ;
        RECT 1564.4400 2034.8400 1566.0400 2035.3200 ;
        RECT 1564.4400 2040.2800 1566.0400 2040.7600 ;
        RECT 1564.4400 2045.7200 1566.0400 2046.2000 ;
        RECT 1576.7800 2023.9600 1579.7800 2024.4400 ;
        RECT 1576.7800 2029.4000 1579.7800 2029.8800 ;
        RECT 1564.4400 2023.9600 1566.0400 2024.4400 ;
        RECT 1564.4400 2029.4000 1566.0400 2029.8800 ;
        RECT 1519.4400 2062.0400 1521.0400 2062.5200 ;
        RECT 1519.4400 2067.4800 1521.0400 2067.9600 ;
        RECT 1519.4400 2072.9200 1521.0400 2073.4000 ;
        RECT 1519.4400 2051.1600 1521.0400 2051.6400 ;
        RECT 1519.4400 2056.6000 1521.0400 2057.0800 ;
        RECT 1519.4400 2034.8400 1521.0400 2035.3200 ;
        RECT 1519.4400 2040.2800 1521.0400 2040.7600 ;
        RECT 1519.4400 2045.7200 1521.0400 2046.2000 ;
        RECT 1519.4400 2023.9600 1521.0400 2024.4400 ;
        RECT 1519.4400 2029.4000 1521.0400 2029.8800 ;
        RECT 1474.4400 2105.5600 1476.0400 2106.0400 ;
        RECT 1474.4400 2111.0000 1476.0400 2111.4800 ;
        RECT 1474.4400 2116.4400 1476.0400 2116.9200 ;
        RECT 1429.4400 2105.5600 1431.0400 2106.0400 ;
        RECT 1429.4400 2111.0000 1431.0400 2111.4800 ;
        RECT 1429.4400 2116.4400 1431.0400 2116.9200 ;
        RECT 1474.4400 2094.6800 1476.0400 2095.1600 ;
        RECT 1474.4400 2100.1200 1476.0400 2100.6000 ;
        RECT 1474.4400 2078.3600 1476.0400 2078.8400 ;
        RECT 1474.4400 2083.8000 1476.0400 2084.2800 ;
        RECT 1474.4400 2089.2400 1476.0400 2089.7200 ;
        RECT 1429.4400 2094.6800 1431.0400 2095.1600 ;
        RECT 1429.4400 2100.1200 1431.0400 2100.6000 ;
        RECT 1429.4400 2078.3600 1431.0400 2078.8400 ;
        RECT 1429.4400 2083.8000 1431.0400 2084.2800 ;
        RECT 1429.4400 2089.2400 1431.0400 2089.7200 ;
        RECT 1384.4400 2105.5600 1386.0400 2106.0400 ;
        RECT 1384.4400 2111.0000 1386.0400 2111.4800 ;
        RECT 1372.6800 2111.0000 1375.6800 2111.4800 ;
        RECT 1372.6800 2105.5600 1375.6800 2106.0400 ;
        RECT 1372.6800 2116.4400 1375.6800 2116.9200 ;
        RECT 1384.4400 2116.4400 1386.0400 2116.9200 ;
        RECT 1384.4400 2094.6800 1386.0400 2095.1600 ;
        RECT 1384.4400 2100.1200 1386.0400 2100.6000 ;
        RECT 1372.6800 2100.1200 1375.6800 2100.6000 ;
        RECT 1372.6800 2094.6800 1375.6800 2095.1600 ;
        RECT 1384.4400 2078.3600 1386.0400 2078.8400 ;
        RECT 1384.4400 2083.8000 1386.0400 2084.2800 ;
        RECT 1372.6800 2083.8000 1375.6800 2084.2800 ;
        RECT 1372.6800 2078.3600 1375.6800 2078.8400 ;
        RECT 1372.6800 2089.2400 1375.6800 2089.7200 ;
        RECT 1384.4400 2089.2400 1386.0400 2089.7200 ;
        RECT 1474.4400 2062.0400 1476.0400 2062.5200 ;
        RECT 1474.4400 2067.4800 1476.0400 2067.9600 ;
        RECT 1474.4400 2072.9200 1476.0400 2073.4000 ;
        RECT 1474.4400 2051.1600 1476.0400 2051.6400 ;
        RECT 1474.4400 2056.6000 1476.0400 2057.0800 ;
        RECT 1429.4400 2062.0400 1431.0400 2062.5200 ;
        RECT 1429.4400 2067.4800 1431.0400 2067.9600 ;
        RECT 1429.4400 2072.9200 1431.0400 2073.4000 ;
        RECT 1429.4400 2051.1600 1431.0400 2051.6400 ;
        RECT 1429.4400 2056.6000 1431.0400 2057.0800 ;
        RECT 1474.4400 2034.8400 1476.0400 2035.3200 ;
        RECT 1474.4400 2040.2800 1476.0400 2040.7600 ;
        RECT 1474.4400 2045.7200 1476.0400 2046.2000 ;
        RECT 1474.4400 2023.9600 1476.0400 2024.4400 ;
        RECT 1474.4400 2029.4000 1476.0400 2029.8800 ;
        RECT 1429.4400 2034.8400 1431.0400 2035.3200 ;
        RECT 1429.4400 2040.2800 1431.0400 2040.7600 ;
        RECT 1429.4400 2045.7200 1431.0400 2046.2000 ;
        RECT 1429.4400 2023.9600 1431.0400 2024.4400 ;
        RECT 1429.4400 2029.4000 1431.0400 2029.8800 ;
        RECT 1384.4400 2062.0400 1386.0400 2062.5200 ;
        RECT 1384.4400 2067.4800 1386.0400 2067.9600 ;
        RECT 1384.4400 2072.9200 1386.0400 2073.4000 ;
        RECT 1372.6800 2062.0400 1375.6800 2062.5200 ;
        RECT 1372.6800 2067.4800 1375.6800 2067.9600 ;
        RECT 1372.6800 2072.9200 1375.6800 2073.4000 ;
        RECT 1384.4400 2051.1600 1386.0400 2051.6400 ;
        RECT 1384.4400 2056.6000 1386.0400 2057.0800 ;
        RECT 1372.6800 2051.1600 1375.6800 2051.6400 ;
        RECT 1372.6800 2056.6000 1375.6800 2057.0800 ;
        RECT 1384.4400 2034.8400 1386.0400 2035.3200 ;
        RECT 1384.4400 2040.2800 1386.0400 2040.7600 ;
        RECT 1384.4400 2045.7200 1386.0400 2046.2000 ;
        RECT 1372.6800 2034.8400 1375.6800 2035.3200 ;
        RECT 1372.6800 2040.2800 1375.6800 2040.7600 ;
        RECT 1372.6800 2045.7200 1375.6800 2046.2000 ;
        RECT 1384.4400 2023.9600 1386.0400 2024.4400 ;
        RECT 1384.4400 2029.4000 1386.0400 2029.8800 ;
        RECT 1372.6800 2023.9600 1375.6800 2024.4400 ;
        RECT 1372.6800 2029.4000 1375.6800 2029.8800 ;
        RECT 1576.7800 2007.6400 1579.7800 2008.1200 ;
        RECT 1576.7800 2013.0800 1579.7800 2013.5600 ;
        RECT 1576.7800 2018.5200 1579.7800 2019.0000 ;
        RECT 1564.4400 2007.6400 1566.0400 2008.1200 ;
        RECT 1564.4400 2013.0800 1566.0400 2013.5600 ;
        RECT 1564.4400 2018.5200 1566.0400 2019.0000 ;
        RECT 1576.7800 1996.7600 1579.7800 1997.2400 ;
        RECT 1576.7800 2002.2000 1579.7800 2002.6800 ;
        RECT 1564.4400 1996.7600 1566.0400 1997.2400 ;
        RECT 1564.4400 2002.2000 1566.0400 2002.6800 ;
        RECT 1576.7800 1980.4400 1579.7800 1980.9200 ;
        RECT 1576.7800 1985.8800 1579.7800 1986.3600 ;
        RECT 1576.7800 1991.3200 1579.7800 1991.8000 ;
        RECT 1564.4400 1980.4400 1566.0400 1980.9200 ;
        RECT 1564.4400 1985.8800 1566.0400 1986.3600 ;
        RECT 1564.4400 1991.3200 1566.0400 1991.8000 ;
        RECT 1576.7800 1969.5600 1579.7800 1970.0400 ;
        RECT 1576.7800 1975.0000 1579.7800 1975.4800 ;
        RECT 1564.4400 1969.5600 1566.0400 1970.0400 ;
        RECT 1564.4400 1975.0000 1566.0400 1975.4800 ;
        RECT 1519.4400 2007.6400 1521.0400 2008.1200 ;
        RECT 1519.4400 2013.0800 1521.0400 2013.5600 ;
        RECT 1519.4400 2018.5200 1521.0400 2019.0000 ;
        RECT 1519.4400 1996.7600 1521.0400 1997.2400 ;
        RECT 1519.4400 2002.2000 1521.0400 2002.6800 ;
        RECT 1519.4400 1980.4400 1521.0400 1980.9200 ;
        RECT 1519.4400 1985.8800 1521.0400 1986.3600 ;
        RECT 1519.4400 1991.3200 1521.0400 1991.8000 ;
        RECT 1519.4400 1969.5600 1521.0400 1970.0400 ;
        RECT 1519.4400 1975.0000 1521.0400 1975.4800 ;
        RECT 1576.7800 1953.2400 1579.7800 1953.7200 ;
        RECT 1576.7800 1958.6800 1579.7800 1959.1600 ;
        RECT 1576.7800 1964.1200 1579.7800 1964.6000 ;
        RECT 1564.4400 1953.2400 1566.0400 1953.7200 ;
        RECT 1564.4400 1958.6800 1566.0400 1959.1600 ;
        RECT 1564.4400 1964.1200 1566.0400 1964.6000 ;
        RECT 1576.7800 1942.3600 1579.7800 1942.8400 ;
        RECT 1576.7800 1947.8000 1579.7800 1948.2800 ;
        RECT 1564.4400 1942.3600 1566.0400 1942.8400 ;
        RECT 1564.4400 1947.8000 1566.0400 1948.2800 ;
        RECT 1576.7800 1926.0400 1579.7800 1926.5200 ;
        RECT 1576.7800 1931.4800 1579.7800 1931.9600 ;
        RECT 1576.7800 1936.9200 1579.7800 1937.4000 ;
        RECT 1564.4400 1926.0400 1566.0400 1926.5200 ;
        RECT 1564.4400 1931.4800 1566.0400 1931.9600 ;
        RECT 1564.4400 1936.9200 1566.0400 1937.4000 ;
        RECT 1576.7800 1920.6000 1579.7800 1921.0800 ;
        RECT 1564.4400 1920.6000 1566.0400 1921.0800 ;
        RECT 1519.4400 1953.2400 1521.0400 1953.7200 ;
        RECT 1519.4400 1958.6800 1521.0400 1959.1600 ;
        RECT 1519.4400 1964.1200 1521.0400 1964.6000 ;
        RECT 1519.4400 1942.3600 1521.0400 1942.8400 ;
        RECT 1519.4400 1947.8000 1521.0400 1948.2800 ;
        RECT 1519.4400 1926.0400 1521.0400 1926.5200 ;
        RECT 1519.4400 1931.4800 1521.0400 1931.9600 ;
        RECT 1519.4400 1936.9200 1521.0400 1937.4000 ;
        RECT 1519.4400 1920.6000 1521.0400 1921.0800 ;
        RECT 1474.4400 2007.6400 1476.0400 2008.1200 ;
        RECT 1474.4400 2013.0800 1476.0400 2013.5600 ;
        RECT 1474.4400 2018.5200 1476.0400 2019.0000 ;
        RECT 1474.4400 1996.7600 1476.0400 1997.2400 ;
        RECT 1474.4400 2002.2000 1476.0400 2002.6800 ;
        RECT 1429.4400 2007.6400 1431.0400 2008.1200 ;
        RECT 1429.4400 2013.0800 1431.0400 2013.5600 ;
        RECT 1429.4400 2018.5200 1431.0400 2019.0000 ;
        RECT 1429.4400 1996.7600 1431.0400 1997.2400 ;
        RECT 1429.4400 2002.2000 1431.0400 2002.6800 ;
        RECT 1474.4400 1980.4400 1476.0400 1980.9200 ;
        RECT 1474.4400 1985.8800 1476.0400 1986.3600 ;
        RECT 1474.4400 1991.3200 1476.0400 1991.8000 ;
        RECT 1474.4400 1969.5600 1476.0400 1970.0400 ;
        RECT 1474.4400 1975.0000 1476.0400 1975.4800 ;
        RECT 1429.4400 1980.4400 1431.0400 1980.9200 ;
        RECT 1429.4400 1985.8800 1431.0400 1986.3600 ;
        RECT 1429.4400 1991.3200 1431.0400 1991.8000 ;
        RECT 1429.4400 1969.5600 1431.0400 1970.0400 ;
        RECT 1429.4400 1975.0000 1431.0400 1975.4800 ;
        RECT 1384.4400 2007.6400 1386.0400 2008.1200 ;
        RECT 1384.4400 2013.0800 1386.0400 2013.5600 ;
        RECT 1384.4400 2018.5200 1386.0400 2019.0000 ;
        RECT 1372.6800 2007.6400 1375.6800 2008.1200 ;
        RECT 1372.6800 2013.0800 1375.6800 2013.5600 ;
        RECT 1372.6800 2018.5200 1375.6800 2019.0000 ;
        RECT 1384.4400 1996.7600 1386.0400 1997.2400 ;
        RECT 1384.4400 2002.2000 1386.0400 2002.6800 ;
        RECT 1372.6800 1996.7600 1375.6800 1997.2400 ;
        RECT 1372.6800 2002.2000 1375.6800 2002.6800 ;
        RECT 1384.4400 1980.4400 1386.0400 1980.9200 ;
        RECT 1384.4400 1985.8800 1386.0400 1986.3600 ;
        RECT 1384.4400 1991.3200 1386.0400 1991.8000 ;
        RECT 1372.6800 1980.4400 1375.6800 1980.9200 ;
        RECT 1372.6800 1985.8800 1375.6800 1986.3600 ;
        RECT 1372.6800 1991.3200 1375.6800 1991.8000 ;
        RECT 1384.4400 1969.5600 1386.0400 1970.0400 ;
        RECT 1384.4400 1975.0000 1386.0400 1975.4800 ;
        RECT 1372.6800 1969.5600 1375.6800 1970.0400 ;
        RECT 1372.6800 1975.0000 1375.6800 1975.4800 ;
        RECT 1474.4400 1953.2400 1476.0400 1953.7200 ;
        RECT 1474.4400 1958.6800 1476.0400 1959.1600 ;
        RECT 1474.4400 1964.1200 1476.0400 1964.6000 ;
        RECT 1474.4400 1942.3600 1476.0400 1942.8400 ;
        RECT 1474.4400 1947.8000 1476.0400 1948.2800 ;
        RECT 1429.4400 1953.2400 1431.0400 1953.7200 ;
        RECT 1429.4400 1958.6800 1431.0400 1959.1600 ;
        RECT 1429.4400 1964.1200 1431.0400 1964.6000 ;
        RECT 1429.4400 1942.3600 1431.0400 1942.8400 ;
        RECT 1429.4400 1947.8000 1431.0400 1948.2800 ;
        RECT 1474.4400 1926.0400 1476.0400 1926.5200 ;
        RECT 1474.4400 1931.4800 1476.0400 1931.9600 ;
        RECT 1474.4400 1936.9200 1476.0400 1937.4000 ;
        RECT 1474.4400 1920.6000 1476.0400 1921.0800 ;
        RECT 1429.4400 1926.0400 1431.0400 1926.5200 ;
        RECT 1429.4400 1931.4800 1431.0400 1931.9600 ;
        RECT 1429.4400 1936.9200 1431.0400 1937.4000 ;
        RECT 1429.4400 1920.6000 1431.0400 1921.0800 ;
        RECT 1384.4400 1953.2400 1386.0400 1953.7200 ;
        RECT 1384.4400 1958.6800 1386.0400 1959.1600 ;
        RECT 1384.4400 1964.1200 1386.0400 1964.6000 ;
        RECT 1372.6800 1953.2400 1375.6800 1953.7200 ;
        RECT 1372.6800 1958.6800 1375.6800 1959.1600 ;
        RECT 1372.6800 1964.1200 1375.6800 1964.6000 ;
        RECT 1384.4400 1942.3600 1386.0400 1942.8400 ;
        RECT 1384.4400 1947.8000 1386.0400 1948.2800 ;
        RECT 1372.6800 1942.3600 1375.6800 1942.8400 ;
        RECT 1372.6800 1947.8000 1375.6800 1948.2800 ;
        RECT 1384.4400 1926.0400 1386.0400 1926.5200 ;
        RECT 1384.4400 1931.4800 1386.0400 1931.9600 ;
        RECT 1384.4400 1936.9200 1386.0400 1937.4000 ;
        RECT 1372.6800 1926.0400 1375.6800 1926.5200 ;
        RECT 1372.6800 1931.4800 1375.6800 1931.9600 ;
        RECT 1372.6800 1936.9200 1375.6800 1937.4000 ;
        RECT 1372.6800 1920.6000 1375.6800 1921.0800 ;
        RECT 1384.4400 1920.6000 1386.0400 1921.0800 ;
        RECT 1372.6800 2125.5100 1579.7800 2128.5100 ;
        RECT 1372.6800 1912.4100 1579.7800 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 1682.7700 1566.0400 1898.8700 ;
        RECT 1519.4400 1682.7700 1521.0400 1898.8700 ;
        RECT 1474.4400 1682.7700 1476.0400 1898.8700 ;
        RECT 1429.4400 1682.7700 1431.0400 1898.8700 ;
        RECT 1384.4400 1682.7700 1386.0400 1898.8700 ;
        RECT 1576.7800 1682.7700 1579.7800 1898.8700 ;
        RECT 1372.6800 1682.7700 1375.6800 1898.8700 ;
      LAYER met3 ;
        RECT 1576.7800 1875.9200 1579.7800 1876.4000 ;
        RECT 1576.7800 1881.3600 1579.7800 1881.8400 ;
        RECT 1564.4400 1875.9200 1566.0400 1876.4000 ;
        RECT 1564.4400 1881.3600 1566.0400 1881.8400 ;
        RECT 1576.7800 1886.8000 1579.7800 1887.2800 ;
        RECT 1564.4400 1886.8000 1566.0400 1887.2800 ;
        RECT 1576.7800 1865.0400 1579.7800 1865.5200 ;
        RECT 1576.7800 1870.4800 1579.7800 1870.9600 ;
        RECT 1564.4400 1865.0400 1566.0400 1865.5200 ;
        RECT 1564.4400 1870.4800 1566.0400 1870.9600 ;
        RECT 1576.7800 1848.7200 1579.7800 1849.2000 ;
        RECT 1576.7800 1854.1600 1579.7800 1854.6400 ;
        RECT 1564.4400 1848.7200 1566.0400 1849.2000 ;
        RECT 1564.4400 1854.1600 1566.0400 1854.6400 ;
        RECT 1576.7800 1859.6000 1579.7800 1860.0800 ;
        RECT 1564.4400 1859.6000 1566.0400 1860.0800 ;
        RECT 1519.4400 1875.9200 1521.0400 1876.4000 ;
        RECT 1519.4400 1881.3600 1521.0400 1881.8400 ;
        RECT 1519.4400 1886.8000 1521.0400 1887.2800 ;
        RECT 1519.4400 1865.0400 1521.0400 1865.5200 ;
        RECT 1519.4400 1870.4800 1521.0400 1870.9600 ;
        RECT 1519.4400 1848.7200 1521.0400 1849.2000 ;
        RECT 1519.4400 1854.1600 1521.0400 1854.6400 ;
        RECT 1519.4400 1859.6000 1521.0400 1860.0800 ;
        RECT 1576.7800 1832.4000 1579.7800 1832.8800 ;
        RECT 1576.7800 1837.8400 1579.7800 1838.3200 ;
        RECT 1576.7800 1843.2800 1579.7800 1843.7600 ;
        RECT 1564.4400 1832.4000 1566.0400 1832.8800 ;
        RECT 1564.4400 1837.8400 1566.0400 1838.3200 ;
        RECT 1564.4400 1843.2800 1566.0400 1843.7600 ;
        RECT 1576.7800 1821.5200 1579.7800 1822.0000 ;
        RECT 1576.7800 1826.9600 1579.7800 1827.4400 ;
        RECT 1564.4400 1821.5200 1566.0400 1822.0000 ;
        RECT 1564.4400 1826.9600 1566.0400 1827.4400 ;
        RECT 1576.7800 1805.2000 1579.7800 1805.6800 ;
        RECT 1576.7800 1810.6400 1579.7800 1811.1200 ;
        RECT 1576.7800 1816.0800 1579.7800 1816.5600 ;
        RECT 1564.4400 1805.2000 1566.0400 1805.6800 ;
        RECT 1564.4400 1810.6400 1566.0400 1811.1200 ;
        RECT 1564.4400 1816.0800 1566.0400 1816.5600 ;
        RECT 1576.7800 1794.3200 1579.7800 1794.8000 ;
        RECT 1576.7800 1799.7600 1579.7800 1800.2400 ;
        RECT 1564.4400 1794.3200 1566.0400 1794.8000 ;
        RECT 1564.4400 1799.7600 1566.0400 1800.2400 ;
        RECT 1519.4400 1832.4000 1521.0400 1832.8800 ;
        RECT 1519.4400 1837.8400 1521.0400 1838.3200 ;
        RECT 1519.4400 1843.2800 1521.0400 1843.7600 ;
        RECT 1519.4400 1821.5200 1521.0400 1822.0000 ;
        RECT 1519.4400 1826.9600 1521.0400 1827.4400 ;
        RECT 1519.4400 1805.2000 1521.0400 1805.6800 ;
        RECT 1519.4400 1810.6400 1521.0400 1811.1200 ;
        RECT 1519.4400 1816.0800 1521.0400 1816.5600 ;
        RECT 1519.4400 1794.3200 1521.0400 1794.8000 ;
        RECT 1519.4400 1799.7600 1521.0400 1800.2400 ;
        RECT 1474.4400 1875.9200 1476.0400 1876.4000 ;
        RECT 1474.4400 1881.3600 1476.0400 1881.8400 ;
        RECT 1474.4400 1886.8000 1476.0400 1887.2800 ;
        RECT 1429.4400 1875.9200 1431.0400 1876.4000 ;
        RECT 1429.4400 1881.3600 1431.0400 1881.8400 ;
        RECT 1429.4400 1886.8000 1431.0400 1887.2800 ;
        RECT 1474.4400 1865.0400 1476.0400 1865.5200 ;
        RECT 1474.4400 1870.4800 1476.0400 1870.9600 ;
        RECT 1474.4400 1848.7200 1476.0400 1849.2000 ;
        RECT 1474.4400 1854.1600 1476.0400 1854.6400 ;
        RECT 1474.4400 1859.6000 1476.0400 1860.0800 ;
        RECT 1429.4400 1865.0400 1431.0400 1865.5200 ;
        RECT 1429.4400 1870.4800 1431.0400 1870.9600 ;
        RECT 1429.4400 1848.7200 1431.0400 1849.2000 ;
        RECT 1429.4400 1854.1600 1431.0400 1854.6400 ;
        RECT 1429.4400 1859.6000 1431.0400 1860.0800 ;
        RECT 1384.4400 1875.9200 1386.0400 1876.4000 ;
        RECT 1384.4400 1881.3600 1386.0400 1881.8400 ;
        RECT 1372.6800 1881.3600 1375.6800 1881.8400 ;
        RECT 1372.6800 1875.9200 1375.6800 1876.4000 ;
        RECT 1372.6800 1886.8000 1375.6800 1887.2800 ;
        RECT 1384.4400 1886.8000 1386.0400 1887.2800 ;
        RECT 1384.4400 1865.0400 1386.0400 1865.5200 ;
        RECT 1384.4400 1870.4800 1386.0400 1870.9600 ;
        RECT 1372.6800 1870.4800 1375.6800 1870.9600 ;
        RECT 1372.6800 1865.0400 1375.6800 1865.5200 ;
        RECT 1384.4400 1848.7200 1386.0400 1849.2000 ;
        RECT 1384.4400 1854.1600 1386.0400 1854.6400 ;
        RECT 1372.6800 1854.1600 1375.6800 1854.6400 ;
        RECT 1372.6800 1848.7200 1375.6800 1849.2000 ;
        RECT 1372.6800 1859.6000 1375.6800 1860.0800 ;
        RECT 1384.4400 1859.6000 1386.0400 1860.0800 ;
        RECT 1474.4400 1832.4000 1476.0400 1832.8800 ;
        RECT 1474.4400 1837.8400 1476.0400 1838.3200 ;
        RECT 1474.4400 1843.2800 1476.0400 1843.7600 ;
        RECT 1474.4400 1821.5200 1476.0400 1822.0000 ;
        RECT 1474.4400 1826.9600 1476.0400 1827.4400 ;
        RECT 1429.4400 1832.4000 1431.0400 1832.8800 ;
        RECT 1429.4400 1837.8400 1431.0400 1838.3200 ;
        RECT 1429.4400 1843.2800 1431.0400 1843.7600 ;
        RECT 1429.4400 1821.5200 1431.0400 1822.0000 ;
        RECT 1429.4400 1826.9600 1431.0400 1827.4400 ;
        RECT 1474.4400 1805.2000 1476.0400 1805.6800 ;
        RECT 1474.4400 1810.6400 1476.0400 1811.1200 ;
        RECT 1474.4400 1816.0800 1476.0400 1816.5600 ;
        RECT 1474.4400 1794.3200 1476.0400 1794.8000 ;
        RECT 1474.4400 1799.7600 1476.0400 1800.2400 ;
        RECT 1429.4400 1805.2000 1431.0400 1805.6800 ;
        RECT 1429.4400 1810.6400 1431.0400 1811.1200 ;
        RECT 1429.4400 1816.0800 1431.0400 1816.5600 ;
        RECT 1429.4400 1794.3200 1431.0400 1794.8000 ;
        RECT 1429.4400 1799.7600 1431.0400 1800.2400 ;
        RECT 1384.4400 1832.4000 1386.0400 1832.8800 ;
        RECT 1384.4400 1837.8400 1386.0400 1838.3200 ;
        RECT 1384.4400 1843.2800 1386.0400 1843.7600 ;
        RECT 1372.6800 1832.4000 1375.6800 1832.8800 ;
        RECT 1372.6800 1837.8400 1375.6800 1838.3200 ;
        RECT 1372.6800 1843.2800 1375.6800 1843.7600 ;
        RECT 1384.4400 1821.5200 1386.0400 1822.0000 ;
        RECT 1384.4400 1826.9600 1386.0400 1827.4400 ;
        RECT 1372.6800 1821.5200 1375.6800 1822.0000 ;
        RECT 1372.6800 1826.9600 1375.6800 1827.4400 ;
        RECT 1384.4400 1805.2000 1386.0400 1805.6800 ;
        RECT 1384.4400 1810.6400 1386.0400 1811.1200 ;
        RECT 1384.4400 1816.0800 1386.0400 1816.5600 ;
        RECT 1372.6800 1805.2000 1375.6800 1805.6800 ;
        RECT 1372.6800 1810.6400 1375.6800 1811.1200 ;
        RECT 1372.6800 1816.0800 1375.6800 1816.5600 ;
        RECT 1384.4400 1794.3200 1386.0400 1794.8000 ;
        RECT 1384.4400 1799.7600 1386.0400 1800.2400 ;
        RECT 1372.6800 1794.3200 1375.6800 1794.8000 ;
        RECT 1372.6800 1799.7600 1375.6800 1800.2400 ;
        RECT 1576.7800 1778.0000 1579.7800 1778.4800 ;
        RECT 1576.7800 1783.4400 1579.7800 1783.9200 ;
        RECT 1576.7800 1788.8800 1579.7800 1789.3600 ;
        RECT 1564.4400 1778.0000 1566.0400 1778.4800 ;
        RECT 1564.4400 1783.4400 1566.0400 1783.9200 ;
        RECT 1564.4400 1788.8800 1566.0400 1789.3600 ;
        RECT 1576.7800 1767.1200 1579.7800 1767.6000 ;
        RECT 1576.7800 1772.5600 1579.7800 1773.0400 ;
        RECT 1564.4400 1767.1200 1566.0400 1767.6000 ;
        RECT 1564.4400 1772.5600 1566.0400 1773.0400 ;
        RECT 1576.7800 1750.8000 1579.7800 1751.2800 ;
        RECT 1576.7800 1756.2400 1579.7800 1756.7200 ;
        RECT 1576.7800 1761.6800 1579.7800 1762.1600 ;
        RECT 1564.4400 1750.8000 1566.0400 1751.2800 ;
        RECT 1564.4400 1756.2400 1566.0400 1756.7200 ;
        RECT 1564.4400 1761.6800 1566.0400 1762.1600 ;
        RECT 1576.7800 1739.9200 1579.7800 1740.4000 ;
        RECT 1576.7800 1745.3600 1579.7800 1745.8400 ;
        RECT 1564.4400 1739.9200 1566.0400 1740.4000 ;
        RECT 1564.4400 1745.3600 1566.0400 1745.8400 ;
        RECT 1519.4400 1778.0000 1521.0400 1778.4800 ;
        RECT 1519.4400 1783.4400 1521.0400 1783.9200 ;
        RECT 1519.4400 1788.8800 1521.0400 1789.3600 ;
        RECT 1519.4400 1767.1200 1521.0400 1767.6000 ;
        RECT 1519.4400 1772.5600 1521.0400 1773.0400 ;
        RECT 1519.4400 1750.8000 1521.0400 1751.2800 ;
        RECT 1519.4400 1756.2400 1521.0400 1756.7200 ;
        RECT 1519.4400 1761.6800 1521.0400 1762.1600 ;
        RECT 1519.4400 1739.9200 1521.0400 1740.4000 ;
        RECT 1519.4400 1745.3600 1521.0400 1745.8400 ;
        RECT 1576.7800 1723.6000 1579.7800 1724.0800 ;
        RECT 1576.7800 1729.0400 1579.7800 1729.5200 ;
        RECT 1576.7800 1734.4800 1579.7800 1734.9600 ;
        RECT 1564.4400 1723.6000 1566.0400 1724.0800 ;
        RECT 1564.4400 1729.0400 1566.0400 1729.5200 ;
        RECT 1564.4400 1734.4800 1566.0400 1734.9600 ;
        RECT 1576.7800 1712.7200 1579.7800 1713.2000 ;
        RECT 1576.7800 1718.1600 1579.7800 1718.6400 ;
        RECT 1564.4400 1712.7200 1566.0400 1713.2000 ;
        RECT 1564.4400 1718.1600 1566.0400 1718.6400 ;
        RECT 1576.7800 1696.4000 1579.7800 1696.8800 ;
        RECT 1576.7800 1701.8400 1579.7800 1702.3200 ;
        RECT 1576.7800 1707.2800 1579.7800 1707.7600 ;
        RECT 1564.4400 1696.4000 1566.0400 1696.8800 ;
        RECT 1564.4400 1701.8400 1566.0400 1702.3200 ;
        RECT 1564.4400 1707.2800 1566.0400 1707.7600 ;
        RECT 1576.7800 1690.9600 1579.7800 1691.4400 ;
        RECT 1564.4400 1690.9600 1566.0400 1691.4400 ;
        RECT 1519.4400 1723.6000 1521.0400 1724.0800 ;
        RECT 1519.4400 1729.0400 1521.0400 1729.5200 ;
        RECT 1519.4400 1734.4800 1521.0400 1734.9600 ;
        RECT 1519.4400 1712.7200 1521.0400 1713.2000 ;
        RECT 1519.4400 1718.1600 1521.0400 1718.6400 ;
        RECT 1519.4400 1696.4000 1521.0400 1696.8800 ;
        RECT 1519.4400 1701.8400 1521.0400 1702.3200 ;
        RECT 1519.4400 1707.2800 1521.0400 1707.7600 ;
        RECT 1519.4400 1690.9600 1521.0400 1691.4400 ;
        RECT 1474.4400 1778.0000 1476.0400 1778.4800 ;
        RECT 1474.4400 1783.4400 1476.0400 1783.9200 ;
        RECT 1474.4400 1788.8800 1476.0400 1789.3600 ;
        RECT 1474.4400 1767.1200 1476.0400 1767.6000 ;
        RECT 1474.4400 1772.5600 1476.0400 1773.0400 ;
        RECT 1429.4400 1778.0000 1431.0400 1778.4800 ;
        RECT 1429.4400 1783.4400 1431.0400 1783.9200 ;
        RECT 1429.4400 1788.8800 1431.0400 1789.3600 ;
        RECT 1429.4400 1767.1200 1431.0400 1767.6000 ;
        RECT 1429.4400 1772.5600 1431.0400 1773.0400 ;
        RECT 1474.4400 1750.8000 1476.0400 1751.2800 ;
        RECT 1474.4400 1756.2400 1476.0400 1756.7200 ;
        RECT 1474.4400 1761.6800 1476.0400 1762.1600 ;
        RECT 1474.4400 1739.9200 1476.0400 1740.4000 ;
        RECT 1474.4400 1745.3600 1476.0400 1745.8400 ;
        RECT 1429.4400 1750.8000 1431.0400 1751.2800 ;
        RECT 1429.4400 1756.2400 1431.0400 1756.7200 ;
        RECT 1429.4400 1761.6800 1431.0400 1762.1600 ;
        RECT 1429.4400 1739.9200 1431.0400 1740.4000 ;
        RECT 1429.4400 1745.3600 1431.0400 1745.8400 ;
        RECT 1384.4400 1778.0000 1386.0400 1778.4800 ;
        RECT 1384.4400 1783.4400 1386.0400 1783.9200 ;
        RECT 1384.4400 1788.8800 1386.0400 1789.3600 ;
        RECT 1372.6800 1778.0000 1375.6800 1778.4800 ;
        RECT 1372.6800 1783.4400 1375.6800 1783.9200 ;
        RECT 1372.6800 1788.8800 1375.6800 1789.3600 ;
        RECT 1384.4400 1767.1200 1386.0400 1767.6000 ;
        RECT 1384.4400 1772.5600 1386.0400 1773.0400 ;
        RECT 1372.6800 1767.1200 1375.6800 1767.6000 ;
        RECT 1372.6800 1772.5600 1375.6800 1773.0400 ;
        RECT 1384.4400 1750.8000 1386.0400 1751.2800 ;
        RECT 1384.4400 1756.2400 1386.0400 1756.7200 ;
        RECT 1384.4400 1761.6800 1386.0400 1762.1600 ;
        RECT 1372.6800 1750.8000 1375.6800 1751.2800 ;
        RECT 1372.6800 1756.2400 1375.6800 1756.7200 ;
        RECT 1372.6800 1761.6800 1375.6800 1762.1600 ;
        RECT 1384.4400 1739.9200 1386.0400 1740.4000 ;
        RECT 1384.4400 1745.3600 1386.0400 1745.8400 ;
        RECT 1372.6800 1739.9200 1375.6800 1740.4000 ;
        RECT 1372.6800 1745.3600 1375.6800 1745.8400 ;
        RECT 1474.4400 1723.6000 1476.0400 1724.0800 ;
        RECT 1474.4400 1729.0400 1476.0400 1729.5200 ;
        RECT 1474.4400 1734.4800 1476.0400 1734.9600 ;
        RECT 1474.4400 1712.7200 1476.0400 1713.2000 ;
        RECT 1474.4400 1718.1600 1476.0400 1718.6400 ;
        RECT 1429.4400 1723.6000 1431.0400 1724.0800 ;
        RECT 1429.4400 1729.0400 1431.0400 1729.5200 ;
        RECT 1429.4400 1734.4800 1431.0400 1734.9600 ;
        RECT 1429.4400 1712.7200 1431.0400 1713.2000 ;
        RECT 1429.4400 1718.1600 1431.0400 1718.6400 ;
        RECT 1474.4400 1696.4000 1476.0400 1696.8800 ;
        RECT 1474.4400 1701.8400 1476.0400 1702.3200 ;
        RECT 1474.4400 1707.2800 1476.0400 1707.7600 ;
        RECT 1474.4400 1690.9600 1476.0400 1691.4400 ;
        RECT 1429.4400 1696.4000 1431.0400 1696.8800 ;
        RECT 1429.4400 1701.8400 1431.0400 1702.3200 ;
        RECT 1429.4400 1707.2800 1431.0400 1707.7600 ;
        RECT 1429.4400 1690.9600 1431.0400 1691.4400 ;
        RECT 1384.4400 1723.6000 1386.0400 1724.0800 ;
        RECT 1384.4400 1729.0400 1386.0400 1729.5200 ;
        RECT 1384.4400 1734.4800 1386.0400 1734.9600 ;
        RECT 1372.6800 1723.6000 1375.6800 1724.0800 ;
        RECT 1372.6800 1729.0400 1375.6800 1729.5200 ;
        RECT 1372.6800 1734.4800 1375.6800 1734.9600 ;
        RECT 1384.4400 1712.7200 1386.0400 1713.2000 ;
        RECT 1384.4400 1718.1600 1386.0400 1718.6400 ;
        RECT 1372.6800 1712.7200 1375.6800 1713.2000 ;
        RECT 1372.6800 1718.1600 1375.6800 1718.6400 ;
        RECT 1384.4400 1696.4000 1386.0400 1696.8800 ;
        RECT 1384.4400 1701.8400 1386.0400 1702.3200 ;
        RECT 1384.4400 1707.2800 1386.0400 1707.7600 ;
        RECT 1372.6800 1696.4000 1375.6800 1696.8800 ;
        RECT 1372.6800 1701.8400 1375.6800 1702.3200 ;
        RECT 1372.6800 1707.2800 1375.6800 1707.7600 ;
        RECT 1372.6800 1690.9600 1375.6800 1691.4400 ;
        RECT 1384.4400 1690.9600 1386.0400 1691.4400 ;
        RECT 1372.6800 1895.8700 1579.7800 1898.8700 ;
        RECT 1372.6800 1682.7700 1579.7800 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 1453.1300 1566.0400 1669.2300 ;
        RECT 1519.4400 1453.1300 1521.0400 1669.2300 ;
        RECT 1474.4400 1453.1300 1476.0400 1669.2300 ;
        RECT 1429.4400 1453.1300 1431.0400 1669.2300 ;
        RECT 1384.4400 1453.1300 1386.0400 1669.2300 ;
        RECT 1576.7800 1453.1300 1579.7800 1669.2300 ;
        RECT 1372.6800 1453.1300 1375.6800 1669.2300 ;
      LAYER met3 ;
        RECT 1576.7800 1646.2800 1579.7800 1646.7600 ;
        RECT 1576.7800 1651.7200 1579.7800 1652.2000 ;
        RECT 1564.4400 1646.2800 1566.0400 1646.7600 ;
        RECT 1564.4400 1651.7200 1566.0400 1652.2000 ;
        RECT 1576.7800 1657.1600 1579.7800 1657.6400 ;
        RECT 1564.4400 1657.1600 1566.0400 1657.6400 ;
        RECT 1576.7800 1635.4000 1579.7800 1635.8800 ;
        RECT 1576.7800 1640.8400 1579.7800 1641.3200 ;
        RECT 1564.4400 1635.4000 1566.0400 1635.8800 ;
        RECT 1564.4400 1640.8400 1566.0400 1641.3200 ;
        RECT 1576.7800 1619.0800 1579.7800 1619.5600 ;
        RECT 1576.7800 1624.5200 1579.7800 1625.0000 ;
        RECT 1564.4400 1619.0800 1566.0400 1619.5600 ;
        RECT 1564.4400 1624.5200 1566.0400 1625.0000 ;
        RECT 1576.7800 1629.9600 1579.7800 1630.4400 ;
        RECT 1564.4400 1629.9600 1566.0400 1630.4400 ;
        RECT 1519.4400 1646.2800 1521.0400 1646.7600 ;
        RECT 1519.4400 1651.7200 1521.0400 1652.2000 ;
        RECT 1519.4400 1657.1600 1521.0400 1657.6400 ;
        RECT 1519.4400 1635.4000 1521.0400 1635.8800 ;
        RECT 1519.4400 1640.8400 1521.0400 1641.3200 ;
        RECT 1519.4400 1619.0800 1521.0400 1619.5600 ;
        RECT 1519.4400 1624.5200 1521.0400 1625.0000 ;
        RECT 1519.4400 1629.9600 1521.0400 1630.4400 ;
        RECT 1576.7800 1602.7600 1579.7800 1603.2400 ;
        RECT 1576.7800 1608.2000 1579.7800 1608.6800 ;
        RECT 1576.7800 1613.6400 1579.7800 1614.1200 ;
        RECT 1564.4400 1602.7600 1566.0400 1603.2400 ;
        RECT 1564.4400 1608.2000 1566.0400 1608.6800 ;
        RECT 1564.4400 1613.6400 1566.0400 1614.1200 ;
        RECT 1576.7800 1591.8800 1579.7800 1592.3600 ;
        RECT 1576.7800 1597.3200 1579.7800 1597.8000 ;
        RECT 1564.4400 1591.8800 1566.0400 1592.3600 ;
        RECT 1564.4400 1597.3200 1566.0400 1597.8000 ;
        RECT 1576.7800 1575.5600 1579.7800 1576.0400 ;
        RECT 1576.7800 1581.0000 1579.7800 1581.4800 ;
        RECT 1576.7800 1586.4400 1579.7800 1586.9200 ;
        RECT 1564.4400 1575.5600 1566.0400 1576.0400 ;
        RECT 1564.4400 1581.0000 1566.0400 1581.4800 ;
        RECT 1564.4400 1586.4400 1566.0400 1586.9200 ;
        RECT 1576.7800 1564.6800 1579.7800 1565.1600 ;
        RECT 1576.7800 1570.1200 1579.7800 1570.6000 ;
        RECT 1564.4400 1564.6800 1566.0400 1565.1600 ;
        RECT 1564.4400 1570.1200 1566.0400 1570.6000 ;
        RECT 1519.4400 1602.7600 1521.0400 1603.2400 ;
        RECT 1519.4400 1608.2000 1521.0400 1608.6800 ;
        RECT 1519.4400 1613.6400 1521.0400 1614.1200 ;
        RECT 1519.4400 1591.8800 1521.0400 1592.3600 ;
        RECT 1519.4400 1597.3200 1521.0400 1597.8000 ;
        RECT 1519.4400 1575.5600 1521.0400 1576.0400 ;
        RECT 1519.4400 1581.0000 1521.0400 1581.4800 ;
        RECT 1519.4400 1586.4400 1521.0400 1586.9200 ;
        RECT 1519.4400 1564.6800 1521.0400 1565.1600 ;
        RECT 1519.4400 1570.1200 1521.0400 1570.6000 ;
        RECT 1474.4400 1646.2800 1476.0400 1646.7600 ;
        RECT 1474.4400 1651.7200 1476.0400 1652.2000 ;
        RECT 1474.4400 1657.1600 1476.0400 1657.6400 ;
        RECT 1429.4400 1646.2800 1431.0400 1646.7600 ;
        RECT 1429.4400 1651.7200 1431.0400 1652.2000 ;
        RECT 1429.4400 1657.1600 1431.0400 1657.6400 ;
        RECT 1474.4400 1635.4000 1476.0400 1635.8800 ;
        RECT 1474.4400 1640.8400 1476.0400 1641.3200 ;
        RECT 1474.4400 1619.0800 1476.0400 1619.5600 ;
        RECT 1474.4400 1624.5200 1476.0400 1625.0000 ;
        RECT 1474.4400 1629.9600 1476.0400 1630.4400 ;
        RECT 1429.4400 1635.4000 1431.0400 1635.8800 ;
        RECT 1429.4400 1640.8400 1431.0400 1641.3200 ;
        RECT 1429.4400 1619.0800 1431.0400 1619.5600 ;
        RECT 1429.4400 1624.5200 1431.0400 1625.0000 ;
        RECT 1429.4400 1629.9600 1431.0400 1630.4400 ;
        RECT 1384.4400 1646.2800 1386.0400 1646.7600 ;
        RECT 1384.4400 1651.7200 1386.0400 1652.2000 ;
        RECT 1372.6800 1651.7200 1375.6800 1652.2000 ;
        RECT 1372.6800 1646.2800 1375.6800 1646.7600 ;
        RECT 1372.6800 1657.1600 1375.6800 1657.6400 ;
        RECT 1384.4400 1657.1600 1386.0400 1657.6400 ;
        RECT 1384.4400 1635.4000 1386.0400 1635.8800 ;
        RECT 1384.4400 1640.8400 1386.0400 1641.3200 ;
        RECT 1372.6800 1640.8400 1375.6800 1641.3200 ;
        RECT 1372.6800 1635.4000 1375.6800 1635.8800 ;
        RECT 1384.4400 1619.0800 1386.0400 1619.5600 ;
        RECT 1384.4400 1624.5200 1386.0400 1625.0000 ;
        RECT 1372.6800 1624.5200 1375.6800 1625.0000 ;
        RECT 1372.6800 1619.0800 1375.6800 1619.5600 ;
        RECT 1372.6800 1629.9600 1375.6800 1630.4400 ;
        RECT 1384.4400 1629.9600 1386.0400 1630.4400 ;
        RECT 1474.4400 1602.7600 1476.0400 1603.2400 ;
        RECT 1474.4400 1608.2000 1476.0400 1608.6800 ;
        RECT 1474.4400 1613.6400 1476.0400 1614.1200 ;
        RECT 1474.4400 1591.8800 1476.0400 1592.3600 ;
        RECT 1474.4400 1597.3200 1476.0400 1597.8000 ;
        RECT 1429.4400 1602.7600 1431.0400 1603.2400 ;
        RECT 1429.4400 1608.2000 1431.0400 1608.6800 ;
        RECT 1429.4400 1613.6400 1431.0400 1614.1200 ;
        RECT 1429.4400 1591.8800 1431.0400 1592.3600 ;
        RECT 1429.4400 1597.3200 1431.0400 1597.8000 ;
        RECT 1474.4400 1575.5600 1476.0400 1576.0400 ;
        RECT 1474.4400 1581.0000 1476.0400 1581.4800 ;
        RECT 1474.4400 1586.4400 1476.0400 1586.9200 ;
        RECT 1474.4400 1564.6800 1476.0400 1565.1600 ;
        RECT 1474.4400 1570.1200 1476.0400 1570.6000 ;
        RECT 1429.4400 1575.5600 1431.0400 1576.0400 ;
        RECT 1429.4400 1581.0000 1431.0400 1581.4800 ;
        RECT 1429.4400 1586.4400 1431.0400 1586.9200 ;
        RECT 1429.4400 1564.6800 1431.0400 1565.1600 ;
        RECT 1429.4400 1570.1200 1431.0400 1570.6000 ;
        RECT 1384.4400 1602.7600 1386.0400 1603.2400 ;
        RECT 1384.4400 1608.2000 1386.0400 1608.6800 ;
        RECT 1384.4400 1613.6400 1386.0400 1614.1200 ;
        RECT 1372.6800 1602.7600 1375.6800 1603.2400 ;
        RECT 1372.6800 1608.2000 1375.6800 1608.6800 ;
        RECT 1372.6800 1613.6400 1375.6800 1614.1200 ;
        RECT 1384.4400 1591.8800 1386.0400 1592.3600 ;
        RECT 1384.4400 1597.3200 1386.0400 1597.8000 ;
        RECT 1372.6800 1591.8800 1375.6800 1592.3600 ;
        RECT 1372.6800 1597.3200 1375.6800 1597.8000 ;
        RECT 1384.4400 1575.5600 1386.0400 1576.0400 ;
        RECT 1384.4400 1581.0000 1386.0400 1581.4800 ;
        RECT 1384.4400 1586.4400 1386.0400 1586.9200 ;
        RECT 1372.6800 1575.5600 1375.6800 1576.0400 ;
        RECT 1372.6800 1581.0000 1375.6800 1581.4800 ;
        RECT 1372.6800 1586.4400 1375.6800 1586.9200 ;
        RECT 1384.4400 1564.6800 1386.0400 1565.1600 ;
        RECT 1384.4400 1570.1200 1386.0400 1570.6000 ;
        RECT 1372.6800 1564.6800 1375.6800 1565.1600 ;
        RECT 1372.6800 1570.1200 1375.6800 1570.6000 ;
        RECT 1576.7800 1548.3600 1579.7800 1548.8400 ;
        RECT 1576.7800 1553.8000 1579.7800 1554.2800 ;
        RECT 1576.7800 1559.2400 1579.7800 1559.7200 ;
        RECT 1564.4400 1548.3600 1566.0400 1548.8400 ;
        RECT 1564.4400 1553.8000 1566.0400 1554.2800 ;
        RECT 1564.4400 1559.2400 1566.0400 1559.7200 ;
        RECT 1576.7800 1537.4800 1579.7800 1537.9600 ;
        RECT 1576.7800 1542.9200 1579.7800 1543.4000 ;
        RECT 1564.4400 1537.4800 1566.0400 1537.9600 ;
        RECT 1564.4400 1542.9200 1566.0400 1543.4000 ;
        RECT 1576.7800 1521.1600 1579.7800 1521.6400 ;
        RECT 1576.7800 1526.6000 1579.7800 1527.0800 ;
        RECT 1576.7800 1532.0400 1579.7800 1532.5200 ;
        RECT 1564.4400 1521.1600 1566.0400 1521.6400 ;
        RECT 1564.4400 1526.6000 1566.0400 1527.0800 ;
        RECT 1564.4400 1532.0400 1566.0400 1532.5200 ;
        RECT 1576.7800 1510.2800 1579.7800 1510.7600 ;
        RECT 1576.7800 1515.7200 1579.7800 1516.2000 ;
        RECT 1564.4400 1510.2800 1566.0400 1510.7600 ;
        RECT 1564.4400 1515.7200 1566.0400 1516.2000 ;
        RECT 1519.4400 1548.3600 1521.0400 1548.8400 ;
        RECT 1519.4400 1553.8000 1521.0400 1554.2800 ;
        RECT 1519.4400 1559.2400 1521.0400 1559.7200 ;
        RECT 1519.4400 1537.4800 1521.0400 1537.9600 ;
        RECT 1519.4400 1542.9200 1521.0400 1543.4000 ;
        RECT 1519.4400 1521.1600 1521.0400 1521.6400 ;
        RECT 1519.4400 1526.6000 1521.0400 1527.0800 ;
        RECT 1519.4400 1532.0400 1521.0400 1532.5200 ;
        RECT 1519.4400 1510.2800 1521.0400 1510.7600 ;
        RECT 1519.4400 1515.7200 1521.0400 1516.2000 ;
        RECT 1576.7800 1493.9600 1579.7800 1494.4400 ;
        RECT 1576.7800 1499.4000 1579.7800 1499.8800 ;
        RECT 1576.7800 1504.8400 1579.7800 1505.3200 ;
        RECT 1564.4400 1493.9600 1566.0400 1494.4400 ;
        RECT 1564.4400 1499.4000 1566.0400 1499.8800 ;
        RECT 1564.4400 1504.8400 1566.0400 1505.3200 ;
        RECT 1576.7800 1483.0800 1579.7800 1483.5600 ;
        RECT 1576.7800 1488.5200 1579.7800 1489.0000 ;
        RECT 1564.4400 1483.0800 1566.0400 1483.5600 ;
        RECT 1564.4400 1488.5200 1566.0400 1489.0000 ;
        RECT 1576.7800 1466.7600 1579.7800 1467.2400 ;
        RECT 1576.7800 1472.2000 1579.7800 1472.6800 ;
        RECT 1576.7800 1477.6400 1579.7800 1478.1200 ;
        RECT 1564.4400 1466.7600 1566.0400 1467.2400 ;
        RECT 1564.4400 1472.2000 1566.0400 1472.6800 ;
        RECT 1564.4400 1477.6400 1566.0400 1478.1200 ;
        RECT 1576.7800 1461.3200 1579.7800 1461.8000 ;
        RECT 1564.4400 1461.3200 1566.0400 1461.8000 ;
        RECT 1519.4400 1493.9600 1521.0400 1494.4400 ;
        RECT 1519.4400 1499.4000 1521.0400 1499.8800 ;
        RECT 1519.4400 1504.8400 1521.0400 1505.3200 ;
        RECT 1519.4400 1483.0800 1521.0400 1483.5600 ;
        RECT 1519.4400 1488.5200 1521.0400 1489.0000 ;
        RECT 1519.4400 1466.7600 1521.0400 1467.2400 ;
        RECT 1519.4400 1472.2000 1521.0400 1472.6800 ;
        RECT 1519.4400 1477.6400 1521.0400 1478.1200 ;
        RECT 1519.4400 1461.3200 1521.0400 1461.8000 ;
        RECT 1474.4400 1548.3600 1476.0400 1548.8400 ;
        RECT 1474.4400 1553.8000 1476.0400 1554.2800 ;
        RECT 1474.4400 1559.2400 1476.0400 1559.7200 ;
        RECT 1474.4400 1537.4800 1476.0400 1537.9600 ;
        RECT 1474.4400 1542.9200 1476.0400 1543.4000 ;
        RECT 1429.4400 1548.3600 1431.0400 1548.8400 ;
        RECT 1429.4400 1553.8000 1431.0400 1554.2800 ;
        RECT 1429.4400 1559.2400 1431.0400 1559.7200 ;
        RECT 1429.4400 1537.4800 1431.0400 1537.9600 ;
        RECT 1429.4400 1542.9200 1431.0400 1543.4000 ;
        RECT 1474.4400 1521.1600 1476.0400 1521.6400 ;
        RECT 1474.4400 1526.6000 1476.0400 1527.0800 ;
        RECT 1474.4400 1532.0400 1476.0400 1532.5200 ;
        RECT 1474.4400 1510.2800 1476.0400 1510.7600 ;
        RECT 1474.4400 1515.7200 1476.0400 1516.2000 ;
        RECT 1429.4400 1521.1600 1431.0400 1521.6400 ;
        RECT 1429.4400 1526.6000 1431.0400 1527.0800 ;
        RECT 1429.4400 1532.0400 1431.0400 1532.5200 ;
        RECT 1429.4400 1510.2800 1431.0400 1510.7600 ;
        RECT 1429.4400 1515.7200 1431.0400 1516.2000 ;
        RECT 1384.4400 1548.3600 1386.0400 1548.8400 ;
        RECT 1384.4400 1553.8000 1386.0400 1554.2800 ;
        RECT 1384.4400 1559.2400 1386.0400 1559.7200 ;
        RECT 1372.6800 1548.3600 1375.6800 1548.8400 ;
        RECT 1372.6800 1553.8000 1375.6800 1554.2800 ;
        RECT 1372.6800 1559.2400 1375.6800 1559.7200 ;
        RECT 1384.4400 1537.4800 1386.0400 1537.9600 ;
        RECT 1384.4400 1542.9200 1386.0400 1543.4000 ;
        RECT 1372.6800 1537.4800 1375.6800 1537.9600 ;
        RECT 1372.6800 1542.9200 1375.6800 1543.4000 ;
        RECT 1384.4400 1521.1600 1386.0400 1521.6400 ;
        RECT 1384.4400 1526.6000 1386.0400 1527.0800 ;
        RECT 1384.4400 1532.0400 1386.0400 1532.5200 ;
        RECT 1372.6800 1521.1600 1375.6800 1521.6400 ;
        RECT 1372.6800 1526.6000 1375.6800 1527.0800 ;
        RECT 1372.6800 1532.0400 1375.6800 1532.5200 ;
        RECT 1384.4400 1510.2800 1386.0400 1510.7600 ;
        RECT 1384.4400 1515.7200 1386.0400 1516.2000 ;
        RECT 1372.6800 1510.2800 1375.6800 1510.7600 ;
        RECT 1372.6800 1515.7200 1375.6800 1516.2000 ;
        RECT 1474.4400 1493.9600 1476.0400 1494.4400 ;
        RECT 1474.4400 1499.4000 1476.0400 1499.8800 ;
        RECT 1474.4400 1504.8400 1476.0400 1505.3200 ;
        RECT 1474.4400 1483.0800 1476.0400 1483.5600 ;
        RECT 1474.4400 1488.5200 1476.0400 1489.0000 ;
        RECT 1429.4400 1493.9600 1431.0400 1494.4400 ;
        RECT 1429.4400 1499.4000 1431.0400 1499.8800 ;
        RECT 1429.4400 1504.8400 1431.0400 1505.3200 ;
        RECT 1429.4400 1483.0800 1431.0400 1483.5600 ;
        RECT 1429.4400 1488.5200 1431.0400 1489.0000 ;
        RECT 1474.4400 1466.7600 1476.0400 1467.2400 ;
        RECT 1474.4400 1472.2000 1476.0400 1472.6800 ;
        RECT 1474.4400 1477.6400 1476.0400 1478.1200 ;
        RECT 1474.4400 1461.3200 1476.0400 1461.8000 ;
        RECT 1429.4400 1466.7600 1431.0400 1467.2400 ;
        RECT 1429.4400 1472.2000 1431.0400 1472.6800 ;
        RECT 1429.4400 1477.6400 1431.0400 1478.1200 ;
        RECT 1429.4400 1461.3200 1431.0400 1461.8000 ;
        RECT 1384.4400 1493.9600 1386.0400 1494.4400 ;
        RECT 1384.4400 1499.4000 1386.0400 1499.8800 ;
        RECT 1384.4400 1504.8400 1386.0400 1505.3200 ;
        RECT 1372.6800 1493.9600 1375.6800 1494.4400 ;
        RECT 1372.6800 1499.4000 1375.6800 1499.8800 ;
        RECT 1372.6800 1504.8400 1375.6800 1505.3200 ;
        RECT 1384.4400 1483.0800 1386.0400 1483.5600 ;
        RECT 1384.4400 1488.5200 1386.0400 1489.0000 ;
        RECT 1372.6800 1483.0800 1375.6800 1483.5600 ;
        RECT 1372.6800 1488.5200 1375.6800 1489.0000 ;
        RECT 1384.4400 1466.7600 1386.0400 1467.2400 ;
        RECT 1384.4400 1472.2000 1386.0400 1472.6800 ;
        RECT 1384.4400 1477.6400 1386.0400 1478.1200 ;
        RECT 1372.6800 1466.7600 1375.6800 1467.2400 ;
        RECT 1372.6800 1472.2000 1375.6800 1472.6800 ;
        RECT 1372.6800 1477.6400 1375.6800 1478.1200 ;
        RECT 1372.6800 1461.3200 1375.6800 1461.8000 ;
        RECT 1384.4400 1461.3200 1386.0400 1461.8000 ;
        RECT 1372.6800 1666.2300 1579.7800 1669.2300 ;
        RECT 1372.6800 1453.1300 1579.7800 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 1223.4900 1566.0400 1439.5900 ;
        RECT 1519.4400 1223.4900 1521.0400 1439.5900 ;
        RECT 1474.4400 1223.4900 1476.0400 1439.5900 ;
        RECT 1429.4400 1223.4900 1431.0400 1439.5900 ;
        RECT 1384.4400 1223.4900 1386.0400 1439.5900 ;
        RECT 1576.7800 1223.4900 1579.7800 1439.5900 ;
        RECT 1372.6800 1223.4900 1375.6800 1439.5900 ;
      LAYER met3 ;
        RECT 1576.7800 1416.6400 1579.7800 1417.1200 ;
        RECT 1576.7800 1422.0800 1579.7800 1422.5600 ;
        RECT 1564.4400 1416.6400 1566.0400 1417.1200 ;
        RECT 1564.4400 1422.0800 1566.0400 1422.5600 ;
        RECT 1576.7800 1427.5200 1579.7800 1428.0000 ;
        RECT 1564.4400 1427.5200 1566.0400 1428.0000 ;
        RECT 1576.7800 1405.7600 1579.7800 1406.2400 ;
        RECT 1576.7800 1411.2000 1579.7800 1411.6800 ;
        RECT 1564.4400 1405.7600 1566.0400 1406.2400 ;
        RECT 1564.4400 1411.2000 1566.0400 1411.6800 ;
        RECT 1576.7800 1389.4400 1579.7800 1389.9200 ;
        RECT 1576.7800 1394.8800 1579.7800 1395.3600 ;
        RECT 1564.4400 1389.4400 1566.0400 1389.9200 ;
        RECT 1564.4400 1394.8800 1566.0400 1395.3600 ;
        RECT 1576.7800 1400.3200 1579.7800 1400.8000 ;
        RECT 1564.4400 1400.3200 1566.0400 1400.8000 ;
        RECT 1519.4400 1416.6400 1521.0400 1417.1200 ;
        RECT 1519.4400 1422.0800 1521.0400 1422.5600 ;
        RECT 1519.4400 1427.5200 1521.0400 1428.0000 ;
        RECT 1519.4400 1405.7600 1521.0400 1406.2400 ;
        RECT 1519.4400 1411.2000 1521.0400 1411.6800 ;
        RECT 1519.4400 1389.4400 1521.0400 1389.9200 ;
        RECT 1519.4400 1394.8800 1521.0400 1395.3600 ;
        RECT 1519.4400 1400.3200 1521.0400 1400.8000 ;
        RECT 1576.7800 1373.1200 1579.7800 1373.6000 ;
        RECT 1576.7800 1378.5600 1579.7800 1379.0400 ;
        RECT 1576.7800 1384.0000 1579.7800 1384.4800 ;
        RECT 1564.4400 1373.1200 1566.0400 1373.6000 ;
        RECT 1564.4400 1378.5600 1566.0400 1379.0400 ;
        RECT 1564.4400 1384.0000 1566.0400 1384.4800 ;
        RECT 1576.7800 1362.2400 1579.7800 1362.7200 ;
        RECT 1576.7800 1367.6800 1579.7800 1368.1600 ;
        RECT 1564.4400 1362.2400 1566.0400 1362.7200 ;
        RECT 1564.4400 1367.6800 1566.0400 1368.1600 ;
        RECT 1576.7800 1345.9200 1579.7800 1346.4000 ;
        RECT 1576.7800 1351.3600 1579.7800 1351.8400 ;
        RECT 1576.7800 1356.8000 1579.7800 1357.2800 ;
        RECT 1564.4400 1345.9200 1566.0400 1346.4000 ;
        RECT 1564.4400 1351.3600 1566.0400 1351.8400 ;
        RECT 1564.4400 1356.8000 1566.0400 1357.2800 ;
        RECT 1576.7800 1335.0400 1579.7800 1335.5200 ;
        RECT 1576.7800 1340.4800 1579.7800 1340.9600 ;
        RECT 1564.4400 1335.0400 1566.0400 1335.5200 ;
        RECT 1564.4400 1340.4800 1566.0400 1340.9600 ;
        RECT 1519.4400 1373.1200 1521.0400 1373.6000 ;
        RECT 1519.4400 1378.5600 1521.0400 1379.0400 ;
        RECT 1519.4400 1384.0000 1521.0400 1384.4800 ;
        RECT 1519.4400 1362.2400 1521.0400 1362.7200 ;
        RECT 1519.4400 1367.6800 1521.0400 1368.1600 ;
        RECT 1519.4400 1345.9200 1521.0400 1346.4000 ;
        RECT 1519.4400 1351.3600 1521.0400 1351.8400 ;
        RECT 1519.4400 1356.8000 1521.0400 1357.2800 ;
        RECT 1519.4400 1335.0400 1521.0400 1335.5200 ;
        RECT 1519.4400 1340.4800 1521.0400 1340.9600 ;
        RECT 1474.4400 1416.6400 1476.0400 1417.1200 ;
        RECT 1474.4400 1422.0800 1476.0400 1422.5600 ;
        RECT 1474.4400 1427.5200 1476.0400 1428.0000 ;
        RECT 1429.4400 1416.6400 1431.0400 1417.1200 ;
        RECT 1429.4400 1422.0800 1431.0400 1422.5600 ;
        RECT 1429.4400 1427.5200 1431.0400 1428.0000 ;
        RECT 1474.4400 1405.7600 1476.0400 1406.2400 ;
        RECT 1474.4400 1411.2000 1476.0400 1411.6800 ;
        RECT 1474.4400 1389.4400 1476.0400 1389.9200 ;
        RECT 1474.4400 1394.8800 1476.0400 1395.3600 ;
        RECT 1474.4400 1400.3200 1476.0400 1400.8000 ;
        RECT 1429.4400 1405.7600 1431.0400 1406.2400 ;
        RECT 1429.4400 1411.2000 1431.0400 1411.6800 ;
        RECT 1429.4400 1389.4400 1431.0400 1389.9200 ;
        RECT 1429.4400 1394.8800 1431.0400 1395.3600 ;
        RECT 1429.4400 1400.3200 1431.0400 1400.8000 ;
        RECT 1384.4400 1416.6400 1386.0400 1417.1200 ;
        RECT 1384.4400 1422.0800 1386.0400 1422.5600 ;
        RECT 1372.6800 1422.0800 1375.6800 1422.5600 ;
        RECT 1372.6800 1416.6400 1375.6800 1417.1200 ;
        RECT 1372.6800 1427.5200 1375.6800 1428.0000 ;
        RECT 1384.4400 1427.5200 1386.0400 1428.0000 ;
        RECT 1384.4400 1405.7600 1386.0400 1406.2400 ;
        RECT 1384.4400 1411.2000 1386.0400 1411.6800 ;
        RECT 1372.6800 1411.2000 1375.6800 1411.6800 ;
        RECT 1372.6800 1405.7600 1375.6800 1406.2400 ;
        RECT 1384.4400 1389.4400 1386.0400 1389.9200 ;
        RECT 1384.4400 1394.8800 1386.0400 1395.3600 ;
        RECT 1372.6800 1394.8800 1375.6800 1395.3600 ;
        RECT 1372.6800 1389.4400 1375.6800 1389.9200 ;
        RECT 1372.6800 1400.3200 1375.6800 1400.8000 ;
        RECT 1384.4400 1400.3200 1386.0400 1400.8000 ;
        RECT 1474.4400 1373.1200 1476.0400 1373.6000 ;
        RECT 1474.4400 1378.5600 1476.0400 1379.0400 ;
        RECT 1474.4400 1384.0000 1476.0400 1384.4800 ;
        RECT 1474.4400 1362.2400 1476.0400 1362.7200 ;
        RECT 1474.4400 1367.6800 1476.0400 1368.1600 ;
        RECT 1429.4400 1373.1200 1431.0400 1373.6000 ;
        RECT 1429.4400 1378.5600 1431.0400 1379.0400 ;
        RECT 1429.4400 1384.0000 1431.0400 1384.4800 ;
        RECT 1429.4400 1362.2400 1431.0400 1362.7200 ;
        RECT 1429.4400 1367.6800 1431.0400 1368.1600 ;
        RECT 1474.4400 1345.9200 1476.0400 1346.4000 ;
        RECT 1474.4400 1351.3600 1476.0400 1351.8400 ;
        RECT 1474.4400 1356.8000 1476.0400 1357.2800 ;
        RECT 1474.4400 1335.0400 1476.0400 1335.5200 ;
        RECT 1474.4400 1340.4800 1476.0400 1340.9600 ;
        RECT 1429.4400 1345.9200 1431.0400 1346.4000 ;
        RECT 1429.4400 1351.3600 1431.0400 1351.8400 ;
        RECT 1429.4400 1356.8000 1431.0400 1357.2800 ;
        RECT 1429.4400 1335.0400 1431.0400 1335.5200 ;
        RECT 1429.4400 1340.4800 1431.0400 1340.9600 ;
        RECT 1384.4400 1373.1200 1386.0400 1373.6000 ;
        RECT 1384.4400 1378.5600 1386.0400 1379.0400 ;
        RECT 1384.4400 1384.0000 1386.0400 1384.4800 ;
        RECT 1372.6800 1373.1200 1375.6800 1373.6000 ;
        RECT 1372.6800 1378.5600 1375.6800 1379.0400 ;
        RECT 1372.6800 1384.0000 1375.6800 1384.4800 ;
        RECT 1384.4400 1362.2400 1386.0400 1362.7200 ;
        RECT 1384.4400 1367.6800 1386.0400 1368.1600 ;
        RECT 1372.6800 1362.2400 1375.6800 1362.7200 ;
        RECT 1372.6800 1367.6800 1375.6800 1368.1600 ;
        RECT 1384.4400 1345.9200 1386.0400 1346.4000 ;
        RECT 1384.4400 1351.3600 1386.0400 1351.8400 ;
        RECT 1384.4400 1356.8000 1386.0400 1357.2800 ;
        RECT 1372.6800 1345.9200 1375.6800 1346.4000 ;
        RECT 1372.6800 1351.3600 1375.6800 1351.8400 ;
        RECT 1372.6800 1356.8000 1375.6800 1357.2800 ;
        RECT 1384.4400 1335.0400 1386.0400 1335.5200 ;
        RECT 1384.4400 1340.4800 1386.0400 1340.9600 ;
        RECT 1372.6800 1335.0400 1375.6800 1335.5200 ;
        RECT 1372.6800 1340.4800 1375.6800 1340.9600 ;
        RECT 1576.7800 1318.7200 1579.7800 1319.2000 ;
        RECT 1576.7800 1324.1600 1579.7800 1324.6400 ;
        RECT 1576.7800 1329.6000 1579.7800 1330.0800 ;
        RECT 1564.4400 1318.7200 1566.0400 1319.2000 ;
        RECT 1564.4400 1324.1600 1566.0400 1324.6400 ;
        RECT 1564.4400 1329.6000 1566.0400 1330.0800 ;
        RECT 1576.7800 1307.8400 1579.7800 1308.3200 ;
        RECT 1576.7800 1313.2800 1579.7800 1313.7600 ;
        RECT 1564.4400 1307.8400 1566.0400 1308.3200 ;
        RECT 1564.4400 1313.2800 1566.0400 1313.7600 ;
        RECT 1576.7800 1291.5200 1579.7800 1292.0000 ;
        RECT 1576.7800 1296.9600 1579.7800 1297.4400 ;
        RECT 1576.7800 1302.4000 1579.7800 1302.8800 ;
        RECT 1564.4400 1291.5200 1566.0400 1292.0000 ;
        RECT 1564.4400 1296.9600 1566.0400 1297.4400 ;
        RECT 1564.4400 1302.4000 1566.0400 1302.8800 ;
        RECT 1576.7800 1280.6400 1579.7800 1281.1200 ;
        RECT 1576.7800 1286.0800 1579.7800 1286.5600 ;
        RECT 1564.4400 1280.6400 1566.0400 1281.1200 ;
        RECT 1564.4400 1286.0800 1566.0400 1286.5600 ;
        RECT 1519.4400 1318.7200 1521.0400 1319.2000 ;
        RECT 1519.4400 1324.1600 1521.0400 1324.6400 ;
        RECT 1519.4400 1329.6000 1521.0400 1330.0800 ;
        RECT 1519.4400 1307.8400 1521.0400 1308.3200 ;
        RECT 1519.4400 1313.2800 1521.0400 1313.7600 ;
        RECT 1519.4400 1291.5200 1521.0400 1292.0000 ;
        RECT 1519.4400 1296.9600 1521.0400 1297.4400 ;
        RECT 1519.4400 1302.4000 1521.0400 1302.8800 ;
        RECT 1519.4400 1280.6400 1521.0400 1281.1200 ;
        RECT 1519.4400 1286.0800 1521.0400 1286.5600 ;
        RECT 1576.7800 1264.3200 1579.7800 1264.8000 ;
        RECT 1576.7800 1269.7600 1579.7800 1270.2400 ;
        RECT 1576.7800 1275.2000 1579.7800 1275.6800 ;
        RECT 1564.4400 1264.3200 1566.0400 1264.8000 ;
        RECT 1564.4400 1269.7600 1566.0400 1270.2400 ;
        RECT 1564.4400 1275.2000 1566.0400 1275.6800 ;
        RECT 1576.7800 1253.4400 1579.7800 1253.9200 ;
        RECT 1576.7800 1258.8800 1579.7800 1259.3600 ;
        RECT 1564.4400 1253.4400 1566.0400 1253.9200 ;
        RECT 1564.4400 1258.8800 1566.0400 1259.3600 ;
        RECT 1576.7800 1237.1200 1579.7800 1237.6000 ;
        RECT 1576.7800 1242.5600 1579.7800 1243.0400 ;
        RECT 1576.7800 1248.0000 1579.7800 1248.4800 ;
        RECT 1564.4400 1237.1200 1566.0400 1237.6000 ;
        RECT 1564.4400 1242.5600 1566.0400 1243.0400 ;
        RECT 1564.4400 1248.0000 1566.0400 1248.4800 ;
        RECT 1576.7800 1231.6800 1579.7800 1232.1600 ;
        RECT 1564.4400 1231.6800 1566.0400 1232.1600 ;
        RECT 1519.4400 1264.3200 1521.0400 1264.8000 ;
        RECT 1519.4400 1269.7600 1521.0400 1270.2400 ;
        RECT 1519.4400 1275.2000 1521.0400 1275.6800 ;
        RECT 1519.4400 1253.4400 1521.0400 1253.9200 ;
        RECT 1519.4400 1258.8800 1521.0400 1259.3600 ;
        RECT 1519.4400 1237.1200 1521.0400 1237.6000 ;
        RECT 1519.4400 1242.5600 1521.0400 1243.0400 ;
        RECT 1519.4400 1248.0000 1521.0400 1248.4800 ;
        RECT 1519.4400 1231.6800 1521.0400 1232.1600 ;
        RECT 1474.4400 1318.7200 1476.0400 1319.2000 ;
        RECT 1474.4400 1324.1600 1476.0400 1324.6400 ;
        RECT 1474.4400 1329.6000 1476.0400 1330.0800 ;
        RECT 1474.4400 1307.8400 1476.0400 1308.3200 ;
        RECT 1474.4400 1313.2800 1476.0400 1313.7600 ;
        RECT 1429.4400 1318.7200 1431.0400 1319.2000 ;
        RECT 1429.4400 1324.1600 1431.0400 1324.6400 ;
        RECT 1429.4400 1329.6000 1431.0400 1330.0800 ;
        RECT 1429.4400 1307.8400 1431.0400 1308.3200 ;
        RECT 1429.4400 1313.2800 1431.0400 1313.7600 ;
        RECT 1474.4400 1291.5200 1476.0400 1292.0000 ;
        RECT 1474.4400 1296.9600 1476.0400 1297.4400 ;
        RECT 1474.4400 1302.4000 1476.0400 1302.8800 ;
        RECT 1474.4400 1280.6400 1476.0400 1281.1200 ;
        RECT 1474.4400 1286.0800 1476.0400 1286.5600 ;
        RECT 1429.4400 1291.5200 1431.0400 1292.0000 ;
        RECT 1429.4400 1296.9600 1431.0400 1297.4400 ;
        RECT 1429.4400 1302.4000 1431.0400 1302.8800 ;
        RECT 1429.4400 1280.6400 1431.0400 1281.1200 ;
        RECT 1429.4400 1286.0800 1431.0400 1286.5600 ;
        RECT 1384.4400 1318.7200 1386.0400 1319.2000 ;
        RECT 1384.4400 1324.1600 1386.0400 1324.6400 ;
        RECT 1384.4400 1329.6000 1386.0400 1330.0800 ;
        RECT 1372.6800 1318.7200 1375.6800 1319.2000 ;
        RECT 1372.6800 1324.1600 1375.6800 1324.6400 ;
        RECT 1372.6800 1329.6000 1375.6800 1330.0800 ;
        RECT 1384.4400 1307.8400 1386.0400 1308.3200 ;
        RECT 1384.4400 1313.2800 1386.0400 1313.7600 ;
        RECT 1372.6800 1307.8400 1375.6800 1308.3200 ;
        RECT 1372.6800 1313.2800 1375.6800 1313.7600 ;
        RECT 1384.4400 1291.5200 1386.0400 1292.0000 ;
        RECT 1384.4400 1296.9600 1386.0400 1297.4400 ;
        RECT 1384.4400 1302.4000 1386.0400 1302.8800 ;
        RECT 1372.6800 1291.5200 1375.6800 1292.0000 ;
        RECT 1372.6800 1296.9600 1375.6800 1297.4400 ;
        RECT 1372.6800 1302.4000 1375.6800 1302.8800 ;
        RECT 1384.4400 1280.6400 1386.0400 1281.1200 ;
        RECT 1384.4400 1286.0800 1386.0400 1286.5600 ;
        RECT 1372.6800 1280.6400 1375.6800 1281.1200 ;
        RECT 1372.6800 1286.0800 1375.6800 1286.5600 ;
        RECT 1474.4400 1264.3200 1476.0400 1264.8000 ;
        RECT 1474.4400 1269.7600 1476.0400 1270.2400 ;
        RECT 1474.4400 1275.2000 1476.0400 1275.6800 ;
        RECT 1474.4400 1253.4400 1476.0400 1253.9200 ;
        RECT 1474.4400 1258.8800 1476.0400 1259.3600 ;
        RECT 1429.4400 1264.3200 1431.0400 1264.8000 ;
        RECT 1429.4400 1269.7600 1431.0400 1270.2400 ;
        RECT 1429.4400 1275.2000 1431.0400 1275.6800 ;
        RECT 1429.4400 1253.4400 1431.0400 1253.9200 ;
        RECT 1429.4400 1258.8800 1431.0400 1259.3600 ;
        RECT 1474.4400 1237.1200 1476.0400 1237.6000 ;
        RECT 1474.4400 1242.5600 1476.0400 1243.0400 ;
        RECT 1474.4400 1248.0000 1476.0400 1248.4800 ;
        RECT 1474.4400 1231.6800 1476.0400 1232.1600 ;
        RECT 1429.4400 1237.1200 1431.0400 1237.6000 ;
        RECT 1429.4400 1242.5600 1431.0400 1243.0400 ;
        RECT 1429.4400 1248.0000 1431.0400 1248.4800 ;
        RECT 1429.4400 1231.6800 1431.0400 1232.1600 ;
        RECT 1384.4400 1264.3200 1386.0400 1264.8000 ;
        RECT 1384.4400 1269.7600 1386.0400 1270.2400 ;
        RECT 1384.4400 1275.2000 1386.0400 1275.6800 ;
        RECT 1372.6800 1264.3200 1375.6800 1264.8000 ;
        RECT 1372.6800 1269.7600 1375.6800 1270.2400 ;
        RECT 1372.6800 1275.2000 1375.6800 1275.6800 ;
        RECT 1384.4400 1253.4400 1386.0400 1253.9200 ;
        RECT 1384.4400 1258.8800 1386.0400 1259.3600 ;
        RECT 1372.6800 1253.4400 1375.6800 1253.9200 ;
        RECT 1372.6800 1258.8800 1375.6800 1259.3600 ;
        RECT 1384.4400 1237.1200 1386.0400 1237.6000 ;
        RECT 1384.4400 1242.5600 1386.0400 1243.0400 ;
        RECT 1384.4400 1248.0000 1386.0400 1248.4800 ;
        RECT 1372.6800 1237.1200 1375.6800 1237.6000 ;
        RECT 1372.6800 1242.5600 1375.6800 1243.0400 ;
        RECT 1372.6800 1248.0000 1375.6800 1248.4800 ;
        RECT 1372.6800 1231.6800 1375.6800 1232.1600 ;
        RECT 1384.4400 1231.6800 1386.0400 1232.1600 ;
        RECT 1372.6800 1436.5900 1579.7800 1439.5900 ;
        RECT 1372.6800 1223.4900 1579.7800 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 993.8500 1566.0400 1209.9500 ;
        RECT 1519.4400 993.8500 1521.0400 1209.9500 ;
        RECT 1474.4400 993.8500 1476.0400 1209.9500 ;
        RECT 1429.4400 993.8500 1431.0400 1209.9500 ;
        RECT 1384.4400 993.8500 1386.0400 1209.9500 ;
        RECT 1576.7800 993.8500 1579.7800 1209.9500 ;
        RECT 1372.6800 993.8500 1375.6800 1209.9500 ;
      LAYER met3 ;
        RECT 1576.7800 1187.0000 1579.7800 1187.4800 ;
        RECT 1576.7800 1192.4400 1579.7800 1192.9200 ;
        RECT 1564.4400 1187.0000 1566.0400 1187.4800 ;
        RECT 1564.4400 1192.4400 1566.0400 1192.9200 ;
        RECT 1576.7800 1197.8800 1579.7800 1198.3600 ;
        RECT 1564.4400 1197.8800 1566.0400 1198.3600 ;
        RECT 1576.7800 1176.1200 1579.7800 1176.6000 ;
        RECT 1576.7800 1181.5600 1579.7800 1182.0400 ;
        RECT 1564.4400 1176.1200 1566.0400 1176.6000 ;
        RECT 1564.4400 1181.5600 1566.0400 1182.0400 ;
        RECT 1576.7800 1159.8000 1579.7800 1160.2800 ;
        RECT 1576.7800 1165.2400 1579.7800 1165.7200 ;
        RECT 1564.4400 1159.8000 1566.0400 1160.2800 ;
        RECT 1564.4400 1165.2400 1566.0400 1165.7200 ;
        RECT 1576.7800 1170.6800 1579.7800 1171.1600 ;
        RECT 1564.4400 1170.6800 1566.0400 1171.1600 ;
        RECT 1519.4400 1187.0000 1521.0400 1187.4800 ;
        RECT 1519.4400 1192.4400 1521.0400 1192.9200 ;
        RECT 1519.4400 1197.8800 1521.0400 1198.3600 ;
        RECT 1519.4400 1176.1200 1521.0400 1176.6000 ;
        RECT 1519.4400 1181.5600 1521.0400 1182.0400 ;
        RECT 1519.4400 1159.8000 1521.0400 1160.2800 ;
        RECT 1519.4400 1165.2400 1521.0400 1165.7200 ;
        RECT 1519.4400 1170.6800 1521.0400 1171.1600 ;
        RECT 1576.7800 1143.4800 1579.7800 1143.9600 ;
        RECT 1576.7800 1148.9200 1579.7800 1149.4000 ;
        RECT 1576.7800 1154.3600 1579.7800 1154.8400 ;
        RECT 1564.4400 1143.4800 1566.0400 1143.9600 ;
        RECT 1564.4400 1148.9200 1566.0400 1149.4000 ;
        RECT 1564.4400 1154.3600 1566.0400 1154.8400 ;
        RECT 1576.7800 1132.6000 1579.7800 1133.0800 ;
        RECT 1576.7800 1138.0400 1579.7800 1138.5200 ;
        RECT 1564.4400 1132.6000 1566.0400 1133.0800 ;
        RECT 1564.4400 1138.0400 1566.0400 1138.5200 ;
        RECT 1576.7800 1116.2800 1579.7800 1116.7600 ;
        RECT 1576.7800 1121.7200 1579.7800 1122.2000 ;
        RECT 1576.7800 1127.1600 1579.7800 1127.6400 ;
        RECT 1564.4400 1116.2800 1566.0400 1116.7600 ;
        RECT 1564.4400 1121.7200 1566.0400 1122.2000 ;
        RECT 1564.4400 1127.1600 1566.0400 1127.6400 ;
        RECT 1576.7800 1105.4000 1579.7800 1105.8800 ;
        RECT 1576.7800 1110.8400 1579.7800 1111.3200 ;
        RECT 1564.4400 1105.4000 1566.0400 1105.8800 ;
        RECT 1564.4400 1110.8400 1566.0400 1111.3200 ;
        RECT 1519.4400 1143.4800 1521.0400 1143.9600 ;
        RECT 1519.4400 1148.9200 1521.0400 1149.4000 ;
        RECT 1519.4400 1154.3600 1521.0400 1154.8400 ;
        RECT 1519.4400 1132.6000 1521.0400 1133.0800 ;
        RECT 1519.4400 1138.0400 1521.0400 1138.5200 ;
        RECT 1519.4400 1116.2800 1521.0400 1116.7600 ;
        RECT 1519.4400 1121.7200 1521.0400 1122.2000 ;
        RECT 1519.4400 1127.1600 1521.0400 1127.6400 ;
        RECT 1519.4400 1105.4000 1521.0400 1105.8800 ;
        RECT 1519.4400 1110.8400 1521.0400 1111.3200 ;
        RECT 1474.4400 1187.0000 1476.0400 1187.4800 ;
        RECT 1474.4400 1192.4400 1476.0400 1192.9200 ;
        RECT 1474.4400 1197.8800 1476.0400 1198.3600 ;
        RECT 1429.4400 1187.0000 1431.0400 1187.4800 ;
        RECT 1429.4400 1192.4400 1431.0400 1192.9200 ;
        RECT 1429.4400 1197.8800 1431.0400 1198.3600 ;
        RECT 1474.4400 1176.1200 1476.0400 1176.6000 ;
        RECT 1474.4400 1181.5600 1476.0400 1182.0400 ;
        RECT 1474.4400 1159.8000 1476.0400 1160.2800 ;
        RECT 1474.4400 1165.2400 1476.0400 1165.7200 ;
        RECT 1474.4400 1170.6800 1476.0400 1171.1600 ;
        RECT 1429.4400 1176.1200 1431.0400 1176.6000 ;
        RECT 1429.4400 1181.5600 1431.0400 1182.0400 ;
        RECT 1429.4400 1159.8000 1431.0400 1160.2800 ;
        RECT 1429.4400 1165.2400 1431.0400 1165.7200 ;
        RECT 1429.4400 1170.6800 1431.0400 1171.1600 ;
        RECT 1384.4400 1187.0000 1386.0400 1187.4800 ;
        RECT 1384.4400 1192.4400 1386.0400 1192.9200 ;
        RECT 1372.6800 1192.4400 1375.6800 1192.9200 ;
        RECT 1372.6800 1187.0000 1375.6800 1187.4800 ;
        RECT 1372.6800 1197.8800 1375.6800 1198.3600 ;
        RECT 1384.4400 1197.8800 1386.0400 1198.3600 ;
        RECT 1384.4400 1176.1200 1386.0400 1176.6000 ;
        RECT 1384.4400 1181.5600 1386.0400 1182.0400 ;
        RECT 1372.6800 1181.5600 1375.6800 1182.0400 ;
        RECT 1372.6800 1176.1200 1375.6800 1176.6000 ;
        RECT 1384.4400 1159.8000 1386.0400 1160.2800 ;
        RECT 1384.4400 1165.2400 1386.0400 1165.7200 ;
        RECT 1372.6800 1165.2400 1375.6800 1165.7200 ;
        RECT 1372.6800 1159.8000 1375.6800 1160.2800 ;
        RECT 1372.6800 1170.6800 1375.6800 1171.1600 ;
        RECT 1384.4400 1170.6800 1386.0400 1171.1600 ;
        RECT 1474.4400 1143.4800 1476.0400 1143.9600 ;
        RECT 1474.4400 1148.9200 1476.0400 1149.4000 ;
        RECT 1474.4400 1154.3600 1476.0400 1154.8400 ;
        RECT 1474.4400 1132.6000 1476.0400 1133.0800 ;
        RECT 1474.4400 1138.0400 1476.0400 1138.5200 ;
        RECT 1429.4400 1143.4800 1431.0400 1143.9600 ;
        RECT 1429.4400 1148.9200 1431.0400 1149.4000 ;
        RECT 1429.4400 1154.3600 1431.0400 1154.8400 ;
        RECT 1429.4400 1132.6000 1431.0400 1133.0800 ;
        RECT 1429.4400 1138.0400 1431.0400 1138.5200 ;
        RECT 1474.4400 1116.2800 1476.0400 1116.7600 ;
        RECT 1474.4400 1121.7200 1476.0400 1122.2000 ;
        RECT 1474.4400 1127.1600 1476.0400 1127.6400 ;
        RECT 1474.4400 1105.4000 1476.0400 1105.8800 ;
        RECT 1474.4400 1110.8400 1476.0400 1111.3200 ;
        RECT 1429.4400 1116.2800 1431.0400 1116.7600 ;
        RECT 1429.4400 1121.7200 1431.0400 1122.2000 ;
        RECT 1429.4400 1127.1600 1431.0400 1127.6400 ;
        RECT 1429.4400 1105.4000 1431.0400 1105.8800 ;
        RECT 1429.4400 1110.8400 1431.0400 1111.3200 ;
        RECT 1384.4400 1143.4800 1386.0400 1143.9600 ;
        RECT 1384.4400 1148.9200 1386.0400 1149.4000 ;
        RECT 1384.4400 1154.3600 1386.0400 1154.8400 ;
        RECT 1372.6800 1143.4800 1375.6800 1143.9600 ;
        RECT 1372.6800 1148.9200 1375.6800 1149.4000 ;
        RECT 1372.6800 1154.3600 1375.6800 1154.8400 ;
        RECT 1384.4400 1132.6000 1386.0400 1133.0800 ;
        RECT 1384.4400 1138.0400 1386.0400 1138.5200 ;
        RECT 1372.6800 1132.6000 1375.6800 1133.0800 ;
        RECT 1372.6800 1138.0400 1375.6800 1138.5200 ;
        RECT 1384.4400 1116.2800 1386.0400 1116.7600 ;
        RECT 1384.4400 1121.7200 1386.0400 1122.2000 ;
        RECT 1384.4400 1127.1600 1386.0400 1127.6400 ;
        RECT 1372.6800 1116.2800 1375.6800 1116.7600 ;
        RECT 1372.6800 1121.7200 1375.6800 1122.2000 ;
        RECT 1372.6800 1127.1600 1375.6800 1127.6400 ;
        RECT 1384.4400 1105.4000 1386.0400 1105.8800 ;
        RECT 1384.4400 1110.8400 1386.0400 1111.3200 ;
        RECT 1372.6800 1105.4000 1375.6800 1105.8800 ;
        RECT 1372.6800 1110.8400 1375.6800 1111.3200 ;
        RECT 1576.7800 1089.0800 1579.7800 1089.5600 ;
        RECT 1576.7800 1094.5200 1579.7800 1095.0000 ;
        RECT 1576.7800 1099.9600 1579.7800 1100.4400 ;
        RECT 1564.4400 1089.0800 1566.0400 1089.5600 ;
        RECT 1564.4400 1094.5200 1566.0400 1095.0000 ;
        RECT 1564.4400 1099.9600 1566.0400 1100.4400 ;
        RECT 1576.7800 1078.2000 1579.7800 1078.6800 ;
        RECT 1576.7800 1083.6400 1579.7800 1084.1200 ;
        RECT 1564.4400 1078.2000 1566.0400 1078.6800 ;
        RECT 1564.4400 1083.6400 1566.0400 1084.1200 ;
        RECT 1576.7800 1061.8800 1579.7800 1062.3600 ;
        RECT 1576.7800 1067.3200 1579.7800 1067.8000 ;
        RECT 1576.7800 1072.7600 1579.7800 1073.2400 ;
        RECT 1564.4400 1061.8800 1566.0400 1062.3600 ;
        RECT 1564.4400 1067.3200 1566.0400 1067.8000 ;
        RECT 1564.4400 1072.7600 1566.0400 1073.2400 ;
        RECT 1576.7800 1051.0000 1579.7800 1051.4800 ;
        RECT 1576.7800 1056.4400 1579.7800 1056.9200 ;
        RECT 1564.4400 1051.0000 1566.0400 1051.4800 ;
        RECT 1564.4400 1056.4400 1566.0400 1056.9200 ;
        RECT 1519.4400 1089.0800 1521.0400 1089.5600 ;
        RECT 1519.4400 1094.5200 1521.0400 1095.0000 ;
        RECT 1519.4400 1099.9600 1521.0400 1100.4400 ;
        RECT 1519.4400 1078.2000 1521.0400 1078.6800 ;
        RECT 1519.4400 1083.6400 1521.0400 1084.1200 ;
        RECT 1519.4400 1061.8800 1521.0400 1062.3600 ;
        RECT 1519.4400 1067.3200 1521.0400 1067.8000 ;
        RECT 1519.4400 1072.7600 1521.0400 1073.2400 ;
        RECT 1519.4400 1051.0000 1521.0400 1051.4800 ;
        RECT 1519.4400 1056.4400 1521.0400 1056.9200 ;
        RECT 1576.7800 1034.6800 1579.7800 1035.1600 ;
        RECT 1576.7800 1040.1200 1579.7800 1040.6000 ;
        RECT 1576.7800 1045.5600 1579.7800 1046.0400 ;
        RECT 1564.4400 1034.6800 1566.0400 1035.1600 ;
        RECT 1564.4400 1040.1200 1566.0400 1040.6000 ;
        RECT 1564.4400 1045.5600 1566.0400 1046.0400 ;
        RECT 1576.7800 1023.8000 1579.7800 1024.2800 ;
        RECT 1576.7800 1029.2400 1579.7800 1029.7200 ;
        RECT 1564.4400 1023.8000 1566.0400 1024.2800 ;
        RECT 1564.4400 1029.2400 1566.0400 1029.7200 ;
        RECT 1576.7800 1007.4800 1579.7800 1007.9600 ;
        RECT 1576.7800 1012.9200 1579.7800 1013.4000 ;
        RECT 1576.7800 1018.3600 1579.7800 1018.8400 ;
        RECT 1564.4400 1007.4800 1566.0400 1007.9600 ;
        RECT 1564.4400 1012.9200 1566.0400 1013.4000 ;
        RECT 1564.4400 1018.3600 1566.0400 1018.8400 ;
        RECT 1576.7800 1002.0400 1579.7800 1002.5200 ;
        RECT 1564.4400 1002.0400 1566.0400 1002.5200 ;
        RECT 1519.4400 1034.6800 1521.0400 1035.1600 ;
        RECT 1519.4400 1040.1200 1521.0400 1040.6000 ;
        RECT 1519.4400 1045.5600 1521.0400 1046.0400 ;
        RECT 1519.4400 1023.8000 1521.0400 1024.2800 ;
        RECT 1519.4400 1029.2400 1521.0400 1029.7200 ;
        RECT 1519.4400 1007.4800 1521.0400 1007.9600 ;
        RECT 1519.4400 1012.9200 1521.0400 1013.4000 ;
        RECT 1519.4400 1018.3600 1521.0400 1018.8400 ;
        RECT 1519.4400 1002.0400 1521.0400 1002.5200 ;
        RECT 1474.4400 1089.0800 1476.0400 1089.5600 ;
        RECT 1474.4400 1094.5200 1476.0400 1095.0000 ;
        RECT 1474.4400 1099.9600 1476.0400 1100.4400 ;
        RECT 1474.4400 1078.2000 1476.0400 1078.6800 ;
        RECT 1474.4400 1083.6400 1476.0400 1084.1200 ;
        RECT 1429.4400 1089.0800 1431.0400 1089.5600 ;
        RECT 1429.4400 1094.5200 1431.0400 1095.0000 ;
        RECT 1429.4400 1099.9600 1431.0400 1100.4400 ;
        RECT 1429.4400 1078.2000 1431.0400 1078.6800 ;
        RECT 1429.4400 1083.6400 1431.0400 1084.1200 ;
        RECT 1474.4400 1061.8800 1476.0400 1062.3600 ;
        RECT 1474.4400 1067.3200 1476.0400 1067.8000 ;
        RECT 1474.4400 1072.7600 1476.0400 1073.2400 ;
        RECT 1474.4400 1051.0000 1476.0400 1051.4800 ;
        RECT 1474.4400 1056.4400 1476.0400 1056.9200 ;
        RECT 1429.4400 1061.8800 1431.0400 1062.3600 ;
        RECT 1429.4400 1067.3200 1431.0400 1067.8000 ;
        RECT 1429.4400 1072.7600 1431.0400 1073.2400 ;
        RECT 1429.4400 1051.0000 1431.0400 1051.4800 ;
        RECT 1429.4400 1056.4400 1431.0400 1056.9200 ;
        RECT 1384.4400 1089.0800 1386.0400 1089.5600 ;
        RECT 1384.4400 1094.5200 1386.0400 1095.0000 ;
        RECT 1384.4400 1099.9600 1386.0400 1100.4400 ;
        RECT 1372.6800 1089.0800 1375.6800 1089.5600 ;
        RECT 1372.6800 1094.5200 1375.6800 1095.0000 ;
        RECT 1372.6800 1099.9600 1375.6800 1100.4400 ;
        RECT 1384.4400 1078.2000 1386.0400 1078.6800 ;
        RECT 1384.4400 1083.6400 1386.0400 1084.1200 ;
        RECT 1372.6800 1078.2000 1375.6800 1078.6800 ;
        RECT 1372.6800 1083.6400 1375.6800 1084.1200 ;
        RECT 1384.4400 1061.8800 1386.0400 1062.3600 ;
        RECT 1384.4400 1067.3200 1386.0400 1067.8000 ;
        RECT 1384.4400 1072.7600 1386.0400 1073.2400 ;
        RECT 1372.6800 1061.8800 1375.6800 1062.3600 ;
        RECT 1372.6800 1067.3200 1375.6800 1067.8000 ;
        RECT 1372.6800 1072.7600 1375.6800 1073.2400 ;
        RECT 1384.4400 1051.0000 1386.0400 1051.4800 ;
        RECT 1384.4400 1056.4400 1386.0400 1056.9200 ;
        RECT 1372.6800 1051.0000 1375.6800 1051.4800 ;
        RECT 1372.6800 1056.4400 1375.6800 1056.9200 ;
        RECT 1474.4400 1034.6800 1476.0400 1035.1600 ;
        RECT 1474.4400 1040.1200 1476.0400 1040.6000 ;
        RECT 1474.4400 1045.5600 1476.0400 1046.0400 ;
        RECT 1474.4400 1023.8000 1476.0400 1024.2800 ;
        RECT 1474.4400 1029.2400 1476.0400 1029.7200 ;
        RECT 1429.4400 1034.6800 1431.0400 1035.1600 ;
        RECT 1429.4400 1040.1200 1431.0400 1040.6000 ;
        RECT 1429.4400 1045.5600 1431.0400 1046.0400 ;
        RECT 1429.4400 1023.8000 1431.0400 1024.2800 ;
        RECT 1429.4400 1029.2400 1431.0400 1029.7200 ;
        RECT 1474.4400 1007.4800 1476.0400 1007.9600 ;
        RECT 1474.4400 1012.9200 1476.0400 1013.4000 ;
        RECT 1474.4400 1018.3600 1476.0400 1018.8400 ;
        RECT 1474.4400 1002.0400 1476.0400 1002.5200 ;
        RECT 1429.4400 1007.4800 1431.0400 1007.9600 ;
        RECT 1429.4400 1012.9200 1431.0400 1013.4000 ;
        RECT 1429.4400 1018.3600 1431.0400 1018.8400 ;
        RECT 1429.4400 1002.0400 1431.0400 1002.5200 ;
        RECT 1384.4400 1034.6800 1386.0400 1035.1600 ;
        RECT 1384.4400 1040.1200 1386.0400 1040.6000 ;
        RECT 1384.4400 1045.5600 1386.0400 1046.0400 ;
        RECT 1372.6800 1034.6800 1375.6800 1035.1600 ;
        RECT 1372.6800 1040.1200 1375.6800 1040.6000 ;
        RECT 1372.6800 1045.5600 1375.6800 1046.0400 ;
        RECT 1384.4400 1023.8000 1386.0400 1024.2800 ;
        RECT 1384.4400 1029.2400 1386.0400 1029.7200 ;
        RECT 1372.6800 1023.8000 1375.6800 1024.2800 ;
        RECT 1372.6800 1029.2400 1375.6800 1029.7200 ;
        RECT 1384.4400 1007.4800 1386.0400 1007.9600 ;
        RECT 1384.4400 1012.9200 1386.0400 1013.4000 ;
        RECT 1384.4400 1018.3600 1386.0400 1018.8400 ;
        RECT 1372.6800 1007.4800 1375.6800 1007.9600 ;
        RECT 1372.6800 1012.9200 1375.6800 1013.4000 ;
        RECT 1372.6800 1018.3600 1375.6800 1018.8400 ;
        RECT 1372.6800 1002.0400 1375.6800 1002.5200 ;
        RECT 1384.4400 1002.0400 1386.0400 1002.5200 ;
        RECT 1372.6800 1206.9500 1579.7800 1209.9500 ;
        RECT 1372.6800 993.8500 1579.7800 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1564.4400 764.2100 1566.0400 980.3100 ;
        RECT 1519.4400 764.2100 1521.0400 980.3100 ;
        RECT 1474.4400 764.2100 1476.0400 980.3100 ;
        RECT 1429.4400 764.2100 1431.0400 980.3100 ;
        RECT 1384.4400 764.2100 1386.0400 980.3100 ;
        RECT 1576.7800 764.2100 1579.7800 980.3100 ;
        RECT 1372.6800 764.2100 1375.6800 980.3100 ;
      LAYER met3 ;
        RECT 1576.7800 957.3600 1579.7800 957.8400 ;
        RECT 1576.7800 962.8000 1579.7800 963.2800 ;
        RECT 1564.4400 957.3600 1566.0400 957.8400 ;
        RECT 1564.4400 962.8000 1566.0400 963.2800 ;
        RECT 1576.7800 968.2400 1579.7800 968.7200 ;
        RECT 1564.4400 968.2400 1566.0400 968.7200 ;
        RECT 1576.7800 946.4800 1579.7800 946.9600 ;
        RECT 1576.7800 951.9200 1579.7800 952.4000 ;
        RECT 1564.4400 946.4800 1566.0400 946.9600 ;
        RECT 1564.4400 951.9200 1566.0400 952.4000 ;
        RECT 1576.7800 930.1600 1579.7800 930.6400 ;
        RECT 1576.7800 935.6000 1579.7800 936.0800 ;
        RECT 1564.4400 930.1600 1566.0400 930.6400 ;
        RECT 1564.4400 935.6000 1566.0400 936.0800 ;
        RECT 1576.7800 941.0400 1579.7800 941.5200 ;
        RECT 1564.4400 941.0400 1566.0400 941.5200 ;
        RECT 1519.4400 957.3600 1521.0400 957.8400 ;
        RECT 1519.4400 962.8000 1521.0400 963.2800 ;
        RECT 1519.4400 968.2400 1521.0400 968.7200 ;
        RECT 1519.4400 946.4800 1521.0400 946.9600 ;
        RECT 1519.4400 951.9200 1521.0400 952.4000 ;
        RECT 1519.4400 930.1600 1521.0400 930.6400 ;
        RECT 1519.4400 935.6000 1521.0400 936.0800 ;
        RECT 1519.4400 941.0400 1521.0400 941.5200 ;
        RECT 1576.7800 913.8400 1579.7800 914.3200 ;
        RECT 1576.7800 919.2800 1579.7800 919.7600 ;
        RECT 1576.7800 924.7200 1579.7800 925.2000 ;
        RECT 1564.4400 913.8400 1566.0400 914.3200 ;
        RECT 1564.4400 919.2800 1566.0400 919.7600 ;
        RECT 1564.4400 924.7200 1566.0400 925.2000 ;
        RECT 1576.7800 902.9600 1579.7800 903.4400 ;
        RECT 1576.7800 908.4000 1579.7800 908.8800 ;
        RECT 1564.4400 902.9600 1566.0400 903.4400 ;
        RECT 1564.4400 908.4000 1566.0400 908.8800 ;
        RECT 1576.7800 886.6400 1579.7800 887.1200 ;
        RECT 1576.7800 892.0800 1579.7800 892.5600 ;
        RECT 1576.7800 897.5200 1579.7800 898.0000 ;
        RECT 1564.4400 886.6400 1566.0400 887.1200 ;
        RECT 1564.4400 892.0800 1566.0400 892.5600 ;
        RECT 1564.4400 897.5200 1566.0400 898.0000 ;
        RECT 1576.7800 875.7600 1579.7800 876.2400 ;
        RECT 1576.7800 881.2000 1579.7800 881.6800 ;
        RECT 1564.4400 875.7600 1566.0400 876.2400 ;
        RECT 1564.4400 881.2000 1566.0400 881.6800 ;
        RECT 1519.4400 913.8400 1521.0400 914.3200 ;
        RECT 1519.4400 919.2800 1521.0400 919.7600 ;
        RECT 1519.4400 924.7200 1521.0400 925.2000 ;
        RECT 1519.4400 902.9600 1521.0400 903.4400 ;
        RECT 1519.4400 908.4000 1521.0400 908.8800 ;
        RECT 1519.4400 886.6400 1521.0400 887.1200 ;
        RECT 1519.4400 892.0800 1521.0400 892.5600 ;
        RECT 1519.4400 897.5200 1521.0400 898.0000 ;
        RECT 1519.4400 875.7600 1521.0400 876.2400 ;
        RECT 1519.4400 881.2000 1521.0400 881.6800 ;
        RECT 1474.4400 957.3600 1476.0400 957.8400 ;
        RECT 1474.4400 962.8000 1476.0400 963.2800 ;
        RECT 1474.4400 968.2400 1476.0400 968.7200 ;
        RECT 1429.4400 957.3600 1431.0400 957.8400 ;
        RECT 1429.4400 962.8000 1431.0400 963.2800 ;
        RECT 1429.4400 968.2400 1431.0400 968.7200 ;
        RECT 1474.4400 946.4800 1476.0400 946.9600 ;
        RECT 1474.4400 951.9200 1476.0400 952.4000 ;
        RECT 1474.4400 930.1600 1476.0400 930.6400 ;
        RECT 1474.4400 935.6000 1476.0400 936.0800 ;
        RECT 1474.4400 941.0400 1476.0400 941.5200 ;
        RECT 1429.4400 946.4800 1431.0400 946.9600 ;
        RECT 1429.4400 951.9200 1431.0400 952.4000 ;
        RECT 1429.4400 930.1600 1431.0400 930.6400 ;
        RECT 1429.4400 935.6000 1431.0400 936.0800 ;
        RECT 1429.4400 941.0400 1431.0400 941.5200 ;
        RECT 1384.4400 957.3600 1386.0400 957.8400 ;
        RECT 1384.4400 962.8000 1386.0400 963.2800 ;
        RECT 1372.6800 962.8000 1375.6800 963.2800 ;
        RECT 1372.6800 957.3600 1375.6800 957.8400 ;
        RECT 1372.6800 968.2400 1375.6800 968.7200 ;
        RECT 1384.4400 968.2400 1386.0400 968.7200 ;
        RECT 1384.4400 946.4800 1386.0400 946.9600 ;
        RECT 1384.4400 951.9200 1386.0400 952.4000 ;
        RECT 1372.6800 951.9200 1375.6800 952.4000 ;
        RECT 1372.6800 946.4800 1375.6800 946.9600 ;
        RECT 1384.4400 930.1600 1386.0400 930.6400 ;
        RECT 1384.4400 935.6000 1386.0400 936.0800 ;
        RECT 1372.6800 935.6000 1375.6800 936.0800 ;
        RECT 1372.6800 930.1600 1375.6800 930.6400 ;
        RECT 1372.6800 941.0400 1375.6800 941.5200 ;
        RECT 1384.4400 941.0400 1386.0400 941.5200 ;
        RECT 1474.4400 913.8400 1476.0400 914.3200 ;
        RECT 1474.4400 919.2800 1476.0400 919.7600 ;
        RECT 1474.4400 924.7200 1476.0400 925.2000 ;
        RECT 1474.4400 902.9600 1476.0400 903.4400 ;
        RECT 1474.4400 908.4000 1476.0400 908.8800 ;
        RECT 1429.4400 913.8400 1431.0400 914.3200 ;
        RECT 1429.4400 919.2800 1431.0400 919.7600 ;
        RECT 1429.4400 924.7200 1431.0400 925.2000 ;
        RECT 1429.4400 902.9600 1431.0400 903.4400 ;
        RECT 1429.4400 908.4000 1431.0400 908.8800 ;
        RECT 1474.4400 886.6400 1476.0400 887.1200 ;
        RECT 1474.4400 892.0800 1476.0400 892.5600 ;
        RECT 1474.4400 897.5200 1476.0400 898.0000 ;
        RECT 1474.4400 875.7600 1476.0400 876.2400 ;
        RECT 1474.4400 881.2000 1476.0400 881.6800 ;
        RECT 1429.4400 886.6400 1431.0400 887.1200 ;
        RECT 1429.4400 892.0800 1431.0400 892.5600 ;
        RECT 1429.4400 897.5200 1431.0400 898.0000 ;
        RECT 1429.4400 875.7600 1431.0400 876.2400 ;
        RECT 1429.4400 881.2000 1431.0400 881.6800 ;
        RECT 1384.4400 913.8400 1386.0400 914.3200 ;
        RECT 1384.4400 919.2800 1386.0400 919.7600 ;
        RECT 1384.4400 924.7200 1386.0400 925.2000 ;
        RECT 1372.6800 913.8400 1375.6800 914.3200 ;
        RECT 1372.6800 919.2800 1375.6800 919.7600 ;
        RECT 1372.6800 924.7200 1375.6800 925.2000 ;
        RECT 1384.4400 902.9600 1386.0400 903.4400 ;
        RECT 1384.4400 908.4000 1386.0400 908.8800 ;
        RECT 1372.6800 902.9600 1375.6800 903.4400 ;
        RECT 1372.6800 908.4000 1375.6800 908.8800 ;
        RECT 1384.4400 886.6400 1386.0400 887.1200 ;
        RECT 1384.4400 892.0800 1386.0400 892.5600 ;
        RECT 1384.4400 897.5200 1386.0400 898.0000 ;
        RECT 1372.6800 886.6400 1375.6800 887.1200 ;
        RECT 1372.6800 892.0800 1375.6800 892.5600 ;
        RECT 1372.6800 897.5200 1375.6800 898.0000 ;
        RECT 1384.4400 875.7600 1386.0400 876.2400 ;
        RECT 1384.4400 881.2000 1386.0400 881.6800 ;
        RECT 1372.6800 875.7600 1375.6800 876.2400 ;
        RECT 1372.6800 881.2000 1375.6800 881.6800 ;
        RECT 1576.7800 859.4400 1579.7800 859.9200 ;
        RECT 1576.7800 864.8800 1579.7800 865.3600 ;
        RECT 1576.7800 870.3200 1579.7800 870.8000 ;
        RECT 1564.4400 859.4400 1566.0400 859.9200 ;
        RECT 1564.4400 864.8800 1566.0400 865.3600 ;
        RECT 1564.4400 870.3200 1566.0400 870.8000 ;
        RECT 1576.7800 848.5600 1579.7800 849.0400 ;
        RECT 1576.7800 854.0000 1579.7800 854.4800 ;
        RECT 1564.4400 848.5600 1566.0400 849.0400 ;
        RECT 1564.4400 854.0000 1566.0400 854.4800 ;
        RECT 1576.7800 832.2400 1579.7800 832.7200 ;
        RECT 1576.7800 837.6800 1579.7800 838.1600 ;
        RECT 1576.7800 843.1200 1579.7800 843.6000 ;
        RECT 1564.4400 832.2400 1566.0400 832.7200 ;
        RECT 1564.4400 837.6800 1566.0400 838.1600 ;
        RECT 1564.4400 843.1200 1566.0400 843.6000 ;
        RECT 1576.7800 821.3600 1579.7800 821.8400 ;
        RECT 1576.7800 826.8000 1579.7800 827.2800 ;
        RECT 1564.4400 821.3600 1566.0400 821.8400 ;
        RECT 1564.4400 826.8000 1566.0400 827.2800 ;
        RECT 1519.4400 859.4400 1521.0400 859.9200 ;
        RECT 1519.4400 864.8800 1521.0400 865.3600 ;
        RECT 1519.4400 870.3200 1521.0400 870.8000 ;
        RECT 1519.4400 848.5600 1521.0400 849.0400 ;
        RECT 1519.4400 854.0000 1521.0400 854.4800 ;
        RECT 1519.4400 832.2400 1521.0400 832.7200 ;
        RECT 1519.4400 837.6800 1521.0400 838.1600 ;
        RECT 1519.4400 843.1200 1521.0400 843.6000 ;
        RECT 1519.4400 821.3600 1521.0400 821.8400 ;
        RECT 1519.4400 826.8000 1521.0400 827.2800 ;
        RECT 1576.7800 805.0400 1579.7800 805.5200 ;
        RECT 1576.7800 810.4800 1579.7800 810.9600 ;
        RECT 1576.7800 815.9200 1579.7800 816.4000 ;
        RECT 1564.4400 805.0400 1566.0400 805.5200 ;
        RECT 1564.4400 810.4800 1566.0400 810.9600 ;
        RECT 1564.4400 815.9200 1566.0400 816.4000 ;
        RECT 1576.7800 794.1600 1579.7800 794.6400 ;
        RECT 1576.7800 799.6000 1579.7800 800.0800 ;
        RECT 1564.4400 794.1600 1566.0400 794.6400 ;
        RECT 1564.4400 799.6000 1566.0400 800.0800 ;
        RECT 1576.7800 777.8400 1579.7800 778.3200 ;
        RECT 1576.7800 783.2800 1579.7800 783.7600 ;
        RECT 1576.7800 788.7200 1579.7800 789.2000 ;
        RECT 1564.4400 777.8400 1566.0400 778.3200 ;
        RECT 1564.4400 783.2800 1566.0400 783.7600 ;
        RECT 1564.4400 788.7200 1566.0400 789.2000 ;
        RECT 1576.7800 772.4000 1579.7800 772.8800 ;
        RECT 1564.4400 772.4000 1566.0400 772.8800 ;
        RECT 1519.4400 805.0400 1521.0400 805.5200 ;
        RECT 1519.4400 810.4800 1521.0400 810.9600 ;
        RECT 1519.4400 815.9200 1521.0400 816.4000 ;
        RECT 1519.4400 794.1600 1521.0400 794.6400 ;
        RECT 1519.4400 799.6000 1521.0400 800.0800 ;
        RECT 1519.4400 777.8400 1521.0400 778.3200 ;
        RECT 1519.4400 783.2800 1521.0400 783.7600 ;
        RECT 1519.4400 788.7200 1521.0400 789.2000 ;
        RECT 1519.4400 772.4000 1521.0400 772.8800 ;
        RECT 1474.4400 859.4400 1476.0400 859.9200 ;
        RECT 1474.4400 864.8800 1476.0400 865.3600 ;
        RECT 1474.4400 870.3200 1476.0400 870.8000 ;
        RECT 1474.4400 848.5600 1476.0400 849.0400 ;
        RECT 1474.4400 854.0000 1476.0400 854.4800 ;
        RECT 1429.4400 859.4400 1431.0400 859.9200 ;
        RECT 1429.4400 864.8800 1431.0400 865.3600 ;
        RECT 1429.4400 870.3200 1431.0400 870.8000 ;
        RECT 1429.4400 848.5600 1431.0400 849.0400 ;
        RECT 1429.4400 854.0000 1431.0400 854.4800 ;
        RECT 1474.4400 832.2400 1476.0400 832.7200 ;
        RECT 1474.4400 837.6800 1476.0400 838.1600 ;
        RECT 1474.4400 843.1200 1476.0400 843.6000 ;
        RECT 1474.4400 821.3600 1476.0400 821.8400 ;
        RECT 1474.4400 826.8000 1476.0400 827.2800 ;
        RECT 1429.4400 832.2400 1431.0400 832.7200 ;
        RECT 1429.4400 837.6800 1431.0400 838.1600 ;
        RECT 1429.4400 843.1200 1431.0400 843.6000 ;
        RECT 1429.4400 821.3600 1431.0400 821.8400 ;
        RECT 1429.4400 826.8000 1431.0400 827.2800 ;
        RECT 1384.4400 859.4400 1386.0400 859.9200 ;
        RECT 1384.4400 864.8800 1386.0400 865.3600 ;
        RECT 1384.4400 870.3200 1386.0400 870.8000 ;
        RECT 1372.6800 859.4400 1375.6800 859.9200 ;
        RECT 1372.6800 864.8800 1375.6800 865.3600 ;
        RECT 1372.6800 870.3200 1375.6800 870.8000 ;
        RECT 1384.4400 848.5600 1386.0400 849.0400 ;
        RECT 1384.4400 854.0000 1386.0400 854.4800 ;
        RECT 1372.6800 848.5600 1375.6800 849.0400 ;
        RECT 1372.6800 854.0000 1375.6800 854.4800 ;
        RECT 1384.4400 832.2400 1386.0400 832.7200 ;
        RECT 1384.4400 837.6800 1386.0400 838.1600 ;
        RECT 1384.4400 843.1200 1386.0400 843.6000 ;
        RECT 1372.6800 832.2400 1375.6800 832.7200 ;
        RECT 1372.6800 837.6800 1375.6800 838.1600 ;
        RECT 1372.6800 843.1200 1375.6800 843.6000 ;
        RECT 1384.4400 821.3600 1386.0400 821.8400 ;
        RECT 1384.4400 826.8000 1386.0400 827.2800 ;
        RECT 1372.6800 821.3600 1375.6800 821.8400 ;
        RECT 1372.6800 826.8000 1375.6800 827.2800 ;
        RECT 1474.4400 805.0400 1476.0400 805.5200 ;
        RECT 1474.4400 810.4800 1476.0400 810.9600 ;
        RECT 1474.4400 815.9200 1476.0400 816.4000 ;
        RECT 1474.4400 794.1600 1476.0400 794.6400 ;
        RECT 1474.4400 799.6000 1476.0400 800.0800 ;
        RECT 1429.4400 805.0400 1431.0400 805.5200 ;
        RECT 1429.4400 810.4800 1431.0400 810.9600 ;
        RECT 1429.4400 815.9200 1431.0400 816.4000 ;
        RECT 1429.4400 794.1600 1431.0400 794.6400 ;
        RECT 1429.4400 799.6000 1431.0400 800.0800 ;
        RECT 1474.4400 777.8400 1476.0400 778.3200 ;
        RECT 1474.4400 783.2800 1476.0400 783.7600 ;
        RECT 1474.4400 788.7200 1476.0400 789.2000 ;
        RECT 1474.4400 772.4000 1476.0400 772.8800 ;
        RECT 1429.4400 777.8400 1431.0400 778.3200 ;
        RECT 1429.4400 783.2800 1431.0400 783.7600 ;
        RECT 1429.4400 788.7200 1431.0400 789.2000 ;
        RECT 1429.4400 772.4000 1431.0400 772.8800 ;
        RECT 1384.4400 805.0400 1386.0400 805.5200 ;
        RECT 1384.4400 810.4800 1386.0400 810.9600 ;
        RECT 1384.4400 815.9200 1386.0400 816.4000 ;
        RECT 1372.6800 805.0400 1375.6800 805.5200 ;
        RECT 1372.6800 810.4800 1375.6800 810.9600 ;
        RECT 1372.6800 815.9200 1375.6800 816.4000 ;
        RECT 1384.4400 794.1600 1386.0400 794.6400 ;
        RECT 1384.4400 799.6000 1386.0400 800.0800 ;
        RECT 1372.6800 794.1600 1375.6800 794.6400 ;
        RECT 1372.6800 799.6000 1375.6800 800.0800 ;
        RECT 1384.4400 777.8400 1386.0400 778.3200 ;
        RECT 1384.4400 783.2800 1386.0400 783.7600 ;
        RECT 1384.4400 788.7200 1386.0400 789.2000 ;
        RECT 1372.6800 777.8400 1375.6800 778.3200 ;
        RECT 1372.6800 783.2800 1375.6800 783.7600 ;
        RECT 1372.6800 788.7200 1375.6800 789.2000 ;
        RECT 1372.6800 772.4000 1375.6800 772.8800 ;
        RECT 1384.4400 772.4000 1386.0400 772.8800 ;
        RECT 1372.6800 977.3100 1579.7800 980.3100 ;
        RECT 1372.6800 764.2100 1579.7800 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1593.9000 2830.6100 1595.9000 2857.5400 ;
        RECT 1797.0000 2830.6100 1799.0000 2857.5400 ;
      LAYER met3 ;
        RECT 1797.0000 2847.3200 1799.0000 2847.8000 ;
        RECT 1593.9000 2847.3200 1595.9000 2847.8000 ;
        RECT 1797.0000 2841.8800 1799.0000 2842.3600 ;
        RECT 1797.0000 2836.4400 1799.0000 2836.9200 ;
        RECT 1593.9000 2841.8800 1595.9000 2842.3600 ;
        RECT 1593.9000 2836.4400 1595.9000 2836.9200 ;
        RECT 1593.9000 2855.5400 1799.0000 2857.5400 ;
        RECT 1593.9000 2830.6100 1799.0000 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 534.5700 1786.2600 750.6700 ;
        RECT 1739.6600 534.5700 1741.2600 750.6700 ;
        RECT 1694.6600 534.5700 1696.2600 750.6700 ;
        RECT 1649.6600 534.5700 1651.2600 750.6700 ;
        RECT 1604.6600 534.5700 1606.2600 750.6700 ;
        RECT 1797.0000 534.5700 1800.0000 750.6700 ;
        RECT 1592.9000 534.5700 1595.9000 750.6700 ;
      LAYER met3 ;
        RECT 1797.0000 727.7200 1800.0000 728.2000 ;
        RECT 1797.0000 733.1600 1800.0000 733.6400 ;
        RECT 1784.6600 727.7200 1786.2600 728.2000 ;
        RECT 1784.6600 733.1600 1786.2600 733.6400 ;
        RECT 1797.0000 738.6000 1800.0000 739.0800 ;
        RECT 1784.6600 738.6000 1786.2600 739.0800 ;
        RECT 1797.0000 716.8400 1800.0000 717.3200 ;
        RECT 1797.0000 722.2800 1800.0000 722.7600 ;
        RECT 1784.6600 716.8400 1786.2600 717.3200 ;
        RECT 1784.6600 722.2800 1786.2600 722.7600 ;
        RECT 1797.0000 700.5200 1800.0000 701.0000 ;
        RECT 1797.0000 705.9600 1800.0000 706.4400 ;
        RECT 1784.6600 700.5200 1786.2600 701.0000 ;
        RECT 1784.6600 705.9600 1786.2600 706.4400 ;
        RECT 1797.0000 711.4000 1800.0000 711.8800 ;
        RECT 1784.6600 711.4000 1786.2600 711.8800 ;
        RECT 1739.6600 727.7200 1741.2600 728.2000 ;
        RECT 1739.6600 733.1600 1741.2600 733.6400 ;
        RECT 1739.6600 738.6000 1741.2600 739.0800 ;
        RECT 1739.6600 716.8400 1741.2600 717.3200 ;
        RECT 1739.6600 722.2800 1741.2600 722.7600 ;
        RECT 1739.6600 700.5200 1741.2600 701.0000 ;
        RECT 1739.6600 705.9600 1741.2600 706.4400 ;
        RECT 1739.6600 711.4000 1741.2600 711.8800 ;
        RECT 1797.0000 684.2000 1800.0000 684.6800 ;
        RECT 1797.0000 689.6400 1800.0000 690.1200 ;
        RECT 1797.0000 695.0800 1800.0000 695.5600 ;
        RECT 1784.6600 684.2000 1786.2600 684.6800 ;
        RECT 1784.6600 689.6400 1786.2600 690.1200 ;
        RECT 1784.6600 695.0800 1786.2600 695.5600 ;
        RECT 1797.0000 673.3200 1800.0000 673.8000 ;
        RECT 1797.0000 678.7600 1800.0000 679.2400 ;
        RECT 1784.6600 673.3200 1786.2600 673.8000 ;
        RECT 1784.6600 678.7600 1786.2600 679.2400 ;
        RECT 1797.0000 657.0000 1800.0000 657.4800 ;
        RECT 1797.0000 662.4400 1800.0000 662.9200 ;
        RECT 1797.0000 667.8800 1800.0000 668.3600 ;
        RECT 1784.6600 657.0000 1786.2600 657.4800 ;
        RECT 1784.6600 662.4400 1786.2600 662.9200 ;
        RECT 1784.6600 667.8800 1786.2600 668.3600 ;
        RECT 1797.0000 646.1200 1800.0000 646.6000 ;
        RECT 1797.0000 651.5600 1800.0000 652.0400 ;
        RECT 1784.6600 646.1200 1786.2600 646.6000 ;
        RECT 1784.6600 651.5600 1786.2600 652.0400 ;
        RECT 1739.6600 684.2000 1741.2600 684.6800 ;
        RECT 1739.6600 689.6400 1741.2600 690.1200 ;
        RECT 1739.6600 695.0800 1741.2600 695.5600 ;
        RECT 1739.6600 673.3200 1741.2600 673.8000 ;
        RECT 1739.6600 678.7600 1741.2600 679.2400 ;
        RECT 1739.6600 657.0000 1741.2600 657.4800 ;
        RECT 1739.6600 662.4400 1741.2600 662.9200 ;
        RECT 1739.6600 667.8800 1741.2600 668.3600 ;
        RECT 1739.6600 646.1200 1741.2600 646.6000 ;
        RECT 1739.6600 651.5600 1741.2600 652.0400 ;
        RECT 1694.6600 727.7200 1696.2600 728.2000 ;
        RECT 1694.6600 733.1600 1696.2600 733.6400 ;
        RECT 1694.6600 738.6000 1696.2600 739.0800 ;
        RECT 1649.6600 727.7200 1651.2600 728.2000 ;
        RECT 1649.6600 733.1600 1651.2600 733.6400 ;
        RECT 1649.6600 738.6000 1651.2600 739.0800 ;
        RECT 1694.6600 716.8400 1696.2600 717.3200 ;
        RECT 1694.6600 722.2800 1696.2600 722.7600 ;
        RECT 1694.6600 700.5200 1696.2600 701.0000 ;
        RECT 1694.6600 705.9600 1696.2600 706.4400 ;
        RECT 1694.6600 711.4000 1696.2600 711.8800 ;
        RECT 1649.6600 716.8400 1651.2600 717.3200 ;
        RECT 1649.6600 722.2800 1651.2600 722.7600 ;
        RECT 1649.6600 700.5200 1651.2600 701.0000 ;
        RECT 1649.6600 705.9600 1651.2600 706.4400 ;
        RECT 1649.6600 711.4000 1651.2600 711.8800 ;
        RECT 1604.6600 727.7200 1606.2600 728.2000 ;
        RECT 1604.6600 733.1600 1606.2600 733.6400 ;
        RECT 1592.9000 733.1600 1595.9000 733.6400 ;
        RECT 1592.9000 727.7200 1595.9000 728.2000 ;
        RECT 1592.9000 738.6000 1595.9000 739.0800 ;
        RECT 1604.6600 738.6000 1606.2600 739.0800 ;
        RECT 1604.6600 716.8400 1606.2600 717.3200 ;
        RECT 1604.6600 722.2800 1606.2600 722.7600 ;
        RECT 1592.9000 722.2800 1595.9000 722.7600 ;
        RECT 1592.9000 716.8400 1595.9000 717.3200 ;
        RECT 1604.6600 700.5200 1606.2600 701.0000 ;
        RECT 1604.6600 705.9600 1606.2600 706.4400 ;
        RECT 1592.9000 705.9600 1595.9000 706.4400 ;
        RECT 1592.9000 700.5200 1595.9000 701.0000 ;
        RECT 1592.9000 711.4000 1595.9000 711.8800 ;
        RECT 1604.6600 711.4000 1606.2600 711.8800 ;
        RECT 1694.6600 684.2000 1696.2600 684.6800 ;
        RECT 1694.6600 689.6400 1696.2600 690.1200 ;
        RECT 1694.6600 695.0800 1696.2600 695.5600 ;
        RECT 1694.6600 673.3200 1696.2600 673.8000 ;
        RECT 1694.6600 678.7600 1696.2600 679.2400 ;
        RECT 1649.6600 684.2000 1651.2600 684.6800 ;
        RECT 1649.6600 689.6400 1651.2600 690.1200 ;
        RECT 1649.6600 695.0800 1651.2600 695.5600 ;
        RECT 1649.6600 673.3200 1651.2600 673.8000 ;
        RECT 1649.6600 678.7600 1651.2600 679.2400 ;
        RECT 1694.6600 657.0000 1696.2600 657.4800 ;
        RECT 1694.6600 662.4400 1696.2600 662.9200 ;
        RECT 1694.6600 667.8800 1696.2600 668.3600 ;
        RECT 1694.6600 646.1200 1696.2600 646.6000 ;
        RECT 1694.6600 651.5600 1696.2600 652.0400 ;
        RECT 1649.6600 657.0000 1651.2600 657.4800 ;
        RECT 1649.6600 662.4400 1651.2600 662.9200 ;
        RECT 1649.6600 667.8800 1651.2600 668.3600 ;
        RECT 1649.6600 646.1200 1651.2600 646.6000 ;
        RECT 1649.6600 651.5600 1651.2600 652.0400 ;
        RECT 1604.6600 684.2000 1606.2600 684.6800 ;
        RECT 1604.6600 689.6400 1606.2600 690.1200 ;
        RECT 1604.6600 695.0800 1606.2600 695.5600 ;
        RECT 1592.9000 684.2000 1595.9000 684.6800 ;
        RECT 1592.9000 689.6400 1595.9000 690.1200 ;
        RECT 1592.9000 695.0800 1595.9000 695.5600 ;
        RECT 1604.6600 673.3200 1606.2600 673.8000 ;
        RECT 1604.6600 678.7600 1606.2600 679.2400 ;
        RECT 1592.9000 673.3200 1595.9000 673.8000 ;
        RECT 1592.9000 678.7600 1595.9000 679.2400 ;
        RECT 1604.6600 657.0000 1606.2600 657.4800 ;
        RECT 1604.6600 662.4400 1606.2600 662.9200 ;
        RECT 1604.6600 667.8800 1606.2600 668.3600 ;
        RECT 1592.9000 657.0000 1595.9000 657.4800 ;
        RECT 1592.9000 662.4400 1595.9000 662.9200 ;
        RECT 1592.9000 667.8800 1595.9000 668.3600 ;
        RECT 1604.6600 646.1200 1606.2600 646.6000 ;
        RECT 1604.6600 651.5600 1606.2600 652.0400 ;
        RECT 1592.9000 646.1200 1595.9000 646.6000 ;
        RECT 1592.9000 651.5600 1595.9000 652.0400 ;
        RECT 1797.0000 629.8000 1800.0000 630.2800 ;
        RECT 1797.0000 635.2400 1800.0000 635.7200 ;
        RECT 1797.0000 640.6800 1800.0000 641.1600 ;
        RECT 1784.6600 629.8000 1786.2600 630.2800 ;
        RECT 1784.6600 635.2400 1786.2600 635.7200 ;
        RECT 1784.6600 640.6800 1786.2600 641.1600 ;
        RECT 1797.0000 618.9200 1800.0000 619.4000 ;
        RECT 1797.0000 624.3600 1800.0000 624.8400 ;
        RECT 1784.6600 618.9200 1786.2600 619.4000 ;
        RECT 1784.6600 624.3600 1786.2600 624.8400 ;
        RECT 1797.0000 602.6000 1800.0000 603.0800 ;
        RECT 1797.0000 608.0400 1800.0000 608.5200 ;
        RECT 1797.0000 613.4800 1800.0000 613.9600 ;
        RECT 1784.6600 602.6000 1786.2600 603.0800 ;
        RECT 1784.6600 608.0400 1786.2600 608.5200 ;
        RECT 1784.6600 613.4800 1786.2600 613.9600 ;
        RECT 1797.0000 591.7200 1800.0000 592.2000 ;
        RECT 1797.0000 597.1600 1800.0000 597.6400 ;
        RECT 1784.6600 591.7200 1786.2600 592.2000 ;
        RECT 1784.6600 597.1600 1786.2600 597.6400 ;
        RECT 1739.6600 629.8000 1741.2600 630.2800 ;
        RECT 1739.6600 635.2400 1741.2600 635.7200 ;
        RECT 1739.6600 640.6800 1741.2600 641.1600 ;
        RECT 1739.6600 618.9200 1741.2600 619.4000 ;
        RECT 1739.6600 624.3600 1741.2600 624.8400 ;
        RECT 1739.6600 602.6000 1741.2600 603.0800 ;
        RECT 1739.6600 608.0400 1741.2600 608.5200 ;
        RECT 1739.6600 613.4800 1741.2600 613.9600 ;
        RECT 1739.6600 591.7200 1741.2600 592.2000 ;
        RECT 1739.6600 597.1600 1741.2600 597.6400 ;
        RECT 1797.0000 575.4000 1800.0000 575.8800 ;
        RECT 1797.0000 580.8400 1800.0000 581.3200 ;
        RECT 1797.0000 586.2800 1800.0000 586.7600 ;
        RECT 1784.6600 575.4000 1786.2600 575.8800 ;
        RECT 1784.6600 580.8400 1786.2600 581.3200 ;
        RECT 1784.6600 586.2800 1786.2600 586.7600 ;
        RECT 1797.0000 564.5200 1800.0000 565.0000 ;
        RECT 1797.0000 569.9600 1800.0000 570.4400 ;
        RECT 1784.6600 564.5200 1786.2600 565.0000 ;
        RECT 1784.6600 569.9600 1786.2600 570.4400 ;
        RECT 1797.0000 548.2000 1800.0000 548.6800 ;
        RECT 1797.0000 553.6400 1800.0000 554.1200 ;
        RECT 1797.0000 559.0800 1800.0000 559.5600 ;
        RECT 1784.6600 548.2000 1786.2600 548.6800 ;
        RECT 1784.6600 553.6400 1786.2600 554.1200 ;
        RECT 1784.6600 559.0800 1786.2600 559.5600 ;
        RECT 1797.0000 542.7600 1800.0000 543.2400 ;
        RECT 1784.6600 542.7600 1786.2600 543.2400 ;
        RECT 1739.6600 575.4000 1741.2600 575.8800 ;
        RECT 1739.6600 580.8400 1741.2600 581.3200 ;
        RECT 1739.6600 586.2800 1741.2600 586.7600 ;
        RECT 1739.6600 564.5200 1741.2600 565.0000 ;
        RECT 1739.6600 569.9600 1741.2600 570.4400 ;
        RECT 1739.6600 548.2000 1741.2600 548.6800 ;
        RECT 1739.6600 553.6400 1741.2600 554.1200 ;
        RECT 1739.6600 559.0800 1741.2600 559.5600 ;
        RECT 1739.6600 542.7600 1741.2600 543.2400 ;
        RECT 1694.6600 629.8000 1696.2600 630.2800 ;
        RECT 1694.6600 635.2400 1696.2600 635.7200 ;
        RECT 1694.6600 640.6800 1696.2600 641.1600 ;
        RECT 1694.6600 618.9200 1696.2600 619.4000 ;
        RECT 1694.6600 624.3600 1696.2600 624.8400 ;
        RECT 1649.6600 629.8000 1651.2600 630.2800 ;
        RECT 1649.6600 635.2400 1651.2600 635.7200 ;
        RECT 1649.6600 640.6800 1651.2600 641.1600 ;
        RECT 1649.6600 618.9200 1651.2600 619.4000 ;
        RECT 1649.6600 624.3600 1651.2600 624.8400 ;
        RECT 1694.6600 602.6000 1696.2600 603.0800 ;
        RECT 1694.6600 608.0400 1696.2600 608.5200 ;
        RECT 1694.6600 613.4800 1696.2600 613.9600 ;
        RECT 1694.6600 591.7200 1696.2600 592.2000 ;
        RECT 1694.6600 597.1600 1696.2600 597.6400 ;
        RECT 1649.6600 602.6000 1651.2600 603.0800 ;
        RECT 1649.6600 608.0400 1651.2600 608.5200 ;
        RECT 1649.6600 613.4800 1651.2600 613.9600 ;
        RECT 1649.6600 591.7200 1651.2600 592.2000 ;
        RECT 1649.6600 597.1600 1651.2600 597.6400 ;
        RECT 1604.6600 629.8000 1606.2600 630.2800 ;
        RECT 1604.6600 635.2400 1606.2600 635.7200 ;
        RECT 1604.6600 640.6800 1606.2600 641.1600 ;
        RECT 1592.9000 629.8000 1595.9000 630.2800 ;
        RECT 1592.9000 635.2400 1595.9000 635.7200 ;
        RECT 1592.9000 640.6800 1595.9000 641.1600 ;
        RECT 1604.6600 618.9200 1606.2600 619.4000 ;
        RECT 1604.6600 624.3600 1606.2600 624.8400 ;
        RECT 1592.9000 618.9200 1595.9000 619.4000 ;
        RECT 1592.9000 624.3600 1595.9000 624.8400 ;
        RECT 1604.6600 602.6000 1606.2600 603.0800 ;
        RECT 1604.6600 608.0400 1606.2600 608.5200 ;
        RECT 1604.6600 613.4800 1606.2600 613.9600 ;
        RECT 1592.9000 602.6000 1595.9000 603.0800 ;
        RECT 1592.9000 608.0400 1595.9000 608.5200 ;
        RECT 1592.9000 613.4800 1595.9000 613.9600 ;
        RECT 1604.6600 591.7200 1606.2600 592.2000 ;
        RECT 1604.6600 597.1600 1606.2600 597.6400 ;
        RECT 1592.9000 591.7200 1595.9000 592.2000 ;
        RECT 1592.9000 597.1600 1595.9000 597.6400 ;
        RECT 1694.6600 575.4000 1696.2600 575.8800 ;
        RECT 1694.6600 580.8400 1696.2600 581.3200 ;
        RECT 1694.6600 586.2800 1696.2600 586.7600 ;
        RECT 1694.6600 564.5200 1696.2600 565.0000 ;
        RECT 1694.6600 569.9600 1696.2600 570.4400 ;
        RECT 1649.6600 575.4000 1651.2600 575.8800 ;
        RECT 1649.6600 580.8400 1651.2600 581.3200 ;
        RECT 1649.6600 586.2800 1651.2600 586.7600 ;
        RECT 1649.6600 564.5200 1651.2600 565.0000 ;
        RECT 1649.6600 569.9600 1651.2600 570.4400 ;
        RECT 1694.6600 548.2000 1696.2600 548.6800 ;
        RECT 1694.6600 553.6400 1696.2600 554.1200 ;
        RECT 1694.6600 559.0800 1696.2600 559.5600 ;
        RECT 1694.6600 542.7600 1696.2600 543.2400 ;
        RECT 1649.6600 548.2000 1651.2600 548.6800 ;
        RECT 1649.6600 553.6400 1651.2600 554.1200 ;
        RECT 1649.6600 559.0800 1651.2600 559.5600 ;
        RECT 1649.6600 542.7600 1651.2600 543.2400 ;
        RECT 1604.6600 575.4000 1606.2600 575.8800 ;
        RECT 1604.6600 580.8400 1606.2600 581.3200 ;
        RECT 1604.6600 586.2800 1606.2600 586.7600 ;
        RECT 1592.9000 575.4000 1595.9000 575.8800 ;
        RECT 1592.9000 580.8400 1595.9000 581.3200 ;
        RECT 1592.9000 586.2800 1595.9000 586.7600 ;
        RECT 1604.6600 564.5200 1606.2600 565.0000 ;
        RECT 1604.6600 569.9600 1606.2600 570.4400 ;
        RECT 1592.9000 564.5200 1595.9000 565.0000 ;
        RECT 1592.9000 569.9600 1595.9000 570.4400 ;
        RECT 1604.6600 548.2000 1606.2600 548.6800 ;
        RECT 1604.6600 553.6400 1606.2600 554.1200 ;
        RECT 1604.6600 559.0800 1606.2600 559.5600 ;
        RECT 1592.9000 548.2000 1595.9000 548.6800 ;
        RECT 1592.9000 553.6400 1595.9000 554.1200 ;
        RECT 1592.9000 559.0800 1595.9000 559.5600 ;
        RECT 1592.9000 542.7600 1595.9000 543.2400 ;
        RECT 1604.6600 542.7600 1606.2600 543.2400 ;
        RECT 1592.9000 747.6700 1800.0000 750.6700 ;
        RECT 1592.9000 534.5700 1800.0000 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 304.9300 1786.2600 521.0300 ;
        RECT 1739.6600 304.9300 1741.2600 521.0300 ;
        RECT 1694.6600 304.9300 1696.2600 521.0300 ;
        RECT 1649.6600 304.9300 1651.2600 521.0300 ;
        RECT 1604.6600 304.9300 1606.2600 521.0300 ;
        RECT 1797.0000 304.9300 1800.0000 521.0300 ;
        RECT 1592.9000 304.9300 1595.9000 521.0300 ;
      LAYER met3 ;
        RECT 1797.0000 498.0800 1800.0000 498.5600 ;
        RECT 1797.0000 503.5200 1800.0000 504.0000 ;
        RECT 1784.6600 498.0800 1786.2600 498.5600 ;
        RECT 1784.6600 503.5200 1786.2600 504.0000 ;
        RECT 1797.0000 508.9600 1800.0000 509.4400 ;
        RECT 1784.6600 508.9600 1786.2600 509.4400 ;
        RECT 1797.0000 487.2000 1800.0000 487.6800 ;
        RECT 1797.0000 492.6400 1800.0000 493.1200 ;
        RECT 1784.6600 487.2000 1786.2600 487.6800 ;
        RECT 1784.6600 492.6400 1786.2600 493.1200 ;
        RECT 1797.0000 470.8800 1800.0000 471.3600 ;
        RECT 1797.0000 476.3200 1800.0000 476.8000 ;
        RECT 1784.6600 470.8800 1786.2600 471.3600 ;
        RECT 1784.6600 476.3200 1786.2600 476.8000 ;
        RECT 1797.0000 481.7600 1800.0000 482.2400 ;
        RECT 1784.6600 481.7600 1786.2600 482.2400 ;
        RECT 1739.6600 498.0800 1741.2600 498.5600 ;
        RECT 1739.6600 503.5200 1741.2600 504.0000 ;
        RECT 1739.6600 508.9600 1741.2600 509.4400 ;
        RECT 1739.6600 487.2000 1741.2600 487.6800 ;
        RECT 1739.6600 492.6400 1741.2600 493.1200 ;
        RECT 1739.6600 470.8800 1741.2600 471.3600 ;
        RECT 1739.6600 476.3200 1741.2600 476.8000 ;
        RECT 1739.6600 481.7600 1741.2600 482.2400 ;
        RECT 1797.0000 454.5600 1800.0000 455.0400 ;
        RECT 1797.0000 460.0000 1800.0000 460.4800 ;
        RECT 1797.0000 465.4400 1800.0000 465.9200 ;
        RECT 1784.6600 454.5600 1786.2600 455.0400 ;
        RECT 1784.6600 460.0000 1786.2600 460.4800 ;
        RECT 1784.6600 465.4400 1786.2600 465.9200 ;
        RECT 1797.0000 443.6800 1800.0000 444.1600 ;
        RECT 1797.0000 449.1200 1800.0000 449.6000 ;
        RECT 1784.6600 443.6800 1786.2600 444.1600 ;
        RECT 1784.6600 449.1200 1786.2600 449.6000 ;
        RECT 1797.0000 427.3600 1800.0000 427.8400 ;
        RECT 1797.0000 432.8000 1800.0000 433.2800 ;
        RECT 1797.0000 438.2400 1800.0000 438.7200 ;
        RECT 1784.6600 427.3600 1786.2600 427.8400 ;
        RECT 1784.6600 432.8000 1786.2600 433.2800 ;
        RECT 1784.6600 438.2400 1786.2600 438.7200 ;
        RECT 1797.0000 416.4800 1800.0000 416.9600 ;
        RECT 1797.0000 421.9200 1800.0000 422.4000 ;
        RECT 1784.6600 416.4800 1786.2600 416.9600 ;
        RECT 1784.6600 421.9200 1786.2600 422.4000 ;
        RECT 1739.6600 454.5600 1741.2600 455.0400 ;
        RECT 1739.6600 460.0000 1741.2600 460.4800 ;
        RECT 1739.6600 465.4400 1741.2600 465.9200 ;
        RECT 1739.6600 443.6800 1741.2600 444.1600 ;
        RECT 1739.6600 449.1200 1741.2600 449.6000 ;
        RECT 1739.6600 427.3600 1741.2600 427.8400 ;
        RECT 1739.6600 432.8000 1741.2600 433.2800 ;
        RECT 1739.6600 438.2400 1741.2600 438.7200 ;
        RECT 1739.6600 416.4800 1741.2600 416.9600 ;
        RECT 1739.6600 421.9200 1741.2600 422.4000 ;
        RECT 1694.6600 498.0800 1696.2600 498.5600 ;
        RECT 1694.6600 503.5200 1696.2600 504.0000 ;
        RECT 1694.6600 508.9600 1696.2600 509.4400 ;
        RECT 1649.6600 498.0800 1651.2600 498.5600 ;
        RECT 1649.6600 503.5200 1651.2600 504.0000 ;
        RECT 1649.6600 508.9600 1651.2600 509.4400 ;
        RECT 1694.6600 487.2000 1696.2600 487.6800 ;
        RECT 1694.6600 492.6400 1696.2600 493.1200 ;
        RECT 1694.6600 470.8800 1696.2600 471.3600 ;
        RECT 1694.6600 476.3200 1696.2600 476.8000 ;
        RECT 1694.6600 481.7600 1696.2600 482.2400 ;
        RECT 1649.6600 487.2000 1651.2600 487.6800 ;
        RECT 1649.6600 492.6400 1651.2600 493.1200 ;
        RECT 1649.6600 470.8800 1651.2600 471.3600 ;
        RECT 1649.6600 476.3200 1651.2600 476.8000 ;
        RECT 1649.6600 481.7600 1651.2600 482.2400 ;
        RECT 1604.6600 498.0800 1606.2600 498.5600 ;
        RECT 1604.6600 503.5200 1606.2600 504.0000 ;
        RECT 1592.9000 503.5200 1595.9000 504.0000 ;
        RECT 1592.9000 498.0800 1595.9000 498.5600 ;
        RECT 1592.9000 508.9600 1595.9000 509.4400 ;
        RECT 1604.6600 508.9600 1606.2600 509.4400 ;
        RECT 1604.6600 487.2000 1606.2600 487.6800 ;
        RECT 1604.6600 492.6400 1606.2600 493.1200 ;
        RECT 1592.9000 492.6400 1595.9000 493.1200 ;
        RECT 1592.9000 487.2000 1595.9000 487.6800 ;
        RECT 1604.6600 470.8800 1606.2600 471.3600 ;
        RECT 1604.6600 476.3200 1606.2600 476.8000 ;
        RECT 1592.9000 476.3200 1595.9000 476.8000 ;
        RECT 1592.9000 470.8800 1595.9000 471.3600 ;
        RECT 1592.9000 481.7600 1595.9000 482.2400 ;
        RECT 1604.6600 481.7600 1606.2600 482.2400 ;
        RECT 1694.6600 454.5600 1696.2600 455.0400 ;
        RECT 1694.6600 460.0000 1696.2600 460.4800 ;
        RECT 1694.6600 465.4400 1696.2600 465.9200 ;
        RECT 1694.6600 443.6800 1696.2600 444.1600 ;
        RECT 1694.6600 449.1200 1696.2600 449.6000 ;
        RECT 1649.6600 454.5600 1651.2600 455.0400 ;
        RECT 1649.6600 460.0000 1651.2600 460.4800 ;
        RECT 1649.6600 465.4400 1651.2600 465.9200 ;
        RECT 1649.6600 443.6800 1651.2600 444.1600 ;
        RECT 1649.6600 449.1200 1651.2600 449.6000 ;
        RECT 1694.6600 427.3600 1696.2600 427.8400 ;
        RECT 1694.6600 432.8000 1696.2600 433.2800 ;
        RECT 1694.6600 438.2400 1696.2600 438.7200 ;
        RECT 1694.6600 416.4800 1696.2600 416.9600 ;
        RECT 1694.6600 421.9200 1696.2600 422.4000 ;
        RECT 1649.6600 427.3600 1651.2600 427.8400 ;
        RECT 1649.6600 432.8000 1651.2600 433.2800 ;
        RECT 1649.6600 438.2400 1651.2600 438.7200 ;
        RECT 1649.6600 416.4800 1651.2600 416.9600 ;
        RECT 1649.6600 421.9200 1651.2600 422.4000 ;
        RECT 1604.6600 454.5600 1606.2600 455.0400 ;
        RECT 1604.6600 460.0000 1606.2600 460.4800 ;
        RECT 1604.6600 465.4400 1606.2600 465.9200 ;
        RECT 1592.9000 454.5600 1595.9000 455.0400 ;
        RECT 1592.9000 460.0000 1595.9000 460.4800 ;
        RECT 1592.9000 465.4400 1595.9000 465.9200 ;
        RECT 1604.6600 443.6800 1606.2600 444.1600 ;
        RECT 1604.6600 449.1200 1606.2600 449.6000 ;
        RECT 1592.9000 443.6800 1595.9000 444.1600 ;
        RECT 1592.9000 449.1200 1595.9000 449.6000 ;
        RECT 1604.6600 427.3600 1606.2600 427.8400 ;
        RECT 1604.6600 432.8000 1606.2600 433.2800 ;
        RECT 1604.6600 438.2400 1606.2600 438.7200 ;
        RECT 1592.9000 427.3600 1595.9000 427.8400 ;
        RECT 1592.9000 432.8000 1595.9000 433.2800 ;
        RECT 1592.9000 438.2400 1595.9000 438.7200 ;
        RECT 1604.6600 416.4800 1606.2600 416.9600 ;
        RECT 1604.6600 421.9200 1606.2600 422.4000 ;
        RECT 1592.9000 416.4800 1595.9000 416.9600 ;
        RECT 1592.9000 421.9200 1595.9000 422.4000 ;
        RECT 1797.0000 400.1600 1800.0000 400.6400 ;
        RECT 1797.0000 405.6000 1800.0000 406.0800 ;
        RECT 1797.0000 411.0400 1800.0000 411.5200 ;
        RECT 1784.6600 400.1600 1786.2600 400.6400 ;
        RECT 1784.6600 405.6000 1786.2600 406.0800 ;
        RECT 1784.6600 411.0400 1786.2600 411.5200 ;
        RECT 1797.0000 389.2800 1800.0000 389.7600 ;
        RECT 1797.0000 394.7200 1800.0000 395.2000 ;
        RECT 1784.6600 389.2800 1786.2600 389.7600 ;
        RECT 1784.6600 394.7200 1786.2600 395.2000 ;
        RECT 1797.0000 372.9600 1800.0000 373.4400 ;
        RECT 1797.0000 378.4000 1800.0000 378.8800 ;
        RECT 1797.0000 383.8400 1800.0000 384.3200 ;
        RECT 1784.6600 372.9600 1786.2600 373.4400 ;
        RECT 1784.6600 378.4000 1786.2600 378.8800 ;
        RECT 1784.6600 383.8400 1786.2600 384.3200 ;
        RECT 1797.0000 362.0800 1800.0000 362.5600 ;
        RECT 1797.0000 367.5200 1800.0000 368.0000 ;
        RECT 1784.6600 362.0800 1786.2600 362.5600 ;
        RECT 1784.6600 367.5200 1786.2600 368.0000 ;
        RECT 1739.6600 400.1600 1741.2600 400.6400 ;
        RECT 1739.6600 405.6000 1741.2600 406.0800 ;
        RECT 1739.6600 411.0400 1741.2600 411.5200 ;
        RECT 1739.6600 389.2800 1741.2600 389.7600 ;
        RECT 1739.6600 394.7200 1741.2600 395.2000 ;
        RECT 1739.6600 372.9600 1741.2600 373.4400 ;
        RECT 1739.6600 378.4000 1741.2600 378.8800 ;
        RECT 1739.6600 383.8400 1741.2600 384.3200 ;
        RECT 1739.6600 362.0800 1741.2600 362.5600 ;
        RECT 1739.6600 367.5200 1741.2600 368.0000 ;
        RECT 1797.0000 345.7600 1800.0000 346.2400 ;
        RECT 1797.0000 351.2000 1800.0000 351.6800 ;
        RECT 1797.0000 356.6400 1800.0000 357.1200 ;
        RECT 1784.6600 345.7600 1786.2600 346.2400 ;
        RECT 1784.6600 351.2000 1786.2600 351.6800 ;
        RECT 1784.6600 356.6400 1786.2600 357.1200 ;
        RECT 1797.0000 334.8800 1800.0000 335.3600 ;
        RECT 1797.0000 340.3200 1800.0000 340.8000 ;
        RECT 1784.6600 334.8800 1786.2600 335.3600 ;
        RECT 1784.6600 340.3200 1786.2600 340.8000 ;
        RECT 1797.0000 318.5600 1800.0000 319.0400 ;
        RECT 1797.0000 324.0000 1800.0000 324.4800 ;
        RECT 1797.0000 329.4400 1800.0000 329.9200 ;
        RECT 1784.6600 318.5600 1786.2600 319.0400 ;
        RECT 1784.6600 324.0000 1786.2600 324.4800 ;
        RECT 1784.6600 329.4400 1786.2600 329.9200 ;
        RECT 1797.0000 313.1200 1800.0000 313.6000 ;
        RECT 1784.6600 313.1200 1786.2600 313.6000 ;
        RECT 1739.6600 345.7600 1741.2600 346.2400 ;
        RECT 1739.6600 351.2000 1741.2600 351.6800 ;
        RECT 1739.6600 356.6400 1741.2600 357.1200 ;
        RECT 1739.6600 334.8800 1741.2600 335.3600 ;
        RECT 1739.6600 340.3200 1741.2600 340.8000 ;
        RECT 1739.6600 318.5600 1741.2600 319.0400 ;
        RECT 1739.6600 324.0000 1741.2600 324.4800 ;
        RECT 1739.6600 329.4400 1741.2600 329.9200 ;
        RECT 1739.6600 313.1200 1741.2600 313.6000 ;
        RECT 1694.6600 400.1600 1696.2600 400.6400 ;
        RECT 1694.6600 405.6000 1696.2600 406.0800 ;
        RECT 1694.6600 411.0400 1696.2600 411.5200 ;
        RECT 1694.6600 389.2800 1696.2600 389.7600 ;
        RECT 1694.6600 394.7200 1696.2600 395.2000 ;
        RECT 1649.6600 400.1600 1651.2600 400.6400 ;
        RECT 1649.6600 405.6000 1651.2600 406.0800 ;
        RECT 1649.6600 411.0400 1651.2600 411.5200 ;
        RECT 1649.6600 389.2800 1651.2600 389.7600 ;
        RECT 1649.6600 394.7200 1651.2600 395.2000 ;
        RECT 1694.6600 372.9600 1696.2600 373.4400 ;
        RECT 1694.6600 378.4000 1696.2600 378.8800 ;
        RECT 1694.6600 383.8400 1696.2600 384.3200 ;
        RECT 1694.6600 362.0800 1696.2600 362.5600 ;
        RECT 1694.6600 367.5200 1696.2600 368.0000 ;
        RECT 1649.6600 372.9600 1651.2600 373.4400 ;
        RECT 1649.6600 378.4000 1651.2600 378.8800 ;
        RECT 1649.6600 383.8400 1651.2600 384.3200 ;
        RECT 1649.6600 362.0800 1651.2600 362.5600 ;
        RECT 1649.6600 367.5200 1651.2600 368.0000 ;
        RECT 1604.6600 400.1600 1606.2600 400.6400 ;
        RECT 1604.6600 405.6000 1606.2600 406.0800 ;
        RECT 1604.6600 411.0400 1606.2600 411.5200 ;
        RECT 1592.9000 400.1600 1595.9000 400.6400 ;
        RECT 1592.9000 405.6000 1595.9000 406.0800 ;
        RECT 1592.9000 411.0400 1595.9000 411.5200 ;
        RECT 1604.6600 389.2800 1606.2600 389.7600 ;
        RECT 1604.6600 394.7200 1606.2600 395.2000 ;
        RECT 1592.9000 389.2800 1595.9000 389.7600 ;
        RECT 1592.9000 394.7200 1595.9000 395.2000 ;
        RECT 1604.6600 372.9600 1606.2600 373.4400 ;
        RECT 1604.6600 378.4000 1606.2600 378.8800 ;
        RECT 1604.6600 383.8400 1606.2600 384.3200 ;
        RECT 1592.9000 372.9600 1595.9000 373.4400 ;
        RECT 1592.9000 378.4000 1595.9000 378.8800 ;
        RECT 1592.9000 383.8400 1595.9000 384.3200 ;
        RECT 1604.6600 362.0800 1606.2600 362.5600 ;
        RECT 1604.6600 367.5200 1606.2600 368.0000 ;
        RECT 1592.9000 362.0800 1595.9000 362.5600 ;
        RECT 1592.9000 367.5200 1595.9000 368.0000 ;
        RECT 1694.6600 345.7600 1696.2600 346.2400 ;
        RECT 1694.6600 351.2000 1696.2600 351.6800 ;
        RECT 1694.6600 356.6400 1696.2600 357.1200 ;
        RECT 1694.6600 334.8800 1696.2600 335.3600 ;
        RECT 1694.6600 340.3200 1696.2600 340.8000 ;
        RECT 1649.6600 345.7600 1651.2600 346.2400 ;
        RECT 1649.6600 351.2000 1651.2600 351.6800 ;
        RECT 1649.6600 356.6400 1651.2600 357.1200 ;
        RECT 1649.6600 334.8800 1651.2600 335.3600 ;
        RECT 1649.6600 340.3200 1651.2600 340.8000 ;
        RECT 1694.6600 318.5600 1696.2600 319.0400 ;
        RECT 1694.6600 324.0000 1696.2600 324.4800 ;
        RECT 1694.6600 329.4400 1696.2600 329.9200 ;
        RECT 1694.6600 313.1200 1696.2600 313.6000 ;
        RECT 1649.6600 318.5600 1651.2600 319.0400 ;
        RECT 1649.6600 324.0000 1651.2600 324.4800 ;
        RECT 1649.6600 329.4400 1651.2600 329.9200 ;
        RECT 1649.6600 313.1200 1651.2600 313.6000 ;
        RECT 1604.6600 345.7600 1606.2600 346.2400 ;
        RECT 1604.6600 351.2000 1606.2600 351.6800 ;
        RECT 1604.6600 356.6400 1606.2600 357.1200 ;
        RECT 1592.9000 345.7600 1595.9000 346.2400 ;
        RECT 1592.9000 351.2000 1595.9000 351.6800 ;
        RECT 1592.9000 356.6400 1595.9000 357.1200 ;
        RECT 1604.6600 334.8800 1606.2600 335.3600 ;
        RECT 1604.6600 340.3200 1606.2600 340.8000 ;
        RECT 1592.9000 334.8800 1595.9000 335.3600 ;
        RECT 1592.9000 340.3200 1595.9000 340.8000 ;
        RECT 1604.6600 318.5600 1606.2600 319.0400 ;
        RECT 1604.6600 324.0000 1606.2600 324.4800 ;
        RECT 1604.6600 329.4400 1606.2600 329.9200 ;
        RECT 1592.9000 318.5600 1595.9000 319.0400 ;
        RECT 1592.9000 324.0000 1595.9000 324.4800 ;
        RECT 1592.9000 329.4400 1595.9000 329.9200 ;
        RECT 1592.9000 313.1200 1595.9000 313.6000 ;
        RECT 1604.6600 313.1200 1606.2600 313.6000 ;
        RECT 1592.9000 518.0300 1800.0000 521.0300 ;
        RECT 1592.9000 304.9300 1800.0000 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 75.2900 1786.2600 291.3900 ;
        RECT 1739.6600 75.2900 1741.2600 291.3900 ;
        RECT 1694.6600 75.2900 1696.2600 291.3900 ;
        RECT 1649.6600 75.2900 1651.2600 291.3900 ;
        RECT 1604.6600 75.2900 1606.2600 291.3900 ;
        RECT 1797.0000 75.2900 1800.0000 291.3900 ;
        RECT 1592.9000 75.2900 1595.9000 291.3900 ;
      LAYER met3 ;
        RECT 1797.0000 268.4400 1800.0000 268.9200 ;
        RECT 1797.0000 273.8800 1800.0000 274.3600 ;
        RECT 1784.6600 268.4400 1786.2600 268.9200 ;
        RECT 1784.6600 273.8800 1786.2600 274.3600 ;
        RECT 1797.0000 279.3200 1800.0000 279.8000 ;
        RECT 1784.6600 279.3200 1786.2600 279.8000 ;
        RECT 1797.0000 257.5600 1800.0000 258.0400 ;
        RECT 1797.0000 263.0000 1800.0000 263.4800 ;
        RECT 1784.6600 257.5600 1786.2600 258.0400 ;
        RECT 1784.6600 263.0000 1786.2600 263.4800 ;
        RECT 1797.0000 241.2400 1800.0000 241.7200 ;
        RECT 1797.0000 246.6800 1800.0000 247.1600 ;
        RECT 1784.6600 241.2400 1786.2600 241.7200 ;
        RECT 1784.6600 246.6800 1786.2600 247.1600 ;
        RECT 1797.0000 252.1200 1800.0000 252.6000 ;
        RECT 1784.6600 252.1200 1786.2600 252.6000 ;
        RECT 1739.6600 268.4400 1741.2600 268.9200 ;
        RECT 1739.6600 273.8800 1741.2600 274.3600 ;
        RECT 1739.6600 279.3200 1741.2600 279.8000 ;
        RECT 1739.6600 257.5600 1741.2600 258.0400 ;
        RECT 1739.6600 263.0000 1741.2600 263.4800 ;
        RECT 1739.6600 241.2400 1741.2600 241.7200 ;
        RECT 1739.6600 246.6800 1741.2600 247.1600 ;
        RECT 1739.6600 252.1200 1741.2600 252.6000 ;
        RECT 1797.0000 224.9200 1800.0000 225.4000 ;
        RECT 1797.0000 230.3600 1800.0000 230.8400 ;
        RECT 1797.0000 235.8000 1800.0000 236.2800 ;
        RECT 1784.6600 224.9200 1786.2600 225.4000 ;
        RECT 1784.6600 230.3600 1786.2600 230.8400 ;
        RECT 1784.6600 235.8000 1786.2600 236.2800 ;
        RECT 1797.0000 214.0400 1800.0000 214.5200 ;
        RECT 1797.0000 219.4800 1800.0000 219.9600 ;
        RECT 1784.6600 214.0400 1786.2600 214.5200 ;
        RECT 1784.6600 219.4800 1786.2600 219.9600 ;
        RECT 1797.0000 197.7200 1800.0000 198.2000 ;
        RECT 1797.0000 203.1600 1800.0000 203.6400 ;
        RECT 1797.0000 208.6000 1800.0000 209.0800 ;
        RECT 1784.6600 197.7200 1786.2600 198.2000 ;
        RECT 1784.6600 203.1600 1786.2600 203.6400 ;
        RECT 1784.6600 208.6000 1786.2600 209.0800 ;
        RECT 1797.0000 186.8400 1800.0000 187.3200 ;
        RECT 1797.0000 192.2800 1800.0000 192.7600 ;
        RECT 1784.6600 186.8400 1786.2600 187.3200 ;
        RECT 1784.6600 192.2800 1786.2600 192.7600 ;
        RECT 1739.6600 224.9200 1741.2600 225.4000 ;
        RECT 1739.6600 230.3600 1741.2600 230.8400 ;
        RECT 1739.6600 235.8000 1741.2600 236.2800 ;
        RECT 1739.6600 214.0400 1741.2600 214.5200 ;
        RECT 1739.6600 219.4800 1741.2600 219.9600 ;
        RECT 1739.6600 197.7200 1741.2600 198.2000 ;
        RECT 1739.6600 203.1600 1741.2600 203.6400 ;
        RECT 1739.6600 208.6000 1741.2600 209.0800 ;
        RECT 1739.6600 186.8400 1741.2600 187.3200 ;
        RECT 1739.6600 192.2800 1741.2600 192.7600 ;
        RECT 1694.6600 268.4400 1696.2600 268.9200 ;
        RECT 1694.6600 273.8800 1696.2600 274.3600 ;
        RECT 1694.6600 279.3200 1696.2600 279.8000 ;
        RECT 1649.6600 268.4400 1651.2600 268.9200 ;
        RECT 1649.6600 273.8800 1651.2600 274.3600 ;
        RECT 1649.6600 279.3200 1651.2600 279.8000 ;
        RECT 1694.6600 257.5600 1696.2600 258.0400 ;
        RECT 1694.6600 263.0000 1696.2600 263.4800 ;
        RECT 1694.6600 241.2400 1696.2600 241.7200 ;
        RECT 1694.6600 246.6800 1696.2600 247.1600 ;
        RECT 1694.6600 252.1200 1696.2600 252.6000 ;
        RECT 1649.6600 257.5600 1651.2600 258.0400 ;
        RECT 1649.6600 263.0000 1651.2600 263.4800 ;
        RECT 1649.6600 241.2400 1651.2600 241.7200 ;
        RECT 1649.6600 246.6800 1651.2600 247.1600 ;
        RECT 1649.6600 252.1200 1651.2600 252.6000 ;
        RECT 1604.6600 268.4400 1606.2600 268.9200 ;
        RECT 1604.6600 273.8800 1606.2600 274.3600 ;
        RECT 1592.9000 273.8800 1595.9000 274.3600 ;
        RECT 1592.9000 268.4400 1595.9000 268.9200 ;
        RECT 1592.9000 279.3200 1595.9000 279.8000 ;
        RECT 1604.6600 279.3200 1606.2600 279.8000 ;
        RECT 1604.6600 257.5600 1606.2600 258.0400 ;
        RECT 1604.6600 263.0000 1606.2600 263.4800 ;
        RECT 1592.9000 263.0000 1595.9000 263.4800 ;
        RECT 1592.9000 257.5600 1595.9000 258.0400 ;
        RECT 1604.6600 241.2400 1606.2600 241.7200 ;
        RECT 1604.6600 246.6800 1606.2600 247.1600 ;
        RECT 1592.9000 246.6800 1595.9000 247.1600 ;
        RECT 1592.9000 241.2400 1595.9000 241.7200 ;
        RECT 1592.9000 252.1200 1595.9000 252.6000 ;
        RECT 1604.6600 252.1200 1606.2600 252.6000 ;
        RECT 1694.6600 224.9200 1696.2600 225.4000 ;
        RECT 1694.6600 230.3600 1696.2600 230.8400 ;
        RECT 1694.6600 235.8000 1696.2600 236.2800 ;
        RECT 1694.6600 214.0400 1696.2600 214.5200 ;
        RECT 1694.6600 219.4800 1696.2600 219.9600 ;
        RECT 1649.6600 224.9200 1651.2600 225.4000 ;
        RECT 1649.6600 230.3600 1651.2600 230.8400 ;
        RECT 1649.6600 235.8000 1651.2600 236.2800 ;
        RECT 1649.6600 214.0400 1651.2600 214.5200 ;
        RECT 1649.6600 219.4800 1651.2600 219.9600 ;
        RECT 1694.6600 197.7200 1696.2600 198.2000 ;
        RECT 1694.6600 203.1600 1696.2600 203.6400 ;
        RECT 1694.6600 208.6000 1696.2600 209.0800 ;
        RECT 1694.6600 186.8400 1696.2600 187.3200 ;
        RECT 1694.6600 192.2800 1696.2600 192.7600 ;
        RECT 1649.6600 197.7200 1651.2600 198.2000 ;
        RECT 1649.6600 203.1600 1651.2600 203.6400 ;
        RECT 1649.6600 208.6000 1651.2600 209.0800 ;
        RECT 1649.6600 186.8400 1651.2600 187.3200 ;
        RECT 1649.6600 192.2800 1651.2600 192.7600 ;
        RECT 1604.6600 224.9200 1606.2600 225.4000 ;
        RECT 1604.6600 230.3600 1606.2600 230.8400 ;
        RECT 1604.6600 235.8000 1606.2600 236.2800 ;
        RECT 1592.9000 224.9200 1595.9000 225.4000 ;
        RECT 1592.9000 230.3600 1595.9000 230.8400 ;
        RECT 1592.9000 235.8000 1595.9000 236.2800 ;
        RECT 1604.6600 214.0400 1606.2600 214.5200 ;
        RECT 1604.6600 219.4800 1606.2600 219.9600 ;
        RECT 1592.9000 214.0400 1595.9000 214.5200 ;
        RECT 1592.9000 219.4800 1595.9000 219.9600 ;
        RECT 1604.6600 197.7200 1606.2600 198.2000 ;
        RECT 1604.6600 203.1600 1606.2600 203.6400 ;
        RECT 1604.6600 208.6000 1606.2600 209.0800 ;
        RECT 1592.9000 197.7200 1595.9000 198.2000 ;
        RECT 1592.9000 203.1600 1595.9000 203.6400 ;
        RECT 1592.9000 208.6000 1595.9000 209.0800 ;
        RECT 1604.6600 186.8400 1606.2600 187.3200 ;
        RECT 1604.6600 192.2800 1606.2600 192.7600 ;
        RECT 1592.9000 186.8400 1595.9000 187.3200 ;
        RECT 1592.9000 192.2800 1595.9000 192.7600 ;
        RECT 1797.0000 170.5200 1800.0000 171.0000 ;
        RECT 1797.0000 175.9600 1800.0000 176.4400 ;
        RECT 1797.0000 181.4000 1800.0000 181.8800 ;
        RECT 1784.6600 170.5200 1786.2600 171.0000 ;
        RECT 1784.6600 175.9600 1786.2600 176.4400 ;
        RECT 1784.6600 181.4000 1786.2600 181.8800 ;
        RECT 1797.0000 159.6400 1800.0000 160.1200 ;
        RECT 1797.0000 165.0800 1800.0000 165.5600 ;
        RECT 1784.6600 159.6400 1786.2600 160.1200 ;
        RECT 1784.6600 165.0800 1786.2600 165.5600 ;
        RECT 1797.0000 143.3200 1800.0000 143.8000 ;
        RECT 1797.0000 148.7600 1800.0000 149.2400 ;
        RECT 1797.0000 154.2000 1800.0000 154.6800 ;
        RECT 1784.6600 143.3200 1786.2600 143.8000 ;
        RECT 1784.6600 148.7600 1786.2600 149.2400 ;
        RECT 1784.6600 154.2000 1786.2600 154.6800 ;
        RECT 1797.0000 132.4400 1800.0000 132.9200 ;
        RECT 1797.0000 137.8800 1800.0000 138.3600 ;
        RECT 1784.6600 132.4400 1786.2600 132.9200 ;
        RECT 1784.6600 137.8800 1786.2600 138.3600 ;
        RECT 1739.6600 170.5200 1741.2600 171.0000 ;
        RECT 1739.6600 175.9600 1741.2600 176.4400 ;
        RECT 1739.6600 181.4000 1741.2600 181.8800 ;
        RECT 1739.6600 159.6400 1741.2600 160.1200 ;
        RECT 1739.6600 165.0800 1741.2600 165.5600 ;
        RECT 1739.6600 143.3200 1741.2600 143.8000 ;
        RECT 1739.6600 148.7600 1741.2600 149.2400 ;
        RECT 1739.6600 154.2000 1741.2600 154.6800 ;
        RECT 1739.6600 132.4400 1741.2600 132.9200 ;
        RECT 1739.6600 137.8800 1741.2600 138.3600 ;
        RECT 1797.0000 116.1200 1800.0000 116.6000 ;
        RECT 1797.0000 121.5600 1800.0000 122.0400 ;
        RECT 1797.0000 127.0000 1800.0000 127.4800 ;
        RECT 1784.6600 116.1200 1786.2600 116.6000 ;
        RECT 1784.6600 121.5600 1786.2600 122.0400 ;
        RECT 1784.6600 127.0000 1786.2600 127.4800 ;
        RECT 1797.0000 105.2400 1800.0000 105.7200 ;
        RECT 1797.0000 110.6800 1800.0000 111.1600 ;
        RECT 1784.6600 105.2400 1786.2600 105.7200 ;
        RECT 1784.6600 110.6800 1786.2600 111.1600 ;
        RECT 1797.0000 88.9200 1800.0000 89.4000 ;
        RECT 1797.0000 94.3600 1800.0000 94.8400 ;
        RECT 1797.0000 99.8000 1800.0000 100.2800 ;
        RECT 1784.6600 88.9200 1786.2600 89.4000 ;
        RECT 1784.6600 94.3600 1786.2600 94.8400 ;
        RECT 1784.6600 99.8000 1786.2600 100.2800 ;
        RECT 1797.0000 83.4800 1800.0000 83.9600 ;
        RECT 1784.6600 83.4800 1786.2600 83.9600 ;
        RECT 1739.6600 116.1200 1741.2600 116.6000 ;
        RECT 1739.6600 121.5600 1741.2600 122.0400 ;
        RECT 1739.6600 127.0000 1741.2600 127.4800 ;
        RECT 1739.6600 105.2400 1741.2600 105.7200 ;
        RECT 1739.6600 110.6800 1741.2600 111.1600 ;
        RECT 1739.6600 88.9200 1741.2600 89.4000 ;
        RECT 1739.6600 94.3600 1741.2600 94.8400 ;
        RECT 1739.6600 99.8000 1741.2600 100.2800 ;
        RECT 1739.6600 83.4800 1741.2600 83.9600 ;
        RECT 1694.6600 170.5200 1696.2600 171.0000 ;
        RECT 1694.6600 175.9600 1696.2600 176.4400 ;
        RECT 1694.6600 181.4000 1696.2600 181.8800 ;
        RECT 1694.6600 159.6400 1696.2600 160.1200 ;
        RECT 1694.6600 165.0800 1696.2600 165.5600 ;
        RECT 1649.6600 170.5200 1651.2600 171.0000 ;
        RECT 1649.6600 175.9600 1651.2600 176.4400 ;
        RECT 1649.6600 181.4000 1651.2600 181.8800 ;
        RECT 1649.6600 159.6400 1651.2600 160.1200 ;
        RECT 1649.6600 165.0800 1651.2600 165.5600 ;
        RECT 1694.6600 143.3200 1696.2600 143.8000 ;
        RECT 1694.6600 148.7600 1696.2600 149.2400 ;
        RECT 1694.6600 154.2000 1696.2600 154.6800 ;
        RECT 1694.6600 132.4400 1696.2600 132.9200 ;
        RECT 1694.6600 137.8800 1696.2600 138.3600 ;
        RECT 1649.6600 143.3200 1651.2600 143.8000 ;
        RECT 1649.6600 148.7600 1651.2600 149.2400 ;
        RECT 1649.6600 154.2000 1651.2600 154.6800 ;
        RECT 1649.6600 132.4400 1651.2600 132.9200 ;
        RECT 1649.6600 137.8800 1651.2600 138.3600 ;
        RECT 1604.6600 170.5200 1606.2600 171.0000 ;
        RECT 1604.6600 175.9600 1606.2600 176.4400 ;
        RECT 1604.6600 181.4000 1606.2600 181.8800 ;
        RECT 1592.9000 170.5200 1595.9000 171.0000 ;
        RECT 1592.9000 175.9600 1595.9000 176.4400 ;
        RECT 1592.9000 181.4000 1595.9000 181.8800 ;
        RECT 1604.6600 159.6400 1606.2600 160.1200 ;
        RECT 1604.6600 165.0800 1606.2600 165.5600 ;
        RECT 1592.9000 159.6400 1595.9000 160.1200 ;
        RECT 1592.9000 165.0800 1595.9000 165.5600 ;
        RECT 1604.6600 143.3200 1606.2600 143.8000 ;
        RECT 1604.6600 148.7600 1606.2600 149.2400 ;
        RECT 1604.6600 154.2000 1606.2600 154.6800 ;
        RECT 1592.9000 143.3200 1595.9000 143.8000 ;
        RECT 1592.9000 148.7600 1595.9000 149.2400 ;
        RECT 1592.9000 154.2000 1595.9000 154.6800 ;
        RECT 1604.6600 132.4400 1606.2600 132.9200 ;
        RECT 1604.6600 137.8800 1606.2600 138.3600 ;
        RECT 1592.9000 132.4400 1595.9000 132.9200 ;
        RECT 1592.9000 137.8800 1595.9000 138.3600 ;
        RECT 1694.6600 116.1200 1696.2600 116.6000 ;
        RECT 1694.6600 121.5600 1696.2600 122.0400 ;
        RECT 1694.6600 127.0000 1696.2600 127.4800 ;
        RECT 1694.6600 105.2400 1696.2600 105.7200 ;
        RECT 1694.6600 110.6800 1696.2600 111.1600 ;
        RECT 1649.6600 116.1200 1651.2600 116.6000 ;
        RECT 1649.6600 121.5600 1651.2600 122.0400 ;
        RECT 1649.6600 127.0000 1651.2600 127.4800 ;
        RECT 1649.6600 105.2400 1651.2600 105.7200 ;
        RECT 1649.6600 110.6800 1651.2600 111.1600 ;
        RECT 1694.6600 88.9200 1696.2600 89.4000 ;
        RECT 1694.6600 94.3600 1696.2600 94.8400 ;
        RECT 1694.6600 99.8000 1696.2600 100.2800 ;
        RECT 1694.6600 83.4800 1696.2600 83.9600 ;
        RECT 1649.6600 88.9200 1651.2600 89.4000 ;
        RECT 1649.6600 94.3600 1651.2600 94.8400 ;
        RECT 1649.6600 99.8000 1651.2600 100.2800 ;
        RECT 1649.6600 83.4800 1651.2600 83.9600 ;
        RECT 1604.6600 116.1200 1606.2600 116.6000 ;
        RECT 1604.6600 121.5600 1606.2600 122.0400 ;
        RECT 1604.6600 127.0000 1606.2600 127.4800 ;
        RECT 1592.9000 116.1200 1595.9000 116.6000 ;
        RECT 1592.9000 121.5600 1595.9000 122.0400 ;
        RECT 1592.9000 127.0000 1595.9000 127.4800 ;
        RECT 1604.6600 105.2400 1606.2600 105.7200 ;
        RECT 1604.6600 110.6800 1606.2600 111.1600 ;
        RECT 1592.9000 105.2400 1595.9000 105.7200 ;
        RECT 1592.9000 110.6800 1595.9000 111.1600 ;
        RECT 1604.6600 88.9200 1606.2600 89.4000 ;
        RECT 1604.6600 94.3600 1606.2600 94.8400 ;
        RECT 1604.6600 99.8000 1606.2600 100.2800 ;
        RECT 1592.9000 88.9200 1595.9000 89.4000 ;
        RECT 1592.9000 94.3600 1595.9000 94.8400 ;
        RECT 1592.9000 99.8000 1595.9000 100.2800 ;
        RECT 1592.9000 83.4800 1595.9000 83.9600 ;
        RECT 1604.6600 83.4800 1606.2600 83.9600 ;
        RECT 1592.9000 288.3900 1800.0000 291.3900 ;
        RECT 1592.9000 75.2900 1800.0000 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1593.9000 34.6700 1595.9000 61.6000 ;
        RECT 1797.0000 34.6700 1799.0000 61.6000 ;
      LAYER met3 ;
        RECT 1797.0000 51.3800 1799.0000 51.8600 ;
        RECT 1593.9000 51.3800 1595.9000 51.8600 ;
        RECT 1797.0000 45.9400 1799.0000 46.4200 ;
        RECT 1797.0000 40.5000 1799.0000 40.9800 ;
        RECT 1593.9000 45.9400 1595.9000 46.4200 ;
        RECT 1593.9000 40.5000 1595.9000 40.9800 ;
        RECT 1593.9000 59.6000 1799.0000 61.6000 ;
        RECT 1593.9000 34.6700 1799.0000 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 2601.3300 1786.2600 2817.4300 ;
        RECT 1739.6600 2601.3300 1741.2600 2817.4300 ;
        RECT 1694.6600 2601.3300 1696.2600 2817.4300 ;
        RECT 1649.6600 2601.3300 1651.2600 2817.4300 ;
        RECT 1604.6600 2601.3300 1606.2600 2817.4300 ;
        RECT 1797.0000 2601.3300 1800.0000 2817.4300 ;
        RECT 1592.9000 2601.3300 1595.9000 2817.4300 ;
      LAYER met3 ;
        RECT 1797.0000 2794.4800 1800.0000 2794.9600 ;
        RECT 1797.0000 2799.9200 1800.0000 2800.4000 ;
        RECT 1784.6600 2794.4800 1786.2600 2794.9600 ;
        RECT 1784.6600 2799.9200 1786.2600 2800.4000 ;
        RECT 1797.0000 2805.3600 1800.0000 2805.8400 ;
        RECT 1784.6600 2805.3600 1786.2600 2805.8400 ;
        RECT 1797.0000 2783.6000 1800.0000 2784.0800 ;
        RECT 1797.0000 2789.0400 1800.0000 2789.5200 ;
        RECT 1784.6600 2783.6000 1786.2600 2784.0800 ;
        RECT 1784.6600 2789.0400 1786.2600 2789.5200 ;
        RECT 1797.0000 2767.2800 1800.0000 2767.7600 ;
        RECT 1797.0000 2772.7200 1800.0000 2773.2000 ;
        RECT 1784.6600 2767.2800 1786.2600 2767.7600 ;
        RECT 1784.6600 2772.7200 1786.2600 2773.2000 ;
        RECT 1797.0000 2778.1600 1800.0000 2778.6400 ;
        RECT 1784.6600 2778.1600 1786.2600 2778.6400 ;
        RECT 1739.6600 2794.4800 1741.2600 2794.9600 ;
        RECT 1739.6600 2799.9200 1741.2600 2800.4000 ;
        RECT 1739.6600 2805.3600 1741.2600 2805.8400 ;
        RECT 1739.6600 2783.6000 1741.2600 2784.0800 ;
        RECT 1739.6600 2789.0400 1741.2600 2789.5200 ;
        RECT 1739.6600 2767.2800 1741.2600 2767.7600 ;
        RECT 1739.6600 2772.7200 1741.2600 2773.2000 ;
        RECT 1739.6600 2778.1600 1741.2600 2778.6400 ;
        RECT 1797.0000 2750.9600 1800.0000 2751.4400 ;
        RECT 1797.0000 2756.4000 1800.0000 2756.8800 ;
        RECT 1797.0000 2761.8400 1800.0000 2762.3200 ;
        RECT 1784.6600 2750.9600 1786.2600 2751.4400 ;
        RECT 1784.6600 2756.4000 1786.2600 2756.8800 ;
        RECT 1784.6600 2761.8400 1786.2600 2762.3200 ;
        RECT 1797.0000 2740.0800 1800.0000 2740.5600 ;
        RECT 1797.0000 2745.5200 1800.0000 2746.0000 ;
        RECT 1784.6600 2740.0800 1786.2600 2740.5600 ;
        RECT 1784.6600 2745.5200 1786.2600 2746.0000 ;
        RECT 1797.0000 2723.7600 1800.0000 2724.2400 ;
        RECT 1797.0000 2729.2000 1800.0000 2729.6800 ;
        RECT 1797.0000 2734.6400 1800.0000 2735.1200 ;
        RECT 1784.6600 2723.7600 1786.2600 2724.2400 ;
        RECT 1784.6600 2729.2000 1786.2600 2729.6800 ;
        RECT 1784.6600 2734.6400 1786.2600 2735.1200 ;
        RECT 1797.0000 2712.8800 1800.0000 2713.3600 ;
        RECT 1797.0000 2718.3200 1800.0000 2718.8000 ;
        RECT 1784.6600 2712.8800 1786.2600 2713.3600 ;
        RECT 1784.6600 2718.3200 1786.2600 2718.8000 ;
        RECT 1739.6600 2750.9600 1741.2600 2751.4400 ;
        RECT 1739.6600 2756.4000 1741.2600 2756.8800 ;
        RECT 1739.6600 2761.8400 1741.2600 2762.3200 ;
        RECT 1739.6600 2740.0800 1741.2600 2740.5600 ;
        RECT 1739.6600 2745.5200 1741.2600 2746.0000 ;
        RECT 1739.6600 2723.7600 1741.2600 2724.2400 ;
        RECT 1739.6600 2729.2000 1741.2600 2729.6800 ;
        RECT 1739.6600 2734.6400 1741.2600 2735.1200 ;
        RECT 1739.6600 2712.8800 1741.2600 2713.3600 ;
        RECT 1739.6600 2718.3200 1741.2600 2718.8000 ;
        RECT 1694.6600 2794.4800 1696.2600 2794.9600 ;
        RECT 1694.6600 2799.9200 1696.2600 2800.4000 ;
        RECT 1694.6600 2805.3600 1696.2600 2805.8400 ;
        RECT 1649.6600 2794.4800 1651.2600 2794.9600 ;
        RECT 1649.6600 2799.9200 1651.2600 2800.4000 ;
        RECT 1649.6600 2805.3600 1651.2600 2805.8400 ;
        RECT 1694.6600 2783.6000 1696.2600 2784.0800 ;
        RECT 1694.6600 2789.0400 1696.2600 2789.5200 ;
        RECT 1694.6600 2767.2800 1696.2600 2767.7600 ;
        RECT 1694.6600 2772.7200 1696.2600 2773.2000 ;
        RECT 1694.6600 2778.1600 1696.2600 2778.6400 ;
        RECT 1649.6600 2783.6000 1651.2600 2784.0800 ;
        RECT 1649.6600 2789.0400 1651.2600 2789.5200 ;
        RECT 1649.6600 2767.2800 1651.2600 2767.7600 ;
        RECT 1649.6600 2772.7200 1651.2600 2773.2000 ;
        RECT 1649.6600 2778.1600 1651.2600 2778.6400 ;
        RECT 1604.6600 2794.4800 1606.2600 2794.9600 ;
        RECT 1604.6600 2799.9200 1606.2600 2800.4000 ;
        RECT 1592.9000 2799.9200 1595.9000 2800.4000 ;
        RECT 1592.9000 2794.4800 1595.9000 2794.9600 ;
        RECT 1592.9000 2805.3600 1595.9000 2805.8400 ;
        RECT 1604.6600 2805.3600 1606.2600 2805.8400 ;
        RECT 1604.6600 2783.6000 1606.2600 2784.0800 ;
        RECT 1604.6600 2789.0400 1606.2600 2789.5200 ;
        RECT 1592.9000 2789.0400 1595.9000 2789.5200 ;
        RECT 1592.9000 2783.6000 1595.9000 2784.0800 ;
        RECT 1604.6600 2767.2800 1606.2600 2767.7600 ;
        RECT 1604.6600 2772.7200 1606.2600 2773.2000 ;
        RECT 1592.9000 2772.7200 1595.9000 2773.2000 ;
        RECT 1592.9000 2767.2800 1595.9000 2767.7600 ;
        RECT 1592.9000 2778.1600 1595.9000 2778.6400 ;
        RECT 1604.6600 2778.1600 1606.2600 2778.6400 ;
        RECT 1694.6600 2750.9600 1696.2600 2751.4400 ;
        RECT 1694.6600 2756.4000 1696.2600 2756.8800 ;
        RECT 1694.6600 2761.8400 1696.2600 2762.3200 ;
        RECT 1694.6600 2740.0800 1696.2600 2740.5600 ;
        RECT 1694.6600 2745.5200 1696.2600 2746.0000 ;
        RECT 1649.6600 2750.9600 1651.2600 2751.4400 ;
        RECT 1649.6600 2756.4000 1651.2600 2756.8800 ;
        RECT 1649.6600 2761.8400 1651.2600 2762.3200 ;
        RECT 1649.6600 2740.0800 1651.2600 2740.5600 ;
        RECT 1649.6600 2745.5200 1651.2600 2746.0000 ;
        RECT 1694.6600 2723.7600 1696.2600 2724.2400 ;
        RECT 1694.6600 2729.2000 1696.2600 2729.6800 ;
        RECT 1694.6600 2734.6400 1696.2600 2735.1200 ;
        RECT 1694.6600 2712.8800 1696.2600 2713.3600 ;
        RECT 1694.6600 2718.3200 1696.2600 2718.8000 ;
        RECT 1649.6600 2723.7600 1651.2600 2724.2400 ;
        RECT 1649.6600 2729.2000 1651.2600 2729.6800 ;
        RECT 1649.6600 2734.6400 1651.2600 2735.1200 ;
        RECT 1649.6600 2712.8800 1651.2600 2713.3600 ;
        RECT 1649.6600 2718.3200 1651.2600 2718.8000 ;
        RECT 1604.6600 2750.9600 1606.2600 2751.4400 ;
        RECT 1604.6600 2756.4000 1606.2600 2756.8800 ;
        RECT 1604.6600 2761.8400 1606.2600 2762.3200 ;
        RECT 1592.9000 2750.9600 1595.9000 2751.4400 ;
        RECT 1592.9000 2756.4000 1595.9000 2756.8800 ;
        RECT 1592.9000 2761.8400 1595.9000 2762.3200 ;
        RECT 1604.6600 2740.0800 1606.2600 2740.5600 ;
        RECT 1604.6600 2745.5200 1606.2600 2746.0000 ;
        RECT 1592.9000 2740.0800 1595.9000 2740.5600 ;
        RECT 1592.9000 2745.5200 1595.9000 2746.0000 ;
        RECT 1604.6600 2723.7600 1606.2600 2724.2400 ;
        RECT 1604.6600 2729.2000 1606.2600 2729.6800 ;
        RECT 1604.6600 2734.6400 1606.2600 2735.1200 ;
        RECT 1592.9000 2723.7600 1595.9000 2724.2400 ;
        RECT 1592.9000 2729.2000 1595.9000 2729.6800 ;
        RECT 1592.9000 2734.6400 1595.9000 2735.1200 ;
        RECT 1604.6600 2712.8800 1606.2600 2713.3600 ;
        RECT 1604.6600 2718.3200 1606.2600 2718.8000 ;
        RECT 1592.9000 2712.8800 1595.9000 2713.3600 ;
        RECT 1592.9000 2718.3200 1595.9000 2718.8000 ;
        RECT 1797.0000 2696.5600 1800.0000 2697.0400 ;
        RECT 1797.0000 2702.0000 1800.0000 2702.4800 ;
        RECT 1797.0000 2707.4400 1800.0000 2707.9200 ;
        RECT 1784.6600 2696.5600 1786.2600 2697.0400 ;
        RECT 1784.6600 2702.0000 1786.2600 2702.4800 ;
        RECT 1784.6600 2707.4400 1786.2600 2707.9200 ;
        RECT 1797.0000 2685.6800 1800.0000 2686.1600 ;
        RECT 1797.0000 2691.1200 1800.0000 2691.6000 ;
        RECT 1784.6600 2685.6800 1786.2600 2686.1600 ;
        RECT 1784.6600 2691.1200 1786.2600 2691.6000 ;
        RECT 1797.0000 2669.3600 1800.0000 2669.8400 ;
        RECT 1797.0000 2674.8000 1800.0000 2675.2800 ;
        RECT 1797.0000 2680.2400 1800.0000 2680.7200 ;
        RECT 1784.6600 2669.3600 1786.2600 2669.8400 ;
        RECT 1784.6600 2674.8000 1786.2600 2675.2800 ;
        RECT 1784.6600 2680.2400 1786.2600 2680.7200 ;
        RECT 1797.0000 2658.4800 1800.0000 2658.9600 ;
        RECT 1797.0000 2663.9200 1800.0000 2664.4000 ;
        RECT 1784.6600 2658.4800 1786.2600 2658.9600 ;
        RECT 1784.6600 2663.9200 1786.2600 2664.4000 ;
        RECT 1739.6600 2696.5600 1741.2600 2697.0400 ;
        RECT 1739.6600 2702.0000 1741.2600 2702.4800 ;
        RECT 1739.6600 2707.4400 1741.2600 2707.9200 ;
        RECT 1739.6600 2685.6800 1741.2600 2686.1600 ;
        RECT 1739.6600 2691.1200 1741.2600 2691.6000 ;
        RECT 1739.6600 2669.3600 1741.2600 2669.8400 ;
        RECT 1739.6600 2674.8000 1741.2600 2675.2800 ;
        RECT 1739.6600 2680.2400 1741.2600 2680.7200 ;
        RECT 1739.6600 2658.4800 1741.2600 2658.9600 ;
        RECT 1739.6600 2663.9200 1741.2600 2664.4000 ;
        RECT 1797.0000 2642.1600 1800.0000 2642.6400 ;
        RECT 1797.0000 2647.6000 1800.0000 2648.0800 ;
        RECT 1797.0000 2653.0400 1800.0000 2653.5200 ;
        RECT 1784.6600 2642.1600 1786.2600 2642.6400 ;
        RECT 1784.6600 2647.6000 1786.2600 2648.0800 ;
        RECT 1784.6600 2653.0400 1786.2600 2653.5200 ;
        RECT 1797.0000 2631.2800 1800.0000 2631.7600 ;
        RECT 1797.0000 2636.7200 1800.0000 2637.2000 ;
        RECT 1784.6600 2631.2800 1786.2600 2631.7600 ;
        RECT 1784.6600 2636.7200 1786.2600 2637.2000 ;
        RECT 1797.0000 2614.9600 1800.0000 2615.4400 ;
        RECT 1797.0000 2620.4000 1800.0000 2620.8800 ;
        RECT 1797.0000 2625.8400 1800.0000 2626.3200 ;
        RECT 1784.6600 2614.9600 1786.2600 2615.4400 ;
        RECT 1784.6600 2620.4000 1786.2600 2620.8800 ;
        RECT 1784.6600 2625.8400 1786.2600 2626.3200 ;
        RECT 1797.0000 2609.5200 1800.0000 2610.0000 ;
        RECT 1784.6600 2609.5200 1786.2600 2610.0000 ;
        RECT 1739.6600 2642.1600 1741.2600 2642.6400 ;
        RECT 1739.6600 2647.6000 1741.2600 2648.0800 ;
        RECT 1739.6600 2653.0400 1741.2600 2653.5200 ;
        RECT 1739.6600 2631.2800 1741.2600 2631.7600 ;
        RECT 1739.6600 2636.7200 1741.2600 2637.2000 ;
        RECT 1739.6600 2614.9600 1741.2600 2615.4400 ;
        RECT 1739.6600 2620.4000 1741.2600 2620.8800 ;
        RECT 1739.6600 2625.8400 1741.2600 2626.3200 ;
        RECT 1739.6600 2609.5200 1741.2600 2610.0000 ;
        RECT 1694.6600 2696.5600 1696.2600 2697.0400 ;
        RECT 1694.6600 2702.0000 1696.2600 2702.4800 ;
        RECT 1694.6600 2707.4400 1696.2600 2707.9200 ;
        RECT 1694.6600 2685.6800 1696.2600 2686.1600 ;
        RECT 1694.6600 2691.1200 1696.2600 2691.6000 ;
        RECT 1649.6600 2696.5600 1651.2600 2697.0400 ;
        RECT 1649.6600 2702.0000 1651.2600 2702.4800 ;
        RECT 1649.6600 2707.4400 1651.2600 2707.9200 ;
        RECT 1649.6600 2685.6800 1651.2600 2686.1600 ;
        RECT 1649.6600 2691.1200 1651.2600 2691.6000 ;
        RECT 1694.6600 2669.3600 1696.2600 2669.8400 ;
        RECT 1694.6600 2674.8000 1696.2600 2675.2800 ;
        RECT 1694.6600 2680.2400 1696.2600 2680.7200 ;
        RECT 1694.6600 2658.4800 1696.2600 2658.9600 ;
        RECT 1694.6600 2663.9200 1696.2600 2664.4000 ;
        RECT 1649.6600 2669.3600 1651.2600 2669.8400 ;
        RECT 1649.6600 2674.8000 1651.2600 2675.2800 ;
        RECT 1649.6600 2680.2400 1651.2600 2680.7200 ;
        RECT 1649.6600 2658.4800 1651.2600 2658.9600 ;
        RECT 1649.6600 2663.9200 1651.2600 2664.4000 ;
        RECT 1604.6600 2696.5600 1606.2600 2697.0400 ;
        RECT 1604.6600 2702.0000 1606.2600 2702.4800 ;
        RECT 1604.6600 2707.4400 1606.2600 2707.9200 ;
        RECT 1592.9000 2696.5600 1595.9000 2697.0400 ;
        RECT 1592.9000 2702.0000 1595.9000 2702.4800 ;
        RECT 1592.9000 2707.4400 1595.9000 2707.9200 ;
        RECT 1604.6600 2685.6800 1606.2600 2686.1600 ;
        RECT 1604.6600 2691.1200 1606.2600 2691.6000 ;
        RECT 1592.9000 2685.6800 1595.9000 2686.1600 ;
        RECT 1592.9000 2691.1200 1595.9000 2691.6000 ;
        RECT 1604.6600 2669.3600 1606.2600 2669.8400 ;
        RECT 1604.6600 2674.8000 1606.2600 2675.2800 ;
        RECT 1604.6600 2680.2400 1606.2600 2680.7200 ;
        RECT 1592.9000 2669.3600 1595.9000 2669.8400 ;
        RECT 1592.9000 2674.8000 1595.9000 2675.2800 ;
        RECT 1592.9000 2680.2400 1595.9000 2680.7200 ;
        RECT 1604.6600 2658.4800 1606.2600 2658.9600 ;
        RECT 1604.6600 2663.9200 1606.2600 2664.4000 ;
        RECT 1592.9000 2658.4800 1595.9000 2658.9600 ;
        RECT 1592.9000 2663.9200 1595.9000 2664.4000 ;
        RECT 1694.6600 2642.1600 1696.2600 2642.6400 ;
        RECT 1694.6600 2647.6000 1696.2600 2648.0800 ;
        RECT 1694.6600 2653.0400 1696.2600 2653.5200 ;
        RECT 1694.6600 2631.2800 1696.2600 2631.7600 ;
        RECT 1694.6600 2636.7200 1696.2600 2637.2000 ;
        RECT 1649.6600 2642.1600 1651.2600 2642.6400 ;
        RECT 1649.6600 2647.6000 1651.2600 2648.0800 ;
        RECT 1649.6600 2653.0400 1651.2600 2653.5200 ;
        RECT 1649.6600 2631.2800 1651.2600 2631.7600 ;
        RECT 1649.6600 2636.7200 1651.2600 2637.2000 ;
        RECT 1694.6600 2614.9600 1696.2600 2615.4400 ;
        RECT 1694.6600 2620.4000 1696.2600 2620.8800 ;
        RECT 1694.6600 2625.8400 1696.2600 2626.3200 ;
        RECT 1694.6600 2609.5200 1696.2600 2610.0000 ;
        RECT 1649.6600 2614.9600 1651.2600 2615.4400 ;
        RECT 1649.6600 2620.4000 1651.2600 2620.8800 ;
        RECT 1649.6600 2625.8400 1651.2600 2626.3200 ;
        RECT 1649.6600 2609.5200 1651.2600 2610.0000 ;
        RECT 1604.6600 2642.1600 1606.2600 2642.6400 ;
        RECT 1604.6600 2647.6000 1606.2600 2648.0800 ;
        RECT 1604.6600 2653.0400 1606.2600 2653.5200 ;
        RECT 1592.9000 2642.1600 1595.9000 2642.6400 ;
        RECT 1592.9000 2647.6000 1595.9000 2648.0800 ;
        RECT 1592.9000 2653.0400 1595.9000 2653.5200 ;
        RECT 1604.6600 2631.2800 1606.2600 2631.7600 ;
        RECT 1604.6600 2636.7200 1606.2600 2637.2000 ;
        RECT 1592.9000 2631.2800 1595.9000 2631.7600 ;
        RECT 1592.9000 2636.7200 1595.9000 2637.2000 ;
        RECT 1604.6600 2614.9600 1606.2600 2615.4400 ;
        RECT 1604.6600 2620.4000 1606.2600 2620.8800 ;
        RECT 1604.6600 2625.8400 1606.2600 2626.3200 ;
        RECT 1592.9000 2614.9600 1595.9000 2615.4400 ;
        RECT 1592.9000 2620.4000 1595.9000 2620.8800 ;
        RECT 1592.9000 2625.8400 1595.9000 2626.3200 ;
        RECT 1592.9000 2609.5200 1595.9000 2610.0000 ;
        RECT 1604.6600 2609.5200 1606.2600 2610.0000 ;
        RECT 1592.9000 2814.4300 1800.0000 2817.4300 ;
        RECT 1592.9000 2601.3300 1800.0000 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 2371.6900 1786.2600 2587.7900 ;
        RECT 1739.6600 2371.6900 1741.2600 2587.7900 ;
        RECT 1694.6600 2371.6900 1696.2600 2587.7900 ;
        RECT 1649.6600 2371.6900 1651.2600 2587.7900 ;
        RECT 1604.6600 2371.6900 1606.2600 2587.7900 ;
        RECT 1797.0000 2371.6900 1800.0000 2587.7900 ;
        RECT 1592.9000 2371.6900 1595.9000 2587.7900 ;
      LAYER met3 ;
        RECT 1797.0000 2564.8400 1800.0000 2565.3200 ;
        RECT 1797.0000 2570.2800 1800.0000 2570.7600 ;
        RECT 1784.6600 2564.8400 1786.2600 2565.3200 ;
        RECT 1784.6600 2570.2800 1786.2600 2570.7600 ;
        RECT 1797.0000 2575.7200 1800.0000 2576.2000 ;
        RECT 1784.6600 2575.7200 1786.2600 2576.2000 ;
        RECT 1797.0000 2553.9600 1800.0000 2554.4400 ;
        RECT 1797.0000 2559.4000 1800.0000 2559.8800 ;
        RECT 1784.6600 2553.9600 1786.2600 2554.4400 ;
        RECT 1784.6600 2559.4000 1786.2600 2559.8800 ;
        RECT 1797.0000 2537.6400 1800.0000 2538.1200 ;
        RECT 1797.0000 2543.0800 1800.0000 2543.5600 ;
        RECT 1784.6600 2537.6400 1786.2600 2538.1200 ;
        RECT 1784.6600 2543.0800 1786.2600 2543.5600 ;
        RECT 1797.0000 2548.5200 1800.0000 2549.0000 ;
        RECT 1784.6600 2548.5200 1786.2600 2549.0000 ;
        RECT 1739.6600 2564.8400 1741.2600 2565.3200 ;
        RECT 1739.6600 2570.2800 1741.2600 2570.7600 ;
        RECT 1739.6600 2575.7200 1741.2600 2576.2000 ;
        RECT 1739.6600 2553.9600 1741.2600 2554.4400 ;
        RECT 1739.6600 2559.4000 1741.2600 2559.8800 ;
        RECT 1739.6600 2537.6400 1741.2600 2538.1200 ;
        RECT 1739.6600 2543.0800 1741.2600 2543.5600 ;
        RECT 1739.6600 2548.5200 1741.2600 2549.0000 ;
        RECT 1797.0000 2521.3200 1800.0000 2521.8000 ;
        RECT 1797.0000 2526.7600 1800.0000 2527.2400 ;
        RECT 1797.0000 2532.2000 1800.0000 2532.6800 ;
        RECT 1784.6600 2521.3200 1786.2600 2521.8000 ;
        RECT 1784.6600 2526.7600 1786.2600 2527.2400 ;
        RECT 1784.6600 2532.2000 1786.2600 2532.6800 ;
        RECT 1797.0000 2510.4400 1800.0000 2510.9200 ;
        RECT 1797.0000 2515.8800 1800.0000 2516.3600 ;
        RECT 1784.6600 2510.4400 1786.2600 2510.9200 ;
        RECT 1784.6600 2515.8800 1786.2600 2516.3600 ;
        RECT 1797.0000 2494.1200 1800.0000 2494.6000 ;
        RECT 1797.0000 2499.5600 1800.0000 2500.0400 ;
        RECT 1797.0000 2505.0000 1800.0000 2505.4800 ;
        RECT 1784.6600 2494.1200 1786.2600 2494.6000 ;
        RECT 1784.6600 2499.5600 1786.2600 2500.0400 ;
        RECT 1784.6600 2505.0000 1786.2600 2505.4800 ;
        RECT 1797.0000 2483.2400 1800.0000 2483.7200 ;
        RECT 1797.0000 2488.6800 1800.0000 2489.1600 ;
        RECT 1784.6600 2483.2400 1786.2600 2483.7200 ;
        RECT 1784.6600 2488.6800 1786.2600 2489.1600 ;
        RECT 1739.6600 2521.3200 1741.2600 2521.8000 ;
        RECT 1739.6600 2526.7600 1741.2600 2527.2400 ;
        RECT 1739.6600 2532.2000 1741.2600 2532.6800 ;
        RECT 1739.6600 2510.4400 1741.2600 2510.9200 ;
        RECT 1739.6600 2515.8800 1741.2600 2516.3600 ;
        RECT 1739.6600 2494.1200 1741.2600 2494.6000 ;
        RECT 1739.6600 2499.5600 1741.2600 2500.0400 ;
        RECT 1739.6600 2505.0000 1741.2600 2505.4800 ;
        RECT 1739.6600 2483.2400 1741.2600 2483.7200 ;
        RECT 1739.6600 2488.6800 1741.2600 2489.1600 ;
        RECT 1694.6600 2564.8400 1696.2600 2565.3200 ;
        RECT 1694.6600 2570.2800 1696.2600 2570.7600 ;
        RECT 1694.6600 2575.7200 1696.2600 2576.2000 ;
        RECT 1649.6600 2564.8400 1651.2600 2565.3200 ;
        RECT 1649.6600 2570.2800 1651.2600 2570.7600 ;
        RECT 1649.6600 2575.7200 1651.2600 2576.2000 ;
        RECT 1694.6600 2553.9600 1696.2600 2554.4400 ;
        RECT 1694.6600 2559.4000 1696.2600 2559.8800 ;
        RECT 1694.6600 2537.6400 1696.2600 2538.1200 ;
        RECT 1694.6600 2543.0800 1696.2600 2543.5600 ;
        RECT 1694.6600 2548.5200 1696.2600 2549.0000 ;
        RECT 1649.6600 2553.9600 1651.2600 2554.4400 ;
        RECT 1649.6600 2559.4000 1651.2600 2559.8800 ;
        RECT 1649.6600 2537.6400 1651.2600 2538.1200 ;
        RECT 1649.6600 2543.0800 1651.2600 2543.5600 ;
        RECT 1649.6600 2548.5200 1651.2600 2549.0000 ;
        RECT 1604.6600 2564.8400 1606.2600 2565.3200 ;
        RECT 1604.6600 2570.2800 1606.2600 2570.7600 ;
        RECT 1592.9000 2570.2800 1595.9000 2570.7600 ;
        RECT 1592.9000 2564.8400 1595.9000 2565.3200 ;
        RECT 1592.9000 2575.7200 1595.9000 2576.2000 ;
        RECT 1604.6600 2575.7200 1606.2600 2576.2000 ;
        RECT 1604.6600 2553.9600 1606.2600 2554.4400 ;
        RECT 1604.6600 2559.4000 1606.2600 2559.8800 ;
        RECT 1592.9000 2559.4000 1595.9000 2559.8800 ;
        RECT 1592.9000 2553.9600 1595.9000 2554.4400 ;
        RECT 1604.6600 2537.6400 1606.2600 2538.1200 ;
        RECT 1604.6600 2543.0800 1606.2600 2543.5600 ;
        RECT 1592.9000 2543.0800 1595.9000 2543.5600 ;
        RECT 1592.9000 2537.6400 1595.9000 2538.1200 ;
        RECT 1592.9000 2548.5200 1595.9000 2549.0000 ;
        RECT 1604.6600 2548.5200 1606.2600 2549.0000 ;
        RECT 1694.6600 2521.3200 1696.2600 2521.8000 ;
        RECT 1694.6600 2526.7600 1696.2600 2527.2400 ;
        RECT 1694.6600 2532.2000 1696.2600 2532.6800 ;
        RECT 1694.6600 2510.4400 1696.2600 2510.9200 ;
        RECT 1694.6600 2515.8800 1696.2600 2516.3600 ;
        RECT 1649.6600 2521.3200 1651.2600 2521.8000 ;
        RECT 1649.6600 2526.7600 1651.2600 2527.2400 ;
        RECT 1649.6600 2532.2000 1651.2600 2532.6800 ;
        RECT 1649.6600 2510.4400 1651.2600 2510.9200 ;
        RECT 1649.6600 2515.8800 1651.2600 2516.3600 ;
        RECT 1694.6600 2494.1200 1696.2600 2494.6000 ;
        RECT 1694.6600 2499.5600 1696.2600 2500.0400 ;
        RECT 1694.6600 2505.0000 1696.2600 2505.4800 ;
        RECT 1694.6600 2483.2400 1696.2600 2483.7200 ;
        RECT 1694.6600 2488.6800 1696.2600 2489.1600 ;
        RECT 1649.6600 2494.1200 1651.2600 2494.6000 ;
        RECT 1649.6600 2499.5600 1651.2600 2500.0400 ;
        RECT 1649.6600 2505.0000 1651.2600 2505.4800 ;
        RECT 1649.6600 2483.2400 1651.2600 2483.7200 ;
        RECT 1649.6600 2488.6800 1651.2600 2489.1600 ;
        RECT 1604.6600 2521.3200 1606.2600 2521.8000 ;
        RECT 1604.6600 2526.7600 1606.2600 2527.2400 ;
        RECT 1604.6600 2532.2000 1606.2600 2532.6800 ;
        RECT 1592.9000 2521.3200 1595.9000 2521.8000 ;
        RECT 1592.9000 2526.7600 1595.9000 2527.2400 ;
        RECT 1592.9000 2532.2000 1595.9000 2532.6800 ;
        RECT 1604.6600 2510.4400 1606.2600 2510.9200 ;
        RECT 1604.6600 2515.8800 1606.2600 2516.3600 ;
        RECT 1592.9000 2510.4400 1595.9000 2510.9200 ;
        RECT 1592.9000 2515.8800 1595.9000 2516.3600 ;
        RECT 1604.6600 2494.1200 1606.2600 2494.6000 ;
        RECT 1604.6600 2499.5600 1606.2600 2500.0400 ;
        RECT 1604.6600 2505.0000 1606.2600 2505.4800 ;
        RECT 1592.9000 2494.1200 1595.9000 2494.6000 ;
        RECT 1592.9000 2499.5600 1595.9000 2500.0400 ;
        RECT 1592.9000 2505.0000 1595.9000 2505.4800 ;
        RECT 1604.6600 2483.2400 1606.2600 2483.7200 ;
        RECT 1604.6600 2488.6800 1606.2600 2489.1600 ;
        RECT 1592.9000 2483.2400 1595.9000 2483.7200 ;
        RECT 1592.9000 2488.6800 1595.9000 2489.1600 ;
        RECT 1797.0000 2466.9200 1800.0000 2467.4000 ;
        RECT 1797.0000 2472.3600 1800.0000 2472.8400 ;
        RECT 1797.0000 2477.8000 1800.0000 2478.2800 ;
        RECT 1784.6600 2466.9200 1786.2600 2467.4000 ;
        RECT 1784.6600 2472.3600 1786.2600 2472.8400 ;
        RECT 1784.6600 2477.8000 1786.2600 2478.2800 ;
        RECT 1797.0000 2456.0400 1800.0000 2456.5200 ;
        RECT 1797.0000 2461.4800 1800.0000 2461.9600 ;
        RECT 1784.6600 2456.0400 1786.2600 2456.5200 ;
        RECT 1784.6600 2461.4800 1786.2600 2461.9600 ;
        RECT 1797.0000 2439.7200 1800.0000 2440.2000 ;
        RECT 1797.0000 2445.1600 1800.0000 2445.6400 ;
        RECT 1797.0000 2450.6000 1800.0000 2451.0800 ;
        RECT 1784.6600 2439.7200 1786.2600 2440.2000 ;
        RECT 1784.6600 2445.1600 1786.2600 2445.6400 ;
        RECT 1784.6600 2450.6000 1786.2600 2451.0800 ;
        RECT 1797.0000 2428.8400 1800.0000 2429.3200 ;
        RECT 1797.0000 2434.2800 1800.0000 2434.7600 ;
        RECT 1784.6600 2428.8400 1786.2600 2429.3200 ;
        RECT 1784.6600 2434.2800 1786.2600 2434.7600 ;
        RECT 1739.6600 2466.9200 1741.2600 2467.4000 ;
        RECT 1739.6600 2472.3600 1741.2600 2472.8400 ;
        RECT 1739.6600 2477.8000 1741.2600 2478.2800 ;
        RECT 1739.6600 2456.0400 1741.2600 2456.5200 ;
        RECT 1739.6600 2461.4800 1741.2600 2461.9600 ;
        RECT 1739.6600 2439.7200 1741.2600 2440.2000 ;
        RECT 1739.6600 2445.1600 1741.2600 2445.6400 ;
        RECT 1739.6600 2450.6000 1741.2600 2451.0800 ;
        RECT 1739.6600 2428.8400 1741.2600 2429.3200 ;
        RECT 1739.6600 2434.2800 1741.2600 2434.7600 ;
        RECT 1797.0000 2412.5200 1800.0000 2413.0000 ;
        RECT 1797.0000 2417.9600 1800.0000 2418.4400 ;
        RECT 1797.0000 2423.4000 1800.0000 2423.8800 ;
        RECT 1784.6600 2412.5200 1786.2600 2413.0000 ;
        RECT 1784.6600 2417.9600 1786.2600 2418.4400 ;
        RECT 1784.6600 2423.4000 1786.2600 2423.8800 ;
        RECT 1797.0000 2401.6400 1800.0000 2402.1200 ;
        RECT 1797.0000 2407.0800 1800.0000 2407.5600 ;
        RECT 1784.6600 2401.6400 1786.2600 2402.1200 ;
        RECT 1784.6600 2407.0800 1786.2600 2407.5600 ;
        RECT 1797.0000 2385.3200 1800.0000 2385.8000 ;
        RECT 1797.0000 2390.7600 1800.0000 2391.2400 ;
        RECT 1797.0000 2396.2000 1800.0000 2396.6800 ;
        RECT 1784.6600 2385.3200 1786.2600 2385.8000 ;
        RECT 1784.6600 2390.7600 1786.2600 2391.2400 ;
        RECT 1784.6600 2396.2000 1786.2600 2396.6800 ;
        RECT 1797.0000 2379.8800 1800.0000 2380.3600 ;
        RECT 1784.6600 2379.8800 1786.2600 2380.3600 ;
        RECT 1739.6600 2412.5200 1741.2600 2413.0000 ;
        RECT 1739.6600 2417.9600 1741.2600 2418.4400 ;
        RECT 1739.6600 2423.4000 1741.2600 2423.8800 ;
        RECT 1739.6600 2401.6400 1741.2600 2402.1200 ;
        RECT 1739.6600 2407.0800 1741.2600 2407.5600 ;
        RECT 1739.6600 2385.3200 1741.2600 2385.8000 ;
        RECT 1739.6600 2390.7600 1741.2600 2391.2400 ;
        RECT 1739.6600 2396.2000 1741.2600 2396.6800 ;
        RECT 1739.6600 2379.8800 1741.2600 2380.3600 ;
        RECT 1694.6600 2466.9200 1696.2600 2467.4000 ;
        RECT 1694.6600 2472.3600 1696.2600 2472.8400 ;
        RECT 1694.6600 2477.8000 1696.2600 2478.2800 ;
        RECT 1694.6600 2456.0400 1696.2600 2456.5200 ;
        RECT 1694.6600 2461.4800 1696.2600 2461.9600 ;
        RECT 1649.6600 2466.9200 1651.2600 2467.4000 ;
        RECT 1649.6600 2472.3600 1651.2600 2472.8400 ;
        RECT 1649.6600 2477.8000 1651.2600 2478.2800 ;
        RECT 1649.6600 2456.0400 1651.2600 2456.5200 ;
        RECT 1649.6600 2461.4800 1651.2600 2461.9600 ;
        RECT 1694.6600 2439.7200 1696.2600 2440.2000 ;
        RECT 1694.6600 2445.1600 1696.2600 2445.6400 ;
        RECT 1694.6600 2450.6000 1696.2600 2451.0800 ;
        RECT 1694.6600 2428.8400 1696.2600 2429.3200 ;
        RECT 1694.6600 2434.2800 1696.2600 2434.7600 ;
        RECT 1649.6600 2439.7200 1651.2600 2440.2000 ;
        RECT 1649.6600 2445.1600 1651.2600 2445.6400 ;
        RECT 1649.6600 2450.6000 1651.2600 2451.0800 ;
        RECT 1649.6600 2428.8400 1651.2600 2429.3200 ;
        RECT 1649.6600 2434.2800 1651.2600 2434.7600 ;
        RECT 1604.6600 2466.9200 1606.2600 2467.4000 ;
        RECT 1604.6600 2472.3600 1606.2600 2472.8400 ;
        RECT 1604.6600 2477.8000 1606.2600 2478.2800 ;
        RECT 1592.9000 2466.9200 1595.9000 2467.4000 ;
        RECT 1592.9000 2472.3600 1595.9000 2472.8400 ;
        RECT 1592.9000 2477.8000 1595.9000 2478.2800 ;
        RECT 1604.6600 2456.0400 1606.2600 2456.5200 ;
        RECT 1604.6600 2461.4800 1606.2600 2461.9600 ;
        RECT 1592.9000 2456.0400 1595.9000 2456.5200 ;
        RECT 1592.9000 2461.4800 1595.9000 2461.9600 ;
        RECT 1604.6600 2439.7200 1606.2600 2440.2000 ;
        RECT 1604.6600 2445.1600 1606.2600 2445.6400 ;
        RECT 1604.6600 2450.6000 1606.2600 2451.0800 ;
        RECT 1592.9000 2439.7200 1595.9000 2440.2000 ;
        RECT 1592.9000 2445.1600 1595.9000 2445.6400 ;
        RECT 1592.9000 2450.6000 1595.9000 2451.0800 ;
        RECT 1604.6600 2428.8400 1606.2600 2429.3200 ;
        RECT 1604.6600 2434.2800 1606.2600 2434.7600 ;
        RECT 1592.9000 2428.8400 1595.9000 2429.3200 ;
        RECT 1592.9000 2434.2800 1595.9000 2434.7600 ;
        RECT 1694.6600 2412.5200 1696.2600 2413.0000 ;
        RECT 1694.6600 2417.9600 1696.2600 2418.4400 ;
        RECT 1694.6600 2423.4000 1696.2600 2423.8800 ;
        RECT 1694.6600 2401.6400 1696.2600 2402.1200 ;
        RECT 1694.6600 2407.0800 1696.2600 2407.5600 ;
        RECT 1649.6600 2412.5200 1651.2600 2413.0000 ;
        RECT 1649.6600 2417.9600 1651.2600 2418.4400 ;
        RECT 1649.6600 2423.4000 1651.2600 2423.8800 ;
        RECT 1649.6600 2401.6400 1651.2600 2402.1200 ;
        RECT 1649.6600 2407.0800 1651.2600 2407.5600 ;
        RECT 1694.6600 2385.3200 1696.2600 2385.8000 ;
        RECT 1694.6600 2390.7600 1696.2600 2391.2400 ;
        RECT 1694.6600 2396.2000 1696.2600 2396.6800 ;
        RECT 1694.6600 2379.8800 1696.2600 2380.3600 ;
        RECT 1649.6600 2385.3200 1651.2600 2385.8000 ;
        RECT 1649.6600 2390.7600 1651.2600 2391.2400 ;
        RECT 1649.6600 2396.2000 1651.2600 2396.6800 ;
        RECT 1649.6600 2379.8800 1651.2600 2380.3600 ;
        RECT 1604.6600 2412.5200 1606.2600 2413.0000 ;
        RECT 1604.6600 2417.9600 1606.2600 2418.4400 ;
        RECT 1604.6600 2423.4000 1606.2600 2423.8800 ;
        RECT 1592.9000 2412.5200 1595.9000 2413.0000 ;
        RECT 1592.9000 2417.9600 1595.9000 2418.4400 ;
        RECT 1592.9000 2423.4000 1595.9000 2423.8800 ;
        RECT 1604.6600 2401.6400 1606.2600 2402.1200 ;
        RECT 1604.6600 2407.0800 1606.2600 2407.5600 ;
        RECT 1592.9000 2401.6400 1595.9000 2402.1200 ;
        RECT 1592.9000 2407.0800 1595.9000 2407.5600 ;
        RECT 1604.6600 2385.3200 1606.2600 2385.8000 ;
        RECT 1604.6600 2390.7600 1606.2600 2391.2400 ;
        RECT 1604.6600 2396.2000 1606.2600 2396.6800 ;
        RECT 1592.9000 2385.3200 1595.9000 2385.8000 ;
        RECT 1592.9000 2390.7600 1595.9000 2391.2400 ;
        RECT 1592.9000 2396.2000 1595.9000 2396.6800 ;
        RECT 1592.9000 2379.8800 1595.9000 2380.3600 ;
        RECT 1604.6600 2379.8800 1606.2600 2380.3600 ;
        RECT 1592.9000 2584.7900 1800.0000 2587.7900 ;
        RECT 1592.9000 2371.6900 1800.0000 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 2142.0500 1786.2600 2358.1500 ;
        RECT 1739.6600 2142.0500 1741.2600 2358.1500 ;
        RECT 1694.6600 2142.0500 1696.2600 2358.1500 ;
        RECT 1649.6600 2142.0500 1651.2600 2358.1500 ;
        RECT 1604.6600 2142.0500 1606.2600 2358.1500 ;
        RECT 1797.0000 2142.0500 1800.0000 2358.1500 ;
        RECT 1592.9000 2142.0500 1595.9000 2358.1500 ;
      LAYER met3 ;
        RECT 1797.0000 2335.2000 1800.0000 2335.6800 ;
        RECT 1797.0000 2340.6400 1800.0000 2341.1200 ;
        RECT 1784.6600 2335.2000 1786.2600 2335.6800 ;
        RECT 1784.6600 2340.6400 1786.2600 2341.1200 ;
        RECT 1797.0000 2346.0800 1800.0000 2346.5600 ;
        RECT 1784.6600 2346.0800 1786.2600 2346.5600 ;
        RECT 1797.0000 2324.3200 1800.0000 2324.8000 ;
        RECT 1797.0000 2329.7600 1800.0000 2330.2400 ;
        RECT 1784.6600 2324.3200 1786.2600 2324.8000 ;
        RECT 1784.6600 2329.7600 1786.2600 2330.2400 ;
        RECT 1797.0000 2308.0000 1800.0000 2308.4800 ;
        RECT 1797.0000 2313.4400 1800.0000 2313.9200 ;
        RECT 1784.6600 2308.0000 1786.2600 2308.4800 ;
        RECT 1784.6600 2313.4400 1786.2600 2313.9200 ;
        RECT 1797.0000 2318.8800 1800.0000 2319.3600 ;
        RECT 1784.6600 2318.8800 1786.2600 2319.3600 ;
        RECT 1739.6600 2335.2000 1741.2600 2335.6800 ;
        RECT 1739.6600 2340.6400 1741.2600 2341.1200 ;
        RECT 1739.6600 2346.0800 1741.2600 2346.5600 ;
        RECT 1739.6600 2324.3200 1741.2600 2324.8000 ;
        RECT 1739.6600 2329.7600 1741.2600 2330.2400 ;
        RECT 1739.6600 2308.0000 1741.2600 2308.4800 ;
        RECT 1739.6600 2313.4400 1741.2600 2313.9200 ;
        RECT 1739.6600 2318.8800 1741.2600 2319.3600 ;
        RECT 1797.0000 2291.6800 1800.0000 2292.1600 ;
        RECT 1797.0000 2297.1200 1800.0000 2297.6000 ;
        RECT 1797.0000 2302.5600 1800.0000 2303.0400 ;
        RECT 1784.6600 2291.6800 1786.2600 2292.1600 ;
        RECT 1784.6600 2297.1200 1786.2600 2297.6000 ;
        RECT 1784.6600 2302.5600 1786.2600 2303.0400 ;
        RECT 1797.0000 2280.8000 1800.0000 2281.2800 ;
        RECT 1797.0000 2286.2400 1800.0000 2286.7200 ;
        RECT 1784.6600 2280.8000 1786.2600 2281.2800 ;
        RECT 1784.6600 2286.2400 1786.2600 2286.7200 ;
        RECT 1797.0000 2264.4800 1800.0000 2264.9600 ;
        RECT 1797.0000 2269.9200 1800.0000 2270.4000 ;
        RECT 1797.0000 2275.3600 1800.0000 2275.8400 ;
        RECT 1784.6600 2264.4800 1786.2600 2264.9600 ;
        RECT 1784.6600 2269.9200 1786.2600 2270.4000 ;
        RECT 1784.6600 2275.3600 1786.2600 2275.8400 ;
        RECT 1797.0000 2253.6000 1800.0000 2254.0800 ;
        RECT 1797.0000 2259.0400 1800.0000 2259.5200 ;
        RECT 1784.6600 2253.6000 1786.2600 2254.0800 ;
        RECT 1784.6600 2259.0400 1786.2600 2259.5200 ;
        RECT 1739.6600 2291.6800 1741.2600 2292.1600 ;
        RECT 1739.6600 2297.1200 1741.2600 2297.6000 ;
        RECT 1739.6600 2302.5600 1741.2600 2303.0400 ;
        RECT 1739.6600 2280.8000 1741.2600 2281.2800 ;
        RECT 1739.6600 2286.2400 1741.2600 2286.7200 ;
        RECT 1739.6600 2264.4800 1741.2600 2264.9600 ;
        RECT 1739.6600 2269.9200 1741.2600 2270.4000 ;
        RECT 1739.6600 2275.3600 1741.2600 2275.8400 ;
        RECT 1739.6600 2253.6000 1741.2600 2254.0800 ;
        RECT 1739.6600 2259.0400 1741.2600 2259.5200 ;
        RECT 1694.6600 2335.2000 1696.2600 2335.6800 ;
        RECT 1694.6600 2340.6400 1696.2600 2341.1200 ;
        RECT 1694.6600 2346.0800 1696.2600 2346.5600 ;
        RECT 1649.6600 2335.2000 1651.2600 2335.6800 ;
        RECT 1649.6600 2340.6400 1651.2600 2341.1200 ;
        RECT 1649.6600 2346.0800 1651.2600 2346.5600 ;
        RECT 1694.6600 2324.3200 1696.2600 2324.8000 ;
        RECT 1694.6600 2329.7600 1696.2600 2330.2400 ;
        RECT 1694.6600 2308.0000 1696.2600 2308.4800 ;
        RECT 1694.6600 2313.4400 1696.2600 2313.9200 ;
        RECT 1694.6600 2318.8800 1696.2600 2319.3600 ;
        RECT 1649.6600 2324.3200 1651.2600 2324.8000 ;
        RECT 1649.6600 2329.7600 1651.2600 2330.2400 ;
        RECT 1649.6600 2308.0000 1651.2600 2308.4800 ;
        RECT 1649.6600 2313.4400 1651.2600 2313.9200 ;
        RECT 1649.6600 2318.8800 1651.2600 2319.3600 ;
        RECT 1604.6600 2335.2000 1606.2600 2335.6800 ;
        RECT 1604.6600 2340.6400 1606.2600 2341.1200 ;
        RECT 1592.9000 2340.6400 1595.9000 2341.1200 ;
        RECT 1592.9000 2335.2000 1595.9000 2335.6800 ;
        RECT 1592.9000 2346.0800 1595.9000 2346.5600 ;
        RECT 1604.6600 2346.0800 1606.2600 2346.5600 ;
        RECT 1604.6600 2324.3200 1606.2600 2324.8000 ;
        RECT 1604.6600 2329.7600 1606.2600 2330.2400 ;
        RECT 1592.9000 2329.7600 1595.9000 2330.2400 ;
        RECT 1592.9000 2324.3200 1595.9000 2324.8000 ;
        RECT 1604.6600 2308.0000 1606.2600 2308.4800 ;
        RECT 1604.6600 2313.4400 1606.2600 2313.9200 ;
        RECT 1592.9000 2313.4400 1595.9000 2313.9200 ;
        RECT 1592.9000 2308.0000 1595.9000 2308.4800 ;
        RECT 1592.9000 2318.8800 1595.9000 2319.3600 ;
        RECT 1604.6600 2318.8800 1606.2600 2319.3600 ;
        RECT 1694.6600 2291.6800 1696.2600 2292.1600 ;
        RECT 1694.6600 2297.1200 1696.2600 2297.6000 ;
        RECT 1694.6600 2302.5600 1696.2600 2303.0400 ;
        RECT 1694.6600 2280.8000 1696.2600 2281.2800 ;
        RECT 1694.6600 2286.2400 1696.2600 2286.7200 ;
        RECT 1649.6600 2291.6800 1651.2600 2292.1600 ;
        RECT 1649.6600 2297.1200 1651.2600 2297.6000 ;
        RECT 1649.6600 2302.5600 1651.2600 2303.0400 ;
        RECT 1649.6600 2280.8000 1651.2600 2281.2800 ;
        RECT 1649.6600 2286.2400 1651.2600 2286.7200 ;
        RECT 1694.6600 2264.4800 1696.2600 2264.9600 ;
        RECT 1694.6600 2269.9200 1696.2600 2270.4000 ;
        RECT 1694.6600 2275.3600 1696.2600 2275.8400 ;
        RECT 1694.6600 2253.6000 1696.2600 2254.0800 ;
        RECT 1694.6600 2259.0400 1696.2600 2259.5200 ;
        RECT 1649.6600 2264.4800 1651.2600 2264.9600 ;
        RECT 1649.6600 2269.9200 1651.2600 2270.4000 ;
        RECT 1649.6600 2275.3600 1651.2600 2275.8400 ;
        RECT 1649.6600 2253.6000 1651.2600 2254.0800 ;
        RECT 1649.6600 2259.0400 1651.2600 2259.5200 ;
        RECT 1604.6600 2291.6800 1606.2600 2292.1600 ;
        RECT 1604.6600 2297.1200 1606.2600 2297.6000 ;
        RECT 1604.6600 2302.5600 1606.2600 2303.0400 ;
        RECT 1592.9000 2291.6800 1595.9000 2292.1600 ;
        RECT 1592.9000 2297.1200 1595.9000 2297.6000 ;
        RECT 1592.9000 2302.5600 1595.9000 2303.0400 ;
        RECT 1604.6600 2280.8000 1606.2600 2281.2800 ;
        RECT 1604.6600 2286.2400 1606.2600 2286.7200 ;
        RECT 1592.9000 2280.8000 1595.9000 2281.2800 ;
        RECT 1592.9000 2286.2400 1595.9000 2286.7200 ;
        RECT 1604.6600 2264.4800 1606.2600 2264.9600 ;
        RECT 1604.6600 2269.9200 1606.2600 2270.4000 ;
        RECT 1604.6600 2275.3600 1606.2600 2275.8400 ;
        RECT 1592.9000 2264.4800 1595.9000 2264.9600 ;
        RECT 1592.9000 2269.9200 1595.9000 2270.4000 ;
        RECT 1592.9000 2275.3600 1595.9000 2275.8400 ;
        RECT 1604.6600 2253.6000 1606.2600 2254.0800 ;
        RECT 1604.6600 2259.0400 1606.2600 2259.5200 ;
        RECT 1592.9000 2253.6000 1595.9000 2254.0800 ;
        RECT 1592.9000 2259.0400 1595.9000 2259.5200 ;
        RECT 1797.0000 2237.2800 1800.0000 2237.7600 ;
        RECT 1797.0000 2242.7200 1800.0000 2243.2000 ;
        RECT 1797.0000 2248.1600 1800.0000 2248.6400 ;
        RECT 1784.6600 2237.2800 1786.2600 2237.7600 ;
        RECT 1784.6600 2242.7200 1786.2600 2243.2000 ;
        RECT 1784.6600 2248.1600 1786.2600 2248.6400 ;
        RECT 1797.0000 2226.4000 1800.0000 2226.8800 ;
        RECT 1797.0000 2231.8400 1800.0000 2232.3200 ;
        RECT 1784.6600 2226.4000 1786.2600 2226.8800 ;
        RECT 1784.6600 2231.8400 1786.2600 2232.3200 ;
        RECT 1797.0000 2210.0800 1800.0000 2210.5600 ;
        RECT 1797.0000 2215.5200 1800.0000 2216.0000 ;
        RECT 1797.0000 2220.9600 1800.0000 2221.4400 ;
        RECT 1784.6600 2210.0800 1786.2600 2210.5600 ;
        RECT 1784.6600 2215.5200 1786.2600 2216.0000 ;
        RECT 1784.6600 2220.9600 1786.2600 2221.4400 ;
        RECT 1797.0000 2199.2000 1800.0000 2199.6800 ;
        RECT 1797.0000 2204.6400 1800.0000 2205.1200 ;
        RECT 1784.6600 2199.2000 1786.2600 2199.6800 ;
        RECT 1784.6600 2204.6400 1786.2600 2205.1200 ;
        RECT 1739.6600 2237.2800 1741.2600 2237.7600 ;
        RECT 1739.6600 2242.7200 1741.2600 2243.2000 ;
        RECT 1739.6600 2248.1600 1741.2600 2248.6400 ;
        RECT 1739.6600 2226.4000 1741.2600 2226.8800 ;
        RECT 1739.6600 2231.8400 1741.2600 2232.3200 ;
        RECT 1739.6600 2210.0800 1741.2600 2210.5600 ;
        RECT 1739.6600 2215.5200 1741.2600 2216.0000 ;
        RECT 1739.6600 2220.9600 1741.2600 2221.4400 ;
        RECT 1739.6600 2199.2000 1741.2600 2199.6800 ;
        RECT 1739.6600 2204.6400 1741.2600 2205.1200 ;
        RECT 1797.0000 2182.8800 1800.0000 2183.3600 ;
        RECT 1797.0000 2188.3200 1800.0000 2188.8000 ;
        RECT 1797.0000 2193.7600 1800.0000 2194.2400 ;
        RECT 1784.6600 2182.8800 1786.2600 2183.3600 ;
        RECT 1784.6600 2188.3200 1786.2600 2188.8000 ;
        RECT 1784.6600 2193.7600 1786.2600 2194.2400 ;
        RECT 1797.0000 2172.0000 1800.0000 2172.4800 ;
        RECT 1797.0000 2177.4400 1800.0000 2177.9200 ;
        RECT 1784.6600 2172.0000 1786.2600 2172.4800 ;
        RECT 1784.6600 2177.4400 1786.2600 2177.9200 ;
        RECT 1797.0000 2155.6800 1800.0000 2156.1600 ;
        RECT 1797.0000 2161.1200 1800.0000 2161.6000 ;
        RECT 1797.0000 2166.5600 1800.0000 2167.0400 ;
        RECT 1784.6600 2155.6800 1786.2600 2156.1600 ;
        RECT 1784.6600 2161.1200 1786.2600 2161.6000 ;
        RECT 1784.6600 2166.5600 1786.2600 2167.0400 ;
        RECT 1797.0000 2150.2400 1800.0000 2150.7200 ;
        RECT 1784.6600 2150.2400 1786.2600 2150.7200 ;
        RECT 1739.6600 2182.8800 1741.2600 2183.3600 ;
        RECT 1739.6600 2188.3200 1741.2600 2188.8000 ;
        RECT 1739.6600 2193.7600 1741.2600 2194.2400 ;
        RECT 1739.6600 2172.0000 1741.2600 2172.4800 ;
        RECT 1739.6600 2177.4400 1741.2600 2177.9200 ;
        RECT 1739.6600 2155.6800 1741.2600 2156.1600 ;
        RECT 1739.6600 2161.1200 1741.2600 2161.6000 ;
        RECT 1739.6600 2166.5600 1741.2600 2167.0400 ;
        RECT 1739.6600 2150.2400 1741.2600 2150.7200 ;
        RECT 1694.6600 2237.2800 1696.2600 2237.7600 ;
        RECT 1694.6600 2242.7200 1696.2600 2243.2000 ;
        RECT 1694.6600 2248.1600 1696.2600 2248.6400 ;
        RECT 1694.6600 2226.4000 1696.2600 2226.8800 ;
        RECT 1694.6600 2231.8400 1696.2600 2232.3200 ;
        RECT 1649.6600 2237.2800 1651.2600 2237.7600 ;
        RECT 1649.6600 2242.7200 1651.2600 2243.2000 ;
        RECT 1649.6600 2248.1600 1651.2600 2248.6400 ;
        RECT 1649.6600 2226.4000 1651.2600 2226.8800 ;
        RECT 1649.6600 2231.8400 1651.2600 2232.3200 ;
        RECT 1694.6600 2210.0800 1696.2600 2210.5600 ;
        RECT 1694.6600 2215.5200 1696.2600 2216.0000 ;
        RECT 1694.6600 2220.9600 1696.2600 2221.4400 ;
        RECT 1694.6600 2199.2000 1696.2600 2199.6800 ;
        RECT 1694.6600 2204.6400 1696.2600 2205.1200 ;
        RECT 1649.6600 2210.0800 1651.2600 2210.5600 ;
        RECT 1649.6600 2215.5200 1651.2600 2216.0000 ;
        RECT 1649.6600 2220.9600 1651.2600 2221.4400 ;
        RECT 1649.6600 2199.2000 1651.2600 2199.6800 ;
        RECT 1649.6600 2204.6400 1651.2600 2205.1200 ;
        RECT 1604.6600 2237.2800 1606.2600 2237.7600 ;
        RECT 1604.6600 2242.7200 1606.2600 2243.2000 ;
        RECT 1604.6600 2248.1600 1606.2600 2248.6400 ;
        RECT 1592.9000 2237.2800 1595.9000 2237.7600 ;
        RECT 1592.9000 2242.7200 1595.9000 2243.2000 ;
        RECT 1592.9000 2248.1600 1595.9000 2248.6400 ;
        RECT 1604.6600 2226.4000 1606.2600 2226.8800 ;
        RECT 1604.6600 2231.8400 1606.2600 2232.3200 ;
        RECT 1592.9000 2226.4000 1595.9000 2226.8800 ;
        RECT 1592.9000 2231.8400 1595.9000 2232.3200 ;
        RECT 1604.6600 2210.0800 1606.2600 2210.5600 ;
        RECT 1604.6600 2215.5200 1606.2600 2216.0000 ;
        RECT 1604.6600 2220.9600 1606.2600 2221.4400 ;
        RECT 1592.9000 2210.0800 1595.9000 2210.5600 ;
        RECT 1592.9000 2215.5200 1595.9000 2216.0000 ;
        RECT 1592.9000 2220.9600 1595.9000 2221.4400 ;
        RECT 1604.6600 2199.2000 1606.2600 2199.6800 ;
        RECT 1604.6600 2204.6400 1606.2600 2205.1200 ;
        RECT 1592.9000 2199.2000 1595.9000 2199.6800 ;
        RECT 1592.9000 2204.6400 1595.9000 2205.1200 ;
        RECT 1694.6600 2182.8800 1696.2600 2183.3600 ;
        RECT 1694.6600 2188.3200 1696.2600 2188.8000 ;
        RECT 1694.6600 2193.7600 1696.2600 2194.2400 ;
        RECT 1694.6600 2172.0000 1696.2600 2172.4800 ;
        RECT 1694.6600 2177.4400 1696.2600 2177.9200 ;
        RECT 1649.6600 2182.8800 1651.2600 2183.3600 ;
        RECT 1649.6600 2188.3200 1651.2600 2188.8000 ;
        RECT 1649.6600 2193.7600 1651.2600 2194.2400 ;
        RECT 1649.6600 2172.0000 1651.2600 2172.4800 ;
        RECT 1649.6600 2177.4400 1651.2600 2177.9200 ;
        RECT 1694.6600 2155.6800 1696.2600 2156.1600 ;
        RECT 1694.6600 2161.1200 1696.2600 2161.6000 ;
        RECT 1694.6600 2166.5600 1696.2600 2167.0400 ;
        RECT 1694.6600 2150.2400 1696.2600 2150.7200 ;
        RECT 1649.6600 2155.6800 1651.2600 2156.1600 ;
        RECT 1649.6600 2161.1200 1651.2600 2161.6000 ;
        RECT 1649.6600 2166.5600 1651.2600 2167.0400 ;
        RECT 1649.6600 2150.2400 1651.2600 2150.7200 ;
        RECT 1604.6600 2182.8800 1606.2600 2183.3600 ;
        RECT 1604.6600 2188.3200 1606.2600 2188.8000 ;
        RECT 1604.6600 2193.7600 1606.2600 2194.2400 ;
        RECT 1592.9000 2182.8800 1595.9000 2183.3600 ;
        RECT 1592.9000 2188.3200 1595.9000 2188.8000 ;
        RECT 1592.9000 2193.7600 1595.9000 2194.2400 ;
        RECT 1604.6600 2172.0000 1606.2600 2172.4800 ;
        RECT 1604.6600 2177.4400 1606.2600 2177.9200 ;
        RECT 1592.9000 2172.0000 1595.9000 2172.4800 ;
        RECT 1592.9000 2177.4400 1595.9000 2177.9200 ;
        RECT 1604.6600 2155.6800 1606.2600 2156.1600 ;
        RECT 1604.6600 2161.1200 1606.2600 2161.6000 ;
        RECT 1604.6600 2166.5600 1606.2600 2167.0400 ;
        RECT 1592.9000 2155.6800 1595.9000 2156.1600 ;
        RECT 1592.9000 2161.1200 1595.9000 2161.6000 ;
        RECT 1592.9000 2166.5600 1595.9000 2167.0400 ;
        RECT 1592.9000 2150.2400 1595.9000 2150.7200 ;
        RECT 1604.6600 2150.2400 1606.2600 2150.7200 ;
        RECT 1592.9000 2355.1500 1800.0000 2358.1500 ;
        RECT 1592.9000 2142.0500 1800.0000 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 1912.4100 1786.2600 2128.5100 ;
        RECT 1739.6600 1912.4100 1741.2600 2128.5100 ;
        RECT 1694.6600 1912.4100 1696.2600 2128.5100 ;
        RECT 1649.6600 1912.4100 1651.2600 2128.5100 ;
        RECT 1604.6600 1912.4100 1606.2600 2128.5100 ;
        RECT 1797.0000 1912.4100 1800.0000 2128.5100 ;
        RECT 1592.9000 1912.4100 1595.9000 2128.5100 ;
      LAYER met3 ;
        RECT 1797.0000 2105.5600 1800.0000 2106.0400 ;
        RECT 1797.0000 2111.0000 1800.0000 2111.4800 ;
        RECT 1784.6600 2105.5600 1786.2600 2106.0400 ;
        RECT 1784.6600 2111.0000 1786.2600 2111.4800 ;
        RECT 1797.0000 2116.4400 1800.0000 2116.9200 ;
        RECT 1784.6600 2116.4400 1786.2600 2116.9200 ;
        RECT 1797.0000 2094.6800 1800.0000 2095.1600 ;
        RECT 1797.0000 2100.1200 1800.0000 2100.6000 ;
        RECT 1784.6600 2094.6800 1786.2600 2095.1600 ;
        RECT 1784.6600 2100.1200 1786.2600 2100.6000 ;
        RECT 1797.0000 2078.3600 1800.0000 2078.8400 ;
        RECT 1797.0000 2083.8000 1800.0000 2084.2800 ;
        RECT 1784.6600 2078.3600 1786.2600 2078.8400 ;
        RECT 1784.6600 2083.8000 1786.2600 2084.2800 ;
        RECT 1797.0000 2089.2400 1800.0000 2089.7200 ;
        RECT 1784.6600 2089.2400 1786.2600 2089.7200 ;
        RECT 1739.6600 2105.5600 1741.2600 2106.0400 ;
        RECT 1739.6600 2111.0000 1741.2600 2111.4800 ;
        RECT 1739.6600 2116.4400 1741.2600 2116.9200 ;
        RECT 1739.6600 2094.6800 1741.2600 2095.1600 ;
        RECT 1739.6600 2100.1200 1741.2600 2100.6000 ;
        RECT 1739.6600 2078.3600 1741.2600 2078.8400 ;
        RECT 1739.6600 2083.8000 1741.2600 2084.2800 ;
        RECT 1739.6600 2089.2400 1741.2600 2089.7200 ;
        RECT 1797.0000 2062.0400 1800.0000 2062.5200 ;
        RECT 1797.0000 2067.4800 1800.0000 2067.9600 ;
        RECT 1797.0000 2072.9200 1800.0000 2073.4000 ;
        RECT 1784.6600 2062.0400 1786.2600 2062.5200 ;
        RECT 1784.6600 2067.4800 1786.2600 2067.9600 ;
        RECT 1784.6600 2072.9200 1786.2600 2073.4000 ;
        RECT 1797.0000 2051.1600 1800.0000 2051.6400 ;
        RECT 1797.0000 2056.6000 1800.0000 2057.0800 ;
        RECT 1784.6600 2051.1600 1786.2600 2051.6400 ;
        RECT 1784.6600 2056.6000 1786.2600 2057.0800 ;
        RECT 1797.0000 2034.8400 1800.0000 2035.3200 ;
        RECT 1797.0000 2040.2800 1800.0000 2040.7600 ;
        RECT 1797.0000 2045.7200 1800.0000 2046.2000 ;
        RECT 1784.6600 2034.8400 1786.2600 2035.3200 ;
        RECT 1784.6600 2040.2800 1786.2600 2040.7600 ;
        RECT 1784.6600 2045.7200 1786.2600 2046.2000 ;
        RECT 1797.0000 2023.9600 1800.0000 2024.4400 ;
        RECT 1797.0000 2029.4000 1800.0000 2029.8800 ;
        RECT 1784.6600 2023.9600 1786.2600 2024.4400 ;
        RECT 1784.6600 2029.4000 1786.2600 2029.8800 ;
        RECT 1739.6600 2062.0400 1741.2600 2062.5200 ;
        RECT 1739.6600 2067.4800 1741.2600 2067.9600 ;
        RECT 1739.6600 2072.9200 1741.2600 2073.4000 ;
        RECT 1739.6600 2051.1600 1741.2600 2051.6400 ;
        RECT 1739.6600 2056.6000 1741.2600 2057.0800 ;
        RECT 1739.6600 2034.8400 1741.2600 2035.3200 ;
        RECT 1739.6600 2040.2800 1741.2600 2040.7600 ;
        RECT 1739.6600 2045.7200 1741.2600 2046.2000 ;
        RECT 1739.6600 2023.9600 1741.2600 2024.4400 ;
        RECT 1739.6600 2029.4000 1741.2600 2029.8800 ;
        RECT 1694.6600 2105.5600 1696.2600 2106.0400 ;
        RECT 1694.6600 2111.0000 1696.2600 2111.4800 ;
        RECT 1694.6600 2116.4400 1696.2600 2116.9200 ;
        RECT 1649.6600 2105.5600 1651.2600 2106.0400 ;
        RECT 1649.6600 2111.0000 1651.2600 2111.4800 ;
        RECT 1649.6600 2116.4400 1651.2600 2116.9200 ;
        RECT 1694.6600 2094.6800 1696.2600 2095.1600 ;
        RECT 1694.6600 2100.1200 1696.2600 2100.6000 ;
        RECT 1694.6600 2078.3600 1696.2600 2078.8400 ;
        RECT 1694.6600 2083.8000 1696.2600 2084.2800 ;
        RECT 1694.6600 2089.2400 1696.2600 2089.7200 ;
        RECT 1649.6600 2094.6800 1651.2600 2095.1600 ;
        RECT 1649.6600 2100.1200 1651.2600 2100.6000 ;
        RECT 1649.6600 2078.3600 1651.2600 2078.8400 ;
        RECT 1649.6600 2083.8000 1651.2600 2084.2800 ;
        RECT 1649.6600 2089.2400 1651.2600 2089.7200 ;
        RECT 1604.6600 2105.5600 1606.2600 2106.0400 ;
        RECT 1604.6600 2111.0000 1606.2600 2111.4800 ;
        RECT 1592.9000 2111.0000 1595.9000 2111.4800 ;
        RECT 1592.9000 2105.5600 1595.9000 2106.0400 ;
        RECT 1592.9000 2116.4400 1595.9000 2116.9200 ;
        RECT 1604.6600 2116.4400 1606.2600 2116.9200 ;
        RECT 1604.6600 2094.6800 1606.2600 2095.1600 ;
        RECT 1604.6600 2100.1200 1606.2600 2100.6000 ;
        RECT 1592.9000 2100.1200 1595.9000 2100.6000 ;
        RECT 1592.9000 2094.6800 1595.9000 2095.1600 ;
        RECT 1604.6600 2078.3600 1606.2600 2078.8400 ;
        RECT 1604.6600 2083.8000 1606.2600 2084.2800 ;
        RECT 1592.9000 2083.8000 1595.9000 2084.2800 ;
        RECT 1592.9000 2078.3600 1595.9000 2078.8400 ;
        RECT 1592.9000 2089.2400 1595.9000 2089.7200 ;
        RECT 1604.6600 2089.2400 1606.2600 2089.7200 ;
        RECT 1694.6600 2062.0400 1696.2600 2062.5200 ;
        RECT 1694.6600 2067.4800 1696.2600 2067.9600 ;
        RECT 1694.6600 2072.9200 1696.2600 2073.4000 ;
        RECT 1694.6600 2051.1600 1696.2600 2051.6400 ;
        RECT 1694.6600 2056.6000 1696.2600 2057.0800 ;
        RECT 1649.6600 2062.0400 1651.2600 2062.5200 ;
        RECT 1649.6600 2067.4800 1651.2600 2067.9600 ;
        RECT 1649.6600 2072.9200 1651.2600 2073.4000 ;
        RECT 1649.6600 2051.1600 1651.2600 2051.6400 ;
        RECT 1649.6600 2056.6000 1651.2600 2057.0800 ;
        RECT 1694.6600 2034.8400 1696.2600 2035.3200 ;
        RECT 1694.6600 2040.2800 1696.2600 2040.7600 ;
        RECT 1694.6600 2045.7200 1696.2600 2046.2000 ;
        RECT 1694.6600 2023.9600 1696.2600 2024.4400 ;
        RECT 1694.6600 2029.4000 1696.2600 2029.8800 ;
        RECT 1649.6600 2034.8400 1651.2600 2035.3200 ;
        RECT 1649.6600 2040.2800 1651.2600 2040.7600 ;
        RECT 1649.6600 2045.7200 1651.2600 2046.2000 ;
        RECT 1649.6600 2023.9600 1651.2600 2024.4400 ;
        RECT 1649.6600 2029.4000 1651.2600 2029.8800 ;
        RECT 1604.6600 2062.0400 1606.2600 2062.5200 ;
        RECT 1604.6600 2067.4800 1606.2600 2067.9600 ;
        RECT 1604.6600 2072.9200 1606.2600 2073.4000 ;
        RECT 1592.9000 2062.0400 1595.9000 2062.5200 ;
        RECT 1592.9000 2067.4800 1595.9000 2067.9600 ;
        RECT 1592.9000 2072.9200 1595.9000 2073.4000 ;
        RECT 1604.6600 2051.1600 1606.2600 2051.6400 ;
        RECT 1604.6600 2056.6000 1606.2600 2057.0800 ;
        RECT 1592.9000 2051.1600 1595.9000 2051.6400 ;
        RECT 1592.9000 2056.6000 1595.9000 2057.0800 ;
        RECT 1604.6600 2034.8400 1606.2600 2035.3200 ;
        RECT 1604.6600 2040.2800 1606.2600 2040.7600 ;
        RECT 1604.6600 2045.7200 1606.2600 2046.2000 ;
        RECT 1592.9000 2034.8400 1595.9000 2035.3200 ;
        RECT 1592.9000 2040.2800 1595.9000 2040.7600 ;
        RECT 1592.9000 2045.7200 1595.9000 2046.2000 ;
        RECT 1604.6600 2023.9600 1606.2600 2024.4400 ;
        RECT 1604.6600 2029.4000 1606.2600 2029.8800 ;
        RECT 1592.9000 2023.9600 1595.9000 2024.4400 ;
        RECT 1592.9000 2029.4000 1595.9000 2029.8800 ;
        RECT 1797.0000 2007.6400 1800.0000 2008.1200 ;
        RECT 1797.0000 2013.0800 1800.0000 2013.5600 ;
        RECT 1797.0000 2018.5200 1800.0000 2019.0000 ;
        RECT 1784.6600 2007.6400 1786.2600 2008.1200 ;
        RECT 1784.6600 2013.0800 1786.2600 2013.5600 ;
        RECT 1784.6600 2018.5200 1786.2600 2019.0000 ;
        RECT 1797.0000 1996.7600 1800.0000 1997.2400 ;
        RECT 1797.0000 2002.2000 1800.0000 2002.6800 ;
        RECT 1784.6600 1996.7600 1786.2600 1997.2400 ;
        RECT 1784.6600 2002.2000 1786.2600 2002.6800 ;
        RECT 1797.0000 1980.4400 1800.0000 1980.9200 ;
        RECT 1797.0000 1985.8800 1800.0000 1986.3600 ;
        RECT 1797.0000 1991.3200 1800.0000 1991.8000 ;
        RECT 1784.6600 1980.4400 1786.2600 1980.9200 ;
        RECT 1784.6600 1985.8800 1786.2600 1986.3600 ;
        RECT 1784.6600 1991.3200 1786.2600 1991.8000 ;
        RECT 1797.0000 1969.5600 1800.0000 1970.0400 ;
        RECT 1797.0000 1975.0000 1800.0000 1975.4800 ;
        RECT 1784.6600 1969.5600 1786.2600 1970.0400 ;
        RECT 1784.6600 1975.0000 1786.2600 1975.4800 ;
        RECT 1739.6600 2007.6400 1741.2600 2008.1200 ;
        RECT 1739.6600 2013.0800 1741.2600 2013.5600 ;
        RECT 1739.6600 2018.5200 1741.2600 2019.0000 ;
        RECT 1739.6600 1996.7600 1741.2600 1997.2400 ;
        RECT 1739.6600 2002.2000 1741.2600 2002.6800 ;
        RECT 1739.6600 1980.4400 1741.2600 1980.9200 ;
        RECT 1739.6600 1985.8800 1741.2600 1986.3600 ;
        RECT 1739.6600 1991.3200 1741.2600 1991.8000 ;
        RECT 1739.6600 1969.5600 1741.2600 1970.0400 ;
        RECT 1739.6600 1975.0000 1741.2600 1975.4800 ;
        RECT 1797.0000 1953.2400 1800.0000 1953.7200 ;
        RECT 1797.0000 1958.6800 1800.0000 1959.1600 ;
        RECT 1797.0000 1964.1200 1800.0000 1964.6000 ;
        RECT 1784.6600 1953.2400 1786.2600 1953.7200 ;
        RECT 1784.6600 1958.6800 1786.2600 1959.1600 ;
        RECT 1784.6600 1964.1200 1786.2600 1964.6000 ;
        RECT 1797.0000 1942.3600 1800.0000 1942.8400 ;
        RECT 1797.0000 1947.8000 1800.0000 1948.2800 ;
        RECT 1784.6600 1942.3600 1786.2600 1942.8400 ;
        RECT 1784.6600 1947.8000 1786.2600 1948.2800 ;
        RECT 1797.0000 1926.0400 1800.0000 1926.5200 ;
        RECT 1797.0000 1931.4800 1800.0000 1931.9600 ;
        RECT 1797.0000 1936.9200 1800.0000 1937.4000 ;
        RECT 1784.6600 1926.0400 1786.2600 1926.5200 ;
        RECT 1784.6600 1931.4800 1786.2600 1931.9600 ;
        RECT 1784.6600 1936.9200 1786.2600 1937.4000 ;
        RECT 1797.0000 1920.6000 1800.0000 1921.0800 ;
        RECT 1784.6600 1920.6000 1786.2600 1921.0800 ;
        RECT 1739.6600 1953.2400 1741.2600 1953.7200 ;
        RECT 1739.6600 1958.6800 1741.2600 1959.1600 ;
        RECT 1739.6600 1964.1200 1741.2600 1964.6000 ;
        RECT 1739.6600 1942.3600 1741.2600 1942.8400 ;
        RECT 1739.6600 1947.8000 1741.2600 1948.2800 ;
        RECT 1739.6600 1926.0400 1741.2600 1926.5200 ;
        RECT 1739.6600 1931.4800 1741.2600 1931.9600 ;
        RECT 1739.6600 1936.9200 1741.2600 1937.4000 ;
        RECT 1739.6600 1920.6000 1741.2600 1921.0800 ;
        RECT 1694.6600 2007.6400 1696.2600 2008.1200 ;
        RECT 1694.6600 2013.0800 1696.2600 2013.5600 ;
        RECT 1694.6600 2018.5200 1696.2600 2019.0000 ;
        RECT 1694.6600 1996.7600 1696.2600 1997.2400 ;
        RECT 1694.6600 2002.2000 1696.2600 2002.6800 ;
        RECT 1649.6600 2007.6400 1651.2600 2008.1200 ;
        RECT 1649.6600 2013.0800 1651.2600 2013.5600 ;
        RECT 1649.6600 2018.5200 1651.2600 2019.0000 ;
        RECT 1649.6600 1996.7600 1651.2600 1997.2400 ;
        RECT 1649.6600 2002.2000 1651.2600 2002.6800 ;
        RECT 1694.6600 1980.4400 1696.2600 1980.9200 ;
        RECT 1694.6600 1985.8800 1696.2600 1986.3600 ;
        RECT 1694.6600 1991.3200 1696.2600 1991.8000 ;
        RECT 1694.6600 1969.5600 1696.2600 1970.0400 ;
        RECT 1694.6600 1975.0000 1696.2600 1975.4800 ;
        RECT 1649.6600 1980.4400 1651.2600 1980.9200 ;
        RECT 1649.6600 1985.8800 1651.2600 1986.3600 ;
        RECT 1649.6600 1991.3200 1651.2600 1991.8000 ;
        RECT 1649.6600 1969.5600 1651.2600 1970.0400 ;
        RECT 1649.6600 1975.0000 1651.2600 1975.4800 ;
        RECT 1604.6600 2007.6400 1606.2600 2008.1200 ;
        RECT 1604.6600 2013.0800 1606.2600 2013.5600 ;
        RECT 1604.6600 2018.5200 1606.2600 2019.0000 ;
        RECT 1592.9000 2007.6400 1595.9000 2008.1200 ;
        RECT 1592.9000 2013.0800 1595.9000 2013.5600 ;
        RECT 1592.9000 2018.5200 1595.9000 2019.0000 ;
        RECT 1604.6600 1996.7600 1606.2600 1997.2400 ;
        RECT 1604.6600 2002.2000 1606.2600 2002.6800 ;
        RECT 1592.9000 1996.7600 1595.9000 1997.2400 ;
        RECT 1592.9000 2002.2000 1595.9000 2002.6800 ;
        RECT 1604.6600 1980.4400 1606.2600 1980.9200 ;
        RECT 1604.6600 1985.8800 1606.2600 1986.3600 ;
        RECT 1604.6600 1991.3200 1606.2600 1991.8000 ;
        RECT 1592.9000 1980.4400 1595.9000 1980.9200 ;
        RECT 1592.9000 1985.8800 1595.9000 1986.3600 ;
        RECT 1592.9000 1991.3200 1595.9000 1991.8000 ;
        RECT 1604.6600 1969.5600 1606.2600 1970.0400 ;
        RECT 1604.6600 1975.0000 1606.2600 1975.4800 ;
        RECT 1592.9000 1969.5600 1595.9000 1970.0400 ;
        RECT 1592.9000 1975.0000 1595.9000 1975.4800 ;
        RECT 1694.6600 1953.2400 1696.2600 1953.7200 ;
        RECT 1694.6600 1958.6800 1696.2600 1959.1600 ;
        RECT 1694.6600 1964.1200 1696.2600 1964.6000 ;
        RECT 1694.6600 1942.3600 1696.2600 1942.8400 ;
        RECT 1694.6600 1947.8000 1696.2600 1948.2800 ;
        RECT 1649.6600 1953.2400 1651.2600 1953.7200 ;
        RECT 1649.6600 1958.6800 1651.2600 1959.1600 ;
        RECT 1649.6600 1964.1200 1651.2600 1964.6000 ;
        RECT 1649.6600 1942.3600 1651.2600 1942.8400 ;
        RECT 1649.6600 1947.8000 1651.2600 1948.2800 ;
        RECT 1694.6600 1926.0400 1696.2600 1926.5200 ;
        RECT 1694.6600 1931.4800 1696.2600 1931.9600 ;
        RECT 1694.6600 1936.9200 1696.2600 1937.4000 ;
        RECT 1694.6600 1920.6000 1696.2600 1921.0800 ;
        RECT 1649.6600 1926.0400 1651.2600 1926.5200 ;
        RECT 1649.6600 1931.4800 1651.2600 1931.9600 ;
        RECT 1649.6600 1936.9200 1651.2600 1937.4000 ;
        RECT 1649.6600 1920.6000 1651.2600 1921.0800 ;
        RECT 1604.6600 1953.2400 1606.2600 1953.7200 ;
        RECT 1604.6600 1958.6800 1606.2600 1959.1600 ;
        RECT 1604.6600 1964.1200 1606.2600 1964.6000 ;
        RECT 1592.9000 1953.2400 1595.9000 1953.7200 ;
        RECT 1592.9000 1958.6800 1595.9000 1959.1600 ;
        RECT 1592.9000 1964.1200 1595.9000 1964.6000 ;
        RECT 1604.6600 1942.3600 1606.2600 1942.8400 ;
        RECT 1604.6600 1947.8000 1606.2600 1948.2800 ;
        RECT 1592.9000 1942.3600 1595.9000 1942.8400 ;
        RECT 1592.9000 1947.8000 1595.9000 1948.2800 ;
        RECT 1604.6600 1926.0400 1606.2600 1926.5200 ;
        RECT 1604.6600 1931.4800 1606.2600 1931.9600 ;
        RECT 1604.6600 1936.9200 1606.2600 1937.4000 ;
        RECT 1592.9000 1926.0400 1595.9000 1926.5200 ;
        RECT 1592.9000 1931.4800 1595.9000 1931.9600 ;
        RECT 1592.9000 1936.9200 1595.9000 1937.4000 ;
        RECT 1592.9000 1920.6000 1595.9000 1921.0800 ;
        RECT 1604.6600 1920.6000 1606.2600 1921.0800 ;
        RECT 1592.9000 2125.5100 1800.0000 2128.5100 ;
        RECT 1592.9000 1912.4100 1800.0000 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 1682.7700 1786.2600 1898.8700 ;
        RECT 1739.6600 1682.7700 1741.2600 1898.8700 ;
        RECT 1694.6600 1682.7700 1696.2600 1898.8700 ;
        RECT 1649.6600 1682.7700 1651.2600 1898.8700 ;
        RECT 1604.6600 1682.7700 1606.2600 1898.8700 ;
        RECT 1797.0000 1682.7700 1800.0000 1898.8700 ;
        RECT 1592.9000 1682.7700 1595.9000 1898.8700 ;
      LAYER met3 ;
        RECT 1797.0000 1875.9200 1800.0000 1876.4000 ;
        RECT 1797.0000 1881.3600 1800.0000 1881.8400 ;
        RECT 1784.6600 1875.9200 1786.2600 1876.4000 ;
        RECT 1784.6600 1881.3600 1786.2600 1881.8400 ;
        RECT 1797.0000 1886.8000 1800.0000 1887.2800 ;
        RECT 1784.6600 1886.8000 1786.2600 1887.2800 ;
        RECT 1797.0000 1865.0400 1800.0000 1865.5200 ;
        RECT 1797.0000 1870.4800 1800.0000 1870.9600 ;
        RECT 1784.6600 1865.0400 1786.2600 1865.5200 ;
        RECT 1784.6600 1870.4800 1786.2600 1870.9600 ;
        RECT 1797.0000 1848.7200 1800.0000 1849.2000 ;
        RECT 1797.0000 1854.1600 1800.0000 1854.6400 ;
        RECT 1784.6600 1848.7200 1786.2600 1849.2000 ;
        RECT 1784.6600 1854.1600 1786.2600 1854.6400 ;
        RECT 1797.0000 1859.6000 1800.0000 1860.0800 ;
        RECT 1784.6600 1859.6000 1786.2600 1860.0800 ;
        RECT 1739.6600 1875.9200 1741.2600 1876.4000 ;
        RECT 1739.6600 1881.3600 1741.2600 1881.8400 ;
        RECT 1739.6600 1886.8000 1741.2600 1887.2800 ;
        RECT 1739.6600 1865.0400 1741.2600 1865.5200 ;
        RECT 1739.6600 1870.4800 1741.2600 1870.9600 ;
        RECT 1739.6600 1848.7200 1741.2600 1849.2000 ;
        RECT 1739.6600 1854.1600 1741.2600 1854.6400 ;
        RECT 1739.6600 1859.6000 1741.2600 1860.0800 ;
        RECT 1797.0000 1832.4000 1800.0000 1832.8800 ;
        RECT 1797.0000 1837.8400 1800.0000 1838.3200 ;
        RECT 1797.0000 1843.2800 1800.0000 1843.7600 ;
        RECT 1784.6600 1832.4000 1786.2600 1832.8800 ;
        RECT 1784.6600 1837.8400 1786.2600 1838.3200 ;
        RECT 1784.6600 1843.2800 1786.2600 1843.7600 ;
        RECT 1797.0000 1821.5200 1800.0000 1822.0000 ;
        RECT 1797.0000 1826.9600 1800.0000 1827.4400 ;
        RECT 1784.6600 1821.5200 1786.2600 1822.0000 ;
        RECT 1784.6600 1826.9600 1786.2600 1827.4400 ;
        RECT 1797.0000 1805.2000 1800.0000 1805.6800 ;
        RECT 1797.0000 1810.6400 1800.0000 1811.1200 ;
        RECT 1797.0000 1816.0800 1800.0000 1816.5600 ;
        RECT 1784.6600 1805.2000 1786.2600 1805.6800 ;
        RECT 1784.6600 1810.6400 1786.2600 1811.1200 ;
        RECT 1784.6600 1816.0800 1786.2600 1816.5600 ;
        RECT 1797.0000 1794.3200 1800.0000 1794.8000 ;
        RECT 1797.0000 1799.7600 1800.0000 1800.2400 ;
        RECT 1784.6600 1794.3200 1786.2600 1794.8000 ;
        RECT 1784.6600 1799.7600 1786.2600 1800.2400 ;
        RECT 1739.6600 1832.4000 1741.2600 1832.8800 ;
        RECT 1739.6600 1837.8400 1741.2600 1838.3200 ;
        RECT 1739.6600 1843.2800 1741.2600 1843.7600 ;
        RECT 1739.6600 1821.5200 1741.2600 1822.0000 ;
        RECT 1739.6600 1826.9600 1741.2600 1827.4400 ;
        RECT 1739.6600 1805.2000 1741.2600 1805.6800 ;
        RECT 1739.6600 1810.6400 1741.2600 1811.1200 ;
        RECT 1739.6600 1816.0800 1741.2600 1816.5600 ;
        RECT 1739.6600 1794.3200 1741.2600 1794.8000 ;
        RECT 1739.6600 1799.7600 1741.2600 1800.2400 ;
        RECT 1694.6600 1875.9200 1696.2600 1876.4000 ;
        RECT 1694.6600 1881.3600 1696.2600 1881.8400 ;
        RECT 1694.6600 1886.8000 1696.2600 1887.2800 ;
        RECT 1649.6600 1875.9200 1651.2600 1876.4000 ;
        RECT 1649.6600 1881.3600 1651.2600 1881.8400 ;
        RECT 1649.6600 1886.8000 1651.2600 1887.2800 ;
        RECT 1694.6600 1865.0400 1696.2600 1865.5200 ;
        RECT 1694.6600 1870.4800 1696.2600 1870.9600 ;
        RECT 1694.6600 1848.7200 1696.2600 1849.2000 ;
        RECT 1694.6600 1854.1600 1696.2600 1854.6400 ;
        RECT 1694.6600 1859.6000 1696.2600 1860.0800 ;
        RECT 1649.6600 1865.0400 1651.2600 1865.5200 ;
        RECT 1649.6600 1870.4800 1651.2600 1870.9600 ;
        RECT 1649.6600 1848.7200 1651.2600 1849.2000 ;
        RECT 1649.6600 1854.1600 1651.2600 1854.6400 ;
        RECT 1649.6600 1859.6000 1651.2600 1860.0800 ;
        RECT 1604.6600 1875.9200 1606.2600 1876.4000 ;
        RECT 1604.6600 1881.3600 1606.2600 1881.8400 ;
        RECT 1592.9000 1881.3600 1595.9000 1881.8400 ;
        RECT 1592.9000 1875.9200 1595.9000 1876.4000 ;
        RECT 1592.9000 1886.8000 1595.9000 1887.2800 ;
        RECT 1604.6600 1886.8000 1606.2600 1887.2800 ;
        RECT 1604.6600 1865.0400 1606.2600 1865.5200 ;
        RECT 1604.6600 1870.4800 1606.2600 1870.9600 ;
        RECT 1592.9000 1870.4800 1595.9000 1870.9600 ;
        RECT 1592.9000 1865.0400 1595.9000 1865.5200 ;
        RECT 1604.6600 1848.7200 1606.2600 1849.2000 ;
        RECT 1604.6600 1854.1600 1606.2600 1854.6400 ;
        RECT 1592.9000 1854.1600 1595.9000 1854.6400 ;
        RECT 1592.9000 1848.7200 1595.9000 1849.2000 ;
        RECT 1592.9000 1859.6000 1595.9000 1860.0800 ;
        RECT 1604.6600 1859.6000 1606.2600 1860.0800 ;
        RECT 1694.6600 1832.4000 1696.2600 1832.8800 ;
        RECT 1694.6600 1837.8400 1696.2600 1838.3200 ;
        RECT 1694.6600 1843.2800 1696.2600 1843.7600 ;
        RECT 1694.6600 1821.5200 1696.2600 1822.0000 ;
        RECT 1694.6600 1826.9600 1696.2600 1827.4400 ;
        RECT 1649.6600 1832.4000 1651.2600 1832.8800 ;
        RECT 1649.6600 1837.8400 1651.2600 1838.3200 ;
        RECT 1649.6600 1843.2800 1651.2600 1843.7600 ;
        RECT 1649.6600 1821.5200 1651.2600 1822.0000 ;
        RECT 1649.6600 1826.9600 1651.2600 1827.4400 ;
        RECT 1694.6600 1805.2000 1696.2600 1805.6800 ;
        RECT 1694.6600 1810.6400 1696.2600 1811.1200 ;
        RECT 1694.6600 1816.0800 1696.2600 1816.5600 ;
        RECT 1694.6600 1794.3200 1696.2600 1794.8000 ;
        RECT 1694.6600 1799.7600 1696.2600 1800.2400 ;
        RECT 1649.6600 1805.2000 1651.2600 1805.6800 ;
        RECT 1649.6600 1810.6400 1651.2600 1811.1200 ;
        RECT 1649.6600 1816.0800 1651.2600 1816.5600 ;
        RECT 1649.6600 1794.3200 1651.2600 1794.8000 ;
        RECT 1649.6600 1799.7600 1651.2600 1800.2400 ;
        RECT 1604.6600 1832.4000 1606.2600 1832.8800 ;
        RECT 1604.6600 1837.8400 1606.2600 1838.3200 ;
        RECT 1604.6600 1843.2800 1606.2600 1843.7600 ;
        RECT 1592.9000 1832.4000 1595.9000 1832.8800 ;
        RECT 1592.9000 1837.8400 1595.9000 1838.3200 ;
        RECT 1592.9000 1843.2800 1595.9000 1843.7600 ;
        RECT 1604.6600 1821.5200 1606.2600 1822.0000 ;
        RECT 1604.6600 1826.9600 1606.2600 1827.4400 ;
        RECT 1592.9000 1821.5200 1595.9000 1822.0000 ;
        RECT 1592.9000 1826.9600 1595.9000 1827.4400 ;
        RECT 1604.6600 1805.2000 1606.2600 1805.6800 ;
        RECT 1604.6600 1810.6400 1606.2600 1811.1200 ;
        RECT 1604.6600 1816.0800 1606.2600 1816.5600 ;
        RECT 1592.9000 1805.2000 1595.9000 1805.6800 ;
        RECT 1592.9000 1810.6400 1595.9000 1811.1200 ;
        RECT 1592.9000 1816.0800 1595.9000 1816.5600 ;
        RECT 1604.6600 1794.3200 1606.2600 1794.8000 ;
        RECT 1604.6600 1799.7600 1606.2600 1800.2400 ;
        RECT 1592.9000 1794.3200 1595.9000 1794.8000 ;
        RECT 1592.9000 1799.7600 1595.9000 1800.2400 ;
        RECT 1797.0000 1778.0000 1800.0000 1778.4800 ;
        RECT 1797.0000 1783.4400 1800.0000 1783.9200 ;
        RECT 1797.0000 1788.8800 1800.0000 1789.3600 ;
        RECT 1784.6600 1778.0000 1786.2600 1778.4800 ;
        RECT 1784.6600 1783.4400 1786.2600 1783.9200 ;
        RECT 1784.6600 1788.8800 1786.2600 1789.3600 ;
        RECT 1797.0000 1767.1200 1800.0000 1767.6000 ;
        RECT 1797.0000 1772.5600 1800.0000 1773.0400 ;
        RECT 1784.6600 1767.1200 1786.2600 1767.6000 ;
        RECT 1784.6600 1772.5600 1786.2600 1773.0400 ;
        RECT 1797.0000 1750.8000 1800.0000 1751.2800 ;
        RECT 1797.0000 1756.2400 1800.0000 1756.7200 ;
        RECT 1797.0000 1761.6800 1800.0000 1762.1600 ;
        RECT 1784.6600 1750.8000 1786.2600 1751.2800 ;
        RECT 1784.6600 1756.2400 1786.2600 1756.7200 ;
        RECT 1784.6600 1761.6800 1786.2600 1762.1600 ;
        RECT 1797.0000 1739.9200 1800.0000 1740.4000 ;
        RECT 1797.0000 1745.3600 1800.0000 1745.8400 ;
        RECT 1784.6600 1739.9200 1786.2600 1740.4000 ;
        RECT 1784.6600 1745.3600 1786.2600 1745.8400 ;
        RECT 1739.6600 1778.0000 1741.2600 1778.4800 ;
        RECT 1739.6600 1783.4400 1741.2600 1783.9200 ;
        RECT 1739.6600 1788.8800 1741.2600 1789.3600 ;
        RECT 1739.6600 1767.1200 1741.2600 1767.6000 ;
        RECT 1739.6600 1772.5600 1741.2600 1773.0400 ;
        RECT 1739.6600 1750.8000 1741.2600 1751.2800 ;
        RECT 1739.6600 1756.2400 1741.2600 1756.7200 ;
        RECT 1739.6600 1761.6800 1741.2600 1762.1600 ;
        RECT 1739.6600 1739.9200 1741.2600 1740.4000 ;
        RECT 1739.6600 1745.3600 1741.2600 1745.8400 ;
        RECT 1797.0000 1723.6000 1800.0000 1724.0800 ;
        RECT 1797.0000 1729.0400 1800.0000 1729.5200 ;
        RECT 1797.0000 1734.4800 1800.0000 1734.9600 ;
        RECT 1784.6600 1723.6000 1786.2600 1724.0800 ;
        RECT 1784.6600 1729.0400 1786.2600 1729.5200 ;
        RECT 1784.6600 1734.4800 1786.2600 1734.9600 ;
        RECT 1797.0000 1712.7200 1800.0000 1713.2000 ;
        RECT 1797.0000 1718.1600 1800.0000 1718.6400 ;
        RECT 1784.6600 1712.7200 1786.2600 1713.2000 ;
        RECT 1784.6600 1718.1600 1786.2600 1718.6400 ;
        RECT 1797.0000 1696.4000 1800.0000 1696.8800 ;
        RECT 1797.0000 1701.8400 1800.0000 1702.3200 ;
        RECT 1797.0000 1707.2800 1800.0000 1707.7600 ;
        RECT 1784.6600 1696.4000 1786.2600 1696.8800 ;
        RECT 1784.6600 1701.8400 1786.2600 1702.3200 ;
        RECT 1784.6600 1707.2800 1786.2600 1707.7600 ;
        RECT 1797.0000 1690.9600 1800.0000 1691.4400 ;
        RECT 1784.6600 1690.9600 1786.2600 1691.4400 ;
        RECT 1739.6600 1723.6000 1741.2600 1724.0800 ;
        RECT 1739.6600 1729.0400 1741.2600 1729.5200 ;
        RECT 1739.6600 1734.4800 1741.2600 1734.9600 ;
        RECT 1739.6600 1712.7200 1741.2600 1713.2000 ;
        RECT 1739.6600 1718.1600 1741.2600 1718.6400 ;
        RECT 1739.6600 1696.4000 1741.2600 1696.8800 ;
        RECT 1739.6600 1701.8400 1741.2600 1702.3200 ;
        RECT 1739.6600 1707.2800 1741.2600 1707.7600 ;
        RECT 1739.6600 1690.9600 1741.2600 1691.4400 ;
        RECT 1694.6600 1778.0000 1696.2600 1778.4800 ;
        RECT 1694.6600 1783.4400 1696.2600 1783.9200 ;
        RECT 1694.6600 1788.8800 1696.2600 1789.3600 ;
        RECT 1694.6600 1767.1200 1696.2600 1767.6000 ;
        RECT 1694.6600 1772.5600 1696.2600 1773.0400 ;
        RECT 1649.6600 1778.0000 1651.2600 1778.4800 ;
        RECT 1649.6600 1783.4400 1651.2600 1783.9200 ;
        RECT 1649.6600 1788.8800 1651.2600 1789.3600 ;
        RECT 1649.6600 1767.1200 1651.2600 1767.6000 ;
        RECT 1649.6600 1772.5600 1651.2600 1773.0400 ;
        RECT 1694.6600 1750.8000 1696.2600 1751.2800 ;
        RECT 1694.6600 1756.2400 1696.2600 1756.7200 ;
        RECT 1694.6600 1761.6800 1696.2600 1762.1600 ;
        RECT 1694.6600 1739.9200 1696.2600 1740.4000 ;
        RECT 1694.6600 1745.3600 1696.2600 1745.8400 ;
        RECT 1649.6600 1750.8000 1651.2600 1751.2800 ;
        RECT 1649.6600 1756.2400 1651.2600 1756.7200 ;
        RECT 1649.6600 1761.6800 1651.2600 1762.1600 ;
        RECT 1649.6600 1739.9200 1651.2600 1740.4000 ;
        RECT 1649.6600 1745.3600 1651.2600 1745.8400 ;
        RECT 1604.6600 1778.0000 1606.2600 1778.4800 ;
        RECT 1604.6600 1783.4400 1606.2600 1783.9200 ;
        RECT 1604.6600 1788.8800 1606.2600 1789.3600 ;
        RECT 1592.9000 1778.0000 1595.9000 1778.4800 ;
        RECT 1592.9000 1783.4400 1595.9000 1783.9200 ;
        RECT 1592.9000 1788.8800 1595.9000 1789.3600 ;
        RECT 1604.6600 1767.1200 1606.2600 1767.6000 ;
        RECT 1604.6600 1772.5600 1606.2600 1773.0400 ;
        RECT 1592.9000 1767.1200 1595.9000 1767.6000 ;
        RECT 1592.9000 1772.5600 1595.9000 1773.0400 ;
        RECT 1604.6600 1750.8000 1606.2600 1751.2800 ;
        RECT 1604.6600 1756.2400 1606.2600 1756.7200 ;
        RECT 1604.6600 1761.6800 1606.2600 1762.1600 ;
        RECT 1592.9000 1750.8000 1595.9000 1751.2800 ;
        RECT 1592.9000 1756.2400 1595.9000 1756.7200 ;
        RECT 1592.9000 1761.6800 1595.9000 1762.1600 ;
        RECT 1604.6600 1739.9200 1606.2600 1740.4000 ;
        RECT 1604.6600 1745.3600 1606.2600 1745.8400 ;
        RECT 1592.9000 1739.9200 1595.9000 1740.4000 ;
        RECT 1592.9000 1745.3600 1595.9000 1745.8400 ;
        RECT 1694.6600 1723.6000 1696.2600 1724.0800 ;
        RECT 1694.6600 1729.0400 1696.2600 1729.5200 ;
        RECT 1694.6600 1734.4800 1696.2600 1734.9600 ;
        RECT 1694.6600 1712.7200 1696.2600 1713.2000 ;
        RECT 1694.6600 1718.1600 1696.2600 1718.6400 ;
        RECT 1649.6600 1723.6000 1651.2600 1724.0800 ;
        RECT 1649.6600 1729.0400 1651.2600 1729.5200 ;
        RECT 1649.6600 1734.4800 1651.2600 1734.9600 ;
        RECT 1649.6600 1712.7200 1651.2600 1713.2000 ;
        RECT 1649.6600 1718.1600 1651.2600 1718.6400 ;
        RECT 1694.6600 1696.4000 1696.2600 1696.8800 ;
        RECT 1694.6600 1701.8400 1696.2600 1702.3200 ;
        RECT 1694.6600 1707.2800 1696.2600 1707.7600 ;
        RECT 1694.6600 1690.9600 1696.2600 1691.4400 ;
        RECT 1649.6600 1696.4000 1651.2600 1696.8800 ;
        RECT 1649.6600 1701.8400 1651.2600 1702.3200 ;
        RECT 1649.6600 1707.2800 1651.2600 1707.7600 ;
        RECT 1649.6600 1690.9600 1651.2600 1691.4400 ;
        RECT 1604.6600 1723.6000 1606.2600 1724.0800 ;
        RECT 1604.6600 1729.0400 1606.2600 1729.5200 ;
        RECT 1604.6600 1734.4800 1606.2600 1734.9600 ;
        RECT 1592.9000 1723.6000 1595.9000 1724.0800 ;
        RECT 1592.9000 1729.0400 1595.9000 1729.5200 ;
        RECT 1592.9000 1734.4800 1595.9000 1734.9600 ;
        RECT 1604.6600 1712.7200 1606.2600 1713.2000 ;
        RECT 1604.6600 1718.1600 1606.2600 1718.6400 ;
        RECT 1592.9000 1712.7200 1595.9000 1713.2000 ;
        RECT 1592.9000 1718.1600 1595.9000 1718.6400 ;
        RECT 1604.6600 1696.4000 1606.2600 1696.8800 ;
        RECT 1604.6600 1701.8400 1606.2600 1702.3200 ;
        RECT 1604.6600 1707.2800 1606.2600 1707.7600 ;
        RECT 1592.9000 1696.4000 1595.9000 1696.8800 ;
        RECT 1592.9000 1701.8400 1595.9000 1702.3200 ;
        RECT 1592.9000 1707.2800 1595.9000 1707.7600 ;
        RECT 1592.9000 1690.9600 1595.9000 1691.4400 ;
        RECT 1604.6600 1690.9600 1606.2600 1691.4400 ;
        RECT 1592.9000 1895.8700 1800.0000 1898.8700 ;
        RECT 1592.9000 1682.7700 1800.0000 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 1453.1300 1786.2600 1669.2300 ;
        RECT 1739.6600 1453.1300 1741.2600 1669.2300 ;
        RECT 1694.6600 1453.1300 1696.2600 1669.2300 ;
        RECT 1649.6600 1453.1300 1651.2600 1669.2300 ;
        RECT 1604.6600 1453.1300 1606.2600 1669.2300 ;
        RECT 1797.0000 1453.1300 1800.0000 1669.2300 ;
        RECT 1592.9000 1453.1300 1595.9000 1669.2300 ;
      LAYER met3 ;
        RECT 1797.0000 1646.2800 1800.0000 1646.7600 ;
        RECT 1797.0000 1651.7200 1800.0000 1652.2000 ;
        RECT 1784.6600 1646.2800 1786.2600 1646.7600 ;
        RECT 1784.6600 1651.7200 1786.2600 1652.2000 ;
        RECT 1797.0000 1657.1600 1800.0000 1657.6400 ;
        RECT 1784.6600 1657.1600 1786.2600 1657.6400 ;
        RECT 1797.0000 1635.4000 1800.0000 1635.8800 ;
        RECT 1797.0000 1640.8400 1800.0000 1641.3200 ;
        RECT 1784.6600 1635.4000 1786.2600 1635.8800 ;
        RECT 1784.6600 1640.8400 1786.2600 1641.3200 ;
        RECT 1797.0000 1619.0800 1800.0000 1619.5600 ;
        RECT 1797.0000 1624.5200 1800.0000 1625.0000 ;
        RECT 1784.6600 1619.0800 1786.2600 1619.5600 ;
        RECT 1784.6600 1624.5200 1786.2600 1625.0000 ;
        RECT 1797.0000 1629.9600 1800.0000 1630.4400 ;
        RECT 1784.6600 1629.9600 1786.2600 1630.4400 ;
        RECT 1739.6600 1646.2800 1741.2600 1646.7600 ;
        RECT 1739.6600 1651.7200 1741.2600 1652.2000 ;
        RECT 1739.6600 1657.1600 1741.2600 1657.6400 ;
        RECT 1739.6600 1635.4000 1741.2600 1635.8800 ;
        RECT 1739.6600 1640.8400 1741.2600 1641.3200 ;
        RECT 1739.6600 1619.0800 1741.2600 1619.5600 ;
        RECT 1739.6600 1624.5200 1741.2600 1625.0000 ;
        RECT 1739.6600 1629.9600 1741.2600 1630.4400 ;
        RECT 1797.0000 1602.7600 1800.0000 1603.2400 ;
        RECT 1797.0000 1608.2000 1800.0000 1608.6800 ;
        RECT 1797.0000 1613.6400 1800.0000 1614.1200 ;
        RECT 1784.6600 1602.7600 1786.2600 1603.2400 ;
        RECT 1784.6600 1608.2000 1786.2600 1608.6800 ;
        RECT 1784.6600 1613.6400 1786.2600 1614.1200 ;
        RECT 1797.0000 1591.8800 1800.0000 1592.3600 ;
        RECT 1797.0000 1597.3200 1800.0000 1597.8000 ;
        RECT 1784.6600 1591.8800 1786.2600 1592.3600 ;
        RECT 1784.6600 1597.3200 1786.2600 1597.8000 ;
        RECT 1797.0000 1575.5600 1800.0000 1576.0400 ;
        RECT 1797.0000 1581.0000 1800.0000 1581.4800 ;
        RECT 1797.0000 1586.4400 1800.0000 1586.9200 ;
        RECT 1784.6600 1575.5600 1786.2600 1576.0400 ;
        RECT 1784.6600 1581.0000 1786.2600 1581.4800 ;
        RECT 1784.6600 1586.4400 1786.2600 1586.9200 ;
        RECT 1797.0000 1564.6800 1800.0000 1565.1600 ;
        RECT 1797.0000 1570.1200 1800.0000 1570.6000 ;
        RECT 1784.6600 1564.6800 1786.2600 1565.1600 ;
        RECT 1784.6600 1570.1200 1786.2600 1570.6000 ;
        RECT 1739.6600 1602.7600 1741.2600 1603.2400 ;
        RECT 1739.6600 1608.2000 1741.2600 1608.6800 ;
        RECT 1739.6600 1613.6400 1741.2600 1614.1200 ;
        RECT 1739.6600 1591.8800 1741.2600 1592.3600 ;
        RECT 1739.6600 1597.3200 1741.2600 1597.8000 ;
        RECT 1739.6600 1575.5600 1741.2600 1576.0400 ;
        RECT 1739.6600 1581.0000 1741.2600 1581.4800 ;
        RECT 1739.6600 1586.4400 1741.2600 1586.9200 ;
        RECT 1739.6600 1564.6800 1741.2600 1565.1600 ;
        RECT 1739.6600 1570.1200 1741.2600 1570.6000 ;
        RECT 1694.6600 1646.2800 1696.2600 1646.7600 ;
        RECT 1694.6600 1651.7200 1696.2600 1652.2000 ;
        RECT 1694.6600 1657.1600 1696.2600 1657.6400 ;
        RECT 1649.6600 1646.2800 1651.2600 1646.7600 ;
        RECT 1649.6600 1651.7200 1651.2600 1652.2000 ;
        RECT 1649.6600 1657.1600 1651.2600 1657.6400 ;
        RECT 1694.6600 1635.4000 1696.2600 1635.8800 ;
        RECT 1694.6600 1640.8400 1696.2600 1641.3200 ;
        RECT 1694.6600 1619.0800 1696.2600 1619.5600 ;
        RECT 1694.6600 1624.5200 1696.2600 1625.0000 ;
        RECT 1694.6600 1629.9600 1696.2600 1630.4400 ;
        RECT 1649.6600 1635.4000 1651.2600 1635.8800 ;
        RECT 1649.6600 1640.8400 1651.2600 1641.3200 ;
        RECT 1649.6600 1619.0800 1651.2600 1619.5600 ;
        RECT 1649.6600 1624.5200 1651.2600 1625.0000 ;
        RECT 1649.6600 1629.9600 1651.2600 1630.4400 ;
        RECT 1604.6600 1646.2800 1606.2600 1646.7600 ;
        RECT 1604.6600 1651.7200 1606.2600 1652.2000 ;
        RECT 1592.9000 1651.7200 1595.9000 1652.2000 ;
        RECT 1592.9000 1646.2800 1595.9000 1646.7600 ;
        RECT 1592.9000 1657.1600 1595.9000 1657.6400 ;
        RECT 1604.6600 1657.1600 1606.2600 1657.6400 ;
        RECT 1604.6600 1635.4000 1606.2600 1635.8800 ;
        RECT 1604.6600 1640.8400 1606.2600 1641.3200 ;
        RECT 1592.9000 1640.8400 1595.9000 1641.3200 ;
        RECT 1592.9000 1635.4000 1595.9000 1635.8800 ;
        RECT 1604.6600 1619.0800 1606.2600 1619.5600 ;
        RECT 1604.6600 1624.5200 1606.2600 1625.0000 ;
        RECT 1592.9000 1624.5200 1595.9000 1625.0000 ;
        RECT 1592.9000 1619.0800 1595.9000 1619.5600 ;
        RECT 1592.9000 1629.9600 1595.9000 1630.4400 ;
        RECT 1604.6600 1629.9600 1606.2600 1630.4400 ;
        RECT 1694.6600 1602.7600 1696.2600 1603.2400 ;
        RECT 1694.6600 1608.2000 1696.2600 1608.6800 ;
        RECT 1694.6600 1613.6400 1696.2600 1614.1200 ;
        RECT 1694.6600 1591.8800 1696.2600 1592.3600 ;
        RECT 1694.6600 1597.3200 1696.2600 1597.8000 ;
        RECT 1649.6600 1602.7600 1651.2600 1603.2400 ;
        RECT 1649.6600 1608.2000 1651.2600 1608.6800 ;
        RECT 1649.6600 1613.6400 1651.2600 1614.1200 ;
        RECT 1649.6600 1591.8800 1651.2600 1592.3600 ;
        RECT 1649.6600 1597.3200 1651.2600 1597.8000 ;
        RECT 1694.6600 1575.5600 1696.2600 1576.0400 ;
        RECT 1694.6600 1581.0000 1696.2600 1581.4800 ;
        RECT 1694.6600 1586.4400 1696.2600 1586.9200 ;
        RECT 1694.6600 1564.6800 1696.2600 1565.1600 ;
        RECT 1694.6600 1570.1200 1696.2600 1570.6000 ;
        RECT 1649.6600 1575.5600 1651.2600 1576.0400 ;
        RECT 1649.6600 1581.0000 1651.2600 1581.4800 ;
        RECT 1649.6600 1586.4400 1651.2600 1586.9200 ;
        RECT 1649.6600 1564.6800 1651.2600 1565.1600 ;
        RECT 1649.6600 1570.1200 1651.2600 1570.6000 ;
        RECT 1604.6600 1602.7600 1606.2600 1603.2400 ;
        RECT 1604.6600 1608.2000 1606.2600 1608.6800 ;
        RECT 1604.6600 1613.6400 1606.2600 1614.1200 ;
        RECT 1592.9000 1602.7600 1595.9000 1603.2400 ;
        RECT 1592.9000 1608.2000 1595.9000 1608.6800 ;
        RECT 1592.9000 1613.6400 1595.9000 1614.1200 ;
        RECT 1604.6600 1591.8800 1606.2600 1592.3600 ;
        RECT 1604.6600 1597.3200 1606.2600 1597.8000 ;
        RECT 1592.9000 1591.8800 1595.9000 1592.3600 ;
        RECT 1592.9000 1597.3200 1595.9000 1597.8000 ;
        RECT 1604.6600 1575.5600 1606.2600 1576.0400 ;
        RECT 1604.6600 1581.0000 1606.2600 1581.4800 ;
        RECT 1604.6600 1586.4400 1606.2600 1586.9200 ;
        RECT 1592.9000 1575.5600 1595.9000 1576.0400 ;
        RECT 1592.9000 1581.0000 1595.9000 1581.4800 ;
        RECT 1592.9000 1586.4400 1595.9000 1586.9200 ;
        RECT 1604.6600 1564.6800 1606.2600 1565.1600 ;
        RECT 1604.6600 1570.1200 1606.2600 1570.6000 ;
        RECT 1592.9000 1564.6800 1595.9000 1565.1600 ;
        RECT 1592.9000 1570.1200 1595.9000 1570.6000 ;
        RECT 1797.0000 1548.3600 1800.0000 1548.8400 ;
        RECT 1797.0000 1553.8000 1800.0000 1554.2800 ;
        RECT 1797.0000 1559.2400 1800.0000 1559.7200 ;
        RECT 1784.6600 1548.3600 1786.2600 1548.8400 ;
        RECT 1784.6600 1553.8000 1786.2600 1554.2800 ;
        RECT 1784.6600 1559.2400 1786.2600 1559.7200 ;
        RECT 1797.0000 1537.4800 1800.0000 1537.9600 ;
        RECT 1797.0000 1542.9200 1800.0000 1543.4000 ;
        RECT 1784.6600 1537.4800 1786.2600 1537.9600 ;
        RECT 1784.6600 1542.9200 1786.2600 1543.4000 ;
        RECT 1797.0000 1521.1600 1800.0000 1521.6400 ;
        RECT 1797.0000 1526.6000 1800.0000 1527.0800 ;
        RECT 1797.0000 1532.0400 1800.0000 1532.5200 ;
        RECT 1784.6600 1521.1600 1786.2600 1521.6400 ;
        RECT 1784.6600 1526.6000 1786.2600 1527.0800 ;
        RECT 1784.6600 1532.0400 1786.2600 1532.5200 ;
        RECT 1797.0000 1510.2800 1800.0000 1510.7600 ;
        RECT 1797.0000 1515.7200 1800.0000 1516.2000 ;
        RECT 1784.6600 1510.2800 1786.2600 1510.7600 ;
        RECT 1784.6600 1515.7200 1786.2600 1516.2000 ;
        RECT 1739.6600 1548.3600 1741.2600 1548.8400 ;
        RECT 1739.6600 1553.8000 1741.2600 1554.2800 ;
        RECT 1739.6600 1559.2400 1741.2600 1559.7200 ;
        RECT 1739.6600 1537.4800 1741.2600 1537.9600 ;
        RECT 1739.6600 1542.9200 1741.2600 1543.4000 ;
        RECT 1739.6600 1521.1600 1741.2600 1521.6400 ;
        RECT 1739.6600 1526.6000 1741.2600 1527.0800 ;
        RECT 1739.6600 1532.0400 1741.2600 1532.5200 ;
        RECT 1739.6600 1510.2800 1741.2600 1510.7600 ;
        RECT 1739.6600 1515.7200 1741.2600 1516.2000 ;
        RECT 1797.0000 1493.9600 1800.0000 1494.4400 ;
        RECT 1797.0000 1499.4000 1800.0000 1499.8800 ;
        RECT 1797.0000 1504.8400 1800.0000 1505.3200 ;
        RECT 1784.6600 1493.9600 1786.2600 1494.4400 ;
        RECT 1784.6600 1499.4000 1786.2600 1499.8800 ;
        RECT 1784.6600 1504.8400 1786.2600 1505.3200 ;
        RECT 1797.0000 1483.0800 1800.0000 1483.5600 ;
        RECT 1797.0000 1488.5200 1800.0000 1489.0000 ;
        RECT 1784.6600 1483.0800 1786.2600 1483.5600 ;
        RECT 1784.6600 1488.5200 1786.2600 1489.0000 ;
        RECT 1797.0000 1466.7600 1800.0000 1467.2400 ;
        RECT 1797.0000 1472.2000 1800.0000 1472.6800 ;
        RECT 1797.0000 1477.6400 1800.0000 1478.1200 ;
        RECT 1784.6600 1466.7600 1786.2600 1467.2400 ;
        RECT 1784.6600 1472.2000 1786.2600 1472.6800 ;
        RECT 1784.6600 1477.6400 1786.2600 1478.1200 ;
        RECT 1797.0000 1461.3200 1800.0000 1461.8000 ;
        RECT 1784.6600 1461.3200 1786.2600 1461.8000 ;
        RECT 1739.6600 1493.9600 1741.2600 1494.4400 ;
        RECT 1739.6600 1499.4000 1741.2600 1499.8800 ;
        RECT 1739.6600 1504.8400 1741.2600 1505.3200 ;
        RECT 1739.6600 1483.0800 1741.2600 1483.5600 ;
        RECT 1739.6600 1488.5200 1741.2600 1489.0000 ;
        RECT 1739.6600 1466.7600 1741.2600 1467.2400 ;
        RECT 1739.6600 1472.2000 1741.2600 1472.6800 ;
        RECT 1739.6600 1477.6400 1741.2600 1478.1200 ;
        RECT 1739.6600 1461.3200 1741.2600 1461.8000 ;
        RECT 1694.6600 1548.3600 1696.2600 1548.8400 ;
        RECT 1694.6600 1553.8000 1696.2600 1554.2800 ;
        RECT 1694.6600 1559.2400 1696.2600 1559.7200 ;
        RECT 1694.6600 1537.4800 1696.2600 1537.9600 ;
        RECT 1694.6600 1542.9200 1696.2600 1543.4000 ;
        RECT 1649.6600 1548.3600 1651.2600 1548.8400 ;
        RECT 1649.6600 1553.8000 1651.2600 1554.2800 ;
        RECT 1649.6600 1559.2400 1651.2600 1559.7200 ;
        RECT 1649.6600 1537.4800 1651.2600 1537.9600 ;
        RECT 1649.6600 1542.9200 1651.2600 1543.4000 ;
        RECT 1694.6600 1521.1600 1696.2600 1521.6400 ;
        RECT 1694.6600 1526.6000 1696.2600 1527.0800 ;
        RECT 1694.6600 1532.0400 1696.2600 1532.5200 ;
        RECT 1694.6600 1510.2800 1696.2600 1510.7600 ;
        RECT 1694.6600 1515.7200 1696.2600 1516.2000 ;
        RECT 1649.6600 1521.1600 1651.2600 1521.6400 ;
        RECT 1649.6600 1526.6000 1651.2600 1527.0800 ;
        RECT 1649.6600 1532.0400 1651.2600 1532.5200 ;
        RECT 1649.6600 1510.2800 1651.2600 1510.7600 ;
        RECT 1649.6600 1515.7200 1651.2600 1516.2000 ;
        RECT 1604.6600 1548.3600 1606.2600 1548.8400 ;
        RECT 1604.6600 1553.8000 1606.2600 1554.2800 ;
        RECT 1604.6600 1559.2400 1606.2600 1559.7200 ;
        RECT 1592.9000 1548.3600 1595.9000 1548.8400 ;
        RECT 1592.9000 1553.8000 1595.9000 1554.2800 ;
        RECT 1592.9000 1559.2400 1595.9000 1559.7200 ;
        RECT 1604.6600 1537.4800 1606.2600 1537.9600 ;
        RECT 1604.6600 1542.9200 1606.2600 1543.4000 ;
        RECT 1592.9000 1537.4800 1595.9000 1537.9600 ;
        RECT 1592.9000 1542.9200 1595.9000 1543.4000 ;
        RECT 1604.6600 1521.1600 1606.2600 1521.6400 ;
        RECT 1604.6600 1526.6000 1606.2600 1527.0800 ;
        RECT 1604.6600 1532.0400 1606.2600 1532.5200 ;
        RECT 1592.9000 1521.1600 1595.9000 1521.6400 ;
        RECT 1592.9000 1526.6000 1595.9000 1527.0800 ;
        RECT 1592.9000 1532.0400 1595.9000 1532.5200 ;
        RECT 1604.6600 1510.2800 1606.2600 1510.7600 ;
        RECT 1604.6600 1515.7200 1606.2600 1516.2000 ;
        RECT 1592.9000 1510.2800 1595.9000 1510.7600 ;
        RECT 1592.9000 1515.7200 1595.9000 1516.2000 ;
        RECT 1694.6600 1493.9600 1696.2600 1494.4400 ;
        RECT 1694.6600 1499.4000 1696.2600 1499.8800 ;
        RECT 1694.6600 1504.8400 1696.2600 1505.3200 ;
        RECT 1694.6600 1483.0800 1696.2600 1483.5600 ;
        RECT 1694.6600 1488.5200 1696.2600 1489.0000 ;
        RECT 1649.6600 1493.9600 1651.2600 1494.4400 ;
        RECT 1649.6600 1499.4000 1651.2600 1499.8800 ;
        RECT 1649.6600 1504.8400 1651.2600 1505.3200 ;
        RECT 1649.6600 1483.0800 1651.2600 1483.5600 ;
        RECT 1649.6600 1488.5200 1651.2600 1489.0000 ;
        RECT 1694.6600 1466.7600 1696.2600 1467.2400 ;
        RECT 1694.6600 1472.2000 1696.2600 1472.6800 ;
        RECT 1694.6600 1477.6400 1696.2600 1478.1200 ;
        RECT 1694.6600 1461.3200 1696.2600 1461.8000 ;
        RECT 1649.6600 1466.7600 1651.2600 1467.2400 ;
        RECT 1649.6600 1472.2000 1651.2600 1472.6800 ;
        RECT 1649.6600 1477.6400 1651.2600 1478.1200 ;
        RECT 1649.6600 1461.3200 1651.2600 1461.8000 ;
        RECT 1604.6600 1493.9600 1606.2600 1494.4400 ;
        RECT 1604.6600 1499.4000 1606.2600 1499.8800 ;
        RECT 1604.6600 1504.8400 1606.2600 1505.3200 ;
        RECT 1592.9000 1493.9600 1595.9000 1494.4400 ;
        RECT 1592.9000 1499.4000 1595.9000 1499.8800 ;
        RECT 1592.9000 1504.8400 1595.9000 1505.3200 ;
        RECT 1604.6600 1483.0800 1606.2600 1483.5600 ;
        RECT 1604.6600 1488.5200 1606.2600 1489.0000 ;
        RECT 1592.9000 1483.0800 1595.9000 1483.5600 ;
        RECT 1592.9000 1488.5200 1595.9000 1489.0000 ;
        RECT 1604.6600 1466.7600 1606.2600 1467.2400 ;
        RECT 1604.6600 1472.2000 1606.2600 1472.6800 ;
        RECT 1604.6600 1477.6400 1606.2600 1478.1200 ;
        RECT 1592.9000 1466.7600 1595.9000 1467.2400 ;
        RECT 1592.9000 1472.2000 1595.9000 1472.6800 ;
        RECT 1592.9000 1477.6400 1595.9000 1478.1200 ;
        RECT 1592.9000 1461.3200 1595.9000 1461.8000 ;
        RECT 1604.6600 1461.3200 1606.2600 1461.8000 ;
        RECT 1592.9000 1666.2300 1800.0000 1669.2300 ;
        RECT 1592.9000 1453.1300 1800.0000 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 1223.4900 1786.2600 1439.5900 ;
        RECT 1739.6600 1223.4900 1741.2600 1439.5900 ;
        RECT 1694.6600 1223.4900 1696.2600 1439.5900 ;
        RECT 1649.6600 1223.4900 1651.2600 1439.5900 ;
        RECT 1604.6600 1223.4900 1606.2600 1439.5900 ;
        RECT 1797.0000 1223.4900 1800.0000 1439.5900 ;
        RECT 1592.9000 1223.4900 1595.9000 1439.5900 ;
      LAYER met3 ;
        RECT 1797.0000 1416.6400 1800.0000 1417.1200 ;
        RECT 1797.0000 1422.0800 1800.0000 1422.5600 ;
        RECT 1784.6600 1416.6400 1786.2600 1417.1200 ;
        RECT 1784.6600 1422.0800 1786.2600 1422.5600 ;
        RECT 1797.0000 1427.5200 1800.0000 1428.0000 ;
        RECT 1784.6600 1427.5200 1786.2600 1428.0000 ;
        RECT 1797.0000 1405.7600 1800.0000 1406.2400 ;
        RECT 1797.0000 1411.2000 1800.0000 1411.6800 ;
        RECT 1784.6600 1405.7600 1786.2600 1406.2400 ;
        RECT 1784.6600 1411.2000 1786.2600 1411.6800 ;
        RECT 1797.0000 1389.4400 1800.0000 1389.9200 ;
        RECT 1797.0000 1394.8800 1800.0000 1395.3600 ;
        RECT 1784.6600 1389.4400 1786.2600 1389.9200 ;
        RECT 1784.6600 1394.8800 1786.2600 1395.3600 ;
        RECT 1797.0000 1400.3200 1800.0000 1400.8000 ;
        RECT 1784.6600 1400.3200 1786.2600 1400.8000 ;
        RECT 1739.6600 1416.6400 1741.2600 1417.1200 ;
        RECT 1739.6600 1422.0800 1741.2600 1422.5600 ;
        RECT 1739.6600 1427.5200 1741.2600 1428.0000 ;
        RECT 1739.6600 1405.7600 1741.2600 1406.2400 ;
        RECT 1739.6600 1411.2000 1741.2600 1411.6800 ;
        RECT 1739.6600 1389.4400 1741.2600 1389.9200 ;
        RECT 1739.6600 1394.8800 1741.2600 1395.3600 ;
        RECT 1739.6600 1400.3200 1741.2600 1400.8000 ;
        RECT 1797.0000 1373.1200 1800.0000 1373.6000 ;
        RECT 1797.0000 1378.5600 1800.0000 1379.0400 ;
        RECT 1797.0000 1384.0000 1800.0000 1384.4800 ;
        RECT 1784.6600 1373.1200 1786.2600 1373.6000 ;
        RECT 1784.6600 1378.5600 1786.2600 1379.0400 ;
        RECT 1784.6600 1384.0000 1786.2600 1384.4800 ;
        RECT 1797.0000 1362.2400 1800.0000 1362.7200 ;
        RECT 1797.0000 1367.6800 1800.0000 1368.1600 ;
        RECT 1784.6600 1362.2400 1786.2600 1362.7200 ;
        RECT 1784.6600 1367.6800 1786.2600 1368.1600 ;
        RECT 1797.0000 1345.9200 1800.0000 1346.4000 ;
        RECT 1797.0000 1351.3600 1800.0000 1351.8400 ;
        RECT 1797.0000 1356.8000 1800.0000 1357.2800 ;
        RECT 1784.6600 1345.9200 1786.2600 1346.4000 ;
        RECT 1784.6600 1351.3600 1786.2600 1351.8400 ;
        RECT 1784.6600 1356.8000 1786.2600 1357.2800 ;
        RECT 1797.0000 1335.0400 1800.0000 1335.5200 ;
        RECT 1797.0000 1340.4800 1800.0000 1340.9600 ;
        RECT 1784.6600 1335.0400 1786.2600 1335.5200 ;
        RECT 1784.6600 1340.4800 1786.2600 1340.9600 ;
        RECT 1739.6600 1373.1200 1741.2600 1373.6000 ;
        RECT 1739.6600 1378.5600 1741.2600 1379.0400 ;
        RECT 1739.6600 1384.0000 1741.2600 1384.4800 ;
        RECT 1739.6600 1362.2400 1741.2600 1362.7200 ;
        RECT 1739.6600 1367.6800 1741.2600 1368.1600 ;
        RECT 1739.6600 1345.9200 1741.2600 1346.4000 ;
        RECT 1739.6600 1351.3600 1741.2600 1351.8400 ;
        RECT 1739.6600 1356.8000 1741.2600 1357.2800 ;
        RECT 1739.6600 1335.0400 1741.2600 1335.5200 ;
        RECT 1739.6600 1340.4800 1741.2600 1340.9600 ;
        RECT 1694.6600 1416.6400 1696.2600 1417.1200 ;
        RECT 1694.6600 1422.0800 1696.2600 1422.5600 ;
        RECT 1694.6600 1427.5200 1696.2600 1428.0000 ;
        RECT 1649.6600 1416.6400 1651.2600 1417.1200 ;
        RECT 1649.6600 1422.0800 1651.2600 1422.5600 ;
        RECT 1649.6600 1427.5200 1651.2600 1428.0000 ;
        RECT 1694.6600 1405.7600 1696.2600 1406.2400 ;
        RECT 1694.6600 1411.2000 1696.2600 1411.6800 ;
        RECT 1694.6600 1389.4400 1696.2600 1389.9200 ;
        RECT 1694.6600 1394.8800 1696.2600 1395.3600 ;
        RECT 1694.6600 1400.3200 1696.2600 1400.8000 ;
        RECT 1649.6600 1405.7600 1651.2600 1406.2400 ;
        RECT 1649.6600 1411.2000 1651.2600 1411.6800 ;
        RECT 1649.6600 1389.4400 1651.2600 1389.9200 ;
        RECT 1649.6600 1394.8800 1651.2600 1395.3600 ;
        RECT 1649.6600 1400.3200 1651.2600 1400.8000 ;
        RECT 1604.6600 1416.6400 1606.2600 1417.1200 ;
        RECT 1604.6600 1422.0800 1606.2600 1422.5600 ;
        RECT 1592.9000 1422.0800 1595.9000 1422.5600 ;
        RECT 1592.9000 1416.6400 1595.9000 1417.1200 ;
        RECT 1592.9000 1427.5200 1595.9000 1428.0000 ;
        RECT 1604.6600 1427.5200 1606.2600 1428.0000 ;
        RECT 1604.6600 1405.7600 1606.2600 1406.2400 ;
        RECT 1604.6600 1411.2000 1606.2600 1411.6800 ;
        RECT 1592.9000 1411.2000 1595.9000 1411.6800 ;
        RECT 1592.9000 1405.7600 1595.9000 1406.2400 ;
        RECT 1604.6600 1389.4400 1606.2600 1389.9200 ;
        RECT 1604.6600 1394.8800 1606.2600 1395.3600 ;
        RECT 1592.9000 1394.8800 1595.9000 1395.3600 ;
        RECT 1592.9000 1389.4400 1595.9000 1389.9200 ;
        RECT 1592.9000 1400.3200 1595.9000 1400.8000 ;
        RECT 1604.6600 1400.3200 1606.2600 1400.8000 ;
        RECT 1694.6600 1373.1200 1696.2600 1373.6000 ;
        RECT 1694.6600 1378.5600 1696.2600 1379.0400 ;
        RECT 1694.6600 1384.0000 1696.2600 1384.4800 ;
        RECT 1694.6600 1362.2400 1696.2600 1362.7200 ;
        RECT 1694.6600 1367.6800 1696.2600 1368.1600 ;
        RECT 1649.6600 1373.1200 1651.2600 1373.6000 ;
        RECT 1649.6600 1378.5600 1651.2600 1379.0400 ;
        RECT 1649.6600 1384.0000 1651.2600 1384.4800 ;
        RECT 1649.6600 1362.2400 1651.2600 1362.7200 ;
        RECT 1649.6600 1367.6800 1651.2600 1368.1600 ;
        RECT 1694.6600 1345.9200 1696.2600 1346.4000 ;
        RECT 1694.6600 1351.3600 1696.2600 1351.8400 ;
        RECT 1694.6600 1356.8000 1696.2600 1357.2800 ;
        RECT 1694.6600 1335.0400 1696.2600 1335.5200 ;
        RECT 1694.6600 1340.4800 1696.2600 1340.9600 ;
        RECT 1649.6600 1345.9200 1651.2600 1346.4000 ;
        RECT 1649.6600 1351.3600 1651.2600 1351.8400 ;
        RECT 1649.6600 1356.8000 1651.2600 1357.2800 ;
        RECT 1649.6600 1335.0400 1651.2600 1335.5200 ;
        RECT 1649.6600 1340.4800 1651.2600 1340.9600 ;
        RECT 1604.6600 1373.1200 1606.2600 1373.6000 ;
        RECT 1604.6600 1378.5600 1606.2600 1379.0400 ;
        RECT 1604.6600 1384.0000 1606.2600 1384.4800 ;
        RECT 1592.9000 1373.1200 1595.9000 1373.6000 ;
        RECT 1592.9000 1378.5600 1595.9000 1379.0400 ;
        RECT 1592.9000 1384.0000 1595.9000 1384.4800 ;
        RECT 1604.6600 1362.2400 1606.2600 1362.7200 ;
        RECT 1604.6600 1367.6800 1606.2600 1368.1600 ;
        RECT 1592.9000 1362.2400 1595.9000 1362.7200 ;
        RECT 1592.9000 1367.6800 1595.9000 1368.1600 ;
        RECT 1604.6600 1345.9200 1606.2600 1346.4000 ;
        RECT 1604.6600 1351.3600 1606.2600 1351.8400 ;
        RECT 1604.6600 1356.8000 1606.2600 1357.2800 ;
        RECT 1592.9000 1345.9200 1595.9000 1346.4000 ;
        RECT 1592.9000 1351.3600 1595.9000 1351.8400 ;
        RECT 1592.9000 1356.8000 1595.9000 1357.2800 ;
        RECT 1604.6600 1335.0400 1606.2600 1335.5200 ;
        RECT 1604.6600 1340.4800 1606.2600 1340.9600 ;
        RECT 1592.9000 1335.0400 1595.9000 1335.5200 ;
        RECT 1592.9000 1340.4800 1595.9000 1340.9600 ;
        RECT 1797.0000 1318.7200 1800.0000 1319.2000 ;
        RECT 1797.0000 1324.1600 1800.0000 1324.6400 ;
        RECT 1797.0000 1329.6000 1800.0000 1330.0800 ;
        RECT 1784.6600 1318.7200 1786.2600 1319.2000 ;
        RECT 1784.6600 1324.1600 1786.2600 1324.6400 ;
        RECT 1784.6600 1329.6000 1786.2600 1330.0800 ;
        RECT 1797.0000 1307.8400 1800.0000 1308.3200 ;
        RECT 1797.0000 1313.2800 1800.0000 1313.7600 ;
        RECT 1784.6600 1307.8400 1786.2600 1308.3200 ;
        RECT 1784.6600 1313.2800 1786.2600 1313.7600 ;
        RECT 1797.0000 1291.5200 1800.0000 1292.0000 ;
        RECT 1797.0000 1296.9600 1800.0000 1297.4400 ;
        RECT 1797.0000 1302.4000 1800.0000 1302.8800 ;
        RECT 1784.6600 1291.5200 1786.2600 1292.0000 ;
        RECT 1784.6600 1296.9600 1786.2600 1297.4400 ;
        RECT 1784.6600 1302.4000 1786.2600 1302.8800 ;
        RECT 1797.0000 1280.6400 1800.0000 1281.1200 ;
        RECT 1797.0000 1286.0800 1800.0000 1286.5600 ;
        RECT 1784.6600 1280.6400 1786.2600 1281.1200 ;
        RECT 1784.6600 1286.0800 1786.2600 1286.5600 ;
        RECT 1739.6600 1318.7200 1741.2600 1319.2000 ;
        RECT 1739.6600 1324.1600 1741.2600 1324.6400 ;
        RECT 1739.6600 1329.6000 1741.2600 1330.0800 ;
        RECT 1739.6600 1307.8400 1741.2600 1308.3200 ;
        RECT 1739.6600 1313.2800 1741.2600 1313.7600 ;
        RECT 1739.6600 1291.5200 1741.2600 1292.0000 ;
        RECT 1739.6600 1296.9600 1741.2600 1297.4400 ;
        RECT 1739.6600 1302.4000 1741.2600 1302.8800 ;
        RECT 1739.6600 1280.6400 1741.2600 1281.1200 ;
        RECT 1739.6600 1286.0800 1741.2600 1286.5600 ;
        RECT 1797.0000 1264.3200 1800.0000 1264.8000 ;
        RECT 1797.0000 1269.7600 1800.0000 1270.2400 ;
        RECT 1797.0000 1275.2000 1800.0000 1275.6800 ;
        RECT 1784.6600 1264.3200 1786.2600 1264.8000 ;
        RECT 1784.6600 1269.7600 1786.2600 1270.2400 ;
        RECT 1784.6600 1275.2000 1786.2600 1275.6800 ;
        RECT 1797.0000 1253.4400 1800.0000 1253.9200 ;
        RECT 1797.0000 1258.8800 1800.0000 1259.3600 ;
        RECT 1784.6600 1253.4400 1786.2600 1253.9200 ;
        RECT 1784.6600 1258.8800 1786.2600 1259.3600 ;
        RECT 1797.0000 1237.1200 1800.0000 1237.6000 ;
        RECT 1797.0000 1242.5600 1800.0000 1243.0400 ;
        RECT 1797.0000 1248.0000 1800.0000 1248.4800 ;
        RECT 1784.6600 1237.1200 1786.2600 1237.6000 ;
        RECT 1784.6600 1242.5600 1786.2600 1243.0400 ;
        RECT 1784.6600 1248.0000 1786.2600 1248.4800 ;
        RECT 1797.0000 1231.6800 1800.0000 1232.1600 ;
        RECT 1784.6600 1231.6800 1786.2600 1232.1600 ;
        RECT 1739.6600 1264.3200 1741.2600 1264.8000 ;
        RECT 1739.6600 1269.7600 1741.2600 1270.2400 ;
        RECT 1739.6600 1275.2000 1741.2600 1275.6800 ;
        RECT 1739.6600 1253.4400 1741.2600 1253.9200 ;
        RECT 1739.6600 1258.8800 1741.2600 1259.3600 ;
        RECT 1739.6600 1237.1200 1741.2600 1237.6000 ;
        RECT 1739.6600 1242.5600 1741.2600 1243.0400 ;
        RECT 1739.6600 1248.0000 1741.2600 1248.4800 ;
        RECT 1739.6600 1231.6800 1741.2600 1232.1600 ;
        RECT 1694.6600 1318.7200 1696.2600 1319.2000 ;
        RECT 1694.6600 1324.1600 1696.2600 1324.6400 ;
        RECT 1694.6600 1329.6000 1696.2600 1330.0800 ;
        RECT 1694.6600 1307.8400 1696.2600 1308.3200 ;
        RECT 1694.6600 1313.2800 1696.2600 1313.7600 ;
        RECT 1649.6600 1318.7200 1651.2600 1319.2000 ;
        RECT 1649.6600 1324.1600 1651.2600 1324.6400 ;
        RECT 1649.6600 1329.6000 1651.2600 1330.0800 ;
        RECT 1649.6600 1307.8400 1651.2600 1308.3200 ;
        RECT 1649.6600 1313.2800 1651.2600 1313.7600 ;
        RECT 1694.6600 1291.5200 1696.2600 1292.0000 ;
        RECT 1694.6600 1296.9600 1696.2600 1297.4400 ;
        RECT 1694.6600 1302.4000 1696.2600 1302.8800 ;
        RECT 1694.6600 1280.6400 1696.2600 1281.1200 ;
        RECT 1694.6600 1286.0800 1696.2600 1286.5600 ;
        RECT 1649.6600 1291.5200 1651.2600 1292.0000 ;
        RECT 1649.6600 1296.9600 1651.2600 1297.4400 ;
        RECT 1649.6600 1302.4000 1651.2600 1302.8800 ;
        RECT 1649.6600 1280.6400 1651.2600 1281.1200 ;
        RECT 1649.6600 1286.0800 1651.2600 1286.5600 ;
        RECT 1604.6600 1318.7200 1606.2600 1319.2000 ;
        RECT 1604.6600 1324.1600 1606.2600 1324.6400 ;
        RECT 1604.6600 1329.6000 1606.2600 1330.0800 ;
        RECT 1592.9000 1318.7200 1595.9000 1319.2000 ;
        RECT 1592.9000 1324.1600 1595.9000 1324.6400 ;
        RECT 1592.9000 1329.6000 1595.9000 1330.0800 ;
        RECT 1604.6600 1307.8400 1606.2600 1308.3200 ;
        RECT 1604.6600 1313.2800 1606.2600 1313.7600 ;
        RECT 1592.9000 1307.8400 1595.9000 1308.3200 ;
        RECT 1592.9000 1313.2800 1595.9000 1313.7600 ;
        RECT 1604.6600 1291.5200 1606.2600 1292.0000 ;
        RECT 1604.6600 1296.9600 1606.2600 1297.4400 ;
        RECT 1604.6600 1302.4000 1606.2600 1302.8800 ;
        RECT 1592.9000 1291.5200 1595.9000 1292.0000 ;
        RECT 1592.9000 1296.9600 1595.9000 1297.4400 ;
        RECT 1592.9000 1302.4000 1595.9000 1302.8800 ;
        RECT 1604.6600 1280.6400 1606.2600 1281.1200 ;
        RECT 1604.6600 1286.0800 1606.2600 1286.5600 ;
        RECT 1592.9000 1280.6400 1595.9000 1281.1200 ;
        RECT 1592.9000 1286.0800 1595.9000 1286.5600 ;
        RECT 1694.6600 1264.3200 1696.2600 1264.8000 ;
        RECT 1694.6600 1269.7600 1696.2600 1270.2400 ;
        RECT 1694.6600 1275.2000 1696.2600 1275.6800 ;
        RECT 1694.6600 1253.4400 1696.2600 1253.9200 ;
        RECT 1694.6600 1258.8800 1696.2600 1259.3600 ;
        RECT 1649.6600 1264.3200 1651.2600 1264.8000 ;
        RECT 1649.6600 1269.7600 1651.2600 1270.2400 ;
        RECT 1649.6600 1275.2000 1651.2600 1275.6800 ;
        RECT 1649.6600 1253.4400 1651.2600 1253.9200 ;
        RECT 1649.6600 1258.8800 1651.2600 1259.3600 ;
        RECT 1694.6600 1237.1200 1696.2600 1237.6000 ;
        RECT 1694.6600 1242.5600 1696.2600 1243.0400 ;
        RECT 1694.6600 1248.0000 1696.2600 1248.4800 ;
        RECT 1694.6600 1231.6800 1696.2600 1232.1600 ;
        RECT 1649.6600 1237.1200 1651.2600 1237.6000 ;
        RECT 1649.6600 1242.5600 1651.2600 1243.0400 ;
        RECT 1649.6600 1248.0000 1651.2600 1248.4800 ;
        RECT 1649.6600 1231.6800 1651.2600 1232.1600 ;
        RECT 1604.6600 1264.3200 1606.2600 1264.8000 ;
        RECT 1604.6600 1269.7600 1606.2600 1270.2400 ;
        RECT 1604.6600 1275.2000 1606.2600 1275.6800 ;
        RECT 1592.9000 1264.3200 1595.9000 1264.8000 ;
        RECT 1592.9000 1269.7600 1595.9000 1270.2400 ;
        RECT 1592.9000 1275.2000 1595.9000 1275.6800 ;
        RECT 1604.6600 1253.4400 1606.2600 1253.9200 ;
        RECT 1604.6600 1258.8800 1606.2600 1259.3600 ;
        RECT 1592.9000 1253.4400 1595.9000 1253.9200 ;
        RECT 1592.9000 1258.8800 1595.9000 1259.3600 ;
        RECT 1604.6600 1237.1200 1606.2600 1237.6000 ;
        RECT 1604.6600 1242.5600 1606.2600 1243.0400 ;
        RECT 1604.6600 1248.0000 1606.2600 1248.4800 ;
        RECT 1592.9000 1237.1200 1595.9000 1237.6000 ;
        RECT 1592.9000 1242.5600 1595.9000 1243.0400 ;
        RECT 1592.9000 1248.0000 1595.9000 1248.4800 ;
        RECT 1592.9000 1231.6800 1595.9000 1232.1600 ;
        RECT 1604.6600 1231.6800 1606.2600 1232.1600 ;
        RECT 1592.9000 1436.5900 1800.0000 1439.5900 ;
        RECT 1592.9000 1223.4900 1800.0000 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 993.8500 1786.2600 1209.9500 ;
        RECT 1739.6600 993.8500 1741.2600 1209.9500 ;
        RECT 1694.6600 993.8500 1696.2600 1209.9500 ;
        RECT 1649.6600 993.8500 1651.2600 1209.9500 ;
        RECT 1604.6600 993.8500 1606.2600 1209.9500 ;
        RECT 1797.0000 993.8500 1800.0000 1209.9500 ;
        RECT 1592.9000 993.8500 1595.9000 1209.9500 ;
      LAYER met3 ;
        RECT 1797.0000 1187.0000 1800.0000 1187.4800 ;
        RECT 1797.0000 1192.4400 1800.0000 1192.9200 ;
        RECT 1784.6600 1187.0000 1786.2600 1187.4800 ;
        RECT 1784.6600 1192.4400 1786.2600 1192.9200 ;
        RECT 1797.0000 1197.8800 1800.0000 1198.3600 ;
        RECT 1784.6600 1197.8800 1786.2600 1198.3600 ;
        RECT 1797.0000 1176.1200 1800.0000 1176.6000 ;
        RECT 1797.0000 1181.5600 1800.0000 1182.0400 ;
        RECT 1784.6600 1176.1200 1786.2600 1176.6000 ;
        RECT 1784.6600 1181.5600 1786.2600 1182.0400 ;
        RECT 1797.0000 1159.8000 1800.0000 1160.2800 ;
        RECT 1797.0000 1165.2400 1800.0000 1165.7200 ;
        RECT 1784.6600 1159.8000 1786.2600 1160.2800 ;
        RECT 1784.6600 1165.2400 1786.2600 1165.7200 ;
        RECT 1797.0000 1170.6800 1800.0000 1171.1600 ;
        RECT 1784.6600 1170.6800 1786.2600 1171.1600 ;
        RECT 1739.6600 1187.0000 1741.2600 1187.4800 ;
        RECT 1739.6600 1192.4400 1741.2600 1192.9200 ;
        RECT 1739.6600 1197.8800 1741.2600 1198.3600 ;
        RECT 1739.6600 1176.1200 1741.2600 1176.6000 ;
        RECT 1739.6600 1181.5600 1741.2600 1182.0400 ;
        RECT 1739.6600 1159.8000 1741.2600 1160.2800 ;
        RECT 1739.6600 1165.2400 1741.2600 1165.7200 ;
        RECT 1739.6600 1170.6800 1741.2600 1171.1600 ;
        RECT 1797.0000 1143.4800 1800.0000 1143.9600 ;
        RECT 1797.0000 1148.9200 1800.0000 1149.4000 ;
        RECT 1797.0000 1154.3600 1800.0000 1154.8400 ;
        RECT 1784.6600 1143.4800 1786.2600 1143.9600 ;
        RECT 1784.6600 1148.9200 1786.2600 1149.4000 ;
        RECT 1784.6600 1154.3600 1786.2600 1154.8400 ;
        RECT 1797.0000 1132.6000 1800.0000 1133.0800 ;
        RECT 1797.0000 1138.0400 1800.0000 1138.5200 ;
        RECT 1784.6600 1132.6000 1786.2600 1133.0800 ;
        RECT 1784.6600 1138.0400 1786.2600 1138.5200 ;
        RECT 1797.0000 1116.2800 1800.0000 1116.7600 ;
        RECT 1797.0000 1121.7200 1800.0000 1122.2000 ;
        RECT 1797.0000 1127.1600 1800.0000 1127.6400 ;
        RECT 1784.6600 1116.2800 1786.2600 1116.7600 ;
        RECT 1784.6600 1121.7200 1786.2600 1122.2000 ;
        RECT 1784.6600 1127.1600 1786.2600 1127.6400 ;
        RECT 1797.0000 1105.4000 1800.0000 1105.8800 ;
        RECT 1797.0000 1110.8400 1800.0000 1111.3200 ;
        RECT 1784.6600 1105.4000 1786.2600 1105.8800 ;
        RECT 1784.6600 1110.8400 1786.2600 1111.3200 ;
        RECT 1739.6600 1143.4800 1741.2600 1143.9600 ;
        RECT 1739.6600 1148.9200 1741.2600 1149.4000 ;
        RECT 1739.6600 1154.3600 1741.2600 1154.8400 ;
        RECT 1739.6600 1132.6000 1741.2600 1133.0800 ;
        RECT 1739.6600 1138.0400 1741.2600 1138.5200 ;
        RECT 1739.6600 1116.2800 1741.2600 1116.7600 ;
        RECT 1739.6600 1121.7200 1741.2600 1122.2000 ;
        RECT 1739.6600 1127.1600 1741.2600 1127.6400 ;
        RECT 1739.6600 1105.4000 1741.2600 1105.8800 ;
        RECT 1739.6600 1110.8400 1741.2600 1111.3200 ;
        RECT 1694.6600 1187.0000 1696.2600 1187.4800 ;
        RECT 1694.6600 1192.4400 1696.2600 1192.9200 ;
        RECT 1694.6600 1197.8800 1696.2600 1198.3600 ;
        RECT 1649.6600 1187.0000 1651.2600 1187.4800 ;
        RECT 1649.6600 1192.4400 1651.2600 1192.9200 ;
        RECT 1649.6600 1197.8800 1651.2600 1198.3600 ;
        RECT 1694.6600 1176.1200 1696.2600 1176.6000 ;
        RECT 1694.6600 1181.5600 1696.2600 1182.0400 ;
        RECT 1694.6600 1159.8000 1696.2600 1160.2800 ;
        RECT 1694.6600 1165.2400 1696.2600 1165.7200 ;
        RECT 1694.6600 1170.6800 1696.2600 1171.1600 ;
        RECT 1649.6600 1176.1200 1651.2600 1176.6000 ;
        RECT 1649.6600 1181.5600 1651.2600 1182.0400 ;
        RECT 1649.6600 1159.8000 1651.2600 1160.2800 ;
        RECT 1649.6600 1165.2400 1651.2600 1165.7200 ;
        RECT 1649.6600 1170.6800 1651.2600 1171.1600 ;
        RECT 1604.6600 1187.0000 1606.2600 1187.4800 ;
        RECT 1604.6600 1192.4400 1606.2600 1192.9200 ;
        RECT 1592.9000 1192.4400 1595.9000 1192.9200 ;
        RECT 1592.9000 1187.0000 1595.9000 1187.4800 ;
        RECT 1592.9000 1197.8800 1595.9000 1198.3600 ;
        RECT 1604.6600 1197.8800 1606.2600 1198.3600 ;
        RECT 1604.6600 1176.1200 1606.2600 1176.6000 ;
        RECT 1604.6600 1181.5600 1606.2600 1182.0400 ;
        RECT 1592.9000 1181.5600 1595.9000 1182.0400 ;
        RECT 1592.9000 1176.1200 1595.9000 1176.6000 ;
        RECT 1604.6600 1159.8000 1606.2600 1160.2800 ;
        RECT 1604.6600 1165.2400 1606.2600 1165.7200 ;
        RECT 1592.9000 1165.2400 1595.9000 1165.7200 ;
        RECT 1592.9000 1159.8000 1595.9000 1160.2800 ;
        RECT 1592.9000 1170.6800 1595.9000 1171.1600 ;
        RECT 1604.6600 1170.6800 1606.2600 1171.1600 ;
        RECT 1694.6600 1143.4800 1696.2600 1143.9600 ;
        RECT 1694.6600 1148.9200 1696.2600 1149.4000 ;
        RECT 1694.6600 1154.3600 1696.2600 1154.8400 ;
        RECT 1694.6600 1132.6000 1696.2600 1133.0800 ;
        RECT 1694.6600 1138.0400 1696.2600 1138.5200 ;
        RECT 1649.6600 1143.4800 1651.2600 1143.9600 ;
        RECT 1649.6600 1148.9200 1651.2600 1149.4000 ;
        RECT 1649.6600 1154.3600 1651.2600 1154.8400 ;
        RECT 1649.6600 1132.6000 1651.2600 1133.0800 ;
        RECT 1649.6600 1138.0400 1651.2600 1138.5200 ;
        RECT 1694.6600 1116.2800 1696.2600 1116.7600 ;
        RECT 1694.6600 1121.7200 1696.2600 1122.2000 ;
        RECT 1694.6600 1127.1600 1696.2600 1127.6400 ;
        RECT 1694.6600 1105.4000 1696.2600 1105.8800 ;
        RECT 1694.6600 1110.8400 1696.2600 1111.3200 ;
        RECT 1649.6600 1116.2800 1651.2600 1116.7600 ;
        RECT 1649.6600 1121.7200 1651.2600 1122.2000 ;
        RECT 1649.6600 1127.1600 1651.2600 1127.6400 ;
        RECT 1649.6600 1105.4000 1651.2600 1105.8800 ;
        RECT 1649.6600 1110.8400 1651.2600 1111.3200 ;
        RECT 1604.6600 1143.4800 1606.2600 1143.9600 ;
        RECT 1604.6600 1148.9200 1606.2600 1149.4000 ;
        RECT 1604.6600 1154.3600 1606.2600 1154.8400 ;
        RECT 1592.9000 1143.4800 1595.9000 1143.9600 ;
        RECT 1592.9000 1148.9200 1595.9000 1149.4000 ;
        RECT 1592.9000 1154.3600 1595.9000 1154.8400 ;
        RECT 1604.6600 1132.6000 1606.2600 1133.0800 ;
        RECT 1604.6600 1138.0400 1606.2600 1138.5200 ;
        RECT 1592.9000 1132.6000 1595.9000 1133.0800 ;
        RECT 1592.9000 1138.0400 1595.9000 1138.5200 ;
        RECT 1604.6600 1116.2800 1606.2600 1116.7600 ;
        RECT 1604.6600 1121.7200 1606.2600 1122.2000 ;
        RECT 1604.6600 1127.1600 1606.2600 1127.6400 ;
        RECT 1592.9000 1116.2800 1595.9000 1116.7600 ;
        RECT 1592.9000 1121.7200 1595.9000 1122.2000 ;
        RECT 1592.9000 1127.1600 1595.9000 1127.6400 ;
        RECT 1604.6600 1105.4000 1606.2600 1105.8800 ;
        RECT 1604.6600 1110.8400 1606.2600 1111.3200 ;
        RECT 1592.9000 1105.4000 1595.9000 1105.8800 ;
        RECT 1592.9000 1110.8400 1595.9000 1111.3200 ;
        RECT 1797.0000 1089.0800 1800.0000 1089.5600 ;
        RECT 1797.0000 1094.5200 1800.0000 1095.0000 ;
        RECT 1797.0000 1099.9600 1800.0000 1100.4400 ;
        RECT 1784.6600 1089.0800 1786.2600 1089.5600 ;
        RECT 1784.6600 1094.5200 1786.2600 1095.0000 ;
        RECT 1784.6600 1099.9600 1786.2600 1100.4400 ;
        RECT 1797.0000 1078.2000 1800.0000 1078.6800 ;
        RECT 1797.0000 1083.6400 1800.0000 1084.1200 ;
        RECT 1784.6600 1078.2000 1786.2600 1078.6800 ;
        RECT 1784.6600 1083.6400 1786.2600 1084.1200 ;
        RECT 1797.0000 1061.8800 1800.0000 1062.3600 ;
        RECT 1797.0000 1067.3200 1800.0000 1067.8000 ;
        RECT 1797.0000 1072.7600 1800.0000 1073.2400 ;
        RECT 1784.6600 1061.8800 1786.2600 1062.3600 ;
        RECT 1784.6600 1067.3200 1786.2600 1067.8000 ;
        RECT 1784.6600 1072.7600 1786.2600 1073.2400 ;
        RECT 1797.0000 1051.0000 1800.0000 1051.4800 ;
        RECT 1797.0000 1056.4400 1800.0000 1056.9200 ;
        RECT 1784.6600 1051.0000 1786.2600 1051.4800 ;
        RECT 1784.6600 1056.4400 1786.2600 1056.9200 ;
        RECT 1739.6600 1089.0800 1741.2600 1089.5600 ;
        RECT 1739.6600 1094.5200 1741.2600 1095.0000 ;
        RECT 1739.6600 1099.9600 1741.2600 1100.4400 ;
        RECT 1739.6600 1078.2000 1741.2600 1078.6800 ;
        RECT 1739.6600 1083.6400 1741.2600 1084.1200 ;
        RECT 1739.6600 1061.8800 1741.2600 1062.3600 ;
        RECT 1739.6600 1067.3200 1741.2600 1067.8000 ;
        RECT 1739.6600 1072.7600 1741.2600 1073.2400 ;
        RECT 1739.6600 1051.0000 1741.2600 1051.4800 ;
        RECT 1739.6600 1056.4400 1741.2600 1056.9200 ;
        RECT 1797.0000 1034.6800 1800.0000 1035.1600 ;
        RECT 1797.0000 1040.1200 1800.0000 1040.6000 ;
        RECT 1797.0000 1045.5600 1800.0000 1046.0400 ;
        RECT 1784.6600 1034.6800 1786.2600 1035.1600 ;
        RECT 1784.6600 1040.1200 1786.2600 1040.6000 ;
        RECT 1784.6600 1045.5600 1786.2600 1046.0400 ;
        RECT 1797.0000 1023.8000 1800.0000 1024.2800 ;
        RECT 1797.0000 1029.2400 1800.0000 1029.7200 ;
        RECT 1784.6600 1023.8000 1786.2600 1024.2800 ;
        RECT 1784.6600 1029.2400 1786.2600 1029.7200 ;
        RECT 1797.0000 1007.4800 1800.0000 1007.9600 ;
        RECT 1797.0000 1012.9200 1800.0000 1013.4000 ;
        RECT 1797.0000 1018.3600 1800.0000 1018.8400 ;
        RECT 1784.6600 1007.4800 1786.2600 1007.9600 ;
        RECT 1784.6600 1012.9200 1786.2600 1013.4000 ;
        RECT 1784.6600 1018.3600 1786.2600 1018.8400 ;
        RECT 1797.0000 1002.0400 1800.0000 1002.5200 ;
        RECT 1784.6600 1002.0400 1786.2600 1002.5200 ;
        RECT 1739.6600 1034.6800 1741.2600 1035.1600 ;
        RECT 1739.6600 1040.1200 1741.2600 1040.6000 ;
        RECT 1739.6600 1045.5600 1741.2600 1046.0400 ;
        RECT 1739.6600 1023.8000 1741.2600 1024.2800 ;
        RECT 1739.6600 1029.2400 1741.2600 1029.7200 ;
        RECT 1739.6600 1007.4800 1741.2600 1007.9600 ;
        RECT 1739.6600 1012.9200 1741.2600 1013.4000 ;
        RECT 1739.6600 1018.3600 1741.2600 1018.8400 ;
        RECT 1739.6600 1002.0400 1741.2600 1002.5200 ;
        RECT 1694.6600 1089.0800 1696.2600 1089.5600 ;
        RECT 1694.6600 1094.5200 1696.2600 1095.0000 ;
        RECT 1694.6600 1099.9600 1696.2600 1100.4400 ;
        RECT 1694.6600 1078.2000 1696.2600 1078.6800 ;
        RECT 1694.6600 1083.6400 1696.2600 1084.1200 ;
        RECT 1649.6600 1089.0800 1651.2600 1089.5600 ;
        RECT 1649.6600 1094.5200 1651.2600 1095.0000 ;
        RECT 1649.6600 1099.9600 1651.2600 1100.4400 ;
        RECT 1649.6600 1078.2000 1651.2600 1078.6800 ;
        RECT 1649.6600 1083.6400 1651.2600 1084.1200 ;
        RECT 1694.6600 1061.8800 1696.2600 1062.3600 ;
        RECT 1694.6600 1067.3200 1696.2600 1067.8000 ;
        RECT 1694.6600 1072.7600 1696.2600 1073.2400 ;
        RECT 1694.6600 1051.0000 1696.2600 1051.4800 ;
        RECT 1694.6600 1056.4400 1696.2600 1056.9200 ;
        RECT 1649.6600 1061.8800 1651.2600 1062.3600 ;
        RECT 1649.6600 1067.3200 1651.2600 1067.8000 ;
        RECT 1649.6600 1072.7600 1651.2600 1073.2400 ;
        RECT 1649.6600 1051.0000 1651.2600 1051.4800 ;
        RECT 1649.6600 1056.4400 1651.2600 1056.9200 ;
        RECT 1604.6600 1089.0800 1606.2600 1089.5600 ;
        RECT 1604.6600 1094.5200 1606.2600 1095.0000 ;
        RECT 1604.6600 1099.9600 1606.2600 1100.4400 ;
        RECT 1592.9000 1089.0800 1595.9000 1089.5600 ;
        RECT 1592.9000 1094.5200 1595.9000 1095.0000 ;
        RECT 1592.9000 1099.9600 1595.9000 1100.4400 ;
        RECT 1604.6600 1078.2000 1606.2600 1078.6800 ;
        RECT 1604.6600 1083.6400 1606.2600 1084.1200 ;
        RECT 1592.9000 1078.2000 1595.9000 1078.6800 ;
        RECT 1592.9000 1083.6400 1595.9000 1084.1200 ;
        RECT 1604.6600 1061.8800 1606.2600 1062.3600 ;
        RECT 1604.6600 1067.3200 1606.2600 1067.8000 ;
        RECT 1604.6600 1072.7600 1606.2600 1073.2400 ;
        RECT 1592.9000 1061.8800 1595.9000 1062.3600 ;
        RECT 1592.9000 1067.3200 1595.9000 1067.8000 ;
        RECT 1592.9000 1072.7600 1595.9000 1073.2400 ;
        RECT 1604.6600 1051.0000 1606.2600 1051.4800 ;
        RECT 1604.6600 1056.4400 1606.2600 1056.9200 ;
        RECT 1592.9000 1051.0000 1595.9000 1051.4800 ;
        RECT 1592.9000 1056.4400 1595.9000 1056.9200 ;
        RECT 1694.6600 1034.6800 1696.2600 1035.1600 ;
        RECT 1694.6600 1040.1200 1696.2600 1040.6000 ;
        RECT 1694.6600 1045.5600 1696.2600 1046.0400 ;
        RECT 1694.6600 1023.8000 1696.2600 1024.2800 ;
        RECT 1694.6600 1029.2400 1696.2600 1029.7200 ;
        RECT 1649.6600 1034.6800 1651.2600 1035.1600 ;
        RECT 1649.6600 1040.1200 1651.2600 1040.6000 ;
        RECT 1649.6600 1045.5600 1651.2600 1046.0400 ;
        RECT 1649.6600 1023.8000 1651.2600 1024.2800 ;
        RECT 1649.6600 1029.2400 1651.2600 1029.7200 ;
        RECT 1694.6600 1007.4800 1696.2600 1007.9600 ;
        RECT 1694.6600 1012.9200 1696.2600 1013.4000 ;
        RECT 1694.6600 1018.3600 1696.2600 1018.8400 ;
        RECT 1694.6600 1002.0400 1696.2600 1002.5200 ;
        RECT 1649.6600 1007.4800 1651.2600 1007.9600 ;
        RECT 1649.6600 1012.9200 1651.2600 1013.4000 ;
        RECT 1649.6600 1018.3600 1651.2600 1018.8400 ;
        RECT 1649.6600 1002.0400 1651.2600 1002.5200 ;
        RECT 1604.6600 1034.6800 1606.2600 1035.1600 ;
        RECT 1604.6600 1040.1200 1606.2600 1040.6000 ;
        RECT 1604.6600 1045.5600 1606.2600 1046.0400 ;
        RECT 1592.9000 1034.6800 1595.9000 1035.1600 ;
        RECT 1592.9000 1040.1200 1595.9000 1040.6000 ;
        RECT 1592.9000 1045.5600 1595.9000 1046.0400 ;
        RECT 1604.6600 1023.8000 1606.2600 1024.2800 ;
        RECT 1604.6600 1029.2400 1606.2600 1029.7200 ;
        RECT 1592.9000 1023.8000 1595.9000 1024.2800 ;
        RECT 1592.9000 1029.2400 1595.9000 1029.7200 ;
        RECT 1604.6600 1007.4800 1606.2600 1007.9600 ;
        RECT 1604.6600 1012.9200 1606.2600 1013.4000 ;
        RECT 1604.6600 1018.3600 1606.2600 1018.8400 ;
        RECT 1592.9000 1007.4800 1595.9000 1007.9600 ;
        RECT 1592.9000 1012.9200 1595.9000 1013.4000 ;
        RECT 1592.9000 1018.3600 1595.9000 1018.8400 ;
        RECT 1592.9000 1002.0400 1595.9000 1002.5200 ;
        RECT 1604.6600 1002.0400 1606.2600 1002.5200 ;
        RECT 1592.9000 1206.9500 1800.0000 1209.9500 ;
        RECT 1592.9000 993.8500 1800.0000 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1784.6600 764.2100 1786.2600 980.3100 ;
        RECT 1739.6600 764.2100 1741.2600 980.3100 ;
        RECT 1694.6600 764.2100 1696.2600 980.3100 ;
        RECT 1649.6600 764.2100 1651.2600 980.3100 ;
        RECT 1604.6600 764.2100 1606.2600 980.3100 ;
        RECT 1797.0000 764.2100 1800.0000 980.3100 ;
        RECT 1592.9000 764.2100 1595.9000 980.3100 ;
      LAYER met3 ;
        RECT 1797.0000 957.3600 1800.0000 957.8400 ;
        RECT 1797.0000 962.8000 1800.0000 963.2800 ;
        RECT 1784.6600 957.3600 1786.2600 957.8400 ;
        RECT 1784.6600 962.8000 1786.2600 963.2800 ;
        RECT 1797.0000 968.2400 1800.0000 968.7200 ;
        RECT 1784.6600 968.2400 1786.2600 968.7200 ;
        RECT 1797.0000 946.4800 1800.0000 946.9600 ;
        RECT 1797.0000 951.9200 1800.0000 952.4000 ;
        RECT 1784.6600 946.4800 1786.2600 946.9600 ;
        RECT 1784.6600 951.9200 1786.2600 952.4000 ;
        RECT 1797.0000 930.1600 1800.0000 930.6400 ;
        RECT 1797.0000 935.6000 1800.0000 936.0800 ;
        RECT 1784.6600 930.1600 1786.2600 930.6400 ;
        RECT 1784.6600 935.6000 1786.2600 936.0800 ;
        RECT 1797.0000 941.0400 1800.0000 941.5200 ;
        RECT 1784.6600 941.0400 1786.2600 941.5200 ;
        RECT 1739.6600 957.3600 1741.2600 957.8400 ;
        RECT 1739.6600 962.8000 1741.2600 963.2800 ;
        RECT 1739.6600 968.2400 1741.2600 968.7200 ;
        RECT 1739.6600 946.4800 1741.2600 946.9600 ;
        RECT 1739.6600 951.9200 1741.2600 952.4000 ;
        RECT 1739.6600 930.1600 1741.2600 930.6400 ;
        RECT 1739.6600 935.6000 1741.2600 936.0800 ;
        RECT 1739.6600 941.0400 1741.2600 941.5200 ;
        RECT 1797.0000 913.8400 1800.0000 914.3200 ;
        RECT 1797.0000 919.2800 1800.0000 919.7600 ;
        RECT 1797.0000 924.7200 1800.0000 925.2000 ;
        RECT 1784.6600 913.8400 1786.2600 914.3200 ;
        RECT 1784.6600 919.2800 1786.2600 919.7600 ;
        RECT 1784.6600 924.7200 1786.2600 925.2000 ;
        RECT 1797.0000 902.9600 1800.0000 903.4400 ;
        RECT 1797.0000 908.4000 1800.0000 908.8800 ;
        RECT 1784.6600 902.9600 1786.2600 903.4400 ;
        RECT 1784.6600 908.4000 1786.2600 908.8800 ;
        RECT 1797.0000 886.6400 1800.0000 887.1200 ;
        RECT 1797.0000 892.0800 1800.0000 892.5600 ;
        RECT 1797.0000 897.5200 1800.0000 898.0000 ;
        RECT 1784.6600 886.6400 1786.2600 887.1200 ;
        RECT 1784.6600 892.0800 1786.2600 892.5600 ;
        RECT 1784.6600 897.5200 1786.2600 898.0000 ;
        RECT 1797.0000 875.7600 1800.0000 876.2400 ;
        RECT 1797.0000 881.2000 1800.0000 881.6800 ;
        RECT 1784.6600 875.7600 1786.2600 876.2400 ;
        RECT 1784.6600 881.2000 1786.2600 881.6800 ;
        RECT 1739.6600 913.8400 1741.2600 914.3200 ;
        RECT 1739.6600 919.2800 1741.2600 919.7600 ;
        RECT 1739.6600 924.7200 1741.2600 925.2000 ;
        RECT 1739.6600 902.9600 1741.2600 903.4400 ;
        RECT 1739.6600 908.4000 1741.2600 908.8800 ;
        RECT 1739.6600 886.6400 1741.2600 887.1200 ;
        RECT 1739.6600 892.0800 1741.2600 892.5600 ;
        RECT 1739.6600 897.5200 1741.2600 898.0000 ;
        RECT 1739.6600 875.7600 1741.2600 876.2400 ;
        RECT 1739.6600 881.2000 1741.2600 881.6800 ;
        RECT 1694.6600 957.3600 1696.2600 957.8400 ;
        RECT 1694.6600 962.8000 1696.2600 963.2800 ;
        RECT 1694.6600 968.2400 1696.2600 968.7200 ;
        RECT 1649.6600 957.3600 1651.2600 957.8400 ;
        RECT 1649.6600 962.8000 1651.2600 963.2800 ;
        RECT 1649.6600 968.2400 1651.2600 968.7200 ;
        RECT 1694.6600 946.4800 1696.2600 946.9600 ;
        RECT 1694.6600 951.9200 1696.2600 952.4000 ;
        RECT 1694.6600 930.1600 1696.2600 930.6400 ;
        RECT 1694.6600 935.6000 1696.2600 936.0800 ;
        RECT 1694.6600 941.0400 1696.2600 941.5200 ;
        RECT 1649.6600 946.4800 1651.2600 946.9600 ;
        RECT 1649.6600 951.9200 1651.2600 952.4000 ;
        RECT 1649.6600 930.1600 1651.2600 930.6400 ;
        RECT 1649.6600 935.6000 1651.2600 936.0800 ;
        RECT 1649.6600 941.0400 1651.2600 941.5200 ;
        RECT 1604.6600 957.3600 1606.2600 957.8400 ;
        RECT 1604.6600 962.8000 1606.2600 963.2800 ;
        RECT 1592.9000 962.8000 1595.9000 963.2800 ;
        RECT 1592.9000 957.3600 1595.9000 957.8400 ;
        RECT 1592.9000 968.2400 1595.9000 968.7200 ;
        RECT 1604.6600 968.2400 1606.2600 968.7200 ;
        RECT 1604.6600 946.4800 1606.2600 946.9600 ;
        RECT 1604.6600 951.9200 1606.2600 952.4000 ;
        RECT 1592.9000 951.9200 1595.9000 952.4000 ;
        RECT 1592.9000 946.4800 1595.9000 946.9600 ;
        RECT 1604.6600 930.1600 1606.2600 930.6400 ;
        RECT 1604.6600 935.6000 1606.2600 936.0800 ;
        RECT 1592.9000 935.6000 1595.9000 936.0800 ;
        RECT 1592.9000 930.1600 1595.9000 930.6400 ;
        RECT 1592.9000 941.0400 1595.9000 941.5200 ;
        RECT 1604.6600 941.0400 1606.2600 941.5200 ;
        RECT 1694.6600 913.8400 1696.2600 914.3200 ;
        RECT 1694.6600 919.2800 1696.2600 919.7600 ;
        RECT 1694.6600 924.7200 1696.2600 925.2000 ;
        RECT 1694.6600 902.9600 1696.2600 903.4400 ;
        RECT 1694.6600 908.4000 1696.2600 908.8800 ;
        RECT 1649.6600 913.8400 1651.2600 914.3200 ;
        RECT 1649.6600 919.2800 1651.2600 919.7600 ;
        RECT 1649.6600 924.7200 1651.2600 925.2000 ;
        RECT 1649.6600 902.9600 1651.2600 903.4400 ;
        RECT 1649.6600 908.4000 1651.2600 908.8800 ;
        RECT 1694.6600 886.6400 1696.2600 887.1200 ;
        RECT 1694.6600 892.0800 1696.2600 892.5600 ;
        RECT 1694.6600 897.5200 1696.2600 898.0000 ;
        RECT 1694.6600 875.7600 1696.2600 876.2400 ;
        RECT 1694.6600 881.2000 1696.2600 881.6800 ;
        RECT 1649.6600 886.6400 1651.2600 887.1200 ;
        RECT 1649.6600 892.0800 1651.2600 892.5600 ;
        RECT 1649.6600 897.5200 1651.2600 898.0000 ;
        RECT 1649.6600 875.7600 1651.2600 876.2400 ;
        RECT 1649.6600 881.2000 1651.2600 881.6800 ;
        RECT 1604.6600 913.8400 1606.2600 914.3200 ;
        RECT 1604.6600 919.2800 1606.2600 919.7600 ;
        RECT 1604.6600 924.7200 1606.2600 925.2000 ;
        RECT 1592.9000 913.8400 1595.9000 914.3200 ;
        RECT 1592.9000 919.2800 1595.9000 919.7600 ;
        RECT 1592.9000 924.7200 1595.9000 925.2000 ;
        RECT 1604.6600 902.9600 1606.2600 903.4400 ;
        RECT 1604.6600 908.4000 1606.2600 908.8800 ;
        RECT 1592.9000 902.9600 1595.9000 903.4400 ;
        RECT 1592.9000 908.4000 1595.9000 908.8800 ;
        RECT 1604.6600 886.6400 1606.2600 887.1200 ;
        RECT 1604.6600 892.0800 1606.2600 892.5600 ;
        RECT 1604.6600 897.5200 1606.2600 898.0000 ;
        RECT 1592.9000 886.6400 1595.9000 887.1200 ;
        RECT 1592.9000 892.0800 1595.9000 892.5600 ;
        RECT 1592.9000 897.5200 1595.9000 898.0000 ;
        RECT 1604.6600 875.7600 1606.2600 876.2400 ;
        RECT 1604.6600 881.2000 1606.2600 881.6800 ;
        RECT 1592.9000 875.7600 1595.9000 876.2400 ;
        RECT 1592.9000 881.2000 1595.9000 881.6800 ;
        RECT 1797.0000 859.4400 1800.0000 859.9200 ;
        RECT 1797.0000 864.8800 1800.0000 865.3600 ;
        RECT 1797.0000 870.3200 1800.0000 870.8000 ;
        RECT 1784.6600 859.4400 1786.2600 859.9200 ;
        RECT 1784.6600 864.8800 1786.2600 865.3600 ;
        RECT 1784.6600 870.3200 1786.2600 870.8000 ;
        RECT 1797.0000 848.5600 1800.0000 849.0400 ;
        RECT 1797.0000 854.0000 1800.0000 854.4800 ;
        RECT 1784.6600 848.5600 1786.2600 849.0400 ;
        RECT 1784.6600 854.0000 1786.2600 854.4800 ;
        RECT 1797.0000 832.2400 1800.0000 832.7200 ;
        RECT 1797.0000 837.6800 1800.0000 838.1600 ;
        RECT 1797.0000 843.1200 1800.0000 843.6000 ;
        RECT 1784.6600 832.2400 1786.2600 832.7200 ;
        RECT 1784.6600 837.6800 1786.2600 838.1600 ;
        RECT 1784.6600 843.1200 1786.2600 843.6000 ;
        RECT 1797.0000 821.3600 1800.0000 821.8400 ;
        RECT 1797.0000 826.8000 1800.0000 827.2800 ;
        RECT 1784.6600 821.3600 1786.2600 821.8400 ;
        RECT 1784.6600 826.8000 1786.2600 827.2800 ;
        RECT 1739.6600 859.4400 1741.2600 859.9200 ;
        RECT 1739.6600 864.8800 1741.2600 865.3600 ;
        RECT 1739.6600 870.3200 1741.2600 870.8000 ;
        RECT 1739.6600 848.5600 1741.2600 849.0400 ;
        RECT 1739.6600 854.0000 1741.2600 854.4800 ;
        RECT 1739.6600 832.2400 1741.2600 832.7200 ;
        RECT 1739.6600 837.6800 1741.2600 838.1600 ;
        RECT 1739.6600 843.1200 1741.2600 843.6000 ;
        RECT 1739.6600 821.3600 1741.2600 821.8400 ;
        RECT 1739.6600 826.8000 1741.2600 827.2800 ;
        RECT 1797.0000 805.0400 1800.0000 805.5200 ;
        RECT 1797.0000 810.4800 1800.0000 810.9600 ;
        RECT 1797.0000 815.9200 1800.0000 816.4000 ;
        RECT 1784.6600 805.0400 1786.2600 805.5200 ;
        RECT 1784.6600 810.4800 1786.2600 810.9600 ;
        RECT 1784.6600 815.9200 1786.2600 816.4000 ;
        RECT 1797.0000 794.1600 1800.0000 794.6400 ;
        RECT 1797.0000 799.6000 1800.0000 800.0800 ;
        RECT 1784.6600 794.1600 1786.2600 794.6400 ;
        RECT 1784.6600 799.6000 1786.2600 800.0800 ;
        RECT 1797.0000 777.8400 1800.0000 778.3200 ;
        RECT 1797.0000 783.2800 1800.0000 783.7600 ;
        RECT 1797.0000 788.7200 1800.0000 789.2000 ;
        RECT 1784.6600 777.8400 1786.2600 778.3200 ;
        RECT 1784.6600 783.2800 1786.2600 783.7600 ;
        RECT 1784.6600 788.7200 1786.2600 789.2000 ;
        RECT 1797.0000 772.4000 1800.0000 772.8800 ;
        RECT 1784.6600 772.4000 1786.2600 772.8800 ;
        RECT 1739.6600 805.0400 1741.2600 805.5200 ;
        RECT 1739.6600 810.4800 1741.2600 810.9600 ;
        RECT 1739.6600 815.9200 1741.2600 816.4000 ;
        RECT 1739.6600 794.1600 1741.2600 794.6400 ;
        RECT 1739.6600 799.6000 1741.2600 800.0800 ;
        RECT 1739.6600 777.8400 1741.2600 778.3200 ;
        RECT 1739.6600 783.2800 1741.2600 783.7600 ;
        RECT 1739.6600 788.7200 1741.2600 789.2000 ;
        RECT 1739.6600 772.4000 1741.2600 772.8800 ;
        RECT 1694.6600 859.4400 1696.2600 859.9200 ;
        RECT 1694.6600 864.8800 1696.2600 865.3600 ;
        RECT 1694.6600 870.3200 1696.2600 870.8000 ;
        RECT 1694.6600 848.5600 1696.2600 849.0400 ;
        RECT 1694.6600 854.0000 1696.2600 854.4800 ;
        RECT 1649.6600 859.4400 1651.2600 859.9200 ;
        RECT 1649.6600 864.8800 1651.2600 865.3600 ;
        RECT 1649.6600 870.3200 1651.2600 870.8000 ;
        RECT 1649.6600 848.5600 1651.2600 849.0400 ;
        RECT 1649.6600 854.0000 1651.2600 854.4800 ;
        RECT 1694.6600 832.2400 1696.2600 832.7200 ;
        RECT 1694.6600 837.6800 1696.2600 838.1600 ;
        RECT 1694.6600 843.1200 1696.2600 843.6000 ;
        RECT 1694.6600 821.3600 1696.2600 821.8400 ;
        RECT 1694.6600 826.8000 1696.2600 827.2800 ;
        RECT 1649.6600 832.2400 1651.2600 832.7200 ;
        RECT 1649.6600 837.6800 1651.2600 838.1600 ;
        RECT 1649.6600 843.1200 1651.2600 843.6000 ;
        RECT 1649.6600 821.3600 1651.2600 821.8400 ;
        RECT 1649.6600 826.8000 1651.2600 827.2800 ;
        RECT 1604.6600 859.4400 1606.2600 859.9200 ;
        RECT 1604.6600 864.8800 1606.2600 865.3600 ;
        RECT 1604.6600 870.3200 1606.2600 870.8000 ;
        RECT 1592.9000 859.4400 1595.9000 859.9200 ;
        RECT 1592.9000 864.8800 1595.9000 865.3600 ;
        RECT 1592.9000 870.3200 1595.9000 870.8000 ;
        RECT 1604.6600 848.5600 1606.2600 849.0400 ;
        RECT 1604.6600 854.0000 1606.2600 854.4800 ;
        RECT 1592.9000 848.5600 1595.9000 849.0400 ;
        RECT 1592.9000 854.0000 1595.9000 854.4800 ;
        RECT 1604.6600 832.2400 1606.2600 832.7200 ;
        RECT 1604.6600 837.6800 1606.2600 838.1600 ;
        RECT 1604.6600 843.1200 1606.2600 843.6000 ;
        RECT 1592.9000 832.2400 1595.9000 832.7200 ;
        RECT 1592.9000 837.6800 1595.9000 838.1600 ;
        RECT 1592.9000 843.1200 1595.9000 843.6000 ;
        RECT 1604.6600 821.3600 1606.2600 821.8400 ;
        RECT 1604.6600 826.8000 1606.2600 827.2800 ;
        RECT 1592.9000 821.3600 1595.9000 821.8400 ;
        RECT 1592.9000 826.8000 1595.9000 827.2800 ;
        RECT 1694.6600 805.0400 1696.2600 805.5200 ;
        RECT 1694.6600 810.4800 1696.2600 810.9600 ;
        RECT 1694.6600 815.9200 1696.2600 816.4000 ;
        RECT 1694.6600 794.1600 1696.2600 794.6400 ;
        RECT 1694.6600 799.6000 1696.2600 800.0800 ;
        RECT 1649.6600 805.0400 1651.2600 805.5200 ;
        RECT 1649.6600 810.4800 1651.2600 810.9600 ;
        RECT 1649.6600 815.9200 1651.2600 816.4000 ;
        RECT 1649.6600 794.1600 1651.2600 794.6400 ;
        RECT 1649.6600 799.6000 1651.2600 800.0800 ;
        RECT 1694.6600 777.8400 1696.2600 778.3200 ;
        RECT 1694.6600 783.2800 1696.2600 783.7600 ;
        RECT 1694.6600 788.7200 1696.2600 789.2000 ;
        RECT 1694.6600 772.4000 1696.2600 772.8800 ;
        RECT 1649.6600 777.8400 1651.2600 778.3200 ;
        RECT 1649.6600 783.2800 1651.2600 783.7600 ;
        RECT 1649.6600 788.7200 1651.2600 789.2000 ;
        RECT 1649.6600 772.4000 1651.2600 772.8800 ;
        RECT 1604.6600 805.0400 1606.2600 805.5200 ;
        RECT 1604.6600 810.4800 1606.2600 810.9600 ;
        RECT 1604.6600 815.9200 1606.2600 816.4000 ;
        RECT 1592.9000 805.0400 1595.9000 805.5200 ;
        RECT 1592.9000 810.4800 1595.9000 810.9600 ;
        RECT 1592.9000 815.9200 1595.9000 816.4000 ;
        RECT 1604.6600 794.1600 1606.2600 794.6400 ;
        RECT 1604.6600 799.6000 1606.2600 800.0800 ;
        RECT 1592.9000 794.1600 1595.9000 794.6400 ;
        RECT 1592.9000 799.6000 1595.9000 800.0800 ;
        RECT 1604.6600 777.8400 1606.2600 778.3200 ;
        RECT 1604.6600 783.2800 1606.2600 783.7600 ;
        RECT 1604.6600 788.7200 1606.2600 789.2000 ;
        RECT 1592.9000 777.8400 1595.9000 778.3200 ;
        RECT 1592.9000 783.2800 1595.9000 783.7600 ;
        RECT 1592.9000 788.7200 1595.9000 789.2000 ;
        RECT 1592.9000 772.4000 1595.9000 772.8800 ;
        RECT 1604.6600 772.4000 1606.2600 772.8800 ;
        RECT 1592.9000 977.3100 1800.0000 980.3100 ;
        RECT 1592.9000 764.2100 1800.0000 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1814.1200 2830.6100 1816.1200 2857.5400 ;
        RECT 2017.2200 2830.6100 2019.2200 2857.5400 ;
      LAYER met3 ;
        RECT 2017.2200 2847.3200 2019.2200 2847.8000 ;
        RECT 1814.1200 2847.3200 1816.1200 2847.8000 ;
        RECT 2017.2200 2841.8800 2019.2200 2842.3600 ;
        RECT 2017.2200 2836.4400 2019.2200 2836.9200 ;
        RECT 1814.1200 2841.8800 1816.1200 2842.3600 ;
        RECT 1814.1200 2836.4400 1816.1200 2836.9200 ;
        RECT 1814.1200 2855.5400 2019.2200 2857.5400 ;
        RECT 1814.1200 2830.6100 2019.2200 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1814.1200 76.2900 1816.1200 521.0800 ;
        RECT 2017.2200 76.2900 2019.2200 521.0800 ;
        RECT 1824.8800 76.2900 1826.4800 521.0800 ;
        RECT 1869.8800 76.2900 1871.4800 521.0800 ;
        RECT 1914.8800 76.2900 1916.4800 521.0800 ;
        RECT 1959.8800 76.2900 1961.4800 521.0800 ;
        RECT 2004.8800 76.2900 2006.4800 521.0800 ;
      LAYER met3 ;
        RECT 2017.2200 513.2400 2019.2200 513.7200 ;
        RECT 2017.2200 507.8000 2019.2200 508.2800 ;
        RECT 2017.2200 502.3600 2019.2200 502.8400 ;
        RECT 2017.2200 496.9200 2019.2200 497.4000 ;
        RECT 2017.2200 491.4800 2019.2200 491.9600 ;
        RECT 2017.2200 486.0400 2019.2200 486.5200 ;
        RECT 2017.2200 480.6000 2019.2200 481.0800 ;
        RECT 2017.2200 475.1600 2019.2200 475.6400 ;
        RECT 2017.2200 469.7200 2019.2200 470.2000 ;
        RECT 2017.2200 464.2800 2019.2200 464.7600 ;
        RECT 2017.2200 458.8400 2019.2200 459.3200 ;
        RECT 2017.2200 453.4000 2019.2200 453.8800 ;
        RECT 2017.2200 447.9600 2019.2200 448.4400 ;
        RECT 2017.2200 442.5200 2019.2200 443.0000 ;
        RECT 2017.2200 437.0800 2019.2200 437.5600 ;
        RECT 2017.2200 431.6400 2019.2200 432.1200 ;
        RECT 2017.2200 426.2000 2019.2200 426.6800 ;
        RECT 2017.2200 420.7600 2019.2200 421.2400 ;
        RECT 2017.2200 415.3200 2019.2200 415.8000 ;
        RECT 2017.2200 409.8800 2019.2200 410.3600 ;
        RECT 2017.2200 404.4400 2019.2200 404.9200 ;
        RECT 2017.2200 399.0000 2019.2200 399.4800 ;
        RECT 2017.2200 393.5600 2019.2200 394.0400 ;
        RECT 2017.2200 388.1200 2019.2200 388.6000 ;
        RECT 2017.2200 377.2400 2019.2200 377.7200 ;
        RECT 2017.2200 371.8000 2019.2200 372.2800 ;
        RECT 2017.2200 366.3600 2019.2200 366.8400 ;
        RECT 2017.2200 360.9200 2019.2200 361.4000 ;
        RECT 2017.2200 355.4800 2019.2200 355.9600 ;
        RECT 2017.2200 382.6800 2019.2200 383.1600 ;
        RECT 2017.2200 350.0400 2019.2200 350.5200 ;
        RECT 2017.2200 344.6000 2019.2200 345.0800 ;
        RECT 2017.2200 339.1600 2019.2200 339.6400 ;
        RECT 2017.2200 333.7200 2019.2200 334.2000 ;
        RECT 2017.2200 328.2800 2019.2200 328.7600 ;
        RECT 2017.2200 322.8400 2019.2200 323.3200 ;
        RECT 2017.2200 317.4000 2019.2200 317.8800 ;
        RECT 2017.2200 311.9600 2019.2200 312.4400 ;
        RECT 2017.2200 306.5200 2019.2200 307.0000 ;
        RECT 2017.2200 301.0800 2019.2200 301.5600 ;
        RECT 1814.1200 513.2400 1816.1200 513.7200 ;
        RECT 1814.1200 507.8000 1816.1200 508.2800 ;
        RECT 1814.1200 502.3600 1816.1200 502.8400 ;
        RECT 1814.1200 496.9200 1816.1200 497.4000 ;
        RECT 1814.1200 491.4800 1816.1200 491.9600 ;
        RECT 1814.1200 486.0400 1816.1200 486.5200 ;
        RECT 1814.1200 480.6000 1816.1200 481.0800 ;
        RECT 1814.1200 475.1600 1816.1200 475.6400 ;
        RECT 1814.1200 469.7200 1816.1200 470.2000 ;
        RECT 1814.1200 464.2800 1816.1200 464.7600 ;
        RECT 1814.1200 458.8400 1816.1200 459.3200 ;
        RECT 1814.1200 453.4000 1816.1200 453.8800 ;
        RECT 1814.1200 447.9600 1816.1200 448.4400 ;
        RECT 1814.1200 442.5200 1816.1200 443.0000 ;
        RECT 1814.1200 437.0800 1816.1200 437.5600 ;
        RECT 1814.1200 431.6400 1816.1200 432.1200 ;
        RECT 1814.1200 426.2000 1816.1200 426.6800 ;
        RECT 1814.1200 420.7600 1816.1200 421.2400 ;
        RECT 1814.1200 415.3200 1816.1200 415.8000 ;
        RECT 1814.1200 409.8800 1816.1200 410.3600 ;
        RECT 1814.1200 404.4400 1816.1200 404.9200 ;
        RECT 1814.1200 399.0000 1816.1200 399.4800 ;
        RECT 1814.1200 393.5600 1816.1200 394.0400 ;
        RECT 1814.1200 388.1200 1816.1200 388.6000 ;
        RECT 1814.1200 377.2400 1816.1200 377.7200 ;
        RECT 1814.1200 371.8000 1816.1200 372.2800 ;
        RECT 1814.1200 366.3600 1816.1200 366.8400 ;
        RECT 1814.1200 360.9200 1816.1200 361.4000 ;
        RECT 1814.1200 355.4800 1816.1200 355.9600 ;
        RECT 1814.1200 382.6800 1816.1200 383.1600 ;
        RECT 1814.1200 350.0400 1816.1200 350.5200 ;
        RECT 1814.1200 344.6000 1816.1200 345.0800 ;
        RECT 1814.1200 339.1600 1816.1200 339.6400 ;
        RECT 1814.1200 333.7200 1816.1200 334.2000 ;
        RECT 1814.1200 328.2800 1816.1200 328.7600 ;
        RECT 1814.1200 322.8400 1816.1200 323.3200 ;
        RECT 1814.1200 317.4000 1816.1200 317.8800 ;
        RECT 1814.1200 311.9600 1816.1200 312.4400 ;
        RECT 1814.1200 306.5200 1816.1200 307.0000 ;
        RECT 1814.1200 301.0800 1816.1200 301.5600 ;
        RECT 2017.2200 295.6400 2019.2200 296.1200 ;
        RECT 2017.2200 290.2000 2019.2200 290.6800 ;
        RECT 2017.2200 284.7600 2019.2200 285.2400 ;
        RECT 2017.2200 279.3200 2019.2200 279.8000 ;
        RECT 2017.2200 273.8800 2019.2200 274.3600 ;
        RECT 2017.2200 268.4400 2019.2200 268.9200 ;
        RECT 2017.2200 263.0000 2019.2200 263.4800 ;
        RECT 2017.2200 257.5600 2019.2200 258.0400 ;
        RECT 2017.2200 252.1200 2019.2200 252.6000 ;
        RECT 2017.2200 246.6800 2019.2200 247.1600 ;
        RECT 2017.2200 241.2400 2019.2200 241.7200 ;
        RECT 2017.2200 235.8000 2019.2200 236.2800 ;
        RECT 2017.2200 230.3600 2019.2200 230.8400 ;
        RECT 2017.2200 224.9200 2019.2200 225.4000 ;
        RECT 2017.2200 219.4800 2019.2200 219.9600 ;
        RECT 2017.2200 208.6000 2019.2200 209.0800 ;
        RECT 2017.2200 203.1600 2019.2200 203.6400 ;
        RECT 2017.2200 197.7200 2019.2200 198.2000 ;
        RECT 2017.2200 192.2800 2019.2200 192.7600 ;
        RECT 2017.2200 186.8400 2019.2200 187.3200 ;
        RECT 2017.2200 214.0400 2019.2200 214.5200 ;
        RECT 2017.2200 181.4000 2019.2200 181.8800 ;
        RECT 2017.2200 175.9600 2019.2200 176.4400 ;
        RECT 2017.2200 170.5200 2019.2200 171.0000 ;
        RECT 2017.2200 165.0800 2019.2200 165.5600 ;
        RECT 2017.2200 159.6400 2019.2200 160.1200 ;
        RECT 2017.2200 154.2000 2019.2200 154.6800 ;
        RECT 2017.2200 148.7600 2019.2200 149.2400 ;
        RECT 2017.2200 143.3200 2019.2200 143.8000 ;
        RECT 2017.2200 137.8800 2019.2200 138.3600 ;
        RECT 2017.2200 132.4400 2019.2200 132.9200 ;
        RECT 2017.2200 127.0000 2019.2200 127.4800 ;
        RECT 2017.2200 121.5600 2019.2200 122.0400 ;
        RECT 2017.2200 116.1200 2019.2200 116.6000 ;
        RECT 2017.2200 110.6800 2019.2200 111.1600 ;
        RECT 2017.2200 105.2400 2019.2200 105.7200 ;
        RECT 2017.2200 99.8000 2019.2200 100.2800 ;
        RECT 2017.2200 94.3600 2019.2200 94.8400 ;
        RECT 2017.2200 88.9200 2019.2200 89.4000 ;
        RECT 2017.2200 83.4800 2019.2200 83.9600 ;
        RECT 1814.1200 295.6400 1816.1200 296.1200 ;
        RECT 1814.1200 290.2000 1816.1200 290.6800 ;
        RECT 1814.1200 284.7600 1816.1200 285.2400 ;
        RECT 1814.1200 279.3200 1816.1200 279.8000 ;
        RECT 1814.1200 273.8800 1816.1200 274.3600 ;
        RECT 1814.1200 268.4400 1816.1200 268.9200 ;
        RECT 1814.1200 263.0000 1816.1200 263.4800 ;
        RECT 1814.1200 257.5600 1816.1200 258.0400 ;
        RECT 1814.1200 252.1200 1816.1200 252.6000 ;
        RECT 1814.1200 246.6800 1816.1200 247.1600 ;
        RECT 1814.1200 241.2400 1816.1200 241.7200 ;
        RECT 1814.1200 235.8000 1816.1200 236.2800 ;
        RECT 1814.1200 230.3600 1816.1200 230.8400 ;
        RECT 1814.1200 224.9200 1816.1200 225.4000 ;
        RECT 1814.1200 219.4800 1816.1200 219.9600 ;
        RECT 1814.1200 208.6000 1816.1200 209.0800 ;
        RECT 1814.1200 203.1600 1816.1200 203.6400 ;
        RECT 1814.1200 197.7200 1816.1200 198.2000 ;
        RECT 1814.1200 192.2800 1816.1200 192.7600 ;
        RECT 1814.1200 186.8400 1816.1200 187.3200 ;
        RECT 1814.1200 214.0400 1816.1200 214.5200 ;
        RECT 1814.1200 181.4000 1816.1200 181.8800 ;
        RECT 1814.1200 175.9600 1816.1200 176.4400 ;
        RECT 1814.1200 170.5200 1816.1200 171.0000 ;
        RECT 1814.1200 165.0800 1816.1200 165.5600 ;
        RECT 1814.1200 159.6400 1816.1200 160.1200 ;
        RECT 1814.1200 154.2000 1816.1200 154.6800 ;
        RECT 1814.1200 148.7600 1816.1200 149.2400 ;
        RECT 1814.1200 143.3200 1816.1200 143.8000 ;
        RECT 1814.1200 137.8800 1816.1200 138.3600 ;
        RECT 1814.1200 132.4400 1816.1200 132.9200 ;
        RECT 1814.1200 127.0000 1816.1200 127.4800 ;
        RECT 1814.1200 121.5600 1816.1200 122.0400 ;
        RECT 1814.1200 116.1200 1816.1200 116.6000 ;
        RECT 1814.1200 110.6800 1816.1200 111.1600 ;
        RECT 1814.1200 105.2400 1816.1200 105.7200 ;
        RECT 1814.1200 99.8000 1816.1200 100.2800 ;
        RECT 1814.1200 94.3600 1816.1200 94.8400 ;
        RECT 1814.1200 88.9200 1816.1200 89.4000 ;
        RECT 1814.1200 83.4800 1816.1200 83.9600 ;
        RECT 1814.1200 519.0800 2019.2200 521.0800 ;
        RECT 1814.1200 76.2900 2019.2200 78.2900 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'S_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1814.1200 34.6700 1816.1200 61.6000 ;
        RECT 2017.2200 34.6700 2019.2200 61.6000 ;
      LAYER met3 ;
        RECT 2017.2200 51.3800 2019.2200 51.8600 ;
        RECT 1814.1200 51.3800 1816.1200 51.8600 ;
        RECT 2017.2200 45.9400 2019.2200 46.4200 ;
        RECT 2017.2200 40.5000 2019.2200 40.9800 ;
        RECT 1814.1200 45.9400 1816.1200 46.4200 ;
        RECT 1814.1200 40.5000 1816.1200 40.9800 ;
        RECT 1814.1200 59.6000 2019.2200 61.6000 ;
        RECT 1814.1200 34.6700 2019.2200 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1814.1200 2372.6900 1816.1200 2817.4800 ;
        RECT 2017.2200 2372.6900 2019.2200 2817.4800 ;
        RECT 1824.8800 2372.6900 1826.4800 2817.4800 ;
        RECT 1869.8800 2372.6900 1871.4800 2817.4800 ;
        RECT 1914.8800 2372.6900 1916.4800 2817.4800 ;
        RECT 1959.8800 2372.6900 1961.4800 2817.4800 ;
        RECT 2004.8800 2372.6900 2006.4800 2817.4800 ;
      LAYER met3 ;
        RECT 2017.2200 2809.6400 2019.2200 2810.1200 ;
        RECT 2017.2200 2804.2000 2019.2200 2804.6800 ;
        RECT 2017.2200 2798.7600 2019.2200 2799.2400 ;
        RECT 2017.2200 2793.3200 2019.2200 2793.8000 ;
        RECT 2017.2200 2787.8800 2019.2200 2788.3600 ;
        RECT 2017.2200 2782.4400 2019.2200 2782.9200 ;
        RECT 2017.2200 2777.0000 2019.2200 2777.4800 ;
        RECT 2017.2200 2771.5600 2019.2200 2772.0400 ;
        RECT 2017.2200 2766.1200 2019.2200 2766.6000 ;
        RECT 2017.2200 2760.6800 2019.2200 2761.1600 ;
        RECT 2017.2200 2755.2400 2019.2200 2755.7200 ;
        RECT 2017.2200 2749.8000 2019.2200 2750.2800 ;
        RECT 2017.2200 2744.3600 2019.2200 2744.8400 ;
        RECT 2017.2200 2738.9200 2019.2200 2739.4000 ;
        RECT 2017.2200 2733.4800 2019.2200 2733.9600 ;
        RECT 2017.2200 2728.0400 2019.2200 2728.5200 ;
        RECT 2017.2200 2722.6000 2019.2200 2723.0800 ;
        RECT 2017.2200 2717.1600 2019.2200 2717.6400 ;
        RECT 2017.2200 2711.7200 2019.2200 2712.2000 ;
        RECT 2017.2200 2706.2800 2019.2200 2706.7600 ;
        RECT 2017.2200 2700.8400 2019.2200 2701.3200 ;
        RECT 2017.2200 2695.4000 2019.2200 2695.8800 ;
        RECT 2017.2200 2689.9600 2019.2200 2690.4400 ;
        RECT 2017.2200 2684.5200 2019.2200 2685.0000 ;
        RECT 2017.2200 2673.6400 2019.2200 2674.1200 ;
        RECT 2017.2200 2668.2000 2019.2200 2668.6800 ;
        RECT 2017.2200 2662.7600 2019.2200 2663.2400 ;
        RECT 2017.2200 2657.3200 2019.2200 2657.8000 ;
        RECT 2017.2200 2651.8800 2019.2200 2652.3600 ;
        RECT 2017.2200 2679.0800 2019.2200 2679.5600 ;
        RECT 2017.2200 2646.4400 2019.2200 2646.9200 ;
        RECT 2017.2200 2641.0000 2019.2200 2641.4800 ;
        RECT 2017.2200 2635.5600 2019.2200 2636.0400 ;
        RECT 2017.2200 2630.1200 2019.2200 2630.6000 ;
        RECT 2017.2200 2624.6800 2019.2200 2625.1600 ;
        RECT 2017.2200 2619.2400 2019.2200 2619.7200 ;
        RECT 2017.2200 2613.8000 2019.2200 2614.2800 ;
        RECT 2017.2200 2608.3600 2019.2200 2608.8400 ;
        RECT 2017.2200 2602.9200 2019.2200 2603.4000 ;
        RECT 2017.2200 2597.4800 2019.2200 2597.9600 ;
        RECT 1814.1200 2809.6400 1816.1200 2810.1200 ;
        RECT 1814.1200 2804.2000 1816.1200 2804.6800 ;
        RECT 1814.1200 2798.7600 1816.1200 2799.2400 ;
        RECT 1814.1200 2793.3200 1816.1200 2793.8000 ;
        RECT 1814.1200 2787.8800 1816.1200 2788.3600 ;
        RECT 1814.1200 2782.4400 1816.1200 2782.9200 ;
        RECT 1814.1200 2777.0000 1816.1200 2777.4800 ;
        RECT 1814.1200 2771.5600 1816.1200 2772.0400 ;
        RECT 1814.1200 2766.1200 1816.1200 2766.6000 ;
        RECT 1814.1200 2760.6800 1816.1200 2761.1600 ;
        RECT 1814.1200 2755.2400 1816.1200 2755.7200 ;
        RECT 1814.1200 2749.8000 1816.1200 2750.2800 ;
        RECT 1814.1200 2744.3600 1816.1200 2744.8400 ;
        RECT 1814.1200 2738.9200 1816.1200 2739.4000 ;
        RECT 1814.1200 2733.4800 1816.1200 2733.9600 ;
        RECT 1814.1200 2728.0400 1816.1200 2728.5200 ;
        RECT 1814.1200 2722.6000 1816.1200 2723.0800 ;
        RECT 1814.1200 2717.1600 1816.1200 2717.6400 ;
        RECT 1814.1200 2711.7200 1816.1200 2712.2000 ;
        RECT 1814.1200 2706.2800 1816.1200 2706.7600 ;
        RECT 1814.1200 2700.8400 1816.1200 2701.3200 ;
        RECT 1814.1200 2695.4000 1816.1200 2695.8800 ;
        RECT 1814.1200 2689.9600 1816.1200 2690.4400 ;
        RECT 1814.1200 2684.5200 1816.1200 2685.0000 ;
        RECT 1814.1200 2673.6400 1816.1200 2674.1200 ;
        RECT 1814.1200 2668.2000 1816.1200 2668.6800 ;
        RECT 1814.1200 2662.7600 1816.1200 2663.2400 ;
        RECT 1814.1200 2657.3200 1816.1200 2657.8000 ;
        RECT 1814.1200 2651.8800 1816.1200 2652.3600 ;
        RECT 1814.1200 2679.0800 1816.1200 2679.5600 ;
        RECT 1814.1200 2646.4400 1816.1200 2646.9200 ;
        RECT 1814.1200 2641.0000 1816.1200 2641.4800 ;
        RECT 1814.1200 2635.5600 1816.1200 2636.0400 ;
        RECT 1814.1200 2630.1200 1816.1200 2630.6000 ;
        RECT 1814.1200 2624.6800 1816.1200 2625.1600 ;
        RECT 1814.1200 2619.2400 1816.1200 2619.7200 ;
        RECT 1814.1200 2613.8000 1816.1200 2614.2800 ;
        RECT 1814.1200 2608.3600 1816.1200 2608.8400 ;
        RECT 1814.1200 2602.9200 1816.1200 2603.4000 ;
        RECT 1814.1200 2597.4800 1816.1200 2597.9600 ;
        RECT 2017.2200 2592.0400 2019.2200 2592.5200 ;
        RECT 2017.2200 2586.6000 2019.2200 2587.0800 ;
        RECT 2017.2200 2581.1600 2019.2200 2581.6400 ;
        RECT 2017.2200 2575.7200 2019.2200 2576.2000 ;
        RECT 2017.2200 2570.2800 2019.2200 2570.7600 ;
        RECT 2017.2200 2564.8400 2019.2200 2565.3200 ;
        RECT 2017.2200 2559.4000 2019.2200 2559.8800 ;
        RECT 2017.2200 2553.9600 2019.2200 2554.4400 ;
        RECT 2017.2200 2548.5200 2019.2200 2549.0000 ;
        RECT 2017.2200 2543.0800 2019.2200 2543.5600 ;
        RECT 2017.2200 2537.6400 2019.2200 2538.1200 ;
        RECT 2017.2200 2532.2000 2019.2200 2532.6800 ;
        RECT 2017.2200 2526.7600 2019.2200 2527.2400 ;
        RECT 2017.2200 2521.3200 2019.2200 2521.8000 ;
        RECT 2017.2200 2515.8800 2019.2200 2516.3600 ;
        RECT 2017.2200 2505.0000 2019.2200 2505.4800 ;
        RECT 2017.2200 2499.5600 2019.2200 2500.0400 ;
        RECT 2017.2200 2494.1200 2019.2200 2494.6000 ;
        RECT 2017.2200 2488.6800 2019.2200 2489.1600 ;
        RECT 2017.2200 2483.2400 2019.2200 2483.7200 ;
        RECT 2017.2200 2510.4400 2019.2200 2510.9200 ;
        RECT 2017.2200 2477.8000 2019.2200 2478.2800 ;
        RECT 2017.2200 2472.3600 2019.2200 2472.8400 ;
        RECT 2017.2200 2466.9200 2019.2200 2467.4000 ;
        RECT 2017.2200 2461.4800 2019.2200 2461.9600 ;
        RECT 2017.2200 2456.0400 2019.2200 2456.5200 ;
        RECT 2017.2200 2450.6000 2019.2200 2451.0800 ;
        RECT 2017.2200 2445.1600 2019.2200 2445.6400 ;
        RECT 2017.2200 2439.7200 2019.2200 2440.2000 ;
        RECT 2017.2200 2434.2800 2019.2200 2434.7600 ;
        RECT 2017.2200 2428.8400 2019.2200 2429.3200 ;
        RECT 2017.2200 2423.4000 2019.2200 2423.8800 ;
        RECT 2017.2200 2417.9600 2019.2200 2418.4400 ;
        RECT 2017.2200 2412.5200 2019.2200 2413.0000 ;
        RECT 2017.2200 2407.0800 2019.2200 2407.5600 ;
        RECT 2017.2200 2401.6400 2019.2200 2402.1200 ;
        RECT 2017.2200 2396.2000 2019.2200 2396.6800 ;
        RECT 2017.2200 2390.7600 2019.2200 2391.2400 ;
        RECT 2017.2200 2385.3200 2019.2200 2385.8000 ;
        RECT 2017.2200 2379.8800 2019.2200 2380.3600 ;
        RECT 1814.1200 2592.0400 1816.1200 2592.5200 ;
        RECT 1814.1200 2586.6000 1816.1200 2587.0800 ;
        RECT 1814.1200 2581.1600 1816.1200 2581.6400 ;
        RECT 1814.1200 2575.7200 1816.1200 2576.2000 ;
        RECT 1814.1200 2570.2800 1816.1200 2570.7600 ;
        RECT 1814.1200 2564.8400 1816.1200 2565.3200 ;
        RECT 1814.1200 2559.4000 1816.1200 2559.8800 ;
        RECT 1814.1200 2553.9600 1816.1200 2554.4400 ;
        RECT 1814.1200 2548.5200 1816.1200 2549.0000 ;
        RECT 1814.1200 2543.0800 1816.1200 2543.5600 ;
        RECT 1814.1200 2537.6400 1816.1200 2538.1200 ;
        RECT 1814.1200 2532.2000 1816.1200 2532.6800 ;
        RECT 1814.1200 2526.7600 1816.1200 2527.2400 ;
        RECT 1814.1200 2521.3200 1816.1200 2521.8000 ;
        RECT 1814.1200 2515.8800 1816.1200 2516.3600 ;
        RECT 1814.1200 2505.0000 1816.1200 2505.4800 ;
        RECT 1814.1200 2499.5600 1816.1200 2500.0400 ;
        RECT 1814.1200 2494.1200 1816.1200 2494.6000 ;
        RECT 1814.1200 2488.6800 1816.1200 2489.1600 ;
        RECT 1814.1200 2483.2400 1816.1200 2483.7200 ;
        RECT 1814.1200 2510.4400 1816.1200 2510.9200 ;
        RECT 1814.1200 2477.8000 1816.1200 2478.2800 ;
        RECT 1814.1200 2472.3600 1816.1200 2472.8400 ;
        RECT 1814.1200 2466.9200 1816.1200 2467.4000 ;
        RECT 1814.1200 2461.4800 1816.1200 2461.9600 ;
        RECT 1814.1200 2456.0400 1816.1200 2456.5200 ;
        RECT 1814.1200 2450.6000 1816.1200 2451.0800 ;
        RECT 1814.1200 2445.1600 1816.1200 2445.6400 ;
        RECT 1814.1200 2439.7200 1816.1200 2440.2000 ;
        RECT 1814.1200 2434.2800 1816.1200 2434.7600 ;
        RECT 1814.1200 2428.8400 1816.1200 2429.3200 ;
        RECT 1814.1200 2423.4000 1816.1200 2423.8800 ;
        RECT 1814.1200 2417.9600 1816.1200 2418.4400 ;
        RECT 1814.1200 2412.5200 1816.1200 2413.0000 ;
        RECT 1814.1200 2407.0800 1816.1200 2407.5600 ;
        RECT 1814.1200 2401.6400 1816.1200 2402.1200 ;
        RECT 1814.1200 2396.2000 1816.1200 2396.6800 ;
        RECT 1814.1200 2390.7600 1816.1200 2391.2400 ;
        RECT 1814.1200 2385.3200 1816.1200 2385.8000 ;
        RECT 1814.1200 2379.8800 1816.1200 2380.3600 ;
        RECT 1814.1200 2815.4800 2019.2200 2817.4800 ;
        RECT 1814.1200 2372.6900 2019.2200 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1814.1200 1913.4100 1816.1200 2358.2000 ;
        RECT 2017.2200 1913.4100 2019.2200 2358.2000 ;
        RECT 1824.8800 1913.4100 1826.4800 2358.2000 ;
        RECT 1869.8800 1913.4100 1871.4800 2358.2000 ;
        RECT 1914.8800 1913.4100 1916.4800 2358.2000 ;
        RECT 1959.8800 1913.4100 1961.4800 2358.2000 ;
        RECT 2004.8800 1913.4100 2006.4800 2358.2000 ;
      LAYER met3 ;
        RECT 2017.2200 2350.3600 2019.2200 2350.8400 ;
        RECT 2017.2200 2344.9200 2019.2200 2345.4000 ;
        RECT 2017.2200 2339.4800 2019.2200 2339.9600 ;
        RECT 2017.2200 2334.0400 2019.2200 2334.5200 ;
        RECT 2017.2200 2328.6000 2019.2200 2329.0800 ;
        RECT 2017.2200 2323.1600 2019.2200 2323.6400 ;
        RECT 2017.2200 2317.7200 2019.2200 2318.2000 ;
        RECT 2017.2200 2312.2800 2019.2200 2312.7600 ;
        RECT 2017.2200 2306.8400 2019.2200 2307.3200 ;
        RECT 2017.2200 2301.4000 2019.2200 2301.8800 ;
        RECT 2017.2200 2295.9600 2019.2200 2296.4400 ;
        RECT 2017.2200 2290.5200 2019.2200 2291.0000 ;
        RECT 2017.2200 2285.0800 2019.2200 2285.5600 ;
        RECT 2017.2200 2279.6400 2019.2200 2280.1200 ;
        RECT 2017.2200 2274.2000 2019.2200 2274.6800 ;
        RECT 2017.2200 2268.7600 2019.2200 2269.2400 ;
        RECT 2017.2200 2263.3200 2019.2200 2263.8000 ;
        RECT 2017.2200 2257.8800 2019.2200 2258.3600 ;
        RECT 2017.2200 2252.4400 2019.2200 2252.9200 ;
        RECT 2017.2200 2247.0000 2019.2200 2247.4800 ;
        RECT 2017.2200 2241.5600 2019.2200 2242.0400 ;
        RECT 2017.2200 2236.1200 2019.2200 2236.6000 ;
        RECT 2017.2200 2230.6800 2019.2200 2231.1600 ;
        RECT 2017.2200 2225.2400 2019.2200 2225.7200 ;
        RECT 2017.2200 2214.3600 2019.2200 2214.8400 ;
        RECT 2017.2200 2208.9200 2019.2200 2209.4000 ;
        RECT 2017.2200 2203.4800 2019.2200 2203.9600 ;
        RECT 2017.2200 2198.0400 2019.2200 2198.5200 ;
        RECT 2017.2200 2192.6000 2019.2200 2193.0800 ;
        RECT 2017.2200 2219.8000 2019.2200 2220.2800 ;
        RECT 2017.2200 2187.1600 2019.2200 2187.6400 ;
        RECT 2017.2200 2181.7200 2019.2200 2182.2000 ;
        RECT 2017.2200 2176.2800 2019.2200 2176.7600 ;
        RECT 2017.2200 2170.8400 2019.2200 2171.3200 ;
        RECT 2017.2200 2165.4000 2019.2200 2165.8800 ;
        RECT 2017.2200 2159.9600 2019.2200 2160.4400 ;
        RECT 2017.2200 2154.5200 2019.2200 2155.0000 ;
        RECT 2017.2200 2149.0800 2019.2200 2149.5600 ;
        RECT 2017.2200 2143.6400 2019.2200 2144.1200 ;
        RECT 2017.2200 2138.2000 2019.2200 2138.6800 ;
        RECT 1814.1200 2350.3600 1816.1200 2350.8400 ;
        RECT 1814.1200 2344.9200 1816.1200 2345.4000 ;
        RECT 1814.1200 2339.4800 1816.1200 2339.9600 ;
        RECT 1814.1200 2334.0400 1816.1200 2334.5200 ;
        RECT 1814.1200 2328.6000 1816.1200 2329.0800 ;
        RECT 1814.1200 2323.1600 1816.1200 2323.6400 ;
        RECT 1814.1200 2317.7200 1816.1200 2318.2000 ;
        RECT 1814.1200 2312.2800 1816.1200 2312.7600 ;
        RECT 1814.1200 2306.8400 1816.1200 2307.3200 ;
        RECT 1814.1200 2301.4000 1816.1200 2301.8800 ;
        RECT 1814.1200 2295.9600 1816.1200 2296.4400 ;
        RECT 1814.1200 2290.5200 1816.1200 2291.0000 ;
        RECT 1814.1200 2285.0800 1816.1200 2285.5600 ;
        RECT 1814.1200 2279.6400 1816.1200 2280.1200 ;
        RECT 1814.1200 2274.2000 1816.1200 2274.6800 ;
        RECT 1814.1200 2268.7600 1816.1200 2269.2400 ;
        RECT 1814.1200 2263.3200 1816.1200 2263.8000 ;
        RECT 1814.1200 2257.8800 1816.1200 2258.3600 ;
        RECT 1814.1200 2252.4400 1816.1200 2252.9200 ;
        RECT 1814.1200 2247.0000 1816.1200 2247.4800 ;
        RECT 1814.1200 2241.5600 1816.1200 2242.0400 ;
        RECT 1814.1200 2236.1200 1816.1200 2236.6000 ;
        RECT 1814.1200 2230.6800 1816.1200 2231.1600 ;
        RECT 1814.1200 2225.2400 1816.1200 2225.7200 ;
        RECT 1814.1200 2214.3600 1816.1200 2214.8400 ;
        RECT 1814.1200 2208.9200 1816.1200 2209.4000 ;
        RECT 1814.1200 2203.4800 1816.1200 2203.9600 ;
        RECT 1814.1200 2198.0400 1816.1200 2198.5200 ;
        RECT 1814.1200 2192.6000 1816.1200 2193.0800 ;
        RECT 1814.1200 2219.8000 1816.1200 2220.2800 ;
        RECT 1814.1200 2187.1600 1816.1200 2187.6400 ;
        RECT 1814.1200 2181.7200 1816.1200 2182.2000 ;
        RECT 1814.1200 2176.2800 1816.1200 2176.7600 ;
        RECT 1814.1200 2170.8400 1816.1200 2171.3200 ;
        RECT 1814.1200 2165.4000 1816.1200 2165.8800 ;
        RECT 1814.1200 2159.9600 1816.1200 2160.4400 ;
        RECT 1814.1200 2154.5200 1816.1200 2155.0000 ;
        RECT 1814.1200 2149.0800 1816.1200 2149.5600 ;
        RECT 1814.1200 2143.6400 1816.1200 2144.1200 ;
        RECT 1814.1200 2138.2000 1816.1200 2138.6800 ;
        RECT 2017.2200 2132.7600 2019.2200 2133.2400 ;
        RECT 2017.2200 2127.3200 2019.2200 2127.8000 ;
        RECT 2017.2200 2121.8800 2019.2200 2122.3600 ;
        RECT 2017.2200 2116.4400 2019.2200 2116.9200 ;
        RECT 2017.2200 2111.0000 2019.2200 2111.4800 ;
        RECT 2017.2200 2105.5600 2019.2200 2106.0400 ;
        RECT 2017.2200 2100.1200 2019.2200 2100.6000 ;
        RECT 2017.2200 2094.6800 2019.2200 2095.1600 ;
        RECT 2017.2200 2089.2400 2019.2200 2089.7200 ;
        RECT 2017.2200 2083.8000 2019.2200 2084.2800 ;
        RECT 2017.2200 2078.3600 2019.2200 2078.8400 ;
        RECT 2017.2200 2072.9200 2019.2200 2073.4000 ;
        RECT 2017.2200 2067.4800 2019.2200 2067.9600 ;
        RECT 2017.2200 2062.0400 2019.2200 2062.5200 ;
        RECT 2017.2200 2056.6000 2019.2200 2057.0800 ;
        RECT 2017.2200 2045.7200 2019.2200 2046.2000 ;
        RECT 2017.2200 2040.2800 2019.2200 2040.7600 ;
        RECT 2017.2200 2034.8400 2019.2200 2035.3200 ;
        RECT 2017.2200 2029.4000 2019.2200 2029.8800 ;
        RECT 2017.2200 2023.9600 2019.2200 2024.4400 ;
        RECT 2017.2200 2051.1600 2019.2200 2051.6400 ;
        RECT 2017.2200 2018.5200 2019.2200 2019.0000 ;
        RECT 2017.2200 2013.0800 2019.2200 2013.5600 ;
        RECT 2017.2200 2007.6400 2019.2200 2008.1200 ;
        RECT 2017.2200 2002.2000 2019.2200 2002.6800 ;
        RECT 2017.2200 1996.7600 2019.2200 1997.2400 ;
        RECT 2017.2200 1991.3200 2019.2200 1991.8000 ;
        RECT 2017.2200 1985.8800 2019.2200 1986.3600 ;
        RECT 2017.2200 1980.4400 2019.2200 1980.9200 ;
        RECT 2017.2200 1975.0000 2019.2200 1975.4800 ;
        RECT 2017.2200 1969.5600 2019.2200 1970.0400 ;
        RECT 2017.2200 1964.1200 2019.2200 1964.6000 ;
        RECT 2017.2200 1958.6800 2019.2200 1959.1600 ;
        RECT 2017.2200 1953.2400 2019.2200 1953.7200 ;
        RECT 2017.2200 1947.8000 2019.2200 1948.2800 ;
        RECT 2017.2200 1942.3600 2019.2200 1942.8400 ;
        RECT 2017.2200 1936.9200 2019.2200 1937.4000 ;
        RECT 2017.2200 1931.4800 2019.2200 1931.9600 ;
        RECT 2017.2200 1926.0400 2019.2200 1926.5200 ;
        RECT 2017.2200 1920.6000 2019.2200 1921.0800 ;
        RECT 1814.1200 2132.7600 1816.1200 2133.2400 ;
        RECT 1814.1200 2127.3200 1816.1200 2127.8000 ;
        RECT 1814.1200 2121.8800 1816.1200 2122.3600 ;
        RECT 1814.1200 2116.4400 1816.1200 2116.9200 ;
        RECT 1814.1200 2111.0000 1816.1200 2111.4800 ;
        RECT 1814.1200 2105.5600 1816.1200 2106.0400 ;
        RECT 1814.1200 2100.1200 1816.1200 2100.6000 ;
        RECT 1814.1200 2094.6800 1816.1200 2095.1600 ;
        RECT 1814.1200 2089.2400 1816.1200 2089.7200 ;
        RECT 1814.1200 2083.8000 1816.1200 2084.2800 ;
        RECT 1814.1200 2078.3600 1816.1200 2078.8400 ;
        RECT 1814.1200 2072.9200 1816.1200 2073.4000 ;
        RECT 1814.1200 2067.4800 1816.1200 2067.9600 ;
        RECT 1814.1200 2062.0400 1816.1200 2062.5200 ;
        RECT 1814.1200 2056.6000 1816.1200 2057.0800 ;
        RECT 1814.1200 2045.7200 1816.1200 2046.2000 ;
        RECT 1814.1200 2040.2800 1816.1200 2040.7600 ;
        RECT 1814.1200 2034.8400 1816.1200 2035.3200 ;
        RECT 1814.1200 2029.4000 1816.1200 2029.8800 ;
        RECT 1814.1200 2023.9600 1816.1200 2024.4400 ;
        RECT 1814.1200 2051.1600 1816.1200 2051.6400 ;
        RECT 1814.1200 2018.5200 1816.1200 2019.0000 ;
        RECT 1814.1200 2013.0800 1816.1200 2013.5600 ;
        RECT 1814.1200 2007.6400 1816.1200 2008.1200 ;
        RECT 1814.1200 2002.2000 1816.1200 2002.6800 ;
        RECT 1814.1200 1996.7600 1816.1200 1997.2400 ;
        RECT 1814.1200 1991.3200 1816.1200 1991.8000 ;
        RECT 1814.1200 1985.8800 1816.1200 1986.3600 ;
        RECT 1814.1200 1980.4400 1816.1200 1980.9200 ;
        RECT 1814.1200 1975.0000 1816.1200 1975.4800 ;
        RECT 1814.1200 1969.5600 1816.1200 1970.0400 ;
        RECT 1814.1200 1964.1200 1816.1200 1964.6000 ;
        RECT 1814.1200 1958.6800 1816.1200 1959.1600 ;
        RECT 1814.1200 1953.2400 1816.1200 1953.7200 ;
        RECT 1814.1200 1947.8000 1816.1200 1948.2800 ;
        RECT 1814.1200 1942.3600 1816.1200 1942.8400 ;
        RECT 1814.1200 1936.9200 1816.1200 1937.4000 ;
        RECT 1814.1200 1931.4800 1816.1200 1931.9600 ;
        RECT 1814.1200 1926.0400 1816.1200 1926.5200 ;
        RECT 1814.1200 1920.6000 1816.1200 1921.0800 ;
        RECT 1814.1200 2356.2000 2019.2200 2358.2000 ;
        RECT 1814.1200 1913.4100 2019.2200 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1814.1200 1454.1300 1816.1200 1898.9200 ;
        RECT 2017.2200 1454.1300 2019.2200 1898.9200 ;
        RECT 1824.8800 1454.1300 1826.4800 1898.9200 ;
        RECT 1869.8800 1454.1300 1871.4800 1898.9200 ;
        RECT 1914.8800 1454.1300 1916.4800 1898.9200 ;
        RECT 1959.8800 1454.1300 1961.4800 1898.9200 ;
        RECT 2004.8800 1454.1300 2006.4800 1898.9200 ;
      LAYER met3 ;
        RECT 2017.2200 1891.0800 2019.2200 1891.5600 ;
        RECT 2017.2200 1885.6400 2019.2200 1886.1200 ;
        RECT 2017.2200 1880.2000 2019.2200 1880.6800 ;
        RECT 2017.2200 1874.7600 2019.2200 1875.2400 ;
        RECT 2017.2200 1869.3200 2019.2200 1869.8000 ;
        RECT 2017.2200 1863.8800 2019.2200 1864.3600 ;
        RECT 2017.2200 1858.4400 2019.2200 1858.9200 ;
        RECT 2017.2200 1853.0000 2019.2200 1853.4800 ;
        RECT 2017.2200 1847.5600 2019.2200 1848.0400 ;
        RECT 2017.2200 1842.1200 2019.2200 1842.6000 ;
        RECT 2017.2200 1836.6800 2019.2200 1837.1600 ;
        RECT 2017.2200 1831.2400 2019.2200 1831.7200 ;
        RECT 2017.2200 1825.8000 2019.2200 1826.2800 ;
        RECT 2017.2200 1820.3600 2019.2200 1820.8400 ;
        RECT 2017.2200 1814.9200 2019.2200 1815.4000 ;
        RECT 2017.2200 1809.4800 2019.2200 1809.9600 ;
        RECT 2017.2200 1804.0400 2019.2200 1804.5200 ;
        RECT 2017.2200 1798.6000 2019.2200 1799.0800 ;
        RECT 2017.2200 1793.1600 2019.2200 1793.6400 ;
        RECT 2017.2200 1787.7200 2019.2200 1788.2000 ;
        RECT 2017.2200 1782.2800 2019.2200 1782.7600 ;
        RECT 2017.2200 1776.8400 2019.2200 1777.3200 ;
        RECT 2017.2200 1771.4000 2019.2200 1771.8800 ;
        RECT 2017.2200 1765.9600 2019.2200 1766.4400 ;
        RECT 2017.2200 1755.0800 2019.2200 1755.5600 ;
        RECT 2017.2200 1749.6400 2019.2200 1750.1200 ;
        RECT 2017.2200 1744.2000 2019.2200 1744.6800 ;
        RECT 2017.2200 1738.7600 2019.2200 1739.2400 ;
        RECT 2017.2200 1733.3200 2019.2200 1733.8000 ;
        RECT 2017.2200 1760.5200 2019.2200 1761.0000 ;
        RECT 2017.2200 1727.8800 2019.2200 1728.3600 ;
        RECT 2017.2200 1722.4400 2019.2200 1722.9200 ;
        RECT 2017.2200 1717.0000 2019.2200 1717.4800 ;
        RECT 2017.2200 1711.5600 2019.2200 1712.0400 ;
        RECT 2017.2200 1706.1200 2019.2200 1706.6000 ;
        RECT 2017.2200 1700.6800 2019.2200 1701.1600 ;
        RECT 2017.2200 1695.2400 2019.2200 1695.7200 ;
        RECT 2017.2200 1689.8000 2019.2200 1690.2800 ;
        RECT 2017.2200 1684.3600 2019.2200 1684.8400 ;
        RECT 2017.2200 1678.9200 2019.2200 1679.4000 ;
        RECT 1814.1200 1891.0800 1816.1200 1891.5600 ;
        RECT 1814.1200 1885.6400 1816.1200 1886.1200 ;
        RECT 1814.1200 1880.2000 1816.1200 1880.6800 ;
        RECT 1814.1200 1874.7600 1816.1200 1875.2400 ;
        RECT 1814.1200 1869.3200 1816.1200 1869.8000 ;
        RECT 1814.1200 1863.8800 1816.1200 1864.3600 ;
        RECT 1814.1200 1858.4400 1816.1200 1858.9200 ;
        RECT 1814.1200 1853.0000 1816.1200 1853.4800 ;
        RECT 1814.1200 1847.5600 1816.1200 1848.0400 ;
        RECT 1814.1200 1842.1200 1816.1200 1842.6000 ;
        RECT 1814.1200 1836.6800 1816.1200 1837.1600 ;
        RECT 1814.1200 1831.2400 1816.1200 1831.7200 ;
        RECT 1814.1200 1825.8000 1816.1200 1826.2800 ;
        RECT 1814.1200 1820.3600 1816.1200 1820.8400 ;
        RECT 1814.1200 1814.9200 1816.1200 1815.4000 ;
        RECT 1814.1200 1809.4800 1816.1200 1809.9600 ;
        RECT 1814.1200 1804.0400 1816.1200 1804.5200 ;
        RECT 1814.1200 1798.6000 1816.1200 1799.0800 ;
        RECT 1814.1200 1793.1600 1816.1200 1793.6400 ;
        RECT 1814.1200 1787.7200 1816.1200 1788.2000 ;
        RECT 1814.1200 1782.2800 1816.1200 1782.7600 ;
        RECT 1814.1200 1776.8400 1816.1200 1777.3200 ;
        RECT 1814.1200 1771.4000 1816.1200 1771.8800 ;
        RECT 1814.1200 1765.9600 1816.1200 1766.4400 ;
        RECT 1814.1200 1755.0800 1816.1200 1755.5600 ;
        RECT 1814.1200 1749.6400 1816.1200 1750.1200 ;
        RECT 1814.1200 1744.2000 1816.1200 1744.6800 ;
        RECT 1814.1200 1738.7600 1816.1200 1739.2400 ;
        RECT 1814.1200 1733.3200 1816.1200 1733.8000 ;
        RECT 1814.1200 1760.5200 1816.1200 1761.0000 ;
        RECT 1814.1200 1727.8800 1816.1200 1728.3600 ;
        RECT 1814.1200 1722.4400 1816.1200 1722.9200 ;
        RECT 1814.1200 1717.0000 1816.1200 1717.4800 ;
        RECT 1814.1200 1711.5600 1816.1200 1712.0400 ;
        RECT 1814.1200 1706.1200 1816.1200 1706.6000 ;
        RECT 1814.1200 1700.6800 1816.1200 1701.1600 ;
        RECT 1814.1200 1695.2400 1816.1200 1695.7200 ;
        RECT 1814.1200 1689.8000 1816.1200 1690.2800 ;
        RECT 1814.1200 1684.3600 1816.1200 1684.8400 ;
        RECT 1814.1200 1678.9200 1816.1200 1679.4000 ;
        RECT 2017.2200 1673.4800 2019.2200 1673.9600 ;
        RECT 2017.2200 1668.0400 2019.2200 1668.5200 ;
        RECT 2017.2200 1662.6000 2019.2200 1663.0800 ;
        RECT 2017.2200 1657.1600 2019.2200 1657.6400 ;
        RECT 2017.2200 1651.7200 2019.2200 1652.2000 ;
        RECT 2017.2200 1646.2800 2019.2200 1646.7600 ;
        RECT 2017.2200 1640.8400 2019.2200 1641.3200 ;
        RECT 2017.2200 1635.4000 2019.2200 1635.8800 ;
        RECT 2017.2200 1629.9600 2019.2200 1630.4400 ;
        RECT 2017.2200 1624.5200 2019.2200 1625.0000 ;
        RECT 2017.2200 1619.0800 2019.2200 1619.5600 ;
        RECT 2017.2200 1613.6400 2019.2200 1614.1200 ;
        RECT 2017.2200 1608.2000 2019.2200 1608.6800 ;
        RECT 2017.2200 1602.7600 2019.2200 1603.2400 ;
        RECT 2017.2200 1597.3200 2019.2200 1597.8000 ;
        RECT 2017.2200 1586.4400 2019.2200 1586.9200 ;
        RECT 2017.2200 1581.0000 2019.2200 1581.4800 ;
        RECT 2017.2200 1575.5600 2019.2200 1576.0400 ;
        RECT 2017.2200 1570.1200 2019.2200 1570.6000 ;
        RECT 2017.2200 1564.6800 2019.2200 1565.1600 ;
        RECT 2017.2200 1591.8800 2019.2200 1592.3600 ;
        RECT 2017.2200 1559.2400 2019.2200 1559.7200 ;
        RECT 2017.2200 1553.8000 2019.2200 1554.2800 ;
        RECT 2017.2200 1548.3600 2019.2200 1548.8400 ;
        RECT 2017.2200 1542.9200 2019.2200 1543.4000 ;
        RECT 2017.2200 1537.4800 2019.2200 1537.9600 ;
        RECT 2017.2200 1532.0400 2019.2200 1532.5200 ;
        RECT 2017.2200 1526.6000 2019.2200 1527.0800 ;
        RECT 2017.2200 1521.1600 2019.2200 1521.6400 ;
        RECT 2017.2200 1515.7200 2019.2200 1516.2000 ;
        RECT 2017.2200 1510.2800 2019.2200 1510.7600 ;
        RECT 2017.2200 1504.8400 2019.2200 1505.3200 ;
        RECT 2017.2200 1499.4000 2019.2200 1499.8800 ;
        RECT 2017.2200 1493.9600 2019.2200 1494.4400 ;
        RECT 2017.2200 1488.5200 2019.2200 1489.0000 ;
        RECT 2017.2200 1483.0800 2019.2200 1483.5600 ;
        RECT 2017.2200 1477.6400 2019.2200 1478.1200 ;
        RECT 2017.2200 1472.2000 2019.2200 1472.6800 ;
        RECT 2017.2200 1466.7600 2019.2200 1467.2400 ;
        RECT 2017.2200 1461.3200 2019.2200 1461.8000 ;
        RECT 1814.1200 1673.4800 1816.1200 1673.9600 ;
        RECT 1814.1200 1668.0400 1816.1200 1668.5200 ;
        RECT 1814.1200 1662.6000 1816.1200 1663.0800 ;
        RECT 1814.1200 1657.1600 1816.1200 1657.6400 ;
        RECT 1814.1200 1651.7200 1816.1200 1652.2000 ;
        RECT 1814.1200 1646.2800 1816.1200 1646.7600 ;
        RECT 1814.1200 1640.8400 1816.1200 1641.3200 ;
        RECT 1814.1200 1635.4000 1816.1200 1635.8800 ;
        RECT 1814.1200 1629.9600 1816.1200 1630.4400 ;
        RECT 1814.1200 1624.5200 1816.1200 1625.0000 ;
        RECT 1814.1200 1619.0800 1816.1200 1619.5600 ;
        RECT 1814.1200 1613.6400 1816.1200 1614.1200 ;
        RECT 1814.1200 1608.2000 1816.1200 1608.6800 ;
        RECT 1814.1200 1602.7600 1816.1200 1603.2400 ;
        RECT 1814.1200 1597.3200 1816.1200 1597.8000 ;
        RECT 1814.1200 1586.4400 1816.1200 1586.9200 ;
        RECT 1814.1200 1581.0000 1816.1200 1581.4800 ;
        RECT 1814.1200 1575.5600 1816.1200 1576.0400 ;
        RECT 1814.1200 1570.1200 1816.1200 1570.6000 ;
        RECT 1814.1200 1564.6800 1816.1200 1565.1600 ;
        RECT 1814.1200 1591.8800 1816.1200 1592.3600 ;
        RECT 1814.1200 1559.2400 1816.1200 1559.7200 ;
        RECT 1814.1200 1553.8000 1816.1200 1554.2800 ;
        RECT 1814.1200 1548.3600 1816.1200 1548.8400 ;
        RECT 1814.1200 1542.9200 1816.1200 1543.4000 ;
        RECT 1814.1200 1537.4800 1816.1200 1537.9600 ;
        RECT 1814.1200 1532.0400 1816.1200 1532.5200 ;
        RECT 1814.1200 1526.6000 1816.1200 1527.0800 ;
        RECT 1814.1200 1521.1600 1816.1200 1521.6400 ;
        RECT 1814.1200 1515.7200 1816.1200 1516.2000 ;
        RECT 1814.1200 1510.2800 1816.1200 1510.7600 ;
        RECT 1814.1200 1504.8400 1816.1200 1505.3200 ;
        RECT 1814.1200 1499.4000 1816.1200 1499.8800 ;
        RECT 1814.1200 1493.9600 1816.1200 1494.4400 ;
        RECT 1814.1200 1488.5200 1816.1200 1489.0000 ;
        RECT 1814.1200 1483.0800 1816.1200 1483.5600 ;
        RECT 1814.1200 1477.6400 1816.1200 1478.1200 ;
        RECT 1814.1200 1472.2000 1816.1200 1472.6800 ;
        RECT 1814.1200 1466.7600 1816.1200 1467.2400 ;
        RECT 1814.1200 1461.3200 1816.1200 1461.8000 ;
        RECT 1814.1200 1896.9200 2019.2200 1898.9200 ;
        RECT 1814.1200 1454.1300 2019.2200 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1814.1200 994.8500 1816.1200 1439.6400 ;
        RECT 2017.2200 994.8500 2019.2200 1439.6400 ;
        RECT 1824.8800 994.8500 1826.4800 1439.6400 ;
        RECT 1869.8800 994.8500 1871.4800 1439.6400 ;
        RECT 1914.8800 994.8500 1916.4800 1439.6400 ;
        RECT 1959.8800 994.8500 1961.4800 1439.6400 ;
        RECT 2004.8800 994.8500 2006.4800 1439.6400 ;
      LAYER met3 ;
        RECT 2017.2200 1431.8000 2019.2200 1432.2800 ;
        RECT 2017.2200 1426.3600 2019.2200 1426.8400 ;
        RECT 2017.2200 1420.9200 2019.2200 1421.4000 ;
        RECT 2017.2200 1415.4800 2019.2200 1415.9600 ;
        RECT 2017.2200 1410.0400 2019.2200 1410.5200 ;
        RECT 2017.2200 1404.6000 2019.2200 1405.0800 ;
        RECT 2017.2200 1399.1600 2019.2200 1399.6400 ;
        RECT 2017.2200 1393.7200 2019.2200 1394.2000 ;
        RECT 2017.2200 1388.2800 2019.2200 1388.7600 ;
        RECT 2017.2200 1382.8400 2019.2200 1383.3200 ;
        RECT 2017.2200 1377.4000 2019.2200 1377.8800 ;
        RECT 2017.2200 1371.9600 2019.2200 1372.4400 ;
        RECT 2017.2200 1366.5200 2019.2200 1367.0000 ;
        RECT 2017.2200 1361.0800 2019.2200 1361.5600 ;
        RECT 2017.2200 1355.6400 2019.2200 1356.1200 ;
        RECT 2017.2200 1350.2000 2019.2200 1350.6800 ;
        RECT 2017.2200 1344.7600 2019.2200 1345.2400 ;
        RECT 2017.2200 1339.3200 2019.2200 1339.8000 ;
        RECT 2017.2200 1333.8800 2019.2200 1334.3600 ;
        RECT 2017.2200 1328.4400 2019.2200 1328.9200 ;
        RECT 2017.2200 1323.0000 2019.2200 1323.4800 ;
        RECT 2017.2200 1317.5600 2019.2200 1318.0400 ;
        RECT 2017.2200 1312.1200 2019.2200 1312.6000 ;
        RECT 2017.2200 1306.6800 2019.2200 1307.1600 ;
        RECT 2017.2200 1295.8000 2019.2200 1296.2800 ;
        RECT 2017.2200 1290.3600 2019.2200 1290.8400 ;
        RECT 2017.2200 1284.9200 2019.2200 1285.4000 ;
        RECT 2017.2200 1279.4800 2019.2200 1279.9600 ;
        RECT 2017.2200 1274.0400 2019.2200 1274.5200 ;
        RECT 2017.2200 1301.2400 2019.2200 1301.7200 ;
        RECT 2017.2200 1268.6000 2019.2200 1269.0800 ;
        RECT 2017.2200 1263.1600 2019.2200 1263.6400 ;
        RECT 2017.2200 1257.7200 2019.2200 1258.2000 ;
        RECT 2017.2200 1252.2800 2019.2200 1252.7600 ;
        RECT 2017.2200 1246.8400 2019.2200 1247.3200 ;
        RECT 2017.2200 1241.4000 2019.2200 1241.8800 ;
        RECT 2017.2200 1235.9600 2019.2200 1236.4400 ;
        RECT 2017.2200 1230.5200 2019.2200 1231.0000 ;
        RECT 2017.2200 1225.0800 2019.2200 1225.5600 ;
        RECT 2017.2200 1219.6400 2019.2200 1220.1200 ;
        RECT 1814.1200 1431.8000 1816.1200 1432.2800 ;
        RECT 1814.1200 1426.3600 1816.1200 1426.8400 ;
        RECT 1814.1200 1420.9200 1816.1200 1421.4000 ;
        RECT 1814.1200 1415.4800 1816.1200 1415.9600 ;
        RECT 1814.1200 1410.0400 1816.1200 1410.5200 ;
        RECT 1814.1200 1404.6000 1816.1200 1405.0800 ;
        RECT 1814.1200 1399.1600 1816.1200 1399.6400 ;
        RECT 1814.1200 1393.7200 1816.1200 1394.2000 ;
        RECT 1814.1200 1388.2800 1816.1200 1388.7600 ;
        RECT 1814.1200 1382.8400 1816.1200 1383.3200 ;
        RECT 1814.1200 1377.4000 1816.1200 1377.8800 ;
        RECT 1814.1200 1371.9600 1816.1200 1372.4400 ;
        RECT 1814.1200 1366.5200 1816.1200 1367.0000 ;
        RECT 1814.1200 1361.0800 1816.1200 1361.5600 ;
        RECT 1814.1200 1355.6400 1816.1200 1356.1200 ;
        RECT 1814.1200 1350.2000 1816.1200 1350.6800 ;
        RECT 1814.1200 1344.7600 1816.1200 1345.2400 ;
        RECT 1814.1200 1339.3200 1816.1200 1339.8000 ;
        RECT 1814.1200 1333.8800 1816.1200 1334.3600 ;
        RECT 1814.1200 1328.4400 1816.1200 1328.9200 ;
        RECT 1814.1200 1323.0000 1816.1200 1323.4800 ;
        RECT 1814.1200 1317.5600 1816.1200 1318.0400 ;
        RECT 1814.1200 1312.1200 1816.1200 1312.6000 ;
        RECT 1814.1200 1306.6800 1816.1200 1307.1600 ;
        RECT 1814.1200 1295.8000 1816.1200 1296.2800 ;
        RECT 1814.1200 1290.3600 1816.1200 1290.8400 ;
        RECT 1814.1200 1284.9200 1816.1200 1285.4000 ;
        RECT 1814.1200 1279.4800 1816.1200 1279.9600 ;
        RECT 1814.1200 1274.0400 1816.1200 1274.5200 ;
        RECT 1814.1200 1301.2400 1816.1200 1301.7200 ;
        RECT 1814.1200 1268.6000 1816.1200 1269.0800 ;
        RECT 1814.1200 1263.1600 1816.1200 1263.6400 ;
        RECT 1814.1200 1257.7200 1816.1200 1258.2000 ;
        RECT 1814.1200 1252.2800 1816.1200 1252.7600 ;
        RECT 1814.1200 1246.8400 1816.1200 1247.3200 ;
        RECT 1814.1200 1241.4000 1816.1200 1241.8800 ;
        RECT 1814.1200 1235.9600 1816.1200 1236.4400 ;
        RECT 1814.1200 1230.5200 1816.1200 1231.0000 ;
        RECT 1814.1200 1225.0800 1816.1200 1225.5600 ;
        RECT 1814.1200 1219.6400 1816.1200 1220.1200 ;
        RECT 2017.2200 1214.2000 2019.2200 1214.6800 ;
        RECT 2017.2200 1208.7600 2019.2200 1209.2400 ;
        RECT 2017.2200 1203.3200 2019.2200 1203.8000 ;
        RECT 2017.2200 1197.8800 2019.2200 1198.3600 ;
        RECT 2017.2200 1192.4400 2019.2200 1192.9200 ;
        RECT 2017.2200 1187.0000 2019.2200 1187.4800 ;
        RECT 2017.2200 1181.5600 2019.2200 1182.0400 ;
        RECT 2017.2200 1176.1200 2019.2200 1176.6000 ;
        RECT 2017.2200 1170.6800 2019.2200 1171.1600 ;
        RECT 2017.2200 1165.2400 2019.2200 1165.7200 ;
        RECT 2017.2200 1159.8000 2019.2200 1160.2800 ;
        RECT 2017.2200 1154.3600 2019.2200 1154.8400 ;
        RECT 2017.2200 1148.9200 2019.2200 1149.4000 ;
        RECT 2017.2200 1143.4800 2019.2200 1143.9600 ;
        RECT 2017.2200 1138.0400 2019.2200 1138.5200 ;
        RECT 2017.2200 1127.1600 2019.2200 1127.6400 ;
        RECT 2017.2200 1121.7200 2019.2200 1122.2000 ;
        RECT 2017.2200 1116.2800 2019.2200 1116.7600 ;
        RECT 2017.2200 1110.8400 2019.2200 1111.3200 ;
        RECT 2017.2200 1105.4000 2019.2200 1105.8800 ;
        RECT 2017.2200 1132.6000 2019.2200 1133.0800 ;
        RECT 2017.2200 1099.9600 2019.2200 1100.4400 ;
        RECT 2017.2200 1094.5200 2019.2200 1095.0000 ;
        RECT 2017.2200 1089.0800 2019.2200 1089.5600 ;
        RECT 2017.2200 1083.6400 2019.2200 1084.1200 ;
        RECT 2017.2200 1078.2000 2019.2200 1078.6800 ;
        RECT 2017.2200 1072.7600 2019.2200 1073.2400 ;
        RECT 2017.2200 1067.3200 2019.2200 1067.8000 ;
        RECT 2017.2200 1061.8800 2019.2200 1062.3600 ;
        RECT 2017.2200 1056.4400 2019.2200 1056.9200 ;
        RECT 2017.2200 1051.0000 2019.2200 1051.4800 ;
        RECT 2017.2200 1045.5600 2019.2200 1046.0400 ;
        RECT 2017.2200 1040.1200 2019.2200 1040.6000 ;
        RECT 2017.2200 1034.6800 2019.2200 1035.1600 ;
        RECT 2017.2200 1029.2400 2019.2200 1029.7200 ;
        RECT 2017.2200 1023.8000 2019.2200 1024.2800 ;
        RECT 2017.2200 1018.3600 2019.2200 1018.8400 ;
        RECT 2017.2200 1012.9200 2019.2200 1013.4000 ;
        RECT 2017.2200 1007.4800 2019.2200 1007.9600 ;
        RECT 2017.2200 1002.0400 2019.2200 1002.5200 ;
        RECT 1814.1200 1214.2000 1816.1200 1214.6800 ;
        RECT 1814.1200 1208.7600 1816.1200 1209.2400 ;
        RECT 1814.1200 1203.3200 1816.1200 1203.8000 ;
        RECT 1814.1200 1197.8800 1816.1200 1198.3600 ;
        RECT 1814.1200 1192.4400 1816.1200 1192.9200 ;
        RECT 1814.1200 1187.0000 1816.1200 1187.4800 ;
        RECT 1814.1200 1181.5600 1816.1200 1182.0400 ;
        RECT 1814.1200 1176.1200 1816.1200 1176.6000 ;
        RECT 1814.1200 1170.6800 1816.1200 1171.1600 ;
        RECT 1814.1200 1165.2400 1816.1200 1165.7200 ;
        RECT 1814.1200 1159.8000 1816.1200 1160.2800 ;
        RECT 1814.1200 1154.3600 1816.1200 1154.8400 ;
        RECT 1814.1200 1148.9200 1816.1200 1149.4000 ;
        RECT 1814.1200 1143.4800 1816.1200 1143.9600 ;
        RECT 1814.1200 1138.0400 1816.1200 1138.5200 ;
        RECT 1814.1200 1127.1600 1816.1200 1127.6400 ;
        RECT 1814.1200 1121.7200 1816.1200 1122.2000 ;
        RECT 1814.1200 1116.2800 1816.1200 1116.7600 ;
        RECT 1814.1200 1110.8400 1816.1200 1111.3200 ;
        RECT 1814.1200 1105.4000 1816.1200 1105.8800 ;
        RECT 1814.1200 1132.6000 1816.1200 1133.0800 ;
        RECT 1814.1200 1099.9600 1816.1200 1100.4400 ;
        RECT 1814.1200 1094.5200 1816.1200 1095.0000 ;
        RECT 1814.1200 1089.0800 1816.1200 1089.5600 ;
        RECT 1814.1200 1083.6400 1816.1200 1084.1200 ;
        RECT 1814.1200 1078.2000 1816.1200 1078.6800 ;
        RECT 1814.1200 1072.7600 1816.1200 1073.2400 ;
        RECT 1814.1200 1067.3200 1816.1200 1067.8000 ;
        RECT 1814.1200 1061.8800 1816.1200 1062.3600 ;
        RECT 1814.1200 1056.4400 1816.1200 1056.9200 ;
        RECT 1814.1200 1051.0000 1816.1200 1051.4800 ;
        RECT 1814.1200 1045.5600 1816.1200 1046.0400 ;
        RECT 1814.1200 1040.1200 1816.1200 1040.6000 ;
        RECT 1814.1200 1034.6800 1816.1200 1035.1600 ;
        RECT 1814.1200 1029.2400 1816.1200 1029.7200 ;
        RECT 1814.1200 1023.8000 1816.1200 1024.2800 ;
        RECT 1814.1200 1018.3600 1816.1200 1018.8400 ;
        RECT 1814.1200 1012.9200 1816.1200 1013.4000 ;
        RECT 1814.1200 1007.4800 1816.1200 1007.9600 ;
        RECT 1814.1200 1002.0400 1816.1200 1002.5200 ;
        RECT 1814.1200 1437.6400 2019.2200 1439.6400 ;
        RECT 1814.1200 994.8500 2019.2200 996.8500 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1814.1200 535.5700 1816.1200 980.3600 ;
        RECT 2017.2200 535.5700 2019.2200 980.3600 ;
        RECT 1824.8800 535.5700 1826.4800 980.3600 ;
        RECT 1869.8800 535.5700 1871.4800 980.3600 ;
        RECT 1914.8800 535.5700 1916.4800 980.3600 ;
        RECT 1959.8800 535.5700 1961.4800 980.3600 ;
        RECT 2004.8800 535.5700 2006.4800 980.3600 ;
      LAYER met3 ;
        RECT 2017.2200 972.5200 2019.2200 973.0000 ;
        RECT 2017.2200 967.0800 2019.2200 967.5600 ;
        RECT 2017.2200 961.6400 2019.2200 962.1200 ;
        RECT 2017.2200 956.2000 2019.2200 956.6800 ;
        RECT 2017.2200 950.7600 2019.2200 951.2400 ;
        RECT 2017.2200 945.3200 2019.2200 945.8000 ;
        RECT 2017.2200 939.8800 2019.2200 940.3600 ;
        RECT 2017.2200 934.4400 2019.2200 934.9200 ;
        RECT 2017.2200 929.0000 2019.2200 929.4800 ;
        RECT 2017.2200 923.5600 2019.2200 924.0400 ;
        RECT 2017.2200 918.1200 2019.2200 918.6000 ;
        RECT 2017.2200 912.6800 2019.2200 913.1600 ;
        RECT 2017.2200 907.2400 2019.2200 907.7200 ;
        RECT 2017.2200 901.8000 2019.2200 902.2800 ;
        RECT 2017.2200 896.3600 2019.2200 896.8400 ;
        RECT 2017.2200 890.9200 2019.2200 891.4000 ;
        RECT 2017.2200 885.4800 2019.2200 885.9600 ;
        RECT 2017.2200 880.0400 2019.2200 880.5200 ;
        RECT 2017.2200 874.6000 2019.2200 875.0800 ;
        RECT 2017.2200 869.1600 2019.2200 869.6400 ;
        RECT 2017.2200 863.7200 2019.2200 864.2000 ;
        RECT 2017.2200 858.2800 2019.2200 858.7600 ;
        RECT 2017.2200 852.8400 2019.2200 853.3200 ;
        RECT 2017.2200 847.4000 2019.2200 847.8800 ;
        RECT 2017.2200 836.5200 2019.2200 837.0000 ;
        RECT 2017.2200 831.0800 2019.2200 831.5600 ;
        RECT 2017.2200 825.6400 2019.2200 826.1200 ;
        RECT 2017.2200 820.2000 2019.2200 820.6800 ;
        RECT 2017.2200 814.7600 2019.2200 815.2400 ;
        RECT 2017.2200 841.9600 2019.2200 842.4400 ;
        RECT 2017.2200 809.3200 2019.2200 809.8000 ;
        RECT 2017.2200 803.8800 2019.2200 804.3600 ;
        RECT 2017.2200 798.4400 2019.2200 798.9200 ;
        RECT 2017.2200 793.0000 2019.2200 793.4800 ;
        RECT 2017.2200 787.5600 2019.2200 788.0400 ;
        RECT 2017.2200 782.1200 2019.2200 782.6000 ;
        RECT 2017.2200 776.6800 2019.2200 777.1600 ;
        RECT 2017.2200 771.2400 2019.2200 771.7200 ;
        RECT 2017.2200 765.8000 2019.2200 766.2800 ;
        RECT 2017.2200 760.3600 2019.2200 760.8400 ;
        RECT 1814.1200 972.5200 1816.1200 973.0000 ;
        RECT 1814.1200 967.0800 1816.1200 967.5600 ;
        RECT 1814.1200 961.6400 1816.1200 962.1200 ;
        RECT 1814.1200 956.2000 1816.1200 956.6800 ;
        RECT 1814.1200 950.7600 1816.1200 951.2400 ;
        RECT 1814.1200 945.3200 1816.1200 945.8000 ;
        RECT 1814.1200 939.8800 1816.1200 940.3600 ;
        RECT 1814.1200 934.4400 1816.1200 934.9200 ;
        RECT 1814.1200 929.0000 1816.1200 929.4800 ;
        RECT 1814.1200 923.5600 1816.1200 924.0400 ;
        RECT 1814.1200 918.1200 1816.1200 918.6000 ;
        RECT 1814.1200 912.6800 1816.1200 913.1600 ;
        RECT 1814.1200 907.2400 1816.1200 907.7200 ;
        RECT 1814.1200 901.8000 1816.1200 902.2800 ;
        RECT 1814.1200 896.3600 1816.1200 896.8400 ;
        RECT 1814.1200 890.9200 1816.1200 891.4000 ;
        RECT 1814.1200 885.4800 1816.1200 885.9600 ;
        RECT 1814.1200 880.0400 1816.1200 880.5200 ;
        RECT 1814.1200 874.6000 1816.1200 875.0800 ;
        RECT 1814.1200 869.1600 1816.1200 869.6400 ;
        RECT 1814.1200 863.7200 1816.1200 864.2000 ;
        RECT 1814.1200 858.2800 1816.1200 858.7600 ;
        RECT 1814.1200 852.8400 1816.1200 853.3200 ;
        RECT 1814.1200 847.4000 1816.1200 847.8800 ;
        RECT 1814.1200 836.5200 1816.1200 837.0000 ;
        RECT 1814.1200 831.0800 1816.1200 831.5600 ;
        RECT 1814.1200 825.6400 1816.1200 826.1200 ;
        RECT 1814.1200 820.2000 1816.1200 820.6800 ;
        RECT 1814.1200 814.7600 1816.1200 815.2400 ;
        RECT 1814.1200 841.9600 1816.1200 842.4400 ;
        RECT 1814.1200 809.3200 1816.1200 809.8000 ;
        RECT 1814.1200 803.8800 1816.1200 804.3600 ;
        RECT 1814.1200 798.4400 1816.1200 798.9200 ;
        RECT 1814.1200 793.0000 1816.1200 793.4800 ;
        RECT 1814.1200 787.5600 1816.1200 788.0400 ;
        RECT 1814.1200 782.1200 1816.1200 782.6000 ;
        RECT 1814.1200 776.6800 1816.1200 777.1600 ;
        RECT 1814.1200 771.2400 1816.1200 771.7200 ;
        RECT 1814.1200 765.8000 1816.1200 766.2800 ;
        RECT 1814.1200 760.3600 1816.1200 760.8400 ;
        RECT 2017.2200 754.9200 2019.2200 755.4000 ;
        RECT 2017.2200 749.4800 2019.2200 749.9600 ;
        RECT 2017.2200 744.0400 2019.2200 744.5200 ;
        RECT 2017.2200 738.6000 2019.2200 739.0800 ;
        RECT 2017.2200 733.1600 2019.2200 733.6400 ;
        RECT 2017.2200 727.7200 2019.2200 728.2000 ;
        RECT 2017.2200 722.2800 2019.2200 722.7600 ;
        RECT 2017.2200 716.8400 2019.2200 717.3200 ;
        RECT 2017.2200 711.4000 2019.2200 711.8800 ;
        RECT 2017.2200 705.9600 2019.2200 706.4400 ;
        RECT 2017.2200 700.5200 2019.2200 701.0000 ;
        RECT 2017.2200 695.0800 2019.2200 695.5600 ;
        RECT 2017.2200 689.6400 2019.2200 690.1200 ;
        RECT 2017.2200 684.2000 2019.2200 684.6800 ;
        RECT 2017.2200 678.7600 2019.2200 679.2400 ;
        RECT 2017.2200 667.8800 2019.2200 668.3600 ;
        RECT 2017.2200 662.4400 2019.2200 662.9200 ;
        RECT 2017.2200 657.0000 2019.2200 657.4800 ;
        RECT 2017.2200 651.5600 2019.2200 652.0400 ;
        RECT 2017.2200 646.1200 2019.2200 646.6000 ;
        RECT 2017.2200 673.3200 2019.2200 673.8000 ;
        RECT 2017.2200 640.6800 2019.2200 641.1600 ;
        RECT 2017.2200 635.2400 2019.2200 635.7200 ;
        RECT 2017.2200 629.8000 2019.2200 630.2800 ;
        RECT 2017.2200 624.3600 2019.2200 624.8400 ;
        RECT 2017.2200 618.9200 2019.2200 619.4000 ;
        RECT 2017.2200 613.4800 2019.2200 613.9600 ;
        RECT 2017.2200 608.0400 2019.2200 608.5200 ;
        RECT 2017.2200 602.6000 2019.2200 603.0800 ;
        RECT 2017.2200 597.1600 2019.2200 597.6400 ;
        RECT 2017.2200 591.7200 2019.2200 592.2000 ;
        RECT 2017.2200 586.2800 2019.2200 586.7600 ;
        RECT 2017.2200 580.8400 2019.2200 581.3200 ;
        RECT 2017.2200 575.4000 2019.2200 575.8800 ;
        RECT 2017.2200 569.9600 2019.2200 570.4400 ;
        RECT 2017.2200 564.5200 2019.2200 565.0000 ;
        RECT 2017.2200 559.0800 2019.2200 559.5600 ;
        RECT 2017.2200 553.6400 2019.2200 554.1200 ;
        RECT 2017.2200 548.2000 2019.2200 548.6800 ;
        RECT 2017.2200 542.7600 2019.2200 543.2400 ;
        RECT 1814.1200 754.9200 1816.1200 755.4000 ;
        RECT 1814.1200 749.4800 1816.1200 749.9600 ;
        RECT 1814.1200 744.0400 1816.1200 744.5200 ;
        RECT 1814.1200 738.6000 1816.1200 739.0800 ;
        RECT 1814.1200 733.1600 1816.1200 733.6400 ;
        RECT 1814.1200 727.7200 1816.1200 728.2000 ;
        RECT 1814.1200 722.2800 1816.1200 722.7600 ;
        RECT 1814.1200 716.8400 1816.1200 717.3200 ;
        RECT 1814.1200 711.4000 1816.1200 711.8800 ;
        RECT 1814.1200 705.9600 1816.1200 706.4400 ;
        RECT 1814.1200 700.5200 1816.1200 701.0000 ;
        RECT 1814.1200 695.0800 1816.1200 695.5600 ;
        RECT 1814.1200 689.6400 1816.1200 690.1200 ;
        RECT 1814.1200 684.2000 1816.1200 684.6800 ;
        RECT 1814.1200 678.7600 1816.1200 679.2400 ;
        RECT 1814.1200 667.8800 1816.1200 668.3600 ;
        RECT 1814.1200 662.4400 1816.1200 662.9200 ;
        RECT 1814.1200 657.0000 1816.1200 657.4800 ;
        RECT 1814.1200 651.5600 1816.1200 652.0400 ;
        RECT 1814.1200 646.1200 1816.1200 646.6000 ;
        RECT 1814.1200 673.3200 1816.1200 673.8000 ;
        RECT 1814.1200 640.6800 1816.1200 641.1600 ;
        RECT 1814.1200 635.2400 1816.1200 635.7200 ;
        RECT 1814.1200 629.8000 1816.1200 630.2800 ;
        RECT 1814.1200 624.3600 1816.1200 624.8400 ;
        RECT 1814.1200 618.9200 1816.1200 619.4000 ;
        RECT 1814.1200 613.4800 1816.1200 613.9600 ;
        RECT 1814.1200 608.0400 1816.1200 608.5200 ;
        RECT 1814.1200 602.6000 1816.1200 603.0800 ;
        RECT 1814.1200 597.1600 1816.1200 597.6400 ;
        RECT 1814.1200 591.7200 1816.1200 592.2000 ;
        RECT 1814.1200 586.2800 1816.1200 586.7600 ;
        RECT 1814.1200 580.8400 1816.1200 581.3200 ;
        RECT 1814.1200 575.4000 1816.1200 575.8800 ;
        RECT 1814.1200 569.9600 1816.1200 570.4400 ;
        RECT 1814.1200 564.5200 1816.1200 565.0000 ;
        RECT 1814.1200 559.0800 1816.1200 559.5600 ;
        RECT 1814.1200 553.6400 1816.1200 554.1200 ;
        RECT 1814.1200 548.2000 1816.1200 548.6800 ;
        RECT 1814.1200 542.7600 1816.1200 543.2400 ;
        RECT 1814.1200 978.3600 2019.2200 980.3600 ;
        RECT 1814.1200 535.5700 2019.2200 537.5700 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 2034.3400 2830.6100 2036.3400 2857.5400 ;
        RECT 2237.4400 2830.6100 2239.4400 2857.5400 ;
      LAYER met3 ;
        RECT 2237.4400 2847.3200 2239.4400 2847.8000 ;
        RECT 2034.3400 2847.3200 2036.3400 2847.8000 ;
        RECT 2237.4400 2841.8800 2239.4400 2842.3600 ;
        RECT 2237.4400 2836.4400 2239.4400 2836.9200 ;
        RECT 2034.3400 2841.8800 2036.3400 2842.3600 ;
        RECT 2034.3400 2836.4400 2036.3400 2836.9200 ;
        RECT 2034.3400 2855.5400 2239.4400 2857.5400 ;
        RECT 2034.3400 2830.6100 2239.4400 2832.6100 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 534.5700 2226.7000 750.6700 ;
        RECT 2180.1000 534.5700 2181.7000 750.6700 ;
        RECT 2135.1000 534.5700 2136.7000 750.6700 ;
        RECT 2090.1000 534.5700 2091.7000 750.6700 ;
        RECT 2045.1000 534.5700 2046.7000 750.6700 ;
        RECT 2237.4400 534.5700 2240.4400 750.6700 ;
        RECT 2033.3400 534.5700 2036.3400 750.6700 ;
      LAYER met3 ;
        RECT 2237.4400 727.7200 2240.4400 728.2000 ;
        RECT 2237.4400 733.1600 2240.4400 733.6400 ;
        RECT 2225.1000 727.7200 2226.7000 728.2000 ;
        RECT 2225.1000 733.1600 2226.7000 733.6400 ;
        RECT 2237.4400 738.6000 2240.4400 739.0800 ;
        RECT 2225.1000 738.6000 2226.7000 739.0800 ;
        RECT 2237.4400 716.8400 2240.4400 717.3200 ;
        RECT 2237.4400 722.2800 2240.4400 722.7600 ;
        RECT 2225.1000 716.8400 2226.7000 717.3200 ;
        RECT 2225.1000 722.2800 2226.7000 722.7600 ;
        RECT 2237.4400 700.5200 2240.4400 701.0000 ;
        RECT 2237.4400 705.9600 2240.4400 706.4400 ;
        RECT 2225.1000 700.5200 2226.7000 701.0000 ;
        RECT 2225.1000 705.9600 2226.7000 706.4400 ;
        RECT 2237.4400 711.4000 2240.4400 711.8800 ;
        RECT 2225.1000 711.4000 2226.7000 711.8800 ;
        RECT 2180.1000 727.7200 2181.7000 728.2000 ;
        RECT 2180.1000 733.1600 2181.7000 733.6400 ;
        RECT 2180.1000 738.6000 2181.7000 739.0800 ;
        RECT 2180.1000 716.8400 2181.7000 717.3200 ;
        RECT 2180.1000 722.2800 2181.7000 722.7600 ;
        RECT 2180.1000 700.5200 2181.7000 701.0000 ;
        RECT 2180.1000 705.9600 2181.7000 706.4400 ;
        RECT 2180.1000 711.4000 2181.7000 711.8800 ;
        RECT 2237.4400 684.2000 2240.4400 684.6800 ;
        RECT 2237.4400 689.6400 2240.4400 690.1200 ;
        RECT 2237.4400 695.0800 2240.4400 695.5600 ;
        RECT 2225.1000 684.2000 2226.7000 684.6800 ;
        RECT 2225.1000 689.6400 2226.7000 690.1200 ;
        RECT 2225.1000 695.0800 2226.7000 695.5600 ;
        RECT 2237.4400 673.3200 2240.4400 673.8000 ;
        RECT 2237.4400 678.7600 2240.4400 679.2400 ;
        RECT 2225.1000 673.3200 2226.7000 673.8000 ;
        RECT 2225.1000 678.7600 2226.7000 679.2400 ;
        RECT 2237.4400 657.0000 2240.4400 657.4800 ;
        RECT 2237.4400 662.4400 2240.4400 662.9200 ;
        RECT 2237.4400 667.8800 2240.4400 668.3600 ;
        RECT 2225.1000 657.0000 2226.7000 657.4800 ;
        RECT 2225.1000 662.4400 2226.7000 662.9200 ;
        RECT 2225.1000 667.8800 2226.7000 668.3600 ;
        RECT 2237.4400 646.1200 2240.4400 646.6000 ;
        RECT 2237.4400 651.5600 2240.4400 652.0400 ;
        RECT 2225.1000 646.1200 2226.7000 646.6000 ;
        RECT 2225.1000 651.5600 2226.7000 652.0400 ;
        RECT 2180.1000 684.2000 2181.7000 684.6800 ;
        RECT 2180.1000 689.6400 2181.7000 690.1200 ;
        RECT 2180.1000 695.0800 2181.7000 695.5600 ;
        RECT 2180.1000 673.3200 2181.7000 673.8000 ;
        RECT 2180.1000 678.7600 2181.7000 679.2400 ;
        RECT 2180.1000 657.0000 2181.7000 657.4800 ;
        RECT 2180.1000 662.4400 2181.7000 662.9200 ;
        RECT 2180.1000 667.8800 2181.7000 668.3600 ;
        RECT 2180.1000 646.1200 2181.7000 646.6000 ;
        RECT 2180.1000 651.5600 2181.7000 652.0400 ;
        RECT 2135.1000 727.7200 2136.7000 728.2000 ;
        RECT 2135.1000 733.1600 2136.7000 733.6400 ;
        RECT 2135.1000 738.6000 2136.7000 739.0800 ;
        RECT 2090.1000 727.7200 2091.7000 728.2000 ;
        RECT 2090.1000 733.1600 2091.7000 733.6400 ;
        RECT 2090.1000 738.6000 2091.7000 739.0800 ;
        RECT 2135.1000 716.8400 2136.7000 717.3200 ;
        RECT 2135.1000 722.2800 2136.7000 722.7600 ;
        RECT 2135.1000 700.5200 2136.7000 701.0000 ;
        RECT 2135.1000 705.9600 2136.7000 706.4400 ;
        RECT 2135.1000 711.4000 2136.7000 711.8800 ;
        RECT 2090.1000 716.8400 2091.7000 717.3200 ;
        RECT 2090.1000 722.2800 2091.7000 722.7600 ;
        RECT 2090.1000 700.5200 2091.7000 701.0000 ;
        RECT 2090.1000 705.9600 2091.7000 706.4400 ;
        RECT 2090.1000 711.4000 2091.7000 711.8800 ;
        RECT 2045.1000 727.7200 2046.7000 728.2000 ;
        RECT 2045.1000 733.1600 2046.7000 733.6400 ;
        RECT 2033.3400 733.1600 2036.3400 733.6400 ;
        RECT 2033.3400 727.7200 2036.3400 728.2000 ;
        RECT 2033.3400 738.6000 2036.3400 739.0800 ;
        RECT 2045.1000 738.6000 2046.7000 739.0800 ;
        RECT 2045.1000 716.8400 2046.7000 717.3200 ;
        RECT 2045.1000 722.2800 2046.7000 722.7600 ;
        RECT 2033.3400 722.2800 2036.3400 722.7600 ;
        RECT 2033.3400 716.8400 2036.3400 717.3200 ;
        RECT 2045.1000 700.5200 2046.7000 701.0000 ;
        RECT 2045.1000 705.9600 2046.7000 706.4400 ;
        RECT 2033.3400 705.9600 2036.3400 706.4400 ;
        RECT 2033.3400 700.5200 2036.3400 701.0000 ;
        RECT 2033.3400 711.4000 2036.3400 711.8800 ;
        RECT 2045.1000 711.4000 2046.7000 711.8800 ;
        RECT 2135.1000 684.2000 2136.7000 684.6800 ;
        RECT 2135.1000 689.6400 2136.7000 690.1200 ;
        RECT 2135.1000 695.0800 2136.7000 695.5600 ;
        RECT 2135.1000 673.3200 2136.7000 673.8000 ;
        RECT 2135.1000 678.7600 2136.7000 679.2400 ;
        RECT 2090.1000 684.2000 2091.7000 684.6800 ;
        RECT 2090.1000 689.6400 2091.7000 690.1200 ;
        RECT 2090.1000 695.0800 2091.7000 695.5600 ;
        RECT 2090.1000 673.3200 2091.7000 673.8000 ;
        RECT 2090.1000 678.7600 2091.7000 679.2400 ;
        RECT 2135.1000 657.0000 2136.7000 657.4800 ;
        RECT 2135.1000 662.4400 2136.7000 662.9200 ;
        RECT 2135.1000 667.8800 2136.7000 668.3600 ;
        RECT 2135.1000 646.1200 2136.7000 646.6000 ;
        RECT 2135.1000 651.5600 2136.7000 652.0400 ;
        RECT 2090.1000 657.0000 2091.7000 657.4800 ;
        RECT 2090.1000 662.4400 2091.7000 662.9200 ;
        RECT 2090.1000 667.8800 2091.7000 668.3600 ;
        RECT 2090.1000 646.1200 2091.7000 646.6000 ;
        RECT 2090.1000 651.5600 2091.7000 652.0400 ;
        RECT 2045.1000 684.2000 2046.7000 684.6800 ;
        RECT 2045.1000 689.6400 2046.7000 690.1200 ;
        RECT 2045.1000 695.0800 2046.7000 695.5600 ;
        RECT 2033.3400 684.2000 2036.3400 684.6800 ;
        RECT 2033.3400 689.6400 2036.3400 690.1200 ;
        RECT 2033.3400 695.0800 2036.3400 695.5600 ;
        RECT 2045.1000 673.3200 2046.7000 673.8000 ;
        RECT 2045.1000 678.7600 2046.7000 679.2400 ;
        RECT 2033.3400 673.3200 2036.3400 673.8000 ;
        RECT 2033.3400 678.7600 2036.3400 679.2400 ;
        RECT 2045.1000 657.0000 2046.7000 657.4800 ;
        RECT 2045.1000 662.4400 2046.7000 662.9200 ;
        RECT 2045.1000 667.8800 2046.7000 668.3600 ;
        RECT 2033.3400 657.0000 2036.3400 657.4800 ;
        RECT 2033.3400 662.4400 2036.3400 662.9200 ;
        RECT 2033.3400 667.8800 2036.3400 668.3600 ;
        RECT 2045.1000 646.1200 2046.7000 646.6000 ;
        RECT 2045.1000 651.5600 2046.7000 652.0400 ;
        RECT 2033.3400 646.1200 2036.3400 646.6000 ;
        RECT 2033.3400 651.5600 2036.3400 652.0400 ;
        RECT 2237.4400 629.8000 2240.4400 630.2800 ;
        RECT 2237.4400 635.2400 2240.4400 635.7200 ;
        RECT 2237.4400 640.6800 2240.4400 641.1600 ;
        RECT 2225.1000 629.8000 2226.7000 630.2800 ;
        RECT 2225.1000 635.2400 2226.7000 635.7200 ;
        RECT 2225.1000 640.6800 2226.7000 641.1600 ;
        RECT 2237.4400 618.9200 2240.4400 619.4000 ;
        RECT 2237.4400 624.3600 2240.4400 624.8400 ;
        RECT 2225.1000 618.9200 2226.7000 619.4000 ;
        RECT 2225.1000 624.3600 2226.7000 624.8400 ;
        RECT 2237.4400 602.6000 2240.4400 603.0800 ;
        RECT 2237.4400 608.0400 2240.4400 608.5200 ;
        RECT 2237.4400 613.4800 2240.4400 613.9600 ;
        RECT 2225.1000 602.6000 2226.7000 603.0800 ;
        RECT 2225.1000 608.0400 2226.7000 608.5200 ;
        RECT 2225.1000 613.4800 2226.7000 613.9600 ;
        RECT 2237.4400 591.7200 2240.4400 592.2000 ;
        RECT 2237.4400 597.1600 2240.4400 597.6400 ;
        RECT 2225.1000 591.7200 2226.7000 592.2000 ;
        RECT 2225.1000 597.1600 2226.7000 597.6400 ;
        RECT 2180.1000 629.8000 2181.7000 630.2800 ;
        RECT 2180.1000 635.2400 2181.7000 635.7200 ;
        RECT 2180.1000 640.6800 2181.7000 641.1600 ;
        RECT 2180.1000 618.9200 2181.7000 619.4000 ;
        RECT 2180.1000 624.3600 2181.7000 624.8400 ;
        RECT 2180.1000 602.6000 2181.7000 603.0800 ;
        RECT 2180.1000 608.0400 2181.7000 608.5200 ;
        RECT 2180.1000 613.4800 2181.7000 613.9600 ;
        RECT 2180.1000 591.7200 2181.7000 592.2000 ;
        RECT 2180.1000 597.1600 2181.7000 597.6400 ;
        RECT 2237.4400 575.4000 2240.4400 575.8800 ;
        RECT 2237.4400 580.8400 2240.4400 581.3200 ;
        RECT 2237.4400 586.2800 2240.4400 586.7600 ;
        RECT 2225.1000 575.4000 2226.7000 575.8800 ;
        RECT 2225.1000 580.8400 2226.7000 581.3200 ;
        RECT 2225.1000 586.2800 2226.7000 586.7600 ;
        RECT 2237.4400 564.5200 2240.4400 565.0000 ;
        RECT 2237.4400 569.9600 2240.4400 570.4400 ;
        RECT 2225.1000 564.5200 2226.7000 565.0000 ;
        RECT 2225.1000 569.9600 2226.7000 570.4400 ;
        RECT 2237.4400 548.2000 2240.4400 548.6800 ;
        RECT 2237.4400 553.6400 2240.4400 554.1200 ;
        RECT 2237.4400 559.0800 2240.4400 559.5600 ;
        RECT 2225.1000 548.2000 2226.7000 548.6800 ;
        RECT 2225.1000 553.6400 2226.7000 554.1200 ;
        RECT 2225.1000 559.0800 2226.7000 559.5600 ;
        RECT 2237.4400 542.7600 2240.4400 543.2400 ;
        RECT 2225.1000 542.7600 2226.7000 543.2400 ;
        RECT 2180.1000 575.4000 2181.7000 575.8800 ;
        RECT 2180.1000 580.8400 2181.7000 581.3200 ;
        RECT 2180.1000 586.2800 2181.7000 586.7600 ;
        RECT 2180.1000 564.5200 2181.7000 565.0000 ;
        RECT 2180.1000 569.9600 2181.7000 570.4400 ;
        RECT 2180.1000 548.2000 2181.7000 548.6800 ;
        RECT 2180.1000 553.6400 2181.7000 554.1200 ;
        RECT 2180.1000 559.0800 2181.7000 559.5600 ;
        RECT 2180.1000 542.7600 2181.7000 543.2400 ;
        RECT 2135.1000 629.8000 2136.7000 630.2800 ;
        RECT 2135.1000 635.2400 2136.7000 635.7200 ;
        RECT 2135.1000 640.6800 2136.7000 641.1600 ;
        RECT 2135.1000 618.9200 2136.7000 619.4000 ;
        RECT 2135.1000 624.3600 2136.7000 624.8400 ;
        RECT 2090.1000 629.8000 2091.7000 630.2800 ;
        RECT 2090.1000 635.2400 2091.7000 635.7200 ;
        RECT 2090.1000 640.6800 2091.7000 641.1600 ;
        RECT 2090.1000 618.9200 2091.7000 619.4000 ;
        RECT 2090.1000 624.3600 2091.7000 624.8400 ;
        RECT 2135.1000 602.6000 2136.7000 603.0800 ;
        RECT 2135.1000 608.0400 2136.7000 608.5200 ;
        RECT 2135.1000 613.4800 2136.7000 613.9600 ;
        RECT 2135.1000 591.7200 2136.7000 592.2000 ;
        RECT 2135.1000 597.1600 2136.7000 597.6400 ;
        RECT 2090.1000 602.6000 2091.7000 603.0800 ;
        RECT 2090.1000 608.0400 2091.7000 608.5200 ;
        RECT 2090.1000 613.4800 2091.7000 613.9600 ;
        RECT 2090.1000 591.7200 2091.7000 592.2000 ;
        RECT 2090.1000 597.1600 2091.7000 597.6400 ;
        RECT 2045.1000 629.8000 2046.7000 630.2800 ;
        RECT 2045.1000 635.2400 2046.7000 635.7200 ;
        RECT 2045.1000 640.6800 2046.7000 641.1600 ;
        RECT 2033.3400 629.8000 2036.3400 630.2800 ;
        RECT 2033.3400 635.2400 2036.3400 635.7200 ;
        RECT 2033.3400 640.6800 2036.3400 641.1600 ;
        RECT 2045.1000 618.9200 2046.7000 619.4000 ;
        RECT 2045.1000 624.3600 2046.7000 624.8400 ;
        RECT 2033.3400 618.9200 2036.3400 619.4000 ;
        RECT 2033.3400 624.3600 2036.3400 624.8400 ;
        RECT 2045.1000 602.6000 2046.7000 603.0800 ;
        RECT 2045.1000 608.0400 2046.7000 608.5200 ;
        RECT 2045.1000 613.4800 2046.7000 613.9600 ;
        RECT 2033.3400 602.6000 2036.3400 603.0800 ;
        RECT 2033.3400 608.0400 2036.3400 608.5200 ;
        RECT 2033.3400 613.4800 2036.3400 613.9600 ;
        RECT 2045.1000 591.7200 2046.7000 592.2000 ;
        RECT 2045.1000 597.1600 2046.7000 597.6400 ;
        RECT 2033.3400 591.7200 2036.3400 592.2000 ;
        RECT 2033.3400 597.1600 2036.3400 597.6400 ;
        RECT 2135.1000 575.4000 2136.7000 575.8800 ;
        RECT 2135.1000 580.8400 2136.7000 581.3200 ;
        RECT 2135.1000 586.2800 2136.7000 586.7600 ;
        RECT 2135.1000 564.5200 2136.7000 565.0000 ;
        RECT 2135.1000 569.9600 2136.7000 570.4400 ;
        RECT 2090.1000 575.4000 2091.7000 575.8800 ;
        RECT 2090.1000 580.8400 2091.7000 581.3200 ;
        RECT 2090.1000 586.2800 2091.7000 586.7600 ;
        RECT 2090.1000 564.5200 2091.7000 565.0000 ;
        RECT 2090.1000 569.9600 2091.7000 570.4400 ;
        RECT 2135.1000 548.2000 2136.7000 548.6800 ;
        RECT 2135.1000 553.6400 2136.7000 554.1200 ;
        RECT 2135.1000 559.0800 2136.7000 559.5600 ;
        RECT 2135.1000 542.7600 2136.7000 543.2400 ;
        RECT 2090.1000 548.2000 2091.7000 548.6800 ;
        RECT 2090.1000 553.6400 2091.7000 554.1200 ;
        RECT 2090.1000 559.0800 2091.7000 559.5600 ;
        RECT 2090.1000 542.7600 2091.7000 543.2400 ;
        RECT 2045.1000 575.4000 2046.7000 575.8800 ;
        RECT 2045.1000 580.8400 2046.7000 581.3200 ;
        RECT 2045.1000 586.2800 2046.7000 586.7600 ;
        RECT 2033.3400 575.4000 2036.3400 575.8800 ;
        RECT 2033.3400 580.8400 2036.3400 581.3200 ;
        RECT 2033.3400 586.2800 2036.3400 586.7600 ;
        RECT 2045.1000 564.5200 2046.7000 565.0000 ;
        RECT 2045.1000 569.9600 2046.7000 570.4400 ;
        RECT 2033.3400 564.5200 2036.3400 565.0000 ;
        RECT 2033.3400 569.9600 2036.3400 570.4400 ;
        RECT 2045.1000 548.2000 2046.7000 548.6800 ;
        RECT 2045.1000 553.6400 2046.7000 554.1200 ;
        RECT 2045.1000 559.0800 2046.7000 559.5600 ;
        RECT 2033.3400 548.2000 2036.3400 548.6800 ;
        RECT 2033.3400 553.6400 2036.3400 554.1200 ;
        RECT 2033.3400 559.0800 2036.3400 559.5600 ;
        RECT 2033.3400 542.7600 2036.3400 543.2400 ;
        RECT 2045.1000 542.7600 2046.7000 543.2400 ;
        RECT 2033.3400 747.6700 2240.4400 750.6700 ;
        RECT 2033.3400 534.5700 2240.4400 537.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 304.9300 2226.7000 521.0300 ;
        RECT 2180.1000 304.9300 2181.7000 521.0300 ;
        RECT 2135.1000 304.9300 2136.7000 521.0300 ;
        RECT 2090.1000 304.9300 2091.7000 521.0300 ;
        RECT 2045.1000 304.9300 2046.7000 521.0300 ;
        RECT 2237.4400 304.9300 2240.4400 521.0300 ;
        RECT 2033.3400 304.9300 2036.3400 521.0300 ;
      LAYER met3 ;
        RECT 2237.4400 498.0800 2240.4400 498.5600 ;
        RECT 2237.4400 503.5200 2240.4400 504.0000 ;
        RECT 2225.1000 498.0800 2226.7000 498.5600 ;
        RECT 2225.1000 503.5200 2226.7000 504.0000 ;
        RECT 2237.4400 508.9600 2240.4400 509.4400 ;
        RECT 2225.1000 508.9600 2226.7000 509.4400 ;
        RECT 2237.4400 487.2000 2240.4400 487.6800 ;
        RECT 2237.4400 492.6400 2240.4400 493.1200 ;
        RECT 2225.1000 487.2000 2226.7000 487.6800 ;
        RECT 2225.1000 492.6400 2226.7000 493.1200 ;
        RECT 2237.4400 470.8800 2240.4400 471.3600 ;
        RECT 2237.4400 476.3200 2240.4400 476.8000 ;
        RECT 2225.1000 470.8800 2226.7000 471.3600 ;
        RECT 2225.1000 476.3200 2226.7000 476.8000 ;
        RECT 2237.4400 481.7600 2240.4400 482.2400 ;
        RECT 2225.1000 481.7600 2226.7000 482.2400 ;
        RECT 2180.1000 498.0800 2181.7000 498.5600 ;
        RECT 2180.1000 503.5200 2181.7000 504.0000 ;
        RECT 2180.1000 508.9600 2181.7000 509.4400 ;
        RECT 2180.1000 487.2000 2181.7000 487.6800 ;
        RECT 2180.1000 492.6400 2181.7000 493.1200 ;
        RECT 2180.1000 470.8800 2181.7000 471.3600 ;
        RECT 2180.1000 476.3200 2181.7000 476.8000 ;
        RECT 2180.1000 481.7600 2181.7000 482.2400 ;
        RECT 2237.4400 454.5600 2240.4400 455.0400 ;
        RECT 2237.4400 460.0000 2240.4400 460.4800 ;
        RECT 2237.4400 465.4400 2240.4400 465.9200 ;
        RECT 2225.1000 454.5600 2226.7000 455.0400 ;
        RECT 2225.1000 460.0000 2226.7000 460.4800 ;
        RECT 2225.1000 465.4400 2226.7000 465.9200 ;
        RECT 2237.4400 443.6800 2240.4400 444.1600 ;
        RECT 2237.4400 449.1200 2240.4400 449.6000 ;
        RECT 2225.1000 443.6800 2226.7000 444.1600 ;
        RECT 2225.1000 449.1200 2226.7000 449.6000 ;
        RECT 2237.4400 427.3600 2240.4400 427.8400 ;
        RECT 2237.4400 432.8000 2240.4400 433.2800 ;
        RECT 2237.4400 438.2400 2240.4400 438.7200 ;
        RECT 2225.1000 427.3600 2226.7000 427.8400 ;
        RECT 2225.1000 432.8000 2226.7000 433.2800 ;
        RECT 2225.1000 438.2400 2226.7000 438.7200 ;
        RECT 2237.4400 416.4800 2240.4400 416.9600 ;
        RECT 2237.4400 421.9200 2240.4400 422.4000 ;
        RECT 2225.1000 416.4800 2226.7000 416.9600 ;
        RECT 2225.1000 421.9200 2226.7000 422.4000 ;
        RECT 2180.1000 454.5600 2181.7000 455.0400 ;
        RECT 2180.1000 460.0000 2181.7000 460.4800 ;
        RECT 2180.1000 465.4400 2181.7000 465.9200 ;
        RECT 2180.1000 443.6800 2181.7000 444.1600 ;
        RECT 2180.1000 449.1200 2181.7000 449.6000 ;
        RECT 2180.1000 427.3600 2181.7000 427.8400 ;
        RECT 2180.1000 432.8000 2181.7000 433.2800 ;
        RECT 2180.1000 438.2400 2181.7000 438.7200 ;
        RECT 2180.1000 416.4800 2181.7000 416.9600 ;
        RECT 2180.1000 421.9200 2181.7000 422.4000 ;
        RECT 2135.1000 498.0800 2136.7000 498.5600 ;
        RECT 2135.1000 503.5200 2136.7000 504.0000 ;
        RECT 2135.1000 508.9600 2136.7000 509.4400 ;
        RECT 2090.1000 498.0800 2091.7000 498.5600 ;
        RECT 2090.1000 503.5200 2091.7000 504.0000 ;
        RECT 2090.1000 508.9600 2091.7000 509.4400 ;
        RECT 2135.1000 487.2000 2136.7000 487.6800 ;
        RECT 2135.1000 492.6400 2136.7000 493.1200 ;
        RECT 2135.1000 470.8800 2136.7000 471.3600 ;
        RECT 2135.1000 476.3200 2136.7000 476.8000 ;
        RECT 2135.1000 481.7600 2136.7000 482.2400 ;
        RECT 2090.1000 487.2000 2091.7000 487.6800 ;
        RECT 2090.1000 492.6400 2091.7000 493.1200 ;
        RECT 2090.1000 470.8800 2091.7000 471.3600 ;
        RECT 2090.1000 476.3200 2091.7000 476.8000 ;
        RECT 2090.1000 481.7600 2091.7000 482.2400 ;
        RECT 2045.1000 498.0800 2046.7000 498.5600 ;
        RECT 2045.1000 503.5200 2046.7000 504.0000 ;
        RECT 2033.3400 503.5200 2036.3400 504.0000 ;
        RECT 2033.3400 498.0800 2036.3400 498.5600 ;
        RECT 2033.3400 508.9600 2036.3400 509.4400 ;
        RECT 2045.1000 508.9600 2046.7000 509.4400 ;
        RECT 2045.1000 487.2000 2046.7000 487.6800 ;
        RECT 2045.1000 492.6400 2046.7000 493.1200 ;
        RECT 2033.3400 492.6400 2036.3400 493.1200 ;
        RECT 2033.3400 487.2000 2036.3400 487.6800 ;
        RECT 2045.1000 470.8800 2046.7000 471.3600 ;
        RECT 2045.1000 476.3200 2046.7000 476.8000 ;
        RECT 2033.3400 476.3200 2036.3400 476.8000 ;
        RECT 2033.3400 470.8800 2036.3400 471.3600 ;
        RECT 2033.3400 481.7600 2036.3400 482.2400 ;
        RECT 2045.1000 481.7600 2046.7000 482.2400 ;
        RECT 2135.1000 454.5600 2136.7000 455.0400 ;
        RECT 2135.1000 460.0000 2136.7000 460.4800 ;
        RECT 2135.1000 465.4400 2136.7000 465.9200 ;
        RECT 2135.1000 443.6800 2136.7000 444.1600 ;
        RECT 2135.1000 449.1200 2136.7000 449.6000 ;
        RECT 2090.1000 454.5600 2091.7000 455.0400 ;
        RECT 2090.1000 460.0000 2091.7000 460.4800 ;
        RECT 2090.1000 465.4400 2091.7000 465.9200 ;
        RECT 2090.1000 443.6800 2091.7000 444.1600 ;
        RECT 2090.1000 449.1200 2091.7000 449.6000 ;
        RECT 2135.1000 427.3600 2136.7000 427.8400 ;
        RECT 2135.1000 432.8000 2136.7000 433.2800 ;
        RECT 2135.1000 438.2400 2136.7000 438.7200 ;
        RECT 2135.1000 416.4800 2136.7000 416.9600 ;
        RECT 2135.1000 421.9200 2136.7000 422.4000 ;
        RECT 2090.1000 427.3600 2091.7000 427.8400 ;
        RECT 2090.1000 432.8000 2091.7000 433.2800 ;
        RECT 2090.1000 438.2400 2091.7000 438.7200 ;
        RECT 2090.1000 416.4800 2091.7000 416.9600 ;
        RECT 2090.1000 421.9200 2091.7000 422.4000 ;
        RECT 2045.1000 454.5600 2046.7000 455.0400 ;
        RECT 2045.1000 460.0000 2046.7000 460.4800 ;
        RECT 2045.1000 465.4400 2046.7000 465.9200 ;
        RECT 2033.3400 454.5600 2036.3400 455.0400 ;
        RECT 2033.3400 460.0000 2036.3400 460.4800 ;
        RECT 2033.3400 465.4400 2036.3400 465.9200 ;
        RECT 2045.1000 443.6800 2046.7000 444.1600 ;
        RECT 2045.1000 449.1200 2046.7000 449.6000 ;
        RECT 2033.3400 443.6800 2036.3400 444.1600 ;
        RECT 2033.3400 449.1200 2036.3400 449.6000 ;
        RECT 2045.1000 427.3600 2046.7000 427.8400 ;
        RECT 2045.1000 432.8000 2046.7000 433.2800 ;
        RECT 2045.1000 438.2400 2046.7000 438.7200 ;
        RECT 2033.3400 427.3600 2036.3400 427.8400 ;
        RECT 2033.3400 432.8000 2036.3400 433.2800 ;
        RECT 2033.3400 438.2400 2036.3400 438.7200 ;
        RECT 2045.1000 416.4800 2046.7000 416.9600 ;
        RECT 2045.1000 421.9200 2046.7000 422.4000 ;
        RECT 2033.3400 416.4800 2036.3400 416.9600 ;
        RECT 2033.3400 421.9200 2036.3400 422.4000 ;
        RECT 2237.4400 400.1600 2240.4400 400.6400 ;
        RECT 2237.4400 405.6000 2240.4400 406.0800 ;
        RECT 2237.4400 411.0400 2240.4400 411.5200 ;
        RECT 2225.1000 400.1600 2226.7000 400.6400 ;
        RECT 2225.1000 405.6000 2226.7000 406.0800 ;
        RECT 2225.1000 411.0400 2226.7000 411.5200 ;
        RECT 2237.4400 389.2800 2240.4400 389.7600 ;
        RECT 2237.4400 394.7200 2240.4400 395.2000 ;
        RECT 2225.1000 389.2800 2226.7000 389.7600 ;
        RECT 2225.1000 394.7200 2226.7000 395.2000 ;
        RECT 2237.4400 372.9600 2240.4400 373.4400 ;
        RECT 2237.4400 378.4000 2240.4400 378.8800 ;
        RECT 2237.4400 383.8400 2240.4400 384.3200 ;
        RECT 2225.1000 372.9600 2226.7000 373.4400 ;
        RECT 2225.1000 378.4000 2226.7000 378.8800 ;
        RECT 2225.1000 383.8400 2226.7000 384.3200 ;
        RECT 2237.4400 362.0800 2240.4400 362.5600 ;
        RECT 2237.4400 367.5200 2240.4400 368.0000 ;
        RECT 2225.1000 362.0800 2226.7000 362.5600 ;
        RECT 2225.1000 367.5200 2226.7000 368.0000 ;
        RECT 2180.1000 400.1600 2181.7000 400.6400 ;
        RECT 2180.1000 405.6000 2181.7000 406.0800 ;
        RECT 2180.1000 411.0400 2181.7000 411.5200 ;
        RECT 2180.1000 389.2800 2181.7000 389.7600 ;
        RECT 2180.1000 394.7200 2181.7000 395.2000 ;
        RECT 2180.1000 372.9600 2181.7000 373.4400 ;
        RECT 2180.1000 378.4000 2181.7000 378.8800 ;
        RECT 2180.1000 383.8400 2181.7000 384.3200 ;
        RECT 2180.1000 362.0800 2181.7000 362.5600 ;
        RECT 2180.1000 367.5200 2181.7000 368.0000 ;
        RECT 2237.4400 345.7600 2240.4400 346.2400 ;
        RECT 2237.4400 351.2000 2240.4400 351.6800 ;
        RECT 2237.4400 356.6400 2240.4400 357.1200 ;
        RECT 2225.1000 345.7600 2226.7000 346.2400 ;
        RECT 2225.1000 351.2000 2226.7000 351.6800 ;
        RECT 2225.1000 356.6400 2226.7000 357.1200 ;
        RECT 2237.4400 334.8800 2240.4400 335.3600 ;
        RECT 2237.4400 340.3200 2240.4400 340.8000 ;
        RECT 2225.1000 334.8800 2226.7000 335.3600 ;
        RECT 2225.1000 340.3200 2226.7000 340.8000 ;
        RECT 2237.4400 318.5600 2240.4400 319.0400 ;
        RECT 2237.4400 324.0000 2240.4400 324.4800 ;
        RECT 2237.4400 329.4400 2240.4400 329.9200 ;
        RECT 2225.1000 318.5600 2226.7000 319.0400 ;
        RECT 2225.1000 324.0000 2226.7000 324.4800 ;
        RECT 2225.1000 329.4400 2226.7000 329.9200 ;
        RECT 2237.4400 313.1200 2240.4400 313.6000 ;
        RECT 2225.1000 313.1200 2226.7000 313.6000 ;
        RECT 2180.1000 345.7600 2181.7000 346.2400 ;
        RECT 2180.1000 351.2000 2181.7000 351.6800 ;
        RECT 2180.1000 356.6400 2181.7000 357.1200 ;
        RECT 2180.1000 334.8800 2181.7000 335.3600 ;
        RECT 2180.1000 340.3200 2181.7000 340.8000 ;
        RECT 2180.1000 318.5600 2181.7000 319.0400 ;
        RECT 2180.1000 324.0000 2181.7000 324.4800 ;
        RECT 2180.1000 329.4400 2181.7000 329.9200 ;
        RECT 2180.1000 313.1200 2181.7000 313.6000 ;
        RECT 2135.1000 400.1600 2136.7000 400.6400 ;
        RECT 2135.1000 405.6000 2136.7000 406.0800 ;
        RECT 2135.1000 411.0400 2136.7000 411.5200 ;
        RECT 2135.1000 389.2800 2136.7000 389.7600 ;
        RECT 2135.1000 394.7200 2136.7000 395.2000 ;
        RECT 2090.1000 400.1600 2091.7000 400.6400 ;
        RECT 2090.1000 405.6000 2091.7000 406.0800 ;
        RECT 2090.1000 411.0400 2091.7000 411.5200 ;
        RECT 2090.1000 389.2800 2091.7000 389.7600 ;
        RECT 2090.1000 394.7200 2091.7000 395.2000 ;
        RECT 2135.1000 372.9600 2136.7000 373.4400 ;
        RECT 2135.1000 378.4000 2136.7000 378.8800 ;
        RECT 2135.1000 383.8400 2136.7000 384.3200 ;
        RECT 2135.1000 362.0800 2136.7000 362.5600 ;
        RECT 2135.1000 367.5200 2136.7000 368.0000 ;
        RECT 2090.1000 372.9600 2091.7000 373.4400 ;
        RECT 2090.1000 378.4000 2091.7000 378.8800 ;
        RECT 2090.1000 383.8400 2091.7000 384.3200 ;
        RECT 2090.1000 362.0800 2091.7000 362.5600 ;
        RECT 2090.1000 367.5200 2091.7000 368.0000 ;
        RECT 2045.1000 400.1600 2046.7000 400.6400 ;
        RECT 2045.1000 405.6000 2046.7000 406.0800 ;
        RECT 2045.1000 411.0400 2046.7000 411.5200 ;
        RECT 2033.3400 400.1600 2036.3400 400.6400 ;
        RECT 2033.3400 405.6000 2036.3400 406.0800 ;
        RECT 2033.3400 411.0400 2036.3400 411.5200 ;
        RECT 2045.1000 389.2800 2046.7000 389.7600 ;
        RECT 2045.1000 394.7200 2046.7000 395.2000 ;
        RECT 2033.3400 389.2800 2036.3400 389.7600 ;
        RECT 2033.3400 394.7200 2036.3400 395.2000 ;
        RECT 2045.1000 372.9600 2046.7000 373.4400 ;
        RECT 2045.1000 378.4000 2046.7000 378.8800 ;
        RECT 2045.1000 383.8400 2046.7000 384.3200 ;
        RECT 2033.3400 372.9600 2036.3400 373.4400 ;
        RECT 2033.3400 378.4000 2036.3400 378.8800 ;
        RECT 2033.3400 383.8400 2036.3400 384.3200 ;
        RECT 2045.1000 362.0800 2046.7000 362.5600 ;
        RECT 2045.1000 367.5200 2046.7000 368.0000 ;
        RECT 2033.3400 362.0800 2036.3400 362.5600 ;
        RECT 2033.3400 367.5200 2036.3400 368.0000 ;
        RECT 2135.1000 345.7600 2136.7000 346.2400 ;
        RECT 2135.1000 351.2000 2136.7000 351.6800 ;
        RECT 2135.1000 356.6400 2136.7000 357.1200 ;
        RECT 2135.1000 334.8800 2136.7000 335.3600 ;
        RECT 2135.1000 340.3200 2136.7000 340.8000 ;
        RECT 2090.1000 345.7600 2091.7000 346.2400 ;
        RECT 2090.1000 351.2000 2091.7000 351.6800 ;
        RECT 2090.1000 356.6400 2091.7000 357.1200 ;
        RECT 2090.1000 334.8800 2091.7000 335.3600 ;
        RECT 2090.1000 340.3200 2091.7000 340.8000 ;
        RECT 2135.1000 318.5600 2136.7000 319.0400 ;
        RECT 2135.1000 324.0000 2136.7000 324.4800 ;
        RECT 2135.1000 329.4400 2136.7000 329.9200 ;
        RECT 2135.1000 313.1200 2136.7000 313.6000 ;
        RECT 2090.1000 318.5600 2091.7000 319.0400 ;
        RECT 2090.1000 324.0000 2091.7000 324.4800 ;
        RECT 2090.1000 329.4400 2091.7000 329.9200 ;
        RECT 2090.1000 313.1200 2091.7000 313.6000 ;
        RECT 2045.1000 345.7600 2046.7000 346.2400 ;
        RECT 2045.1000 351.2000 2046.7000 351.6800 ;
        RECT 2045.1000 356.6400 2046.7000 357.1200 ;
        RECT 2033.3400 345.7600 2036.3400 346.2400 ;
        RECT 2033.3400 351.2000 2036.3400 351.6800 ;
        RECT 2033.3400 356.6400 2036.3400 357.1200 ;
        RECT 2045.1000 334.8800 2046.7000 335.3600 ;
        RECT 2045.1000 340.3200 2046.7000 340.8000 ;
        RECT 2033.3400 334.8800 2036.3400 335.3600 ;
        RECT 2033.3400 340.3200 2036.3400 340.8000 ;
        RECT 2045.1000 318.5600 2046.7000 319.0400 ;
        RECT 2045.1000 324.0000 2046.7000 324.4800 ;
        RECT 2045.1000 329.4400 2046.7000 329.9200 ;
        RECT 2033.3400 318.5600 2036.3400 319.0400 ;
        RECT 2033.3400 324.0000 2036.3400 324.4800 ;
        RECT 2033.3400 329.4400 2036.3400 329.9200 ;
        RECT 2033.3400 313.1200 2036.3400 313.6000 ;
        RECT 2045.1000 313.1200 2046.7000 313.6000 ;
        RECT 2033.3400 518.0300 2240.4400 521.0300 ;
        RECT 2033.3400 304.9300 2240.4400 307.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 75.2900 2226.7000 291.3900 ;
        RECT 2180.1000 75.2900 2181.7000 291.3900 ;
        RECT 2135.1000 75.2900 2136.7000 291.3900 ;
        RECT 2090.1000 75.2900 2091.7000 291.3900 ;
        RECT 2045.1000 75.2900 2046.7000 291.3900 ;
        RECT 2237.4400 75.2900 2240.4400 291.3900 ;
        RECT 2033.3400 75.2900 2036.3400 291.3900 ;
      LAYER met3 ;
        RECT 2237.4400 268.4400 2240.4400 268.9200 ;
        RECT 2237.4400 273.8800 2240.4400 274.3600 ;
        RECT 2225.1000 268.4400 2226.7000 268.9200 ;
        RECT 2225.1000 273.8800 2226.7000 274.3600 ;
        RECT 2237.4400 279.3200 2240.4400 279.8000 ;
        RECT 2225.1000 279.3200 2226.7000 279.8000 ;
        RECT 2237.4400 257.5600 2240.4400 258.0400 ;
        RECT 2237.4400 263.0000 2240.4400 263.4800 ;
        RECT 2225.1000 257.5600 2226.7000 258.0400 ;
        RECT 2225.1000 263.0000 2226.7000 263.4800 ;
        RECT 2237.4400 241.2400 2240.4400 241.7200 ;
        RECT 2237.4400 246.6800 2240.4400 247.1600 ;
        RECT 2225.1000 241.2400 2226.7000 241.7200 ;
        RECT 2225.1000 246.6800 2226.7000 247.1600 ;
        RECT 2237.4400 252.1200 2240.4400 252.6000 ;
        RECT 2225.1000 252.1200 2226.7000 252.6000 ;
        RECT 2180.1000 268.4400 2181.7000 268.9200 ;
        RECT 2180.1000 273.8800 2181.7000 274.3600 ;
        RECT 2180.1000 279.3200 2181.7000 279.8000 ;
        RECT 2180.1000 257.5600 2181.7000 258.0400 ;
        RECT 2180.1000 263.0000 2181.7000 263.4800 ;
        RECT 2180.1000 241.2400 2181.7000 241.7200 ;
        RECT 2180.1000 246.6800 2181.7000 247.1600 ;
        RECT 2180.1000 252.1200 2181.7000 252.6000 ;
        RECT 2237.4400 224.9200 2240.4400 225.4000 ;
        RECT 2237.4400 230.3600 2240.4400 230.8400 ;
        RECT 2237.4400 235.8000 2240.4400 236.2800 ;
        RECT 2225.1000 224.9200 2226.7000 225.4000 ;
        RECT 2225.1000 230.3600 2226.7000 230.8400 ;
        RECT 2225.1000 235.8000 2226.7000 236.2800 ;
        RECT 2237.4400 214.0400 2240.4400 214.5200 ;
        RECT 2237.4400 219.4800 2240.4400 219.9600 ;
        RECT 2225.1000 214.0400 2226.7000 214.5200 ;
        RECT 2225.1000 219.4800 2226.7000 219.9600 ;
        RECT 2237.4400 197.7200 2240.4400 198.2000 ;
        RECT 2237.4400 203.1600 2240.4400 203.6400 ;
        RECT 2237.4400 208.6000 2240.4400 209.0800 ;
        RECT 2225.1000 197.7200 2226.7000 198.2000 ;
        RECT 2225.1000 203.1600 2226.7000 203.6400 ;
        RECT 2225.1000 208.6000 2226.7000 209.0800 ;
        RECT 2237.4400 186.8400 2240.4400 187.3200 ;
        RECT 2237.4400 192.2800 2240.4400 192.7600 ;
        RECT 2225.1000 186.8400 2226.7000 187.3200 ;
        RECT 2225.1000 192.2800 2226.7000 192.7600 ;
        RECT 2180.1000 224.9200 2181.7000 225.4000 ;
        RECT 2180.1000 230.3600 2181.7000 230.8400 ;
        RECT 2180.1000 235.8000 2181.7000 236.2800 ;
        RECT 2180.1000 214.0400 2181.7000 214.5200 ;
        RECT 2180.1000 219.4800 2181.7000 219.9600 ;
        RECT 2180.1000 197.7200 2181.7000 198.2000 ;
        RECT 2180.1000 203.1600 2181.7000 203.6400 ;
        RECT 2180.1000 208.6000 2181.7000 209.0800 ;
        RECT 2180.1000 186.8400 2181.7000 187.3200 ;
        RECT 2180.1000 192.2800 2181.7000 192.7600 ;
        RECT 2135.1000 268.4400 2136.7000 268.9200 ;
        RECT 2135.1000 273.8800 2136.7000 274.3600 ;
        RECT 2135.1000 279.3200 2136.7000 279.8000 ;
        RECT 2090.1000 268.4400 2091.7000 268.9200 ;
        RECT 2090.1000 273.8800 2091.7000 274.3600 ;
        RECT 2090.1000 279.3200 2091.7000 279.8000 ;
        RECT 2135.1000 257.5600 2136.7000 258.0400 ;
        RECT 2135.1000 263.0000 2136.7000 263.4800 ;
        RECT 2135.1000 241.2400 2136.7000 241.7200 ;
        RECT 2135.1000 246.6800 2136.7000 247.1600 ;
        RECT 2135.1000 252.1200 2136.7000 252.6000 ;
        RECT 2090.1000 257.5600 2091.7000 258.0400 ;
        RECT 2090.1000 263.0000 2091.7000 263.4800 ;
        RECT 2090.1000 241.2400 2091.7000 241.7200 ;
        RECT 2090.1000 246.6800 2091.7000 247.1600 ;
        RECT 2090.1000 252.1200 2091.7000 252.6000 ;
        RECT 2045.1000 268.4400 2046.7000 268.9200 ;
        RECT 2045.1000 273.8800 2046.7000 274.3600 ;
        RECT 2033.3400 273.8800 2036.3400 274.3600 ;
        RECT 2033.3400 268.4400 2036.3400 268.9200 ;
        RECT 2033.3400 279.3200 2036.3400 279.8000 ;
        RECT 2045.1000 279.3200 2046.7000 279.8000 ;
        RECT 2045.1000 257.5600 2046.7000 258.0400 ;
        RECT 2045.1000 263.0000 2046.7000 263.4800 ;
        RECT 2033.3400 263.0000 2036.3400 263.4800 ;
        RECT 2033.3400 257.5600 2036.3400 258.0400 ;
        RECT 2045.1000 241.2400 2046.7000 241.7200 ;
        RECT 2045.1000 246.6800 2046.7000 247.1600 ;
        RECT 2033.3400 246.6800 2036.3400 247.1600 ;
        RECT 2033.3400 241.2400 2036.3400 241.7200 ;
        RECT 2033.3400 252.1200 2036.3400 252.6000 ;
        RECT 2045.1000 252.1200 2046.7000 252.6000 ;
        RECT 2135.1000 224.9200 2136.7000 225.4000 ;
        RECT 2135.1000 230.3600 2136.7000 230.8400 ;
        RECT 2135.1000 235.8000 2136.7000 236.2800 ;
        RECT 2135.1000 214.0400 2136.7000 214.5200 ;
        RECT 2135.1000 219.4800 2136.7000 219.9600 ;
        RECT 2090.1000 224.9200 2091.7000 225.4000 ;
        RECT 2090.1000 230.3600 2091.7000 230.8400 ;
        RECT 2090.1000 235.8000 2091.7000 236.2800 ;
        RECT 2090.1000 214.0400 2091.7000 214.5200 ;
        RECT 2090.1000 219.4800 2091.7000 219.9600 ;
        RECT 2135.1000 197.7200 2136.7000 198.2000 ;
        RECT 2135.1000 203.1600 2136.7000 203.6400 ;
        RECT 2135.1000 208.6000 2136.7000 209.0800 ;
        RECT 2135.1000 186.8400 2136.7000 187.3200 ;
        RECT 2135.1000 192.2800 2136.7000 192.7600 ;
        RECT 2090.1000 197.7200 2091.7000 198.2000 ;
        RECT 2090.1000 203.1600 2091.7000 203.6400 ;
        RECT 2090.1000 208.6000 2091.7000 209.0800 ;
        RECT 2090.1000 186.8400 2091.7000 187.3200 ;
        RECT 2090.1000 192.2800 2091.7000 192.7600 ;
        RECT 2045.1000 224.9200 2046.7000 225.4000 ;
        RECT 2045.1000 230.3600 2046.7000 230.8400 ;
        RECT 2045.1000 235.8000 2046.7000 236.2800 ;
        RECT 2033.3400 224.9200 2036.3400 225.4000 ;
        RECT 2033.3400 230.3600 2036.3400 230.8400 ;
        RECT 2033.3400 235.8000 2036.3400 236.2800 ;
        RECT 2045.1000 214.0400 2046.7000 214.5200 ;
        RECT 2045.1000 219.4800 2046.7000 219.9600 ;
        RECT 2033.3400 214.0400 2036.3400 214.5200 ;
        RECT 2033.3400 219.4800 2036.3400 219.9600 ;
        RECT 2045.1000 197.7200 2046.7000 198.2000 ;
        RECT 2045.1000 203.1600 2046.7000 203.6400 ;
        RECT 2045.1000 208.6000 2046.7000 209.0800 ;
        RECT 2033.3400 197.7200 2036.3400 198.2000 ;
        RECT 2033.3400 203.1600 2036.3400 203.6400 ;
        RECT 2033.3400 208.6000 2036.3400 209.0800 ;
        RECT 2045.1000 186.8400 2046.7000 187.3200 ;
        RECT 2045.1000 192.2800 2046.7000 192.7600 ;
        RECT 2033.3400 186.8400 2036.3400 187.3200 ;
        RECT 2033.3400 192.2800 2036.3400 192.7600 ;
        RECT 2237.4400 170.5200 2240.4400 171.0000 ;
        RECT 2237.4400 175.9600 2240.4400 176.4400 ;
        RECT 2237.4400 181.4000 2240.4400 181.8800 ;
        RECT 2225.1000 170.5200 2226.7000 171.0000 ;
        RECT 2225.1000 175.9600 2226.7000 176.4400 ;
        RECT 2225.1000 181.4000 2226.7000 181.8800 ;
        RECT 2237.4400 159.6400 2240.4400 160.1200 ;
        RECT 2237.4400 165.0800 2240.4400 165.5600 ;
        RECT 2225.1000 159.6400 2226.7000 160.1200 ;
        RECT 2225.1000 165.0800 2226.7000 165.5600 ;
        RECT 2237.4400 143.3200 2240.4400 143.8000 ;
        RECT 2237.4400 148.7600 2240.4400 149.2400 ;
        RECT 2237.4400 154.2000 2240.4400 154.6800 ;
        RECT 2225.1000 143.3200 2226.7000 143.8000 ;
        RECT 2225.1000 148.7600 2226.7000 149.2400 ;
        RECT 2225.1000 154.2000 2226.7000 154.6800 ;
        RECT 2237.4400 132.4400 2240.4400 132.9200 ;
        RECT 2237.4400 137.8800 2240.4400 138.3600 ;
        RECT 2225.1000 132.4400 2226.7000 132.9200 ;
        RECT 2225.1000 137.8800 2226.7000 138.3600 ;
        RECT 2180.1000 170.5200 2181.7000 171.0000 ;
        RECT 2180.1000 175.9600 2181.7000 176.4400 ;
        RECT 2180.1000 181.4000 2181.7000 181.8800 ;
        RECT 2180.1000 159.6400 2181.7000 160.1200 ;
        RECT 2180.1000 165.0800 2181.7000 165.5600 ;
        RECT 2180.1000 143.3200 2181.7000 143.8000 ;
        RECT 2180.1000 148.7600 2181.7000 149.2400 ;
        RECT 2180.1000 154.2000 2181.7000 154.6800 ;
        RECT 2180.1000 132.4400 2181.7000 132.9200 ;
        RECT 2180.1000 137.8800 2181.7000 138.3600 ;
        RECT 2237.4400 116.1200 2240.4400 116.6000 ;
        RECT 2237.4400 121.5600 2240.4400 122.0400 ;
        RECT 2237.4400 127.0000 2240.4400 127.4800 ;
        RECT 2225.1000 116.1200 2226.7000 116.6000 ;
        RECT 2225.1000 121.5600 2226.7000 122.0400 ;
        RECT 2225.1000 127.0000 2226.7000 127.4800 ;
        RECT 2237.4400 105.2400 2240.4400 105.7200 ;
        RECT 2237.4400 110.6800 2240.4400 111.1600 ;
        RECT 2225.1000 105.2400 2226.7000 105.7200 ;
        RECT 2225.1000 110.6800 2226.7000 111.1600 ;
        RECT 2237.4400 88.9200 2240.4400 89.4000 ;
        RECT 2237.4400 94.3600 2240.4400 94.8400 ;
        RECT 2237.4400 99.8000 2240.4400 100.2800 ;
        RECT 2225.1000 88.9200 2226.7000 89.4000 ;
        RECT 2225.1000 94.3600 2226.7000 94.8400 ;
        RECT 2225.1000 99.8000 2226.7000 100.2800 ;
        RECT 2237.4400 83.4800 2240.4400 83.9600 ;
        RECT 2225.1000 83.4800 2226.7000 83.9600 ;
        RECT 2180.1000 116.1200 2181.7000 116.6000 ;
        RECT 2180.1000 121.5600 2181.7000 122.0400 ;
        RECT 2180.1000 127.0000 2181.7000 127.4800 ;
        RECT 2180.1000 105.2400 2181.7000 105.7200 ;
        RECT 2180.1000 110.6800 2181.7000 111.1600 ;
        RECT 2180.1000 88.9200 2181.7000 89.4000 ;
        RECT 2180.1000 94.3600 2181.7000 94.8400 ;
        RECT 2180.1000 99.8000 2181.7000 100.2800 ;
        RECT 2180.1000 83.4800 2181.7000 83.9600 ;
        RECT 2135.1000 170.5200 2136.7000 171.0000 ;
        RECT 2135.1000 175.9600 2136.7000 176.4400 ;
        RECT 2135.1000 181.4000 2136.7000 181.8800 ;
        RECT 2135.1000 159.6400 2136.7000 160.1200 ;
        RECT 2135.1000 165.0800 2136.7000 165.5600 ;
        RECT 2090.1000 170.5200 2091.7000 171.0000 ;
        RECT 2090.1000 175.9600 2091.7000 176.4400 ;
        RECT 2090.1000 181.4000 2091.7000 181.8800 ;
        RECT 2090.1000 159.6400 2091.7000 160.1200 ;
        RECT 2090.1000 165.0800 2091.7000 165.5600 ;
        RECT 2135.1000 143.3200 2136.7000 143.8000 ;
        RECT 2135.1000 148.7600 2136.7000 149.2400 ;
        RECT 2135.1000 154.2000 2136.7000 154.6800 ;
        RECT 2135.1000 132.4400 2136.7000 132.9200 ;
        RECT 2135.1000 137.8800 2136.7000 138.3600 ;
        RECT 2090.1000 143.3200 2091.7000 143.8000 ;
        RECT 2090.1000 148.7600 2091.7000 149.2400 ;
        RECT 2090.1000 154.2000 2091.7000 154.6800 ;
        RECT 2090.1000 132.4400 2091.7000 132.9200 ;
        RECT 2090.1000 137.8800 2091.7000 138.3600 ;
        RECT 2045.1000 170.5200 2046.7000 171.0000 ;
        RECT 2045.1000 175.9600 2046.7000 176.4400 ;
        RECT 2045.1000 181.4000 2046.7000 181.8800 ;
        RECT 2033.3400 170.5200 2036.3400 171.0000 ;
        RECT 2033.3400 175.9600 2036.3400 176.4400 ;
        RECT 2033.3400 181.4000 2036.3400 181.8800 ;
        RECT 2045.1000 159.6400 2046.7000 160.1200 ;
        RECT 2045.1000 165.0800 2046.7000 165.5600 ;
        RECT 2033.3400 159.6400 2036.3400 160.1200 ;
        RECT 2033.3400 165.0800 2036.3400 165.5600 ;
        RECT 2045.1000 143.3200 2046.7000 143.8000 ;
        RECT 2045.1000 148.7600 2046.7000 149.2400 ;
        RECT 2045.1000 154.2000 2046.7000 154.6800 ;
        RECT 2033.3400 143.3200 2036.3400 143.8000 ;
        RECT 2033.3400 148.7600 2036.3400 149.2400 ;
        RECT 2033.3400 154.2000 2036.3400 154.6800 ;
        RECT 2045.1000 132.4400 2046.7000 132.9200 ;
        RECT 2045.1000 137.8800 2046.7000 138.3600 ;
        RECT 2033.3400 132.4400 2036.3400 132.9200 ;
        RECT 2033.3400 137.8800 2036.3400 138.3600 ;
        RECT 2135.1000 116.1200 2136.7000 116.6000 ;
        RECT 2135.1000 121.5600 2136.7000 122.0400 ;
        RECT 2135.1000 127.0000 2136.7000 127.4800 ;
        RECT 2135.1000 105.2400 2136.7000 105.7200 ;
        RECT 2135.1000 110.6800 2136.7000 111.1600 ;
        RECT 2090.1000 116.1200 2091.7000 116.6000 ;
        RECT 2090.1000 121.5600 2091.7000 122.0400 ;
        RECT 2090.1000 127.0000 2091.7000 127.4800 ;
        RECT 2090.1000 105.2400 2091.7000 105.7200 ;
        RECT 2090.1000 110.6800 2091.7000 111.1600 ;
        RECT 2135.1000 88.9200 2136.7000 89.4000 ;
        RECT 2135.1000 94.3600 2136.7000 94.8400 ;
        RECT 2135.1000 99.8000 2136.7000 100.2800 ;
        RECT 2135.1000 83.4800 2136.7000 83.9600 ;
        RECT 2090.1000 88.9200 2091.7000 89.4000 ;
        RECT 2090.1000 94.3600 2091.7000 94.8400 ;
        RECT 2090.1000 99.8000 2091.7000 100.2800 ;
        RECT 2090.1000 83.4800 2091.7000 83.9600 ;
        RECT 2045.1000 116.1200 2046.7000 116.6000 ;
        RECT 2045.1000 121.5600 2046.7000 122.0400 ;
        RECT 2045.1000 127.0000 2046.7000 127.4800 ;
        RECT 2033.3400 116.1200 2036.3400 116.6000 ;
        RECT 2033.3400 121.5600 2036.3400 122.0400 ;
        RECT 2033.3400 127.0000 2036.3400 127.4800 ;
        RECT 2045.1000 105.2400 2046.7000 105.7200 ;
        RECT 2045.1000 110.6800 2046.7000 111.1600 ;
        RECT 2033.3400 105.2400 2036.3400 105.7200 ;
        RECT 2033.3400 110.6800 2036.3400 111.1600 ;
        RECT 2045.1000 88.9200 2046.7000 89.4000 ;
        RECT 2045.1000 94.3600 2046.7000 94.8400 ;
        RECT 2045.1000 99.8000 2046.7000 100.2800 ;
        RECT 2033.3400 88.9200 2036.3400 89.4000 ;
        RECT 2033.3400 94.3600 2036.3400 94.8400 ;
        RECT 2033.3400 99.8000 2036.3400 100.2800 ;
        RECT 2033.3400 83.4800 2036.3400 83.9600 ;
        RECT 2045.1000 83.4800 2046.7000 83.9600 ;
        RECT 2033.3400 288.3900 2240.4400 291.3900 ;
        RECT 2033.3400 75.2900 2240.4400 78.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 2034.3400 34.6700 2036.3400 61.6000 ;
        RECT 2237.4400 34.6700 2239.4400 61.6000 ;
      LAYER met3 ;
        RECT 2237.4400 51.3800 2239.4400 51.8600 ;
        RECT 2034.3400 51.3800 2036.3400 51.8600 ;
        RECT 2237.4400 45.9400 2239.4400 46.4200 ;
        RECT 2237.4400 40.5000 2239.4400 40.9800 ;
        RECT 2034.3400 45.9400 2036.3400 46.4200 ;
        RECT 2034.3400 40.5000 2036.3400 40.9800 ;
        RECT 2034.3400 59.6000 2239.4400 61.6000 ;
        RECT 2034.3400 34.6700 2239.4400 36.6700 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 2601.3300 2226.7000 2817.4300 ;
        RECT 2180.1000 2601.3300 2181.7000 2817.4300 ;
        RECT 2135.1000 2601.3300 2136.7000 2817.4300 ;
        RECT 2090.1000 2601.3300 2091.7000 2817.4300 ;
        RECT 2045.1000 2601.3300 2046.7000 2817.4300 ;
        RECT 2237.4400 2601.3300 2240.4400 2817.4300 ;
        RECT 2033.3400 2601.3300 2036.3400 2817.4300 ;
      LAYER met3 ;
        RECT 2237.4400 2794.4800 2240.4400 2794.9600 ;
        RECT 2237.4400 2799.9200 2240.4400 2800.4000 ;
        RECT 2225.1000 2794.4800 2226.7000 2794.9600 ;
        RECT 2225.1000 2799.9200 2226.7000 2800.4000 ;
        RECT 2237.4400 2805.3600 2240.4400 2805.8400 ;
        RECT 2225.1000 2805.3600 2226.7000 2805.8400 ;
        RECT 2237.4400 2783.6000 2240.4400 2784.0800 ;
        RECT 2237.4400 2789.0400 2240.4400 2789.5200 ;
        RECT 2225.1000 2783.6000 2226.7000 2784.0800 ;
        RECT 2225.1000 2789.0400 2226.7000 2789.5200 ;
        RECT 2237.4400 2767.2800 2240.4400 2767.7600 ;
        RECT 2237.4400 2772.7200 2240.4400 2773.2000 ;
        RECT 2225.1000 2767.2800 2226.7000 2767.7600 ;
        RECT 2225.1000 2772.7200 2226.7000 2773.2000 ;
        RECT 2237.4400 2778.1600 2240.4400 2778.6400 ;
        RECT 2225.1000 2778.1600 2226.7000 2778.6400 ;
        RECT 2180.1000 2794.4800 2181.7000 2794.9600 ;
        RECT 2180.1000 2799.9200 2181.7000 2800.4000 ;
        RECT 2180.1000 2805.3600 2181.7000 2805.8400 ;
        RECT 2180.1000 2783.6000 2181.7000 2784.0800 ;
        RECT 2180.1000 2789.0400 2181.7000 2789.5200 ;
        RECT 2180.1000 2767.2800 2181.7000 2767.7600 ;
        RECT 2180.1000 2772.7200 2181.7000 2773.2000 ;
        RECT 2180.1000 2778.1600 2181.7000 2778.6400 ;
        RECT 2237.4400 2750.9600 2240.4400 2751.4400 ;
        RECT 2237.4400 2756.4000 2240.4400 2756.8800 ;
        RECT 2237.4400 2761.8400 2240.4400 2762.3200 ;
        RECT 2225.1000 2750.9600 2226.7000 2751.4400 ;
        RECT 2225.1000 2756.4000 2226.7000 2756.8800 ;
        RECT 2225.1000 2761.8400 2226.7000 2762.3200 ;
        RECT 2237.4400 2740.0800 2240.4400 2740.5600 ;
        RECT 2237.4400 2745.5200 2240.4400 2746.0000 ;
        RECT 2225.1000 2740.0800 2226.7000 2740.5600 ;
        RECT 2225.1000 2745.5200 2226.7000 2746.0000 ;
        RECT 2237.4400 2723.7600 2240.4400 2724.2400 ;
        RECT 2237.4400 2729.2000 2240.4400 2729.6800 ;
        RECT 2237.4400 2734.6400 2240.4400 2735.1200 ;
        RECT 2225.1000 2723.7600 2226.7000 2724.2400 ;
        RECT 2225.1000 2729.2000 2226.7000 2729.6800 ;
        RECT 2225.1000 2734.6400 2226.7000 2735.1200 ;
        RECT 2237.4400 2712.8800 2240.4400 2713.3600 ;
        RECT 2237.4400 2718.3200 2240.4400 2718.8000 ;
        RECT 2225.1000 2712.8800 2226.7000 2713.3600 ;
        RECT 2225.1000 2718.3200 2226.7000 2718.8000 ;
        RECT 2180.1000 2750.9600 2181.7000 2751.4400 ;
        RECT 2180.1000 2756.4000 2181.7000 2756.8800 ;
        RECT 2180.1000 2761.8400 2181.7000 2762.3200 ;
        RECT 2180.1000 2740.0800 2181.7000 2740.5600 ;
        RECT 2180.1000 2745.5200 2181.7000 2746.0000 ;
        RECT 2180.1000 2723.7600 2181.7000 2724.2400 ;
        RECT 2180.1000 2729.2000 2181.7000 2729.6800 ;
        RECT 2180.1000 2734.6400 2181.7000 2735.1200 ;
        RECT 2180.1000 2712.8800 2181.7000 2713.3600 ;
        RECT 2180.1000 2718.3200 2181.7000 2718.8000 ;
        RECT 2135.1000 2794.4800 2136.7000 2794.9600 ;
        RECT 2135.1000 2799.9200 2136.7000 2800.4000 ;
        RECT 2135.1000 2805.3600 2136.7000 2805.8400 ;
        RECT 2090.1000 2794.4800 2091.7000 2794.9600 ;
        RECT 2090.1000 2799.9200 2091.7000 2800.4000 ;
        RECT 2090.1000 2805.3600 2091.7000 2805.8400 ;
        RECT 2135.1000 2783.6000 2136.7000 2784.0800 ;
        RECT 2135.1000 2789.0400 2136.7000 2789.5200 ;
        RECT 2135.1000 2767.2800 2136.7000 2767.7600 ;
        RECT 2135.1000 2772.7200 2136.7000 2773.2000 ;
        RECT 2135.1000 2778.1600 2136.7000 2778.6400 ;
        RECT 2090.1000 2783.6000 2091.7000 2784.0800 ;
        RECT 2090.1000 2789.0400 2091.7000 2789.5200 ;
        RECT 2090.1000 2767.2800 2091.7000 2767.7600 ;
        RECT 2090.1000 2772.7200 2091.7000 2773.2000 ;
        RECT 2090.1000 2778.1600 2091.7000 2778.6400 ;
        RECT 2045.1000 2794.4800 2046.7000 2794.9600 ;
        RECT 2045.1000 2799.9200 2046.7000 2800.4000 ;
        RECT 2033.3400 2799.9200 2036.3400 2800.4000 ;
        RECT 2033.3400 2794.4800 2036.3400 2794.9600 ;
        RECT 2033.3400 2805.3600 2036.3400 2805.8400 ;
        RECT 2045.1000 2805.3600 2046.7000 2805.8400 ;
        RECT 2045.1000 2783.6000 2046.7000 2784.0800 ;
        RECT 2045.1000 2789.0400 2046.7000 2789.5200 ;
        RECT 2033.3400 2789.0400 2036.3400 2789.5200 ;
        RECT 2033.3400 2783.6000 2036.3400 2784.0800 ;
        RECT 2045.1000 2767.2800 2046.7000 2767.7600 ;
        RECT 2045.1000 2772.7200 2046.7000 2773.2000 ;
        RECT 2033.3400 2772.7200 2036.3400 2773.2000 ;
        RECT 2033.3400 2767.2800 2036.3400 2767.7600 ;
        RECT 2033.3400 2778.1600 2036.3400 2778.6400 ;
        RECT 2045.1000 2778.1600 2046.7000 2778.6400 ;
        RECT 2135.1000 2750.9600 2136.7000 2751.4400 ;
        RECT 2135.1000 2756.4000 2136.7000 2756.8800 ;
        RECT 2135.1000 2761.8400 2136.7000 2762.3200 ;
        RECT 2135.1000 2740.0800 2136.7000 2740.5600 ;
        RECT 2135.1000 2745.5200 2136.7000 2746.0000 ;
        RECT 2090.1000 2750.9600 2091.7000 2751.4400 ;
        RECT 2090.1000 2756.4000 2091.7000 2756.8800 ;
        RECT 2090.1000 2761.8400 2091.7000 2762.3200 ;
        RECT 2090.1000 2740.0800 2091.7000 2740.5600 ;
        RECT 2090.1000 2745.5200 2091.7000 2746.0000 ;
        RECT 2135.1000 2723.7600 2136.7000 2724.2400 ;
        RECT 2135.1000 2729.2000 2136.7000 2729.6800 ;
        RECT 2135.1000 2734.6400 2136.7000 2735.1200 ;
        RECT 2135.1000 2712.8800 2136.7000 2713.3600 ;
        RECT 2135.1000 2718.3200 2136.7000 2718.8000 ;
        RECT 2090.1000 2723.7600 2091.7000 2724.2400 ;
        RECT 2090.1000 2729.2000 2091.7000 2729.6800 ;
        RECT 2090.1000 2734.6400 2091.7000 2735.1200 ;
        RECT 2090.1000 2712.8800 2091.7000 2713.3600 ;
        RECT 2090.1000 2718.3200 2091.7000 2718.8000 ;
        RECT 2045.1000 2750.9600 2046.7000 2751.4400 ;
        RECT 2045.1000 2756.4000 2046.7000 2756.8800 ;
        RECT 2045.1000 2761.8400 2046.7000 2762.3200 ;
        RECT 2033.3400 2750.9600 2036.3400 2751.4400 ;
        RECT 2033.3400 2756.4000 2036.3400 2756.8800 ;
        RECT 2033.3400 2761.8400 2036.3400 2762.3200 ;
        RECT 2045.1000 2740.0800 2046.7000 2740.5600 ;
        RECT 2045.1000 2745.5200 2046.7000 2746.0000 ;
        RECT 2033.3400 2740.0800 2036.3400 2740.5600 ;
        RECT 2033.3400 2745.5200 2036.3400 2746.0000 ;
        RECT 2045.1000 2723.7600 2046.7000 2724.2400 ;
        RECT 2045.1000 2729.2000 2046.7000 2729.6800 ;
        RECT 2045.1000 2734.6400 2046.7000 2735.1200 ;
        RECT 2033.3400 2723.7600 2036.3400 2724.2400 ;
        RECT 2033.3400 2729.2000 2036.3400 2729.6800 ;
        RECT 2033.3400 2734.6400 2036.3400 2735.1200 ;
        RECT 2045.1000 2712.8800 2046.7000 2713.3600 ;
        RECT 2045.1000 2718.3200 2046.7000 2718.8000 ;
        RECT 2033.3400 2712.8800 2036.3400 2713.3600 ;
        RECT 2033.3400 2718.3200 2036.3400 2718.8000 ;
        RECT 2237.4400 2696.5600 2240.4400 2697.0400 ;
        RECT 2237.4400 2702.0000 2240.4400 2702.4800 ;
        RECT 2237.4400 2707.4400 2240.4400 2707.9200 ;
        RECT 2225.1000 2696.5600 2226.7000 2697.0400 ;
        RECT 2225.1000 2702.0000 2226.7000 2702.4800 ;
        RECT 2225.1000 2707.4400 2226.7000 2707.9200 ;
        RECT 2237.4400 2685.6800 2240.4400 2686.1600 ;
        RECT 2237.4400 2691.1200 2240.4400 2691.6000 ;
        RECT 2225.1000 2685.6800 2226.7000 2686.1600 ;
        RECT 2225.1000 2691.1200 2226.7000 2691.6000 ;
        RECT 2237.4400 2669.3600 2240.4400 2669.8400 ;
        RECT 2237.4400 2674.8000 2240.4400 2675.2800 ;
        RECT 2237.4400 2680.2400 2240.4400 2680.7200 ;
        RECT 2225.1000 2669.3600 2226.7000 2669.8400 ;
        RECT 2225.1000 2674.8000 2226.7000 2675.2800 ;
        RECT 2225.1000 2680.2400 2226.7000 2680.7200 ;
        RECT 2237.4400 2658.4800 2240.4400 2658.9600 ;
        RECT 2237.4400 2663.9200 2240.4400 2664.4000 ;
        RECT 2225.1000 2658.4800 2226.7000 2658.9600 ;
        RECT 2225.1000 2663.9200 2226.7000 2664.4000 ;
        RECT 2180.1000 2696.5600 2181.7000 2697.0400 ;
        RECT 2180.1000 2702.0000 2181.7000 2702.4800 ;
        RECT 2180.1000 2707.4400 2181.7000 2707.9200 ;
        RECT 2180.1000 2685.6800 2181.7000 2686.1600 ;
        RECT 2180.1000 2691.1200 2181.7000 2691.6000 ;
        RECT 2180.1000 2669.3600 2181.7000 2669.8400 ;
        RECT 2180.1000 2674.8000 2181.7000 2675.2800 ;
        RECT 2180.1000 2680.2400 2181.7000 2680.7200 ;
        RECT 2180.1000 2658.4800 2181.7000 2658.9600 ;
        RECT 2180.1000 2663.9200 2181.7000 2664.4000 ;
        RECT 2237.4400 2642.1600 2240.4400 2642.6400 ;
        RECT 2237.4400 2647.6000 2240.4400 2648.0800 ;
        RECT 2237.4400 2653.0400 2240.4400 2653.5200 ;
        RECT 2225.1000 2642.1600 2226.7000 2642.6400 ;
        RECT 2225.1000 2647.6000 2226.7000 2648.0800 ;
        RECT 2225.1000 2653.0400 2226.7000 2653.5200 ;
        RECT 2237.4400 2631.2800 2240.4400 2631.7600 ;
        RECT 2237.4400 2636.7200 2240.4400 2637.2000 ;
        RECT 2225.1000 2631.2800 2226.7000 2631.7600 ;
        RECT 2225.1000 2636.7200 2226.7000 2637.2000 ;
        RECT 2237.4400 2614.9600 2240.4400 2615.4400 ;
        RECT 2237.4400 2620.4000 2240.4400 2620.8800 ;
        RECT 2237.4400 2625.8400 2240.4400 2626.3200 ;
        RECT 2225.1000 2614.9600 2226.7000 2615.4400 ;
        RECT 2225.1000 2620.4000 2226.7000 2620.8800 ;
        RECT 2225.1000 2625.8400 2226.7000 2626.3200 ;
        RECT 2237.4400 2609.5200 2240.4400 2610.0000 ;
        RECT 2225.1000 2609.5200 2226.7000 2610.0000 ;
        RECT 2180.1000 2642.1600 2181.7000 2642.6400 ;
        RECT 2180.1000 2647.6000 2181.7000 2648.0800 ;
        RECT 2180.1000 2653.0400 2181.7000 2653.5200 ;
        RECT 2180.1000 2631.2800 2181.7000 2631.7600 ;
        RECT 2180.1000 2636.7200 2181.7000 2637.2000 ;
        RECT 2180.1000 2614.9600 2181.7000 2615.4400 ;
        RECT 2180.1000 2620.4000 2181.7000 2620.8800 ;
        RECT 2180.1000 2625.8400 2181.7000 2626.3200 ;
        RECT 2180.1000 2609.5200 2181.7000 2610.0000 ;
        RECT 2135.1000 2696.5600 2136.7000 2697.0400 ;
        RECT 2135.1000 2702.0000 2136.7000 2702.4800 ;
        RECT 2135.1000 2707.4400 2136.7000 2707.9200 ;
        RECT 2135.1000 2685.6800 2136.7000 2686.1600 ;
        RECT 2135.1000 2691.1200 2136.7000 2691.6000 ;
        RECT 2090.1000 2696.5600 2091.7000 2697.0400 ;
        RECT 2090.1000 2702.0000 2091.7000 2702.4800 ;
        RECT 2090.1000 2707.4400 2091.7000 2707.9200 ;
        RECT 2090.1000 2685.6800 2091.7000 2686.1600 ;
        RECT 2090.1000 2691.1200 2091.7000 2691.6000 ;
        RECT 2135.1000 2669.3600 2136.7000 2669.8400 ;
        RECT 2135.1000 2674.8000 2136.7000 2675.2800 ;
        RECT 2135.1000 2680.2400 2136.7000 2680.7200 ;
        RECT 2135.1000 2658.4800 2136.7000 2658.9600 ;
        RECT 2135.1000 2663.9200 2136.7000 2664.4000 ;
        RECT 2090.1000 2669.3600 2091.7000 2669.8400 ;
        RECT 2090.1000 2674.8000 2091.7000 2675.2800 ;
        RECT 2090.1000 2680.2400 2091.7000 2680.7200 ;
        RECT 2090.1000 2658.4800 2091.7000 2658.9600 ;
        RECT 2090.1000 2663.9200 2091.7000 2664.4000 ;
        RECT 2045.1000 2696.5600 2046.7000 2697.0400 ;
        RECT 2045.1000 2702.0000 2046.7000 2702.4800 ;
        RECT 2045.1000 2707.4400 2046.7000 2707.9200 ;
        RECT 2033.3400 2696.5600 2036.3400 2697.0400 ;
        RECT 2033.3400 2702.0000 2036.3400 2702.4800 ;
        RECT 2033.3400 2707.4400 2036.3400 2707.9200 ;
        RECT 2045.1000 2685.6800 2046.7000 2686.1600 ;
        RECT 2045.1000 2691.1200 2046.7000 2691.6000 ;
        RECT 2033.3400 2685.6800 2036.3400 2686.1600 ;
        RECT 2033.3400 2691.1200 2036.3400 2691.6000 ;
        RECT 2045.1000 2669.3600 2046.7000 2669.8400 ;
        RECT 2045.1000 2674.8000 2046.7000 2675.2800 ;
        RECT 2045.1000 2680.2400 2046.7000 2680.7200 ;
        RECT 2033.3400 2669.3600 2036.3400 2669.8400 ;
        RECT 2033.3400 2674.8000 2036.3400 2675.2800 ;
        RECT 2033.3400 2680.2400 2036.3400 2680.7200 ;
        RECT 2045.1000 2658.4800 2046.7000 2658.9600 ;
        RECT 2045.1000 2663.9200 2046.7000 2664.4000 ;
        RECT 2033.3400 2658.4800 2036.3400 2658.9600 ;
        RECT 2033.3400 2663.9200 2036.3400 2664.4000 ;
        RECT 2135.1000 2642.1600 2136.7000 2642.6400 ;
        RECT 2135.1000 2647.6000 2136.7000 2648.0800 ;
        RECT 2135.1000 2653.0400 2136.7000 2653.5200 ;
        RECT 2135.1000 2631.2800 2136.7000 2631.7600 ;
        RECT 2135.1000 2636.7200 2136.7000 2637.2000 ;
        RECT 2090.1000 2642.1600 2091.7000 2642.6400 ;
        RECT 2090.1000 2647.6000 2091.7000 2648.0800 ;
        RECT 2090.1000 2653.0400 2091.7000 2653.5200 ;
        RECT 2090.1000 2631.2800 2091.7000 2631.7600 ;
        RECT 2090.1000 2636.7200 2091.7000 2637.2000 ;
        RECT 2135.1000 2614.9600 2136.7000 2615.4400 ;
        RECT 2135.1000 2620.4000 2136.7000 2620.8800 ;
        RECT 2135.1000 2625.8400 2136.7000 2626.3200 ;
        RECT 2135.1000 2609.5200 2136.7000 2610.0000 ;
        RECT 2090.1000 2614.9600 2091.7000 2615.4400 ;
        RECT 2090.1000 2620.4000 2091.7000 2620.8800 ;
        RECT 2090.1000 2625.8400 2091.7000 2626.3200 ;
        RECT 2090.1000 2609.5200 2091.7000 2610.0000 ;
        RECT 2045.1000 2642.1600 2046.7000 2642.6400 ;
        RECT 2045.1000 2647.6000 2046.7000 2648.0800 ;
        RECT 2045.1000 2653.0400 2046.7000 2653.5200 ;
        RECT 2033.3400 2642.1600 2036.3400 2642.6400 ;
        RECT 2033.3400 2647.6000 2036.3400 2648.0800 ;
        RECT 2033.3400 2653.0400 2036.3400 2653.5200 ;
        RECT 2045.1000 2631.2800 2046.7000 2631.7600 ;
        RECT 2045.1000 2636.7200 2046.7000 2637.2000 ;
        RECT 2033.3400 2631.2800 2036.3400 2631.7600 ;
        RECT 2033.3400 2636.7200 2036.3400 2637.2000 ;
        RECT 2045.1000 2614.9600 2046.7000 2615.4400 ;
        RECT 2045.1000 2620.4000 2046.7000 2620.8800 ;
        RECT 2045.1000 2625.8400 2046.7000 2626.3200 ;
        RECT 2033.3400 2614.9600 2036.3400 2615.4400 ;
        RECT 2033.3400 2620.4000 2036.3400 2620.8800 ;
        RECT 2033.3400 2625.8400 2036.3400 2626.3200 ;
        RECT 2033.3400 2609.5200 2036.3400 2610.0000 ;
        RECT 2045.1000 2609.5200 2046.7000 2610.0000 ;
        RECT 2033.3400 2814.4300 2240.4400 2817.4300 ;
        RECT 2033.3400 2601.3300 2240.4400 2604.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 2371.6900 2226.7000 2587.7900 ;
        RECT 2180.1000 2371.6900 2181.7000 2587.7900 ;
        RECT 2135.1000 2371.6900 2136.7000 2587.7900 ;
        RECT 2090.1000 2371.6900 2091.7000 2587.7900 ;
        RECT 2045.1000 2371.6900 2046.7000 2587.7900 ;
        RECT 2237.4400 2371.6900 2240.4400 2587.7900 ;
        RECT 2033.3400 2371.6900 2036.3400 2587.7900 ;
      LAYER met3 ;
        RECT 2237.4400 2564.8400 2240.4400 2565.3200 ;
        RECT 2237.4400 2570.2800 2240.4400 2570.7600 ;
        RECT 2225.1000 2564.8400 2226.7000 2565.3200 ;
        RECT 2225.1000 2570.2800 2226.7000 2570.7600 ;
        RECT 2237.4400 2575.7200 2240.4400 2576.2000 ;
        RECT 2225.1000 2575.7200 2226.7000 2576.2000 ;
        RECT 2237.4400 2553.9600 2240.4400 2554.4400 ;
        RECT 2237.4400 2559.4000 2240.4400 2559.8800 ;
        RECT 2225.1000 2553.9600 2226.7000 2554.4400 ;
        RECT 2225.1000 2559.4000 2226.7000 2559.8800 ;
        RECT 2237.4400 2537.6400 2240.4400 2538.1200 ;
        RECT 2237.4400 2543.0800 2240.4400 2543.5600 ;
        RECT 2225.1000 2537.6400 2226.7000 2538.1200 ;
        RECT 2225.1000 2543.0800 2226.7000 2543.5600 ;
        RECT 2237.4400 2548.5200 2240.4400 2549.0000 ;
        RECT 2225.1000 2548.5200 2226.7000 2549.0000 ;
        RECT 2180.1000 2564.8400 2181.7000 2565.3200 ;
        RECT 2180.1000 2570.2800 2181.7000 2570.7600 ;
        RECT 2180.1000 2575.7200 2181.7000 2576.2000 ;
        RECT 2180.1000 2553.9600 2181.7000 2554.4400 ;
        RECT 2180.1000 2559.4000 2181.7000 2559.8800 ;
        RECT 2180.1000 2537.6400 2181.7000 2538.1200 ;
        RECT 2180.1000 2543.0800 2181.7000 2543.5600 ;
        RECT 2180.1000 2548.5200 2181.7000 2549.0000 ;
        RECT 2237.4400 2521.3200 2240.4400 2521.8000 ;
        RECT 2237.4400 2526.7600 2240.4400 2527.2400 ;
        RECT 2237.4400 2532.2000 2240.4400 2532.6800 ;
        RECT 2225.1000 2521.3200 2226.7000 2521.8000 ;
        RECT 2225.1000 2526.7600 2226.7000 2527.2400 ;
        RECT 2225.1000 2532.2000 2226.7000 2532.6800 ;
        RECT 2237.4400 2510.4400 2240.4400 2510.9200 ;
        RECT 2237.4400 2515.8800 2240.4400 2516.3600 ;
        RECT 2225.1000 2510.4400 2226.7000 2510.9200 ;
        RECT 2225.1000 2515.8800 2226.7000 2516.3600 ;
        RECT 2237.4400 2494.1200 2240.4400 2494.6000 ;
        RECT 2237.4400 2499.5600 2240.4400 2500.0400 ;
        RECT 2237.4400 2505.0000 2240.4400 2505.4800 ;
        RECT 2225.1000 2494.1200 2226.7000 2494.6000 ;
        RECT 2225.1000 2499.5600 2226.7000 2500.0400 ;
        RECT 2225.1000 2505.0000 2226.7000 2505.4800 ;
        RECT 2237.4400 2483.2400 2240.4400 2483.7200 ;
        RECT 2237.4400 2488.6800 2240.4400 2489.1600 ;
        RECT 2225.1000 2483.2400 2226.7000 2483.7200 ;
        RECT 2225.1000 2488.6800 2226.7000 2489.1600 ;
        RECT 2180.1000 2521.3200 2181.7000 2521.8000 ;
        RECT 2180.1000 2526.7600 2181.7000 2527.2400 ;
        RECT 2180.1000 2532.2000 2181.7000 2532.6800 ;
        RECT 2180.1000 2510.4400 2181.7000 2510.9200 ;
        RECT 2180.1000 2515.8800 2181.7000 2516.3600 ;
        RECT 2180.1000 2494.1200 2181.7000 2494.6000 ;
        RECT 2180.1000 2499.5600 2181.7000 2500.0400 ;
        RECT 2180.1000 2505.0000 2181.7000 2505.4800 ;
        RECT 2180.1000 2483.2400 2181.7000 2483.7200 ;
        RECT 2180.1000 2488.6800 2181.7000 2489.1600 ;
        RECT 2135.1000 2564.8400 2136.7000 2565.3200 ;
        RECT 2135.1000 2570.2800 2136.7000 2570.7600 ;
        RECT 2135.1000 2575.7200 2136.7000 2576.2000 ;
        RECT 2090.1000 2564.8400 2091.7000 2565.3200 ;
        RECT 2090.1000 2570.2800 2091.7000 2570.7600 ;
        RECT 2090.1000 2575.7200 2091.7000 2576.2000 ;
        RECT 2135.1000 2553.9600 2136.7000 2554.4400 ;
        RECT 2135.1000 2559.4000 2136.7000 2559.8800 ;
        RECT 2135.1000 2537.6400 2136.7000 2538.1200 ;
        RECT 2135.1000 2543.0800 2136.7000 2543.5600 ;
        RECT 2135.1000 2548.5200 2136.7000 2549.0000 ;
        RECT 2090.1000 2553.9600 2091.7000 2554.4400 ;
        RECT 2090.1000 2559.4000 2091.7000 2559.8800 ;
        RECT 2090.1000 2537.6400 2091.7000 2538.1200 ;
        RECT 2090.1000 2543.0800 2091.7000 2543.5600 ;
        RECT 2090.1000 2548.5200 2091.7000 2549.0000 ;
        RECT 2045.1000 2564.8400 2046.7000 2565.3200 ;
        RECT 2045.1000 2570.2800 2046.7000 2570.7600 ;
        RECT 2033.3400 2570.2800 2036.3400 2570.7600 ;
        RECT 2033.3400 2564.8400 2036.3400 2565.3200 ;
        RECT 2033.3400 2575.7200 2036.3400 2576.2000 ;
        RECT 2045.1000 2575.7200 2046.7000 2576.2000 ;
        RECT 2045.1000 2553.9600 2046.7000 2554.4400 ;
        RECT 2045.1000 2559.4000 2046.7000 2559.8800 ;
        RECT 2033.3400 2559.4000 2036.3400 2559.8800 ;
        RECT 2033.3400 2553.9600 2036.3400 2554.4400 ;
        RECT 2045.1000 2537.6400 2046.7000 2538.1200 ;
        RECT 2045.1000 2543.0800 2046.7000 2543.5600 ;
        RECT 2033.3400 2543.0800 2036.3400 2543.5600 ;
        RECT 2033.3400 2537.6400 2036.3400 2538.1200 ;
        RECT 2033.3400 2548.5200 2036.3400 2549.0000 ;
        RECT 2045.1000 2548.5200 2046.7000 2549.0000 ;
        RECT 2135.1000 2521.3200 2136.7000 2521.8000 ;
        RECT 2135.1000 2526.7600 2136.7000 2527.2400 ;
        RECT 2135.1000 2532.2000 2136.7000 2532.6800 ;
        RECT 2135.1000 2510.4400 2136.7000 2510.9200 ;
        RECT 2135.1000 2515.8800 2136.7000 2516.3600 ;
        RECT 2090.1000 2521.3200 2091.7000 2521.8000 ;
        RECT 2090.1000 2526.7600 2091.7000 2527.2400 ;
        RECT 2090.1000 2532.2000 2091.7000 2532.6800 ;
        RECT 2090.1000 2510.4400 2091.7000 2510.9200 ;
        RECT 2090.1000 2515.8800 2091.7000 2516.3600 ;
        RECT 2135.1000 2494.1200 2136.7000 2494.6000 ;
        RECT 2135.1000 2499.5600 2136.7000 2500.0400 ;
        RECT 2135.1000 2505.0000 2136.7000 2505.4800 ;
        RECT 2135.1000 2483.2400 2136.7000 2483.7200 ;
        RECT 2135.1000 2488.6800 2136.7000 2489.1600 ;
        RECT 2090.1000 2494.1200 2091.7000 2494.6000 ;
        RECT 2090.1000 2499.5600 2091.7000 2500.0400 ;
        RECT 2090.1000 2505.0000 2091.7000 2505.4800 ;
        RECT 2090.1000 2483.2400 2091.7000 2483.7200 ;
        RECT 2090.1000 2488.6800 2091.7000 2489.1600 ;
        RECT 2045.1000 2521.3200 2046.7000 2521.8000 ;
        RECT 2045.1000 2526.7600 2046.7000 2527.2400 ;
        RECT 2045.1000 2532.2000 2046.7000 2532.6800 ;
        RECT 2033.3400 2521.3200 2036.3400 2521.8000 ;
        RECT 2033.3400 2526.7600 2036.3400 2527.2400 ;
        RECT 2033.3400 2532.2000 2036.3400 2532.6800 ;
        RECT 2045.1000 2510.4400 2046.7000 2510.9200 ;
        RECT 2045.1000 2515.8800 2046.7000 2516.3600 ;
        RECT 2033.3400 2510.4400 2036.3400 2510.9200 ;
        RECT 2033.3400 2515.8800 2036.3400 2516.3600 ;
        RECT 2045.1000 2494.1200 2046.7000 2494.6000 ;
        RECT 2045.1000 2499.5600 2046.7000 2500.0400 ;
        RECT 2045.1000 2505.0000 2046.7000 2505.4800 ;
        RECT 2033.3400 2494.1200 2036.3400 2494.6000 ;
        RECT 2033.3400 2499.5600 2036.3400 2500.0400 ;
        RECT 2033.3400 2505.0000 2036.3400 2505.4800 ;
        RECT 2045.1000 2483.2400 2046.7000 2483.7200 ;
        RECT 2045.1000 2488.6800 2046.7000 2489.1600 ;
        RECT 2033.3400 2483.2400 2036.3400 2483.7200 ;
        RECT 2033.3400 2488.6800 2036.3400 2489.1600 ;
        RECT 2237.4400 2466.9200 2240.4400 2467.4000 ;
        RECT 2237.4400 2472.3600 2240.4400 2472.8400 ;
        RECT 2237.4400 2477.8000 2240.4400 2478.2800 ;
        RECT 2225.1000 2466.9200 2226.7000 2467.4000 ;
        RECT 2225.1000 2472.3600 2226.7000 2472.8400 ;
        RECT 2225.1000 2477.8000 2226.7000 2478.2800 ;
        RECT 2237.4400 2456.0400 2240.4400 2456.5200 ;
        RECT 2237.4400 2461.4800 2240.4400 2461.9600 ;
        RECT 2225.1000 2456.0400 2226.7000 2456.5200 ;
        RECT 2225.1000 2461.4800 2226.7000 2461.9600 ;
        RECT 2237.4400 2439.7200 2240.4400 2440.2000 ;
        RECT 2237.4400 2445.1600 2240.4400 2445.6400 ;
        RECT 2237.4400 2450.6000 2240.4400 2451.0800 ;
        RECT 2225.1000 2439.7200 2226.7000 2440.2000 ;
        RECT 2225.1000 2445.1600 2226.7000 2445.6400 ;
        RECT 2225.1000 2450.6000 2226.7000 2451.0800 ;
        RECT 2237.4400 2428.8400 2240.4400 2429.3200 ;
        RECT 2237.4400 2434.2800 2240.4400 2434.7600 ;
        RECT 2225.1000 2428.8400 2226.7000 2429.3200 ;
        RECT 2225.1000 2434.2800 2226.7000 2434.7600 ;
        RECT 2180.1000 2466.9200 2181.7000 2467.4000 ;
        RECT 2180.1000 2472.3600 2181.7000 2472.8400 ;
        RECT 2180.1000 2477.8000 2181.7000 2478.2800 ;
        RECT 2180.1000 2456.0400 2181.7000 2456.5200 ;
        RECT 2180.1000 2461.4800 2181.7000 2461.9600 ;
        RECT 2180.1000 2439.7200 2181.7000 2440.2000 ;
        RECT 2180.1000 2445.1600 2181.7000 2445.6400 ;
        RECT 2180.1000 2450.6000 2181.7000 2451.0800 ;
        RECT 2180.1000 2428.8400 2181.7000 2429.3200 ;
        RECT 2180.1000 2434.2800 2181.7000 2434.7600 ;
        RECT 2237.4400 2412.5200 2240.4400 2413.0000 ;
        RECT 2237.4400 2417.9600 2240.4400 2418.4400 ;
        RECT 2237.4400 2423.4000 2240.4400 2423.8800 ;
        RECT 2225.1000 2412.5200 2226.7000 2413.0000 ;
        RECT 2225.1000 2417.9600 2226.7000 2418.4400 ;
        RECT 2225.1000 2423.4000 2226.7000 2423.8800 ;
        RECT 2237.4400 2401.6400 2240.4400 2402.1200 ;
        RECT 2237.4400 2407.0800 2240.4400 2407.5600 ;
        RECT 2225.1000 2401.6400 2226.7000 2402.1200 ;
        RECT 2225.1000 2407.0800 2226.7000 2407.5600 ;
        RECT 2237.4400 2385.3200 2240.4400 2385.8000 ;
        RECT 2237.4400 2390.7600 2240.4400 2391.2400 ;
        RECT 2237.4400 2396.2000 2240.4400 2396.6800 ;
        RECT 2225.1000 2385.3200 2226.7000 2385.8000 ;
        RECT 2225.1000 2390.7600 2226.7000 2391.2400 ;
        RECT 2225.1000 2396.2000 2226.7000 2396.6800 ;
        RECT 2237.4400 2379.8800 2240.4400 2380.3600 ;
        RECT 2225.1000 2379.8800 2226.7000 2380.3600 ;
        RECT 2180.1000 2412.5200 2181.7000 2413.0000 ;
        RECT 2180.1000 2417.9600 2181.7000 2418.4400 ;
        RECT 2180.1000 2423.4000 2181.7000 2423.8800 ;
        RECT 2180.1000 2401.6400 2181.7000 2402.1200 ;
        RECT 2180.1000 2407.0800 2181.7000 2407.5600 ;
        RECT 2180.1000 2385.3200 2181.7000 2385.8000 ;
        RECT 2180.1000 2390.7600 2181.7000 2391.2400 ;
        RECT 2180.1000 2396.2000 2181.7000 2396.6800 ;
        RECT 2180.1000 2379.8800 2181.7000 2380.3600 ;
        RECT 2135.1000 2466.9200 2136.7000 2467.4000 ;
        RECT 2135.1000 2472.3600 2136.7000 2472.8400 ;
        RECT 2135.1000 2477.8000 2136.7000 2478.2800 ;
        RECT 2135.1000 2456.0400 2136.7000 2456.5200 ;
        RECT 2135.1000 2461.4800 2136.7000 2461.9600 ;
        RECT 2090.1000 2466.9200 2091.7000 2467.4000 ;
        RECT 2090.1000 2472.3600 2091.7000 2472.8400 ;
        RECT 2090.1000 2477.8000 2091.7000 2478.2800 ;
        RECT 2090.1000 2456.0400 2091.7000 2456.5200 ;
        RECT 2090.1000 2461.4800 2091.7000 2461.9600 ;
        RECT 2135.1000 2439.7200 2136.7000 2440.2000 ;
        RECT 2135.1000 2445.1600 2136.7000 2445.6400 ;
        RECT 2135.1000 2450.6000 2136.7000 2451.0800 ;
        RECT 2135.1000 2428.8400 2136.7000 2429.3200 ;
        RECT 2135.1000 2434.2800 2136.7000 2434.7600 ;
        RECT 2090.1000 2439.7200 2091.7000 2440.2000 ;
        RECT 2090.1000 2445.1600 2091.7000 2445.6400 ;
        RECT 2090.1000 2450.6000 2091.7000 2451.0800 ;
        RECT 2090.1000 2428.8400 2091.7000 2429.3200 ;
        RECT 2090.1000 2434.2800 2091.7000 2434.7600 ;
        RECT 2045.1000 2466.9200 2046.7000 2467.4000 ;
        RECT 2045.1000 2472.3600 2046.7000 2472.8400 ;
        RECT 2045.1000 2477.8000 2046.7000 2478.2800 ;
        RECT 2033.3400 2466.9200 2036.3400 2467.4000 ;
        RECT 2033.3400 2472.3600 2036.3400 2472.8400 ;
        RECT 2033.3400 2477.8000 2036.3400 2478.2800 ;
        RECT 2045.1000 2456.0400 2046.7000 2456.5200 ;
        RECT 2045.1000 2461.4800 2046.7000 2461.9600 ;
        RECT 2033.3400 2456.0400 2036.3400 2456.5200 ;
        RECT 2033.3400 2461.4800 2036.3400 2461.9600 ;
        RECT 2045.1000 2439.7200 2046.7000 2440.2000 ;
        RECT 2045.1000 2445.1600 2046.7000 2445.6400 ;
        RECT 2045.1000 2450.6000 2046.7000 2451.0800 ;
        RECT 2033.3400 2439.7200 2036.3400 2440.2000 ;
        RECT 2033.3400 2445.1600 2036.3400 2445.6400 ;
        RECT 2033.3400 2450.6000 2036.3400 2451.0800 ;
        RECT 2045.1000 2428.8400 2046.7000 2429.3200 ;
        RECT 2045.1000 2434.2800 2046.7000 2434.7600 ;
        RECT 2033.3400 2428.8400 2036.3400 2429.3200 ;
        RECT 2033.3400 2434.2800 2036.3400 2434.7600 ;
        RECT 2135.1000 2412.5200 2136.7000 2413.0000 ;
        RECT 2135.1000 2417.9600 2136.7000 2418.4400 ;
        RECT 2135.1000 2423.4000 2136.7000 2423.8800 ;
        RECT 2135.1000 2401.6400 2136.7000 2402.1200 ;
        RECT 2135.1000 2407.0800 2136.7000 2407.5600 ;
        RECT 2090.1000 2412.5200 2091.7000 2413.0000 ;
        RECT 2090.1000 2417.9600 2091.7000 2418.4400 ;
        RECT 2090.1000 2423.4000 2091.7000 2423.8800 ;
        RECT 2090.1000 2401.6400 2091.7000 2402.1200 ;
        RECT 2090.1000 2407.0800 2091.7000 2407.5600 ;
        RECT 2135.1000 2385.3200 2136.7000 2385.8000 ;
        RECT 2135.1000 2390.7600 2136.7000 2391.2400 ;
        RECT 2135.1000 2396.2000 2136.7000 2396.6800 ;
        RECT 2135.1000 2379.8800 2136.7000 2380.3600 ;
        RECT 2090.1000 2385.3200 2091.7000 2385.8000 ;
        RECT 2090.1000 2390.7600 2091.7000 2391.2400 ;
        RECT 2090.1000 2396.2000 2091.7000 2396.6800 ;
        RECT 2090.1000 2379.8800 2091.7000 2380.3600 ;
        RECT 2045.1000 2412.5200 2046.7000 2413.0000 ;
        RECT 2045.1000 2417.9600 2046.7000 2418.4400 ;
        RECT 2045.1000 2423.4000 2046.7000 2423.8800 ;
        RECT 2033.3400 2412.5200 2036.3400 2413.0000 ;
        RECT 2033.3400 2417.9600 2036.3400 2418.4400 ;
        RECT 2033.3400 2423.4000 2036.3400 2423.8800 ;
        RECT 2045.1000 2401.6400 2046.7000 2402.1200 ;
        RECT 2045.1000 2407.0800 2046.7000 2407.5600 ;
        RECT 2033.3400 2401.6400 2036.3400 2402.1200 ;
        RECT 2033.3400 2407.0800 2036.3400 2407.5600 ;
        RECT 2045.1000 2385.3200 2046.7000 2385.8000 ;
        RECT 2045.1000 2390.7600 2046.7000 2391.2400 ;
        RECT 2045.1000 2396.2000 2046.7000 2396.6800 ;
        RECT 2033.3400 2385.3200 2036.3400 2385.8000 ;
        RECT 2033.3400 2390.7600 2036.3400 2391.2400 ;
        RECT 2033.3400 2396.2000 2036.3400 2396.6800 ;
        RECT 2033.3400 2379.8800 2036.3400 2380.3600 ;
        RECT 2045.1000 2379.8800 2046.7000 2380.3600 ;
        RECT 2033.3400 2584.7900 2240.4400 2587.7900 ;
        RECT 2033.3400 2371.6900 2240.4400 2374.6900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 2142.0500 2226.7000 2358.1500 ;
        RECT 2180.1000 2142.0500 2181.7000 2358.1500 ;
        RECT 2135.1000 2142.0500 2136.7000 2358.1500 ;
        RECT 2090.1000 2142.0500 2091.7000 2358.1500 ;
        RECT 2045.1000 2142.0500 2046.7000 2358.1500 ;
        RECT 2237.4400 2142.0500 2240.4400 2358.1500 ;
        RECT 2033.3400 2142.0500 2036.3400 2358.1500 ;
      LAYER met3 ;
        RECT 2237.4400 2335.2000 2240.4400 2335.6800 ;
        RECT 2237.4400 2340.6400 2240.4400 2341.1200 ;
        RECT 2225.1000 2335.2000 2226.7000 2335.6800 ;
        RECT 2225.1000 2340.6400 2226.7000 2341.1200 ;
        RECT 2237.4400 2346.0800 2240.4400 2346.5600 ;
        RECT 2225.1000 2346.0800 2226.7000 2346.5600 ;
        RECT 2237.4400 2324.3200 2240.4400 2324.8000 ;
        RECT 2237.4400 2329.7600 2240.4400 2330.2400 ;
        RECT 2225.1000 2324.3200 2226.7000 2324.8000 ;
        RECT 2225.1000 2329.7600 2226.7000 2330.2400 ;
        RECT 2237.4400 2308.0000 2240.4400 2308.4800 ;
        RECT 2237.4400 2313.4400 2240.4400 2313.9200 ;
        RECT 2225.1000 2308.0000 2226.7000 2308.4800 ;
        RECT 2225.1000 2313.4400 2226.7000 2313.9200 ;
        RECT 2237.4400 2318.8800 2240.4400 2319.3600 ;
        RECT 2225.1000 2318.8800 2226.7000 2319.3600 ;
        RECT 2180.1000 2335.2000 2181.7000 2335.6800 ;
        RECT 2180.1000 2340.6400 2181.7000 2341.1200 ;
        RECT 2180.1000 2346.0800 2181.7000 2346.5600 ;
        RECT 2180.1000 2324.3200 2181.7000 2324.8000 ;
        RECT 2180.1000 2329.7600 2181.7000 2330.2400 ;
        RECT 2180.1000 2308.0000 2181.7000 2308.4800 ;
        RECT 2180.1000 2313.4400 2181.7000 2313.9200 ;
        RECT 2180.1000 2318.8800 2181.7000 2319.3600 ;
        RECT 2237.4400 2291.6800 2240.4400 2292.1600 ;
        RECT 2237.4400 2297.1200 2240.4400 2297.6000 ;
        RECT 2237.4400 2302.5600 2240.4400 2303.0400 ;
        RECT 2225.1000 2291.6800 2226.7000 2292.1600 ;
        RECT 2225.1000 2297.1200 2226.7000 2297.6000 ;
        RECT 2225.1000 2302.5600 2226.7000 2303.0400 ;
        RECT 2237.4400 2280.8000 2240.4400 2281.2800 ;
        RECT 2237.4400 2286.2400 2240.4400 2286.7200 ;
        RECT 2225.1000 2280.8000 2226.7000 2281.2800 ;
        RECT 2225.1000 2286.2400 2226.7000 2286.7200 ;
        RECT 2237.4400 2264.4800 2240.4400 2264.9600 ;
        RECT 2237.4400 2269.9200 2240.4400 2270.4000 ;
        RECT 2237.4400 2275.3600 2240.4400 2275.8400 ;
        RECT 2225.1000 2264.4800 2226.7000 2264.9600 ;
        RECT 2225.1000 2269.9200 2226.7000 2270.4000 ;
        RECT 2225.1000 2275.3600 2226.7000 2275.8400 ;
        RECT 2237.4400 2253.6000 2240.4400 2254.0800 ;
        RECT 2237.4400 2259.0400 2240.4400 2259.5200 ;
        RECT 2225.1000 2253.6000 2226.7000 2254.0800 ;
        RECT 2225.1000 2259.0400 2226.7000 2259.5200 ;
        RECT 2180.1000 2291.6800 2181.7000 2292.1600 ;
        RECT 2180.1000 2297.1200 2181.7000 2297.6000 ;
        RECT 2180.1000 2302.5600 2181.7000 2303.0400 ;
        RECT 2180.1000 2280.8000 2181.7000 2281.2800 ;
        RECT 2180.1000 2286.2400 2181.7000 2286.7200 ;
        RECT 2180.1000 2264.4800 2181.7000 2264.9600 ;
        RECT 2180.1000 2269.9200 2181.7000 2270.4000 ;
        RECT 2180.1000 2275.3600 2181.7000 2275.8400 ;
        RECT 2180.1000 2253.6000 2181.7000 2254.0800 ;
        RECT 2180.1000 2259.0400 2181.7000 2259.5200 ;
        RECT 2135.1000 2335.2000 2136.7000 2335.6800 ;
        RECT 2135.1000 2340.6400 2136.7000 2341.1200 ;
        RECT 2135.1000 2346.0800 2136.7000 2346.5600 ;
        RECT 2090.1000 2335.2000 2091.7000 2335.6800 ;
        RECT 2090.1000 2340.6400 2091.7000 2341.1200 ;
        RECT 2090.1000 2346.0800 2091.7000 2346.5600 ;
        RECT 2135.1000 2324.3200 2136.7000 2324.8000 ;
        RECT 2135.1000 2329.7600 2136.7000 2330.2400 ;
        RECT 2135.1000 2308.0000 2136.7000 2308.4800 ;
        RECT 2135.1000 2313.4400 2136.7000 2313.9200 ;
        RECT 2135.1000 2318.8800 2136.7000 2319.3600 ;
        RECT 2090.1000 2324.3200 2091.7000 2324.8000 ;
        RECT 2090.1000 2329.7600 2091.7000 2330.2400 ;
        RECT 2090.1000 2308.0000 2091.7000 2308.4800 ;
        RECT 2090.1000 2313.4400 2091.7000 2313.9200 ;
        RECT 2090.1000 2318.8800 2091.7000 2319.3600 ;
        RECT 2045.1000 2335.2000 2046.7000 2335.6800 ;
        RECT 2045.1000 2340.6400 2046.7000 2341.1200 ;
        RECT 2033.3400 2340.6400 2036.3400 2341.1200 ;
        RECT 2033.3400 2335.2000 2036.3400 2335.6800 ;
        RECT 2033.3400 2346.0800 2036.3400 2346.5600 ;
        RECT 2045.1000 2346.0800 2046.7000 2346.5600 ;
        RECT 2045.1000 2324.3200 2046.7000 2324.8000 ;
        RECT 2045.1000 2329.7600 2046.7000 2330.2400 ;
        RECT 2033.3400 2329.7600 2036.3400 2330.2400 ;
        RECT 2033.3400 2324.3200 2036.3400 2324.8000 ;
        RECT 2045.1000 2308.0000 2046.7000 2308.4800 ;
        RECT 2045.1000 2313.4400 2046.7000 2313.9200 ;
        RECT 2033.3400 2313.4400 2036.3400 2313.9200 ;
        RECT 2033.3400 2308.0000 2036.3400 2308.4800 ;
        RECT 2033.3400 2318.8800 2036.3400 2319.3600 ;
        RECT 2045.1000 2318.8800 2046.7000 2319.3600 ;
        RECT 2135.1000 2291.6800 2136.7000 2292.1600 ;
        RECT 2135.1000 2297.1200 2136.7000 2297.6000 ;
        RECT 2135.1000 2302.5600 2136.7000 2303.0400 ;
        RECT 2135.1000 2280.8000 2136.7000 2281.2800 ;
        RECT 2135.1000 2286.2400 2136.7000 2286.7200 ;
        RECT 2090.1000 2291.6800 2091.7000 2292.1600 ;
        RECT 2090.1000 2297.1200 2091.7000 2297.6000 ;
        RECT 2090.1000 2302.5600 2091.7000 2303.0400 ;
        RECT 2090.1000 2280.8000 2091.7000 2281.2800 ;
        RECT 2090.1000 2286.2400 2091.7000 2286.7200 ;
        RECT 2135.1000 2264.4800 2136.7000 2264.9600 ;
        RECT 2135.1000 2269.9200 2136.7000 2270.4000 ;
        RECT 2135.1000 2275.3600 2136.7000 2275.8400 ;
        RECT 2135.1000 2253.6000 2136.7000 2254.0800 ;
        RECT 2135.1000 2259.0400 2136.7000 2259.5200 ;
        RECT 2090.1000 2264.4800 2091.7000 2264.9600 ;
        RECT 2090.1000 2269.9200 2091.7000 2270.4000 ;
        RECT 2090.1000 2275.3600 2091.7000 2275.8400 ;
        RECT 2090.1000 2253.6000 2091.7000 2254.0800 ;
        RECT 2090.1000 2259.0400 2091.7000 2259.5200 ;
        RECT 2045.1000 2291.6800 2046.7000 2292.1600 ;
        RECT 2045.1000 2297.1200 2046.7000 2297.6000 ;
        RECT 2045.1000 2302.5600 2046.7000 2303.0400 ;
        RECT 2033.3400 2291.6800 2036.3400 2292.1600 ;
        RECT 2033.3400 2297.1200 2036.3400 2297.6000 ;
        RECT 2033.3400 2302.5600 2036.3400 2303.0400 ;
        RECT 2045.1000 2280.8000 2046.7000 2281.2800 ;
        RECT 2045.1000 2286.2400 2046.7000 2286.7200 ;
        RECT 2033.3400 2280.8000 2036.3400 2281.2800 ;
        RECT 2033.3400 2286.2400 2036.3400 2286.7200 ;
        RECT 2045.1000 2264.4800 2046.7000 2264.9600 ;
        RECT 2045.1000 2269.9200 2046.7000 2270.4000 ;
        RECT 2045.1000 2275.3600 2046.7000 2275.8400 ;
        RECT 2033.3400 2264.4800 2036.3400 2264.9600 ;
        RECT 2033.3400 2269.9200 2036.3400 2270.4000 ;
        RECT 2033.3400 2275.3600 2036.3400 2275.8400 ;
        RECT 2045.1000 2253.6000 2046.7000 2254.0800 ;
        RECT 2045.1000 2259.0400 2046.7000 2259.5200 ;
        RECT 2033.3400 2253.6000 2036.3400 2254.0800 ;
        RECT 2033.3400 2259.0400 2036.3400 2259.5200 ;
        RECT 2237.4400 2237.2800 2240.4400 2237.7600 ;
        RECT 2237.4400 2242.7200 2240.4400 2243.2000 ;
        RECT 2237.4400 2248.1600 2240.4400 2248.6400 ;
        RECT 2225.1000 2237.2800 2226.7000 2237.7600 ;
        RECT 2225.1000 2242.7200 2226.7000 2243.2000 ;
        RECT 2225.1000 2248.1600 2226.7000 2248.6400 ;
        RECT 2237.4400 2226.4000 2240.4400 2226.8800 ;
        RECT 2237.4400 2231.8400 2240.4400 2232.3200 ;
        RECT 2225.1000 2226.4000 2226.7000 2226.8800 ;
        RECT 2225.1000 2231.8400 2226.7000 2232.3200 ;
        RECT 2237.4400 2210.0800 2240.4400 2210.5600 ;
        RECT 2237.4400 2215.5200 2240.4400 2216.0000 ;
        RECT 2237.4400 2220.9600 2240.4400 2221.4400 ;
        RECT 2225.1000 2210.0800 2226.7000 2210.5600 ;
        RECT 2225.1000 2215.5200 2226.7000 2216.0000 ;
        RECT 2225.1000 2220.9600 2226.7000 2221.4400 ;
        RECT 2237.4400 2199.2000 2240.4400 2199.6800 ;
        RECT 2237.4400 2204.6400 2240.4400 2205.1200 ;
        RECT 2225.1000 2199.2000 2226.7000 2199.6800 ;
        RECT 2225.1000 2204.6400 2226.7000 2205.1200 ;
        RECT 2180.1000 2237.2800 2181.7000 2237.7600 ;
        RECT 2180.1000 2242.7200 2181.7000 2243.2000 ;
        RECT 2180.1000 2248.1600 2181.7000 2248.6400 ;
        RECT 2180.1000 2226.4000 2181.7000 2226.8800 ;
        RECT 2180.1000 2231.8400 2181.7000 2232.3200 ;
        RECT 2180.1000 2210.0800 2181.7000 2210.5600 ;
        RECT 2180.1000 2215.5200 2181.7000 2216.0000 ;
        RECT 2180.1000 2220.9600 2181.7000 2221.4400 ;
        RECT 2180.1000 2199.2000 2181.7000 2199.6800 ;
        RECT 2180.1000 2204.6400 2181.7000 2205.1200 ;
        RECT 2237.4400 2182.8800 2240.4400 2183.3600 ;
        RECT 2237.4400 2188.3200 2240.4400 2188.8000 ;
        RECT 2237.4400 2193.7600 2240.4400 2194.2400 ;
        RECT 2225.1000 2182.8800 2226.7000 2183.3600 ;
        RECT 2225.1000 2188.3200 2226.7000 2188.8000 ;
        RECT 2225.1000 2193.7600 2226.7000 2194.2400 ;
        RECT 2237.4400 2172.0000 2240.4400 2172.4800 ;
        RECT 2237.4400 2177.4400 2240.4400 2177.9200 ;
        RECT 2225.1000 2172.0000 2226.7000 2172.4800 ;
        RECT 2225.1000 2177.4400 2226.7000 2177.9200 ;
        RECT 2237.4400 2155.6800 2240.4400 2156.1600 ;
        RECT 2237.4400 2161.1200 2240.4400 2161.6000 ;
        RECT 2237.4400 2166.5600 2240.4400 2167.0400 ;
        RECT 2225.1000 2155.6800 2226.7000 2156.1600 ;
        RECT 2225.1000 2161.1200 2226.7000 2161.6000 ;
        RECT 2225.1000 2166.5600 2226.7000 2167.0400 ;
        RECT 2237.4400 2150.2400 2240.4400 2150.7200 ;
        RECT 2225.1000 2150.2400 2226.7000 2150.7200 ;
        RECT 2180.1000 2182.8800 2181.7000 2183.3600 ;
        RECT 2180.1000 2188.3200 2181.7000 2188.8000 ;
        RECT 2180.1000 2193.7600 2181.7000 2194.2400 ;
        RECT 2180.1000 2172.0000 2181.7000 2172.4800 ;
        RECT 2180.1000 2177.4400 2181.7000 2177.9200 ;
        RECT 2180.1000 2155.6800 2181.7000 2156.1600 ;
        RECT 2180.1000 2161.1200 2181.7000 2161.6000 ;
        RECT 2180.1000 2166.5600 2181.7000 2167.0400 ;
        RECT 2180.1000 2150.2400 2181.7000 2150.7200 ;
        RECT 2135.1000 2237.2800 2136.7000 2237.7600 ;
        RECT 2135.1000 2242.7200 2136.7000 2243.2000 ;
        RECT 2135.1000 2248.1600 2136.7000 2248.6400 ;
        RECT 2135.1000 2226.4000 2136.7000 2226.8800 ;
        RECT 2135.1000 2231.8400 2136.7000 2232.3200 ;
        RECT 2090.1000 2237.2800 2091.7000 2237.7600 ;
        RECT 2090.1000 2242.7200 2091.7000 2243.2000 ;
        RECT 2090.1000 2248.1600 2091.7000 2248.6400 ;
        RECT 2090.1000 2226.4000 2091.7000 2226.8800 ;
        RECT 2090.1000 2231.8400 2091.7000 2232.3200 ;
        RECT 2135.1000 2210.0800 2136.7000 2210.5600 ;
        RECT 2135.1000 2215.5200 2136.7000 2216.0000 ;
        RECT 2135.1000 2220.9600 2136.7000 2221.4400 ;
        RECT 2135.1000 2199.2000 2136.7000 2199.6800 ;
        RECT 2135.1000 2204.6400 2136.7000 2205.1200 ;
        RECT 2090.1000 2210.0800 2091.7000 2210.5600 ;
        RECT 2090.1000 2215.5200 2091.7000 2216.0000 ;
        RECT 2090.1000 2220.9600 2091.7000 2221.4400 ;
        RECT 2090.1000 2199.2000 2091.7000 2199.6800 ;
        RECT 2090.1000 2204.6400 2091.7000 2205.1200 ;
        RECT 2045.1000 2237.2800 2046.7000 2237.7600 ;
        RECT 2045.1000 2242.7200 2046.7000 2243.2000 ;
        RECT 2045.1000 2248.1600 2046.7000 2248.6400 ;
        RECT 2033.3400 2237.2800 2036.3400 2237.7600 ;
        RECT 2033.3400 2242.7200 2036.3400 2243.2000 ;
        RECT 2033.3400 2248.1600 2036.3400 2248.6400 ;
        RECT 2045.1000 2226.4000 2046.7000 2226.8800 ;
        RECT 2045.1000 2231.8400 2046.7000 2232.3200 ;
        RECT 2033.3400 2226.4000 2036.3400 2226.8800 ;
        RECT 2033.3400 2231.8400 2036.3400 2232.3200 ;
        RECT 2045.1000 2210.0800 2046.7000 2210.5600 ;
        RECT 2045.1000 2215.5200 2046.7000 2216.0000 ;
        RECT 2045.1000 2220.9600 2046.7000 2221.4400 ;
        RECT 2033.3400 2210.0800 2036.3400 2210.5600 ;
        RECT 2033.3400 2215.5200 2036.3400 2216.0000 ;
        RECT 2033.3400 2220.9600 2036.3400 2221.4400 ;
        RECT 2045.1000 2199.2000 2046.7000 2199.6800 ;
        RECT 2045.1000 2204.6400 2046.7000 2205.1200 ;
        RECT 2033.3400 2199.2000 2036.3400 2199.6800 ;
        RECT 2033.3400 2204.6400 2036.3400 2205.1200 ;
        RECT 2135.1000 2182.8800 2136.7000 2183.3600 ;
        RECT 2135.1000 2188.3200 2136.7000 2188.8000 ;
        RECT 2135.1000 2193.7600 2136.7000 2194.2400 ;
        RECT 2135.1000 2172.0000 2136.7000 2172.4800 ;
        RECT 2135.1000 2177.4400 2136.7000 2177.9200 ;
        RECT 2090.1000 2182.8800 2091.7000 2183.3600 ;
        RECT 2090.1000 2188.3200 2091.7000 2188.8000 ;
        RECT 2090.1000 2193.7600 2091.7000 2194.2400 ;
        RECT 2090.1000 2172.0000 2091.7000 2172.4800 ;
        RECT 2090.1000 2177.4400 2091.7000 2177.9200 ;
        RECT 2135.1000 2155.6800 2136.7000 2156.1600 ;
        RECT 2135.1000 2161.1200 2136.7000 2161.6000 ;
        RECT 2135.1000 2166.5600 2136.7000 2167.0400 ;
        RECT 2135.1000 2150.2400 2136.7000 2150.7200 ;
        RECT 2090.1000 2155.6800 2091.7000 2156.1600 ;
        RECT 2090.1000 2161.1200 2091.7000 2161.6000 ;
        RECT 2090.1000 2166.5600 2091.7000 2167.0400 ;
        RECT 2090.1000 2150.2400 2091.7000 2150.7200 ;
        RECT 2045.1000 2182.8800 2046.7000 2183.3600 ;
        RECT 2045.1000 2188.3200 2046.7000 2188.8000 ;
        RECT 2045.1000 2193.7600 2046.7000 2194.2400 ;
        RECT 2033.3400 2182.8800 2036.3400 2183.3600 ;
        RECT 2033.3400 2188.3200 2036.3400 2188.8000 ;
        RECT 2033.3400 2193.7600 2036.3400 2194.2400 ;
        RECT 2045.1000 2172.0000 2046.7000 2172.4800 ;
        RECT 2045.1000 2177.4400 2046.7000 2177.9200 ;
        RECT 2033.3400 2172.0000 2036.3400 2172.4800 ;
        RECT 2033.3400 2177.4400 2036.3400 2177.9200 ;
        RECT 2045.1000 2155.6800 2046.7000 2156.1600 ;
        RECT 2045.1000 2161.1200 2046.7000 2161.6000 ;
        RECT 2045.1000 2166.5600 2046.7000 2167.0400 ;
        RECT 2033.3400 2155.6800 2036.3400 2156.1600 ;
        RECT 2033.3400 2161.1200 2036.3400 2161.6000 ;
        RECT 2033.3400 2166.5600 2036.3400 2167.0400 ;
        RECT 2033.3400 2150.2400 2036.3400 2150.7200 ;
        RECT 2045.1000 2150.2400 2046.7000 2150.7200 ;
        RECT 2033.3400 2355.1500 2240.4400 2358.1500 ;
        RECT 2033.3400 2142.0500 2240.4400 2145.0500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 1912.4100 2226.7000 2128.5100 ;
        RECT 2180.1000 1912.4100 2181.7000 2128.5100 ;
        RECT 2135.1000 1912.4100 2136.7000 2128.5100 ;
        RECT 2090.1000 1912.4100 2091.7000 2128.5100 ;
        RECT 2045.1000 1912.4100 2046.7000 2128.5100 ;
        RECT 2237.4400 1912.4100 2240.4400 2128.5100 ;
        RECT 2033.3400 1912.4100 2036.3400 2128.5100 ;
      LAYER met3 ;
        RECT 2237.4400 2105.5600 2240.4400 2106.0400 ;
        RECT 2237.4400 2111.0000 2240.4400 2111.4800 ;
        RECT 2225.1000 2105.5600 2226.7000 2106.0400 ;
        RECT 2225.1000 2111.0000 2226.7000 2111.4800 ;
        RECT 2237.4400 2116.4400 2240.4400 2116.9200 ;
        RECT 2225.1000 2116.4400 2226.7000 2116.9200 ;
        RECT 2237.4400 2094.6800 2240.4400 2095.1600 ;
        RECT 2237.4400 2100.1200 2240.4400 2100.6000 ;
        RECT 2225.1000 2094.6800 2226.7000 2095.1600 ;
        RECT 2225.1000 2100.1200 2226.7000 2100.6000 ;
        RECT 2237.4400 2078.3600 2240.4400 2078.8400 ;
        RECT 2237.4400 2083.8000 2240.4400 2084.2800 ;
        RECT 2225.1000 2078.3600 2226.7000 2078.8400 ;
        RECT 2225.1000 2083.8000 2226.7000 2084.2800 ;
        RECT 2237.4400 2089.2400 2240.4400 2089.7200 ;
        RECT 2225.1000 2089.2400 2226.7000 2089.7200 ;
        RECT 2180.1000 2105.5600 2181.7000 2106.0400 ;
        RECT 2180.1000 2111.0000 2181.7000 2111.4800 ;
        RECT 2180.1000 2116.4400 2181.7000 2116.9200 ;
        RECT 2180.1000 2094.6800 2181.7000 2095.1600 ;
        RECT 2180.1000 2100.1200 2181.7000 2100.6000 ;
        RECT 2180.1000 2078.3600 2181.7000 2078.8400 ;
        RECT 2180.1000 2083.8000 2181.7000 2084.2800 ;
        RECT 2180.1000 2089.2400 2181.7000 2089.7200 ;
        RECT 2237.4400 2062.0400 2240.4400 2062.5200 ;
        RECT 2237.4400 2067.4800 2240.4400 2067.9600 ;
        RECT 2237.4400 2072.9200 2240.4400 2073.4000 ;
        RECT 2225.1000 2062.0400 2226.7000 2062.5200 ;
        RECT 2225.1000 2067.4800 2226.7000 2067.9600 ;
        RECT 2225.1000 2072.9200 2226.7000 2073.4000 ;
        RECT 2237.4400 2051.1600 2240.4400 2051.6400 ;
        RECT 2237.4400 2056.6000 2240.4400 2057.0800 ;
        RECT 2225.1000 2051.1600 2226.7000 2051.6400 ;
        RECT 2225.1000 2056.6000 2226.7000 2057.0800 ;
        RECT 2237.4400 2034.8400 2240.4400 2035.3200 ;
        RECT 2237.4400 2040.2800 2240.4400 2040.7600 ;
        RECT 2237.4400 2045.7200 2240.4400 2046.2000 ;
        RECT 2225.1000 2034.8400 2226.7000 2035.3200 ;
        RECT 2225.1000 2040.2800 2226.7000 2040.7600 ;
        RECT 2225.1000 2045.7200 2226.7000 2046.2000 ;
        RECT 2237.4400 2023.9600 2240.4400 2024.4400 ;
        RECT 2237.4400 2029.4000 2240.4400 2029.8800 ;
        RECT 2225.1000 2023.9600 2226.7000 2024.4400 ;
        RECT 2225.1000 2029.4000 2226.7000 2029.8800 ;
        RECT 2180.1000 2062.0400 2181.7000 2062.5200 ;
        RECT 2180.1000 2067.4800 2181.7000 2067.9600 ;
        RECT 2180.1000 2072.9200 2181.7000 2073.4000 ;
        RECT 2180.1000 2051.1600 2181.7000 2051.6400 ;
        RECT 2180.1000 2056.6000 2181.7000 2057.0800 ;
        RECT 2180.1000 2034.8400 2181.7000 2035.3200 ;
        RECT 2180.1000 2040.2800 2181.7000 2040.7600 ;
        RECT 2180.1000 2045.7200 2181.7000 2046.2000 ;
        RECT 2180.1000 2023.9600 2181.7000 2024.4400 ;
        RECT 2180.1000 2029.4000 2181.7000 2029.8800 ;
        RECT 2135.1000 2105.5600 2136.7000 2106.0400 ;
        RECT 2135.1000 2111.0000 2136.7000 2111.4800 ;
        RECT 2135.1000 2116.4400 2136.7000 2116.9200 ;
        RECT 2090.1000 2105.5600 2091.7000 2106.0400 ;
        RECT 2090.1000 2111.0000 2091.7000 2111.4800 ;
        RECT 2090.1000 2116.4400 2091.7000 2116.9200 ;
        RECT 2135.1000 2094.6800 2136.7000 2095.1600 ;
        RECT 2135.1000 2100.1200 2136.7000 2100.6000 ;
        RECT 2135.1000 2078.3600 2136.7000 2078.8400 ;
        RECT 2135.1000 2083.8000 2136.7000 2084.2800 ;
        RECT 2135.1000 2089.2400 2136.7000 2089.7200 ;
        RECT 2090.1000 2094.6800 2091.7000 2095.1600 ;
        RECT 2090.1000 2100.1200 2091.7000 2100.6000 ;
        RECT 2090.1000 2078.3600 2091.7000 2078.8400 ;
        RECT 2090.1000 2083.8000 2091.7000 2084.2800 ;
        RECT 2090.1000 2089.2400 2091.7000 2089.7200 ;
        RECT 2045.1000 2105.5600 2046.7000 2106.0400 ;
        RECT 2045.1000 2111.0000 2046.7000 2111.4800 ;
        RECT 2033.3400 2111.0000 2036.3400 2111.4800 ;
        RECT 2033.3400 2105.5600 2036.3400 2106.0400 ;
        RECT 2033.3400 2116.4400 2036.3400 2116.9200 ;
        RECT 2045.1000 2116.4400 2046.7000 2116.9200 ;
        RECT 2045.1000 2094.6800 2046.7000 2095.1600 ;
        RECT 2045.1000 2100.1200 2046.7000 2100.6000 ;
        RECT 2033.3400 2100.1200 2036.3400 2100.6000 ;
        RECT 2033.3400 2094.6800 2036.3400 2095.1600 ;
        RECT 2045.1000 2078.3600 2046.7000 2078.8400 ;
        RECT 2045.1000 2083.8000 2046.7000 2084.2800 ;
        RECT 2033.3400 2083.8000 2036.3400 2084.2800 ;
        RECT 2033.3400 2078.3600 2036.3400 2078.8400 ;
        RECT 2033.3400 2089.2400 2036.3400 2089.7200 ;
        RECT 2045.1000 2089.2400 2046.7000 2089.7200 ;
        RECT 2135.1000 2062.0400 2136.7000 2062.5200 ;
        RECT 2135.1000 2067.4800 2136.7000 2067.9600 ;
        RECT 2135.1000 2072.9200 2136.7000 2073.4000 ;
        RECT 2135.1000 2051.1600 2136.7000 2051.6400 ;
        RECT 2135.1000 2056.6000 2136.7000 2057.0800 ;
        RECT 2090.1000 2062.0400 2091.7000 2062.5200 ;
        RECT 2090.1000 2067.4800 2091.7000 2067.9600 ;
        RECT 2090.1000 2072.9200 2091.7000 2073.4000 ;
        RECT 2090.1000 2051.1600 2091.7000 2051.6400 ;
        RECT 2090.1000 2056.6000 2091.7000 2057.0800 ;
        RECT 2135.1000 2034.8400 2136.7000 2035.3200 ;
        RECT 2135.1000 2040.2800 2136.7000 2040.7600 ;
        RECT 2135.1000 2045.7200 2136.7000 2046.2000 ;
        RECT 2135.1000 2023.9600 2136.7000 2024.4400 ;
        RECT 2135.1000 2029.4000 2136.7000 2029.8800 ;
        RECT 2090.1000 2034.8400 2091.7000 2035.3200 ;
        RECT 2090.1000 2040.2800 2091.7000 2040.7600 ;
        RECT 2090.1000 2045.7200 2091.7000 2046.2000 ;
        RECT 2090.1000 2023.9600 2091.7000 2024.4400 ;
        RECT 2090.1000 2029.4000 2091.7000 2029.8800 ;
        RECT 2045.1000 2062.0400 2046.7000 2062.5200 ;
        RECT 2045.1000 2067.4800 2046.7000 2067.9600 ;
        RECT 2045.1000 2072.9200 2046.7000 2073.4000 ;
        RECT 2033.3400 2062.0400 2036.3400 2062.5200 ;
        RECT 2033.3400 2067.4800 2036.3400 2067.9600 ;
        RECT 2033.3400 2072.9200 2036.3400 2073.4000 ;
        RECT 2045.1000 2051.1600 2046.7000 2051.6400 ;
        RECT 2045.1000 2056.6000 2046.7000 2057.0800 ;
        RECT 2033.3400 2051.1600 2036.3400 2051.6400 ;
        RECT 2033.3400 2056.6000 2036.3400 2057.0800 ;
        RECT 2045.1000 2034.8400 2046.7000 2035.3200 ;
        RECT 2045.1000 2040.2800 2046.7000 2040.7600 ;
        RECT 2045.1000 2045.7200 2046.7000 2046.2000 ;
        RECT 2033.3400 2034.8400 2036.3400 2035.3200 ;
        RECT 2033.3400 2040.2800 2036.3400 2040.7600 ;
        RECT 2033.3400 2045.7200 2036.3400 2046.2000 ;
        RECT 2045.1000 2023.9600 2046.7000 2024.4400 ;
        RECT 2045.1000 2029.4000 2046.7000 2029.8800 ;
        RECT 2033.3400 2023.9600 2036.3400 2024.4400 ;
        RECT 2033.3400 2029.4000 2036.3400 2029.8800 ;
        RECT 2237.4400 2007.6400 2240.4400 2008.1200 ;
        RECT 2237.4400 2013.0800 2240.4400 2013.5600 ;
        RECT 2237.4400 2018.5200 2240.4400 2019.0000 ;
        RECT 2225.1000 2007.6400 2226.7000 2008.1200 ;
        RECT 2225.1000 2013.0800 2226.7000 2013.5600 ;
        RECT 2225.1000 2018.5200 2226.7000 2019.0000 ;
        RECT 2237.4400 1996.7600 2240.4400 1997.2400 ;
        RECT 2237.4400 2002.2000 2240.4400 2002.6800 ;
        RECT 2225.1000 1996.7600 2226.7000 1997.2400 ;
        RECT 2225.1000 2002.2000 2226.7000 2002.6800 ;
        RECT 2237.4400 1980.4400 2240.4400 1980.9200 ;
        RECT 2237.4400 1985.8800 2240.4400 1986.3600 ;
        RECT 2237.4400 1991.3200 2240.4400 1991.8000 ;
        RECT 2225.1000 1980.4400 2226.7000 1980.9200 ;
        RECT 2225.1000 1985.8800 2226.7000 1986.3600 ;
        RECT 2225.1000 1991.3200 2226.7000 1991.8000 ;
        RECT 2237.4400 1969.5600 2240.4400 1970.0400 ;
        RECT 2237.4400 1975.0000 2240.4400 1975.4800 ;
        RECT 2225.1000 1969.5600 2226.7000 1970.0400 ;
        RECT 2225.1000 1975.0000 2226.7000 1975.4800 ;
        RECT 2180.1000 2007.6400 2181.7000 2008.1200 ;
        RECT 2180.1000 2013.0800 2181.7000 2013.5600 ;
        RECT 2180.1000 2018.5200 2181.7000 2019.0000 ;
        RECT 2180.1000 1996.7600 2181.7000 1997.2400 ;
        RECT 2180.1000 2002.2000 2181.7000 2002.6800 ;
        RECT 2180.1000 1980.4400 2181.7000 1980.9200 ;
        RECT 2180.1000 1985.8800 2181.7000 1986.3600 ;
        RECT 2180.1000 1991.3200 2181.7000 1991.8000 ;
        RECT 2180.1000 1969.5600 2181.7000 1970.0400 ;
        RECT 2180.1000 1975.0000 2181.7000 1975.4800 ;
        RECT 2237.4400 1953.2400 2240.4400 1953.7200 ;
        RECT 2237.4400 1958.6800 2240.4400 1959.1600 ;
        RECT 2237.4400 1964.1200 2240.4400 1964.6000 ;
        RECT 2225.1000 1953.2400 2226.7000 1953.7200 ;
        RECT 2225.1000 1958.6800 2226.7000 1959.1600 ;
        RECT 2225.1000 1964.1200 2226.7000 1964.6000 ;
        RECT 2237.4400 1942.3600 2240.4400 1942.8400 ;
        RECT 2237.4400 1947.8000 2240.4400 1948.2800 ;
        RECT 2225.1000 1942.3600 2226.7000 1942.8400 ;
        RECT 2225.1000 1947.8000 2226.7000 1948.2800 ;
        RECT 2237.4400 1926.0400 2240.4400 1926.5200 ;
        RECT 2237.4400 1931.4800 2240.4400 1931.9600 ;
        RECT 2237.4400 1936.9200 2240.4400 1937.4000 ;
        RECT 2225.1000 1926.0400 2226.7000 1926.5200 ;
        RECT 2225.1000 1931.4800 2226.7000 1931.9600 ;
        RECT 2225.1000 1936.9200 2226.7000 1937.4000 ;
        RECT 2237.4400 1920.6000 2240.4400 1921.0800 ;
        RECT 2225.1000 1920.6000 2226.7000 1921.0800 ;
        RECT 2180.1000 1953.2400 2181.7000 1953.7200 ;
        RECT 2180.1000 1958.6800 2181.7000 1959.1600 ;
        RECT 2180.1000 1964.1200 2181.7000 1964.6000 ;
        RECT 2180.1000 1942.3600 2181.7000 1942.8400 ;
        RECT 2180.1000 1947.8000 2181.7000 1948.2800 ;
        RECT 2180.1000 1926.0400 2181.7000 1926.5200 ;
        RECT 2180.1000 1931.4800 2181.7000 1931.9600 ;
        RECT 2180.1000 1936.9200 2181.7000 1937.4000 ;
        RECT 2180.1000 1920.6000 2181.7000 1921.0800 ;
        RECT 2135.1000 2007.6400 2136.7000 2008.1200 ;
        RECT 2135.1000 2013.0800 2136.7000 2013.5600 ;
        RECT 2135.1000 2018.5200 2136.7000 2019.0000 ;
        RECT 2135.1000 1996.7600 2136.7000 1997.2400 ;
        RECT 2135.1000 2002.2000 2136.7000 2002.6800 ;
        RECT 2090.1000 2007.6400 2091.7000 2008.1200 ;
        RECT 2090.1000 2013.0800 2091.7000 2013.5600 ;
        RECT 2090.1000 2018.5200 2091.7000 2019.0000 ;
        RECT 2090.1000 1996.7600 2091.7000 1997.2400 ;
        RECT 2090.1000 2002.2000 2091.7000 2002.6800 ;
        RECT 2135.1000 1980.4400 2136.7000 1980.9200 ;
        RECT 2135.1000 1985.8800 2136.7000 1986.3600 ;
        RECT 2135.1000 1991.3200 2136.7000 1991.8000 ;
        RECT 2135.1000 1969.5600 2136.7000 1970.0400 ;
        RECT 2135.1000 1975.0000 2136.7000 1975.4800 ;
        RECT 2090.1000 1980.4400 2091.7000 1980.9200 ;
        RECT 2090.1000 1985.8800 2091.7000 1986.3600 ;
        RECT 2090.1000 1991.3200 2091.7000 1991.8000 ;
        RECT 2090.1000 1969.5600 2091.7000 1970.0400 ;
        RECT 2090.1000 1975.0000 2091.7000 1975.4800 ;
        RECT 2045.1000 2007.6400 2046.7000 2008.1200 ;
        RECT 2045.1000 2013.0800 2046.7000 2013.5600 ;
        RECT 2045.1000 2018.5200 2046.7000 2019.0000 ;
        RECT 2033.3400 2007.6400 2036.3400 2008.1200 ;
        RECT 2033.3400 2013.0800 2036.3400 2013.5600 ;
        RECT 2033.3400 2018.5200 2036.3400 2019.0000 ;
        RECT 2045.1000 1996.7600 2046.7000 1997.2400 ;
        RECT 2045.1000 2002.2000 2046.7000 2002.6800 ;
        RECT 2033.3400 1996.7600 2036.3400 1997.2400 ;
        RECT 2033.3400 2002.2000 2036.3400 2002.6800 ;
        RECT 2045.1000 1980.4400 2046.7000 1980.9200 ;
        RECT 2045.1000 1985.8800 2046.7000 1986.3600 ;
        RECT 2045.1000 1991.3200 2046.7000 1991.8000 ;
        RECT 2033.3400 1980.4400 2036.3400 1980.9200 ;
        RECT 2033.3400 1985.8800 2036.3400 1986.3600 ;
        RECT 2033.3400 1991.3200 2036.3400 1991.8000 ;
        RECT 2045.1000 1969.5600 2046.7000 1970.0400 ;
        RECT 2045.1000 1975.0000 2046.7000 1975.4800 ;
        RECT 2033.3400 1969.5600 2036.3400 1970.0400 ;
        RECT 2033.3400 1975.0000 2036.3400 1975.4800 ;
        RECT 2135.1000 1953.2400 2136.7000 1953.7200 ;
        RECT 2135.1000 1958.6800 2136.7000 1959.1600 ;
        RECT 2135.1000 1964.1200 2136.7000 1964.6000 ;
        RECT 2135.1000 1942.3600 2136.7000 1942.8400 ;
        RECT 2135.1000 1947.8000 2136.7000 1948.2800 ;
        RECT 2090.1000 1953.2400 2091.7000 1953.7200 ;
        RECT 2090.1000 1958.6800 2091.7000 1959.1600 ;
        RECT 2090.1000 1964.1200 2091.7000 1964.6000 ;
        RECT 2090.1000 1942.3600 2091.7000 1942.8400 ;
        RECT 2090.1000 1947.8000 2091.7000 1948.2800 ;
        RECT 2135.1000 1926.0400 2136.7000 1926.5200 ;
        RECT 2135.1000 1931.4800 2136.7000 1931.9600 ;
        RECT 2135.1000 1936.9200 2136.7000 1937.4000 ;
        RECT 2135.1000 1920.6000 2136.7000 1921.0800 ;
        RECT 2090.1000 1926.0400 2091.7000 1926.5200 ;
        RECT 2090.1000 1931.4800 2091.7000 1931.9600 ;
        RECT 2090.1000 1936.9200 2091.7000 1937.4000 ;
        RECT 2090.1000 1920.6000 2091.7000 1921.0800 ;
        RECT 2045.1000 1953.2400 2046.7000 1953.7200 ;
        RECT 2045.1000 1958.6800 2046.7000 1959.1600 ;
        RECT 2045.1000 1964.1200 2046.7000 1964.6000 ;
        RECT 2033.3400 1953.2400 2036.3400 1953.7200 ;
        RECT 2033.3400 1958.6800 2036.3400 1959.1600 ;
        RECT 2033.3400 1964.1200 2036.3400 1964.6000 ;
        RECT 2045.1000 1942.3600 2046.7000 1942.8400 ;
        RECT 2045.1000 1947.8000 2046.7000 1948.2800 ;
        RECT 2033.3400 1942.3600 2036.3400 1942.8400 ;
        RECT 2033.3400 1947.8000 2036.3400 1948.2800 ;
        RECT 2045.1000 1926.0400 2046.7000 1926.5200 ;
        RECT 2045.1000 1931.4800 2046.7000 1931.9600 ;
        RECT 2045.1000 1936.9200 2046.7000 1937.4000 ;
        RECT 2033.3400 1926.0400 2036.3400 1926.5200 ;
        RECT 2033.3400 1931.4800 2036.3400 1931.9600 ;
        RECT 2033.3400 1936.9200 2036.3400 1937.4000 ;
        RECT 2033.3400 1920.6000 2036.3400 1921.0800 ;
        RECT 2045.1000 1920.6000 2046.7000 1921.0800 ;
        RECT 2033.3400 2125.5100 2240.4400 2128.5100 ;
        RECT 2033.3400 1912.4100 2240.4400 1915.4100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 1682.7700 2226.7000 1898.8700 ;
        RECT 2180.1000 1682.7700 2181.7000 1898.8700 ;
        RECT 2135.1000 1682.7700 2136.7000 1898.8700 ;
        RECT 2090.1000 1682.7700 2091.7000 1898.8700 ;
        RECT 2045.1000 1682.7700 2046.7000 1898.8700 ;
        RECT 2237.4400 1682.7700 2240.4400 1898.8700 ;
        RECT 2033.3400 1682.7700 2036.3400 1898.8700 ;
      LAYER met3 ;
        RECT 2237.4400 1875.9200 2240.4400 1876.4000 ;
        RECT 2237.4400 1881.3600 2240.4400 1881.8400 ;
        RECT 2225.1000 1875.9200 2226.7000 1876.4000 ;
        RECT 2225.1000 1881.3600 2226.7000 1881.8400 ;
        RECT 2237.4400 1886.8000 2240.4400 1887.2800 ;
        RECT 2225.1000 1886.8000 2226.7000 1887.2800 ;
        RECT 2237.4400 1865.0400 2240.4400 1865.5200 ;
        RECT 2237.4400 1870.4800 2240.4400 1870.9600 ;
        RECT 2225.1000 1865.0400 2226.7000 1865.5200 ;
        RECT 2225.1000 1870.4800 2226.7000 1870.9600 ;
        RECT 2237.4400 1848.7200 2240.4400 1849.2000 ;
        RECT 2237.4400 1854.1600 2240.4400 1854.6400 ;
        RECT 2225.1000 1848.7200 2226.7000 1849.2000 ;
        RECT 2225.1000 1854.1600 2226.7000 1854.6400 ;
        RECT 2237.4400 1859.6000 2240.4400 1860.0800 ;
        RECT 2225.1000 1859.6000 2226.7000 1860.0800 ;
        RECT 2180.1000 1875.9200 2181.7000 1876.4000 ;
        RECT 2180.1000 1881.3600 2181.7000 1881.8400 ;
        RECT 2180.1000 1886.8000 2181.7000 1887.2800 ;
        RECT 2180.1000 1865.0400 2181.7000 1865.5200 ;
        RECT 2180.1000 1870.4800 2181.7000 1870.9600 ;
        RECT 2180.1000 1848.7200 2181.7000 1849.2000 ;
        RECT 2180.1000 1854.1600 2181.7000 1854.6400 ;
        RECT 2180.1000 1859.6000 2181.7000 1860.0800 ;
        RECT 2237.4400 1832.4000 2240.4400 1832.8800 ;
        RECT 2237.4400 1837.8400 2240.4400 1838.3200 ;
        RECT 2237.4400 1843.2800 2240.4400 1843.7600 ;
        RECT 2225.1000 1832.4000 2226.7000 1832.8800 ;
        RECT 2225.1000 1837.8400 2226.7000 1838.3200 ;
        RECT 2225.1000 1843.2800 2226.7000 1843.7600 ;
        RECT 2237.4400 1821.5200 2240.4400 1822.0000 ;
        RECT 2237.4400 1826.9600 2240.4400 1827.4400 ;
        RECT 2225.1000 1821.5200 2226.7000 1822.0000 ;
        RECT 2225.1000 1826.9600 2226.7000 1827.4400 ;
        RECT 2237.4400 1805.2000 2240.4400 1805.6800 ;
        RECT 2237.4400 1810.6400 2240.4400 1811.1200 ;
        RECT 2237.4400 1816.0800 2240.4400 1816.5600 ;
        RECT 2225.1000 1805.2000 2226.7000 1805.6800 ;
        RECT 2225.1000 1810.6400 2226.7000 1811.1200 ;
        RECT 2225.1000 1816.0800 2226.7000 1816.5600 ;
        RECT 2237.4400 1794.3200 2240.4400 1794.8000 ;
        RECT 2237.4400 1799.7600 2240.4400 1800.2400 ;
        RECT 2225.1000 1794.3200 2226.7000 1794.8000 ;
        RECT 2225.1000 1799.7600 2226.7000 1800.2400 ;
        RECT 2180.1000 1832.4000 2181.7000 1832.8800 ;
        RECT 2180.1000 1837.8400 2181.7000 1838.3200 ;
        RECT 2180.1000 1843.2800 2181.7000 1843.7600 ;
        RECT 2180.1000 1821.5200 2181.7000 1822.0000 ;
        RECT 2180.1000 1826.9600 2181.7000 1827.4400 ;
        RECT 2180.1000 1805.2000 2181.7000 1805.6800 ;
        RECT 2180.1000 1810.6400 2181.7000 1811.1200 ;
        RECT 2180.1000 1816.0800 2181.7000 1816.5600 ;
        RECT 2180.1000 1794.3200 2181.7000 1794.8000 ;
        RECT 2180.1000 1799.7600 2181.7000 1800.2400 ;
        RECT 2135.1000 1875.9200 2136.7000 1876.4000 ;
        RECT 2135.1000 1881.3600 2136.7000 1881.8400 ;
        RECT 2135.1000 1886.8000 2136.7000 1887.2800 ;
        RECT 2090.1000 1875.9200 2091.7000 1876.4000 ;
        RECT 2090.1000 1881.3600 2091.7000 1881.8400 ;
        RECT 2090.1000 1886.8000 2091.7000 1887.2800 ;
        RECT 2135.1000 1865.0400 2136.7000 1865.5200 ;
        RECT 2135.1000 1870.4800 2136.7000 1870.9600 ;
        RECT 2135.1000 1848.7200 2136.7000 1849.2000 ;
        RECT 2135.1000 1854.1600 2136.7000 1854.6400 ;
        RECT 2135.1000 1859.6000 2136.7000 1860.0800 ;
        RECT 2090.1000 1865.0400 2091.7000 1865.5200 ;
        RECT 2090.1000 1870.4800 2091.7000 1870.9600 ;
        RECT 2090.1000 1848.7200 2091.7000 1849.2000 ;
        RECT 2090.1000 1854.1600 2091.7000 1854.6400 ;
        RECT 2090.1000 1859.6000 2091.7000 1860.0800 ;
        RECT 2045.1000 1875.9200 2046.7000 1876.4000 ;
        RECT 2045.1000 1881.3600 2046.7000 1881.8400 ;
        RECT 2033.3400 1881.3600 2036.3400 1881.8400 ;
        RECT 2033.3400 1875.9200 2036.3400 1876.4000 ;
        RECT 2033.3400 1886.8000 2036.3400 1887.2800 ;
        RECT 2045.1000 1886.8000 2046.7000 1887.2800 ;
        RECT 2045.1000 1865.0400 2046.7000 1865.5200 ;
        RECT 2045.1000 1870.4800 2046.7000 1870.9600 ;
        RECT 2033.3400 1870.4800 2036.3400 1870.9600 ;
        RECT 2033.3400 1865.0400 2036.3400 1865.5200 ;
        RECT 2045.1000 1848.7200 2046.7000 1849.2000 ;
        RECT 2045.1000 1854.1600 2046.7000 1854.6400 ;
        RECT 2033.3400 1854.1600 2036.3400 1854.6400 ;
        RECT 2033.3400 1848.7200 2036.3400 1849.2000 ;
        RECT 2033.3400 1859.6000 2036.3400 1860.0800 ;
        RECT 2045.1000 1859.6000 2046.7000 1860.0800 ;
        RECT 2135.1000 1832.4000 2136.7000 1832.8800 ;
        RECT 2135.1000 1837.8400 2136.7000 1838.3200 ;
        RECT 2135.1000 1843.2800 2136.7000 1843.7600 ;
        RECT 2135.1000 1821.5200 2136.7000 1822.0000 ;
        RECT 2135.1000 1826.9600 2136.7000 1827.4400 ;
        RECT 2090.1000 1832.4000 2091.7000 1832.8800 ;
        RECT 2090.1000 1837.8400 2091.7000 1838.3200 ;
        RECT 2090.1000 1843.2800 2091.7000 1843.7600 ;
        RECT 2090.1000 1821.5200 2091.7000 1822.0000 ;
        RECT 2090.1000 1826.9600 2091.7000 1827.4400 ;
        RECT 2135.1000 1805.2000 2136.7000 1805.6800 ;
        RECT 2135.1000 1810.6400 2136.7000 1811.1200 ;
        RECT 2135.1000 1816.0800 2136.7000 1816.5600 ;
        RECT 2135.1000 1794.3200 2136.7000 1794.8000 ;
        RECT 2135.1000 1799.7600 2136.7000 1800.2400 ;
        RECT 2090.1000 1805.2000 2091.7000 1805.6800 ;
        RECT 2090.1000 1810.6400 2091.7000 1811.1200 ;
        RECT 2090.1000 1816.0800 2091.7000 1816.5600 ;
        RECT 2090.1000 1794.3200 2091.7000 1794.8000 ;
        RECT 2090.1000 1799.7600 2091.7000 1800.2400 ;
        RECT 2045.1000 1832.4000 2046.7000 1832.8800 ;
        RECT 2045.1000 1837.8400 2046.7000 1838.3200 ;
        RECT 2045.1000 1843.2800 2046.7000 1843.7600 ;
        RECT 2033.3400 1832.4000 2036.3400 1832.8800 ;
        RECT 2033.3400 1837.8400 2036.3400 1838.3200 ;
        RECT 2033.3400 1843.2800 2036.3400 1843.7600 ;
        RECT 2045.1000 1821.5200 2046.7000 1822.0000 ;
        RECT 2045.1000 1826.9600 2046.7000 1827.4400 ;
        RECT 2033.3400 1821.5200 2036.3400 1822.0000 ;
        RECT 2033.3400 1826.9600 2036.3400 1827.4400 ;
        RECT 2045.1000 1805.2000 2046.7000 1805.6800 ;
        RECT 2045.1000 1810.6400 2046.7000 1811.1200 ;
        RECT 2045.1000 1816.0800 2046.7000 1816.5600 ;
        RECT 2033.3400 1805.2000 2036.3400 1805.6800 ;
        RECT 2033.3400 1810.6400 2036.3400 1811.1200 ;
        RECT 2033.3400 1816.0800 2036.3400 1816.5600 ;
        RECT 2045.1000 1794.3200 2046.7000 1794.8000 ;
        RECT 2045.1000 1799.7600 2046.7000 1800.2400 ;
        RECT 2033.3400 1794.3200 2036.3400 1794.8000 ;
        RECT 2033.3400 1799.7600 2036.3400 1800.2400 ;
        RECT 2237.4400 1778.0000 2240.4400 1778.4800 ;
        RECT 2237.4400 1783.4400 2240.4400 1783.9200 ;
        RECT 2237.4400 1788.8800 2240.4400 1789.3600 ;
        RECT 2225.1000 1778.0000 2226.7000 1778.4800 ;
        RECT 2225.1000 1783.4400 2226.7000 1783.9200 ;
        RECT 2225.1000 1788.8800 2226.7000 1789.3600 ;
        RECT 2237.4400 1767.1200 2240.4400 1767.6000 ;
        RECT 2237.4400 1772.5600 2240.4400 1773.0400 ;
        RECT 2225.1000 1767.1200 2226.7000 1767.6000 ;
        RECT 2225.1000 1772.5600 2226.7000 1773.0400 ;
        RECT 2237.4400 1750.8000 2240.4400 1751.2800 ;
        RECT 2237.4400 1756.2400 2240.4400 1756.7200 ;
        RECT 2237.4400 1761.6800 2240.4400 1762.1600 ;
        RECT 2225.1000 1750.8000 2226.7000 1751.2800 ;
        RECT 2225.1000 1756.2400 2226.7000 1756.7200 ;
        RECT 2225.1000 1761.6800 2226.7000 1762.1600 ;
        RECT 2237.4400 1739.9200 2240.4400 1740.4000 ;
        RECT 2237.4400 1745.3600 2240.4400 1745.8400 ;
        RECT 2225.1000 1739.9200 2226.7000 1740.4000 ;
        RECT 2225.1000 1745.3600 2226.7000 1745.8400 ;
        RECT 2180.1000 1778.0000 2181.7000 1778.4800 ;
        RECT 2180.1000 1783.4400 2181.7000 1783.9200 ;
        RECT 2180.1000 1788.8800 2181.7000 1789.3600 ;
        RECT 2180.1000 1767.1200 2181.7000 1767.6000 ;
        RECT 2180.1000 1772.5600 2181.7000 1773.0400 ;
        RECT 2180.1000 1750.8000 2181.7000 1751.2800 ;
        RECT 2180.1000 1756.2400 2181.7000 1756.7200 ;
        RECT 2180.1000 1761.6800 2181.7000 1762.1600 ;
        RECT 2180.1000 1739.9200 2181.7000 1740.4000 ;
        RECT 2180.1000 1745.3600 2181.7000 1745.8400 ;
        RECT 2237.4400 1723.6000 2240.4400 1724.0800 ;
        RECT 2237.4400 1729.0400 2240.4400 1729.5200 ;
        RECT 2237.4400 1734.4800 2240.4400 1734.9600 ;
        RECT 2225.1000 1723.6000 2226.7000 1724.0800 ;
        RECT 2225.1000 1729.0400 2226.7000 1729.5200 ;
        RECT 2225.1000 1734.4800 2226.7000 1734.9600 ;
        RECT 2237.4400 1712.7200 2240.4400 1713.2000 ;
        RECT 2237.4400 1718.1600 2240.4400 1718.6400 ;
        RECT 2225.1000 1712.7200 2226.7000 1713.2000 ;
        RECT 2225.1000 1718.1600 2226.7000 1718.6400 ;
        RECT 2237.4400 1696.4000 2240.4400 1696.8800 ;
        RECT 2237.4400 1701.8400 2240.4400 1702.3200 ;
        RECT 2237.4400 1707.2800 2240.4400 1707.7600 ;
        RECT 2225.1000 1696.4000 2226.7000 1696.8800 ;
        RECT 2225.1000 1701.8400 2226.7000 1702.3200 ;
        RECT 2225.1000 1707.2800 2226.7000 1707.7600 ;
        RECT 2237.4400 1690.9600 2240.4400 1691.4400 ;
        RECT 2225.1000 1690.9600 2226.7000 1691.4400 ;
        RECT 2180.1000 1723.6000 2181.7000 1724.0800 ;
        RECT 2180.1000 1729.0400 2181.7000 1729.5200 ;
        RECT 2180.1000 1734.4800 2181.7000 1734.9600 ;
        RECT 2180.1000 1712.7200 2181.7000 1713.2000 ;
        RECT 2180.1000 1718.1600 2181.7000 1718.6400 ;
        RECT 2180.1000 1696.4000 2181.7000 1696.8800 ;
        RECT 2180.1000 1701.8400 2181.7000 1702.3200 ;
        RECT 2180.1000 1707.2800 2181.7000 1707.7600 ;
        RECT 2180.1000 1690.9600 2181.7000 1691.4400 ;
        RECT 2135.1000 1778.0000 2136.7000 1778.4800 ;
        RECT 2135.1000 1783.4400 2136.7000 1783.9200 ;
        RECT 2135.1000 1788.8800 2136.7000 1789.3600 ;
        RECT 2135.1000 1767.1200 2136.7000 1767.6000 ;
        RECT 2135.1000 1772.5600 2136.7000 1773.0400 ;
        RECT 2090.1000 1778.0000 2091.7000 1778.4800 ;
        RECT 2090.1000 1783.4400 2091.7000 1783.9200 ;
        RECT 2090.1000 1788.8800 2091.7000 1789.3600 ;
        RECT 2090.1000 1767.1200 2091.7000 1767.6000 ;
        RECT 2090.1000 1772.5600 2091.7000 1773.0400 ;
        RECT 2135.1000 1750.8000 2136.7000 1751.2800 ;
        RECT 2135.1000 1756.2400 2136.7000 1756.7200 ;
        RECT 2135.1000 1761.6800 2136.7000 1762.1600 ;
        RECT 2135.1000 1739.9200 2136.7000 1740.4000 ;
        RECT 2135.1000 1745.3600 2136.7000 1745.8400 ;
        RECT 2090.1000 1750.8000 2091.7000 1751.2800 ;
        RECT 2090.1000 1756.2400 2091.7000 1756.7200 ;
        RECT 2090.1000 1761.6800 2091.7000 1762.1600 ;
        RECT 2090.1000 1739.9200 2091.7000 1740.4000 ;
        RECT 2090.1000 1745.3600 2091.7000 1745.8400 ;
        RECT 2045.1000 1778.0000 2046.7000 1778.4800 ;
        RECT 2045.1000 1783.4400 2046.7000 1783.9200 ;
        RECT 2045.1000 1788.8800 2046.7000 1789.3600 ;
        RECT 2033.3400 1778.0000 2036.3400 1778.4800 ;
        RECT 2033.3400 1783.4400 2036.3400 1783.9200 ;
        RECT 2033.3400 1788.8800 2036.3400 1789.3600 ;
        RECT 2045.1000 1767.1200 2046.7000 1767.6000 ;
        RECT 2045.1000 1772.5600 2046.7000 1773.0400 ;
        RECT 2033.3400 1767.1200 2036.3400 1767.6000 ;
        RECT 2033.3400 1772.5600 2036.3400 1773.0400 ;
        RECT 2045.1000 1750.8000 2046.7000 1751.2800 ;
        RECT 2045.1000 1756.2400 2046.7000 1756.7200 ;
        RECT 2045.1000 1761.6800 2046.7000 1762.1600 ;
        RECT 2033.3400 1750.8000 2036.3400 1751.2800 ;
        RECT 2033.3400 1756.2400 2036.3400 1756.7200 ;
        RECT 2033.3400 1761.6800 2036.3400 1762.1600 ;
        RECT 2045.1000 1739.9200 2046.7000 1740.4000 ;
        RECT 2045.1000 1745.3600 2046.7000 1745.8400 ;
        RECT 2033.3400 1739.9200 2036.3400 1740.4000 ;
        RECT 2033.3400 1745.3600 2036.3400 1745.8400 ;
        RECT 2135.1000 1723.6000 2136.7000 1724.0800 ;
        RECT 2135.1000 1729.0400 2136.7000 1729.5200 ;
        RECT 2135.1000 1734.4800 2136.7000 1734.9600 ;
        RECT 2135.1000 1712.7200 2136.7000 1713.2000 ;
        RECT 2135.1000 1718.1600 2136.7000 1718.6400 ;
        RECT 2090.1000 1723.6000 2091.7000 1724.0800 ;
        RECT 2090.1000 1729.0400 2091.7000 1729.5200 ;
        RECT 2090.1000 1734.4800 2091.7000 1734.9600 ;
        RECT 2090.1000 1712.7200 2091.7000 1713.2000 ;
        RECT 2090.1000 1718.1600 2091.7000 1718.6400 ;
        RECT 2135.1000 1696.4000 2136.7000 1696.8800 ;
        RECT 2135.1000 1701.8400 2136.7000 1702.3200 ;
        RECT 2135.1000 1707.2800 2136.7000 1707.7600 ;
        RECT 2135.1000 1690.9600 2136.7000 1691.4400 ;
        RECT 2090.1000 1696.4000 2091.7000 1696.8800 ;
        RECT 2090.1000 1701.8400 2091.7000 1702.3200 ;
        RECT 2090.1000 1707.2800 2091.7000 1707.7600 ;
        RECT 2090.1000 1690.9600 2091.7000 1691.4400 ;
        RECT 2045.1000 1723.6000 2046.7000 1724.0800 ;
        RECT 2045.1000 1729.0400 2046.7000 1729.5200 ;
        RECT 2045.1000 1734.4800 2046.7000 1734.9600 ;
        RECT 2033.3400 1723.6000 2036.3400 1724.0800 ;
        RECT 2033.3400 1729.0400 2036.3400 1729.5200 ;
        RECT 2033.3400 1734.4800 2036.3400 1734.9600 ;
        RECT 2045.1000 1712.7200 2046.7000 1713.2000 ;
        RECT 2045.1000 1718.1600 2046.7000 1718.6400 ;
        RECT 2033.3400 1712.7200 2036.3400 1713.2000 ;
        RECT 2033.3400 1718.1600 2036.3400 1718.6400 ;
        RECT 2045.1000 1696.4000 2046.7000 1696.8800 ;
        RECT 2045.1000 1701.8400 2046.7000 1702.3200 ;
        RECT 2045.1000 1707.2800 2046.7000 1707.7600 ;
        RECT 2033.3400 1696.4000 2036.3400 1696.8800 ;
        RECT 2033.3400 1701.8400 2036.3400 1702.3200 ;
        RECT 2033.3400 1707.2800 2036.3400 1707.7600 ;
        RECT 2033.3400 1690.9600 2036.3400 1691.4400 ;
        RECT 2045.1000 1690.9600 2046.7000 1691.4400 ;
        RECT 2033.3400 1895.8700 2240.4400 1898.8700 ;
        RECT 2033.3400 1682.7700 2240.4400 1685.7700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 1453.1300 2226.7000 1669.2300 ;
        RECT 2180.1000 1453.1300 2181.7000 1669.2300 ;
        RECT 2135.1000 1453.1300 2136.7000 1669.2300 ;
        RECT 2090.1000 1453.1300 2091.7000 1669.2300 ;
        RECT 2045.1000 1453.1300 2046.7000 1669.2300 ;
        RECT 2237.4400 1453.1300 2240.4400 1669.2300 ;
        RECT 2033.3400 1453.1300 2036.3400 1669.2300 ;
      LAYER met3 ;
        RECT 2237.4400 1646.2800 2240.4400 1646.7600 ;
        RECT 2237.4400 1651.7200 2240.4400 1652.2000 ;
        RECT 2225.1000 1646.2800 2226.7000 1646.7600 ;
        RECT 2225.1000 1651.7200 2226.7000 1652.2000 ;
        RECT 2237.4400 1657.1600 2240.4400 1657.6400 ;
        RECT 2225.1000 1657.1600 2226.7000 1657.6400 ;
        RECT 2237.4400 1635.4000 2240.4400 1635.8800 ;
        RECT 2237.4400 1640.8400 2240.4400 1641.3200 ;
        RECT 2225.1000 1635.4000 2226.7000 1635.8800 ;
        RECT 2225.1000 1640.8400 2226.7000 1641.3200 ;
        RECT 2237.4400 1619.0800 2240.4400 1619.5600 ;
        RECT 2237.4400 1624.5200 2240.4400 1625.0000 ;
        RECT 2225.1000 1619.0800 2226.7000 1619.5600 ;
        RECT 2225.1000 1624.5200 2226.7000 1625.0000 ;
        RECT 2237.4400 1629.9600 2240.4400 1630.4400 ;
        RECT 2225.1000 1629.9600 2226.7000 1630.4400 ;
        RECT 2180.1000 1646.2800 2181.7000 1646.7600 ;
        RECT 2180.1000 1651.7200 2181.7000 1652.2000 ;
        RECT 2180.1000 1657.1600 2181.7000 1657.6400 ;
        RECT 2180.1000 1635.4000 2181.7000 1635.8800 ;
        RECT 2180.1000 1640.8400 2181.7000 1641.3200 ;
        RECT 2180.1000 1619.0800 2181.7000 1619.5600 ;
        RECT 2180.1000 1624.5200 2181.7000 1625.0000 ;
        RECT 2180.1000 1629.9600 2181.7000 1630.4400 ;
        RECT 2237.4400 1602.7600 2240.4400 1603.2400 ;
        RECT 2237.4400 1608.2000 2240.4400 1608.6800 ;
        RECT 2237.4400 1613.6400 2240.4400 1614.1200 ;
        RECT 2225.1000 1602.7600 2226.7000 1603.2400 ;
        RECT 2225.1000 1608.2000 2226.7000 1608.6800 ;
        RECT 2225.1000 1613.6400 2226.7000 1614.1200 ;
        RECT 2237.4400 1591.8800 2240.4400 1592.3600 ;
        RECT 2237.4400 1597.3200 2240.4400 1597.8000 ;
        RECT 2225.1000 1591.8800 2226.7000 1592.3600 ;
        RECT 2225.1000 1597.3200 2226.7000 1597.8000 ;
        RECT 2237.4400 1575.5600 2240.4400 1576.0400 ;
        RECT 2237.4400 1581.0000 2240.4400 1581.4800 ;
        RECT 2237.4400 1586.4400 2240.4400 1586.9200 ;
        RECT 2225.1000 1575.5600 2226.7000 1576.0400 ;
        RECT 2225.1000 1581.0000 2226.7000 1581.4800 ;
        RECT 2225.1000 1586.4400 2226.7000 1586.9200 ;
        RECT 2237.4400 1564.6800 2240.4400 1565.1600 ;
        RECT 2237.4400 1570.1200 2240.4400 1570.6000 ;
        RECT 2225.1000 1564.6800 2226.7000 1565.1600 ;
        RECT 2225.1000 1570.1200 2226.7000 1570.6000 ;
        RECT 2180.1000 1602.7600 2181.7000 1603.2400 ;
        RECT 2180.1000 1608.2000 2181.7000 1608.6800 ;
        RECT 2180.1000 1613.6400 2181.7000 1614.1200 ;
        RECT 2180.1000 1591.8800 2181.7000 1592.3600 ;
        RECT 2180.1000 1597.3200 2181.7000 1597.8000 ;
        RECT 2180.1000 1575.5600 2181.7000 1576.0400 ;
        RECT 2180.1000 1581.0000 2181.7000 1581.4800 ;
        RECT 2180.1000 1586.4400 2181.7000 1586.9200 ;
        RECT 2180.1000 1564.6800 2181.7000 1565.1600 ;
        RECT 2180.1000 1570.1200 2181.7000 1570.6000 ;
        RECT 2135.1000 1646.2800 2136.7000 1646.7600 ;
        RECT 2135.1000 1651.7200 2136.7000 1652.2000 ;
        RECT 2135.1000 1657.1600 2136.7000 1657.6400 ;
        RECT 2090.1000 1646.2800 2091.7000 1646.7600 ;
        RECT 2090.1000 1651.7200 2091.7000 1652.2000 ;
        RECT 2090.1000 1657.1600 2091.7000 1657.6400 ;
        RECT 2135.1000 1635.4000 2136.7000 1635.8800 ;
        RECT 2135.1000 1640.8400 2136.7000 1641.3200 ;
        RECT 2135.1000 1619.0800 2136.7000 1619.5600 ;
        RECT 2135.1000 1624.5200 2136.7000 1625.0000 ;
        RECT 2135.1000 1629.9600 2136.7000 1630.4400 ;
        RECT 2090.1000 1635.4000 2091.7000 1635.8800 ;
        RECT 2090.1000 1640.8400 2091.7000 1641.3200 ;
        RECT 2090.1000 1619.0800 2091.7000 1619.5600 ;
        RECT 2090.1000 1624.5200 2091.7000 1625.0000 ;
        RECT 2090.1000 1629.9600 2091.7000 1630.4400 ;
        RECT 2045.1000 1646.2800 2046.7000 1646.7600 ;
        RECT 2045.1000 1651.7200 2046.7000 1652.2000 ;
        RECT 2033.3400 1651.7200 2036.3400 1652.2000 ;
        RECT 2033.3400 1646.2800 2036.3400 1646.7600 ;
        RECT 2033.3400 1657.1600 2036.3400 1657.6400 ;
        RECT 2045.1000 1657.1600 2046.7000 1657.6400 ;
        RECT 2045.1000 1635.4000 2046.7000 1635.8800 ;
        RECT 2045.1000 1640.8400 2046.7000 1641.3200 ;
        RECT 2033.3400 1640.8400 2036.3400 1641.3200 ;
        RECT 2033.3400 1635.4000 2036.3400 1635.8800 ;
        RECT 2045.1000 1619.0800 2046.7000 1619.5600 ;
        RECT 2045.1000 1624.5200 2046.7000 1625.0000 ;
        RECT 2033.3400 1624.5200 2036.3400 1625.0000 ;
        RECT 2033.3400 1619.0800 2036.3400 1619.5600 ;
        RECT 2033.3400 1629.9600 2036.3400 1630.4400 ;
        RECT 2045.1000 1629.9600 2046.7000 1630.4400 ;
        RECT 2135.1000 1602.7600 2136.7000 1603.2400 ;
        RECT 2135.1000 1608.2000 2136.7000 1608.6800 ;
        RECT 2135.1000 1613.6400 2136.7000 1614.1200 ;
        RECT 2135.1000 1591.8800 2136.7000 1592.3600 ;
        RECT 2135.1000 1597.3200 2136.7000 1597.8000 ;
        RECT 2090.1000 1602.7600 2091.7000 1603.2400 ;
        RECT 2090.1000 1608.2000 2091.7000 1608.6800 ;
        RECT 2090.1000 1613.6400 2091.7000 1614.1200 ;
        RECT 2090.1000 1591.8800 2091.7000 1592.3600 ;
        RECT 2090.1000 1597.3200 2091.7000 1597.8000 ;
        RECT 2135.1000 1575.5600 2136.7000 1576.0400 ;
        RECT 2135.1000 1581.0000 2136.7000 1581.4800 ;
        RECT 2135.1000 1586.4400 2136.7000 1586.9200 ;
        RECT 2135.1000 1564.6800 2136.7000 1565.1600 ;
        RECT 2135.1000 1570.1200 2136.7000 1570.6000 ;
        RECT 2090.1000 1575.5600 2091.7000 1576.0400 ;
        RECT 2090.1000 1581.0000 2091.7000 1581.4800 ;
        RECT 2090.1000 1586.4400 2091.7000 1586.9200 ;
        RECT 2090.1000 1564.6800 2091.7000 1565.1600 ;
        RECT 2090.1000 1570.1200 2091.7000 1570.6000 ;
        RECT 2045.1000 1602.7600 2046.7000 1603.2400 ;
        RECT 2045.1000 1608.2000 2046.7000 1608.6800 ;
        RECT 2045.1000 1613.6400 2046.7000 1614.1200 ;
        RECT 2033.3400 1602.7600 2036.3400 1603.2400 ;
        RECT 2033.3400 1608.2000 2036.3400 1608.6800 ;
        RECT 2033.3400 1613.6400 2036.3400 1614.1200 ;
        RECT 2045.1000 1591.8800 2046.7000 1592.3600 ;
        RECT 2045.1000 1597.3200 2046.7000 1597.8000 ;
        RECT 2033.3400 1591.8800 2036.3400 1592.3600 ;
        RECT 2033.3400 1597.3200 2036.3400 1597.8000 ;
        RECT 2045.1000 1575.5600 2046.7000 1576.0400 ;
        RECT 2045.1000 1581.0000 2046.7000 1581.4800 ;
        RECT 2045.1000 1586.4400 2046.7000 1586.9200 ;
        RECT 2033.3400 1575.5600 2036.3400 1576.0400 ;
        RECT 2033.3400 1581.0000 2036.3400 1581.4800 ;
        RECT 2033.3400 1586.4400 2036.3400 1586.9200 ;
        RECT 2045.1000 1564.6800 2046.7000 1565.1600 ;
        RECT 2045.1000 1570.1200 2046.7000 1570.6000 ;
        RECT 2033.3400 1564.6800 2036.3400 1565.1600 ;
        RECT 2033.3400 1570.1200 2036.3400 1570.6000 ;
        RECT 2237.4400 1548.3600 2240.4400 1548.8400 ;
        RECT 2237.4400 1553.8000 2240.4400 1554.2800 ;
        RECT 2237.4400 1559.2400 2240.4400 1559.7200 ;
        RECT 2225.1000 1548.3600 2226.7000 1548.8400 ;
        RECT 2225.1000 1553.8000 2226.7000 1554.2800 ;
        RECT 2225.1000 1559.2400 2226.7000 1559.7200 ;
        RECT 2237.4400 1537.4800 2240.4400 1537.9600 ;
        RECT 2237.4400 1542.9200 2240.4400 1543.4000 ;
        RECT 2225.1000 1537.4800 2226.7000 1537.9600 ;
        RECT 2225.1000 1542.9200 2226.7000 1543.4000 ;
        RECT 2237.4400 1521.1600 2240.4400 1521.6400 ;
        RECT 2237.4400 1526.6000 2240.4400 1527.0800 ;
        RECT 2237.4400 1532.0400 2240.4400 1532.5200 ;
        RECT 2225.1000 1521.1600 2226.7000 1521.6400 ;
        RECT 2225.1000 1526.6000 2226.7000 1527.0800 ;
        RECT 2225.1000 1532.0400 2226.7000 1532.5200 ;
        RECT 2237.4400 1510.2800 2240.4400 1510.7600 ;
        RECT 2237.4400 1515.7200 2240.4400 1516.2000 ;
        RECT 2225.1000 1510.2800 2226.7000 1510.7600 ;
        RECT 2225.1000 1515.7200 2226.7000 1516.2000 ;
        RECT 2180.1000 1548.3600 2181.7000 1548.8400 ;
        RECT 2180.1000 1553.8000 2181.7000 1554.2800 ;
        RECT 2180.1000 1559.2400 2181.7000 1559.7200 ;
        RECT 2180.1000 1537.4800 2181.7000 1537.9600 ;
        RECT 2180.1000 1542.9200 2181.7000 1543.4000 ;
        RECT 2180.1000 1521.1600 2181.7000 1521.6400 ;
        RECT 2180.1000 1526.6000 2181.7000 1527.0800 ;
        RECT 2180.1000 1532.0400 2181.7000 1532.5200 ;
        RECT 2180.1000 1510.2800 2181.7000 1510.7600 ;
        RECT 2180.1000 1515.7200 2181.7000 1516.2000 ;
        RECT 2237.4400 1493.9600 2240.4400 1494.4400 ;
        RECT 2237.4400 1499.4000 2240.4400 1499.8800 ;
        RECT 2237.4400 1504.8400 2240.4400 1505.3200 ;
        RECT 2225.1000 1493.9600 2226.7000 1494.4400 ;
        RECT 2225.1000 1499.4000 2226.7000 1499.8800 ;
        RECT 2225.1000 1504.8400 2226.7000 1505.3200 ;
        RECT 2237.4400 1483.0800 2240.4400 1483.5600 ;
        RECT 2237.4400 1488.5200 2240.4400 1489.0000 ;
        RECT 2225.1000 1483.0800 2226.7000 1483.5600 ;
        RECT 2225.1000 1488.5200 2226.7000 1489.0000 ;
        RECT 2237.4400 1466.7600 2240.4400 1467.2400 ;
        RECT 2237.4400 1472.2000 2240.4400 1472.6800 ;
        RECT 2237.4400 1477.6400 2240.4400 1478.1200 ;
        RECT 2225.1000 1466.7600 2226.7000 1467.2400 ;
        RECT 2225.1000 1472.2000 2226.7000 1472.6800 ;
        RECT 2225.1000 1477.6400 2226.7000 1478.1200 ;
        RECT 2237.4400 1461.3200 2240.4400 1461.8000 ;
        RECT 2225.1000 1461.3200 2226.7000 1461.8000 ;
        RECT 2180.1000 1493.9600 2181.7000 1494.4400 ;
        RECT 2180.1000 1499.4000 2181.7000 1499.8800 ;
        RECT 2180.1000 1504.8400 2181.7000 1505.3200 ;
        RECT 2180.1000 1483.0800 2181.7000 1483.5600 ;
        RECT 2180.1000 1488.5200 2181.7000 1489.0000 ;
        RECT 2180.1000 1466.7600 2181.7000 1467.2400 ;
        RECT 2180.1000 1472.2000 2181.7000 1472.6800 ;
        RECT 2180.1000 1477.6400 2181.7000 1478.1200 ;
        RECT 2180.1000 1461.3200 2181.7000 1461.8000 ;
        RECT 2135.1000 1548.3600 2136.7000 1548.8400 ;
        RECT 2135.1000 1553.8000 2136.7000 1554.2800 ;
        RECT 2135.1000 1559.2400 2136.7000 1559.7200 ;
        RECT 2135.1000 1537.4800 2136.7000 1537.9600 ;
        RECT 2135.1000 1542.9200 2136.7000 1543.4000 ;
        RECT 2090.1000 1548.3600 2091.7000 1548.8400 ;
        RECT 2090.1000 1553.8000 2091.7000 1554.2800 ;
        RECT 2090.1000 1559.2400 2091.7000 1559.7200 ;
        RECT 2090.1000 1537.4800 2091.7000 1537.9600 ;
        RECT 2090.1000 1542.9200 2091.7000 1543.4000 ;
        RECT 2135.1000 1521.1600 2136.7000 1521.6400 ;
        RECT 2135.1000 1526.6000 2136.7000 1527.0800 ;
        RECT 2135.1000 1532.0400 2136.7000 1532.5200 ;
        RECT 2135.1000 1510.2800 2136.7000 1510.7600 ;
        RECT 2135.1000 1515.7200 2136.7000 1516.2000 ;
        RECT 2090.1000 1521.1600 2091.7000 1521.6400 ;
        RECT 2090.1000 1526.6000 2091.7000 1527.0800 ;
        RECT 2090.1000 1532.0400 2091.7000 1532.5200 ;
        RECT 2090.1000 1510.2800 2091.7000 1510.7600 ;
        RECT 2090.1000 1515.7200 2091.7000 1516.2000 ;
        RECT 2045.1000 1548.3600 2046.7000 1548.8400 ;
        RECT 2045.1000 1553.8000 2046.7000 1554.2800 ;
        RECT 2045.1000 1559.2400 2046.7000 1559.7200 ;
        RECT 2033.3400 1548.3600 2036.3400 1548.8400 ;
        RECT 2033.3400 1553.8000 2036.3400 1554.2800 ;
        RECT 2033.3400 1559.2400 2036.3400 1559.7200 ;
        RECT 2045.1000 1537.4800 2046.7000 1537.9600 ;
        RECT 2045.1000 1542.9200 2046.7000 1543.4000 ;
        RECT 2033.3400 1537.4800 2036.3400 1537.9600 ;
        RECT 2033.3400 1542.9200 2036.3400 1543.4000 ;
        RECT 2045.1000 1521.1600 2046.7000 1521.6400 ;
        RECT 2045.1000 1526.6000 2046.7000 1527.0800 ;
        RECT 2045.1000 1532.0400 2046.7000 1532.5200 ;
        RECT 2033.3400 1521.1600 2036.3400 1521.6400 ;
        RECT 2033.3400 1526.6000 2036.3400 1527.0800 ;
        RECT 2033.3400 1532.0400 2036.3400 1532.5200 ;
        RECT 2045.1000 1510.2800 2046.7000 1510.7600 ;
        RECT 2045.1000 1515.7200 2046.7000 1516.2000 ;
        RECT 2033.3400 1510.2800 2036.3400 1510.7600 ;
        RECT 2033.3400 1515.7200 2036.3400 1516.2000 ;
        RECT 2135.1000 1493.9600 2136.7000 1494.4400 ;
        RECT 2135.1000 1499.4000 2136.7000 1499.8800 ;
        RECT 2135.1000 1504.8400 2136.7000 1505.3200 ;
        RECT 2135.1000 1483.0800 2136.7000 1483.5600 ;
        RECT 2135.1000 1488.5200 2136.7000 1489.0000 ;
        RECT 2090.1000 1493.9600 2091.7000 1494.4400 ;
        RECT 2090.1000 1499.4000 2091.7000 1499.8800 ;
        RECT 2090.1000 1504.8400 2091.7000 1505.3200 ;
        RECT 2090.1000 1483.0800 2091.7000 1483.5600 ;
        RECT 2090.1000 1488.5200 2091.7000 1489.0000 ;
        RECT 2135.1000 1466.7600 2136.7000 1467.2400 ;
        RECT 2135.1000 1472.2000 2136.7000 1472.6800 ;
        RECT 2135.1000 1477.6400 2136.7000 1478.1200 ;
        RECT 2135.1000 1461.3200 2136.7000 1461.8000 ;
        RECT 2090.1000 1466.7600 2091.7000 1467.2400 ;
        RECT 2090.1000 1472.2000 2091.7000 1472.6800 ;
        RECT 2090.1000 1477.6400 2091.7000 1478.1200 ;
        RECT 2090.1000 1461.3200 2091.7000 1461.8000 ;
        RECT 2045.1000 1493.9600 2046.7000 1494.4400 ;
        RECT 2045.1000 1499.4000 2046.7000 1499.8800 ;
        RECT 2045.1000 1504.8400 2046.7000 1505.3200 ;
        RECT 2033.3400 1493.9600 2036.3400 1494.4400 ;
        RECT 2033.3400 1499.4000 2036.3400 1499.8800 ;
        RECT 2033.3400 1504.8400 2036.3400 1505.3200 ;
        RECT 2045.1000 1483.0800 2046.7000 1483.5600 ;
        RECT 2045.1000 1488.5200 2046.7000 1489.0000 ;
        RECT 2033.3400 1483.0800 2036.3400 1483.5600 ;
        RECT 2033.3400 1488.5200 2036.3400 1489.0000 ;
        RECT 2045.1000 1466.7600 2046.7000 1467.2400 ;
        RECT 2045.1000 1472.2000 2046.7000 1472.6800 ;
        RECT 2045.1000 1477.6400 2046.7000 1478.1200 ;
        RECT 2033.3400 1466.7600 2036.3400 1467.2400 ;
        RECT 2033.3400 1472.2000 2036.3400 1472.6800 ;
        RECT 2033.3400 1477.6400 2036.3400 1478.1200 ;
        RECT 2033.3400 1461.3200 2036.3400 1461.8000 ;
        RECT 2045.1000 1461.3200 2046.7000 1461.8000 ;
        RECT 2033.3400 1666.2300 2240.4400 1669.2300 ;
        RECT 2033.3400 1453.1300 2240.4400 1456.1300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 1223.4900 2226.7000 1439.5900 ;
        RECT 2180.1000 1223.4900 2181.7000 1439.5900 ;
        RECT 2135.1000 1223.4900 2136.7000 1439.5900 ;
        RECT 2090.1000 1223.4900 2091.7000 1439.5900 ;
        RECT 2045.1000 1223.4900 2046.7000 1439.5900 ;
        RECT 2237.4400 1223.4900 2240.4400 1439.5900 ;
        RECT 2033.3400 1223.4900 2036.3400 1439.5900 ;
      LAYER met3 ;
        RECT 2237.4400 1416.6400 2240.4400 1417.1200 ;
        RECT 2237.4400 1422.0800 2240.4400 1422.5600 ;
        RECT 2225.1000 1416.6400 2226.7000 1417.1200 ;
        RECT 2225.1000 1422.0800 2226.7000 1422.5600 ;
        RECT 2237.4400 1427.5200 2240.4400 1428.0000 ;
        RECT 2225.1000 1427.5200 2226.7000 1428.0000 ;
        RECT 2237.4400 1405.7600 2240.4400 1406.2400 ;
        RECT 2237.4400 1411.2000 2240.4400 1411.6800 ;
        RECT 2225.1000 1405.7600 2226.7000 1406.2400 ;
        RECT 2225.1000 1411.2000 2226.7000 1411.6800 ;
        RECT 2237.4400 1389.4400 2240.4400 1389.9200 ;
        RECT 2237.4400 1394.8800 2240.4400 1395.3600 ;
        RECT 2225.1000 1389.4400 2226.7000 1389.9200 ;
        RECT 2225.1000 1394.8800 2226.7000 1395.3600 ;
        RECT 2237.4400 1400.3200 2240.4400 1400.8000 ;
        RECT 2225.1000 1400.3200 2226.7000 1400.8000 ;
        RECT 2180.1000 1416.6400 2181.7000 1417.1200 ;
        RECT 2180.1000 1422.0800 2181.7000 1422.5600 ;
        RECT 2180.1000 1427.5200 2181.7000 1428.0000 ;
        RECT 2180.1000 1405.7600 2181.7000 1406.2400 ;
        RECT 2180.1000 1411.2000 2181.7000 1411.6800 ;
        RECT 2180.1000 1389.4400 2181.7000 1389.9200 ;
        RECT 2180.1000 1394.8800 2181.7000 1395.3600 ;
        RECT 2180.1000 1400.3200 2181.7000 1400.8000 ;
        RECT 2237.4400 1373.1200 2240.4400 1373.6000 ;
        RECT 2237.4400 1378.5600 2240.4400 1379.0400 ;
        RECT 2237.4400 1384.0000 2240.4400 1384.4800 ;
        RECT 2225.1000 1373.1200 2226.7000 1373.6000 ;
        RECT 2225.1000 1378.5600 2226.7000 1379.0400 ;
        RECT 2225.1000 1384.0000 2226.7000 1384.4800 ;
        RECT 2237.4400 1362.2400 2240.4400 1362.7200 ;
        RECT 2237.4400 1367.6800 2240.4400 1368.1600 ;
        RECT 2225.1000 1362.2400 2226.7000 1362.7200 ;
        RECT 2225.1000 1367.6800 2226.7000 1368.1600 ;
        RECT 2237.4400 1345.9200 2240.4400 1346.4000 ;
        RECT 2237.4400 1351.3600 2240.4400 1351.8400 ;
        RECT 2237.4400 1356.8000 2240.4400 1357.2800 ;
        RECT 2225.1000 1345.9200 2226.7000 1346.4000 ;
        RECT 2225.1000 1351.3600 2226.7000 1351.8400 ;
        RECT 2225.1000 1356.8000 2226.7000 1357.2800 ;
        RECT 2237.4400 1335.0400 2240.4400 1335.5200 ;
        RECT 2237.4400 1340.4800 2240.4400 1340.9600 ;
        RECT 2225.1000 1335.0400 2226.7000 1335.5200 ;
        RECT 2225.1000 1340.4800 2226.7000 1340.9600 ;
        RECT 2180.1000 1373.1200 2181.7000 1373.6000 ;
        RECT 2180.1000 1378.5600 2181.7000 1379.0400 ;
        RECT 2180.1000 1384.0000 2181.7000 1384.4800 ;
        RECT 2180.1000 1362.2400 2181.7000 1362.7200 ;
        RECT 2180.1000 1367.6800 2181.7000 1368.1600 ;
        RECT 2180.1000 1345.9200 2181.7000 1346.4000 ;
        RECT 2180.1000 1351.3600 2181.7000 1351.8400 ;
        RECT 2180.1000 1356.8000 2181.7000 1357.2800 ;
        RECT 2180.1000 1335.0400 2181.7000 1335.5200 ;
        RECT 2180.1000 1340.4800 2181.7000 1340.9600 ;
        RECT 2135.1000 1416.6400 2136.7000 1417.1200 ;
        RECT 2135.1000 1422.0800 2136.7000 1422.5600 ;
        RECT 2135.1000 1427.5200 2136.7000 1428.0000 ;
        RECT 2090.1000 1416.6400 2091.7000 1417.1200 ;
        RECT 2090.1000 1422.0800 2091.7000 1422.5600 ;
        RECT 2090.1000 1427.5200 2091.7000 1428.0000 ;
        RECT 2135.1000 1405.7600 2136.7000 1406.2400 ;
        RECT 2135.1000 1411.2000 2136.7000 1411.6800 ;
        RECT 2135.1000 1389.4400 2136.7000 1389.9200 ;
        RECT 2135.1000 1394.8800 2136.7000 1395.3600 ;
        RECT 2135.1000 1400.3200 2136.7000 1400.8000 ;
        RECT 2090.1000 1405.7600 2091.7000 1406.2400 ;
        RECT 2090.1000 1411.2000 2091.7000 1411.6800 ;
        RECT 2090.1000 1389.4400 2091.7000 1389.9200 ;
        RECT 2090.1000 1394.8800 2091.7000 1395.3600 ;
        RECT 2090.1000 1400.3200 2091.7000 1400.8000 ;
        RECT 2045.1000 1416.6400 2046.7000 1417.1200 ;
        RECT 2045.1000 1422.0800 2046.7000 1422.5600 ;
        RECT 2033.3400 1422.0800 2036.3400 1422.5600 ;
        RECT 2033.3400 1416.6400 2036.3400 1417.1200 ;
        RECT 2033.3400 1427.5200 2036.3400 1428.0000 ;
        RECT 2045.1000 1427.5200 2046.7000 1428.0000 ;
        RECT 2045.1000 1405.7600 2046.7000 1406.2400 ;
        RECT 2045.1000 1411.2000 2046.7000 1411.6800 ;
        RECT 2033.3400 1411.2000 2036.3400 1411.6800 ;
        RECT 2033.3400 1405.7600 2036.3400 1406.2400 ;
        RECT 2045.1000 1389.4400 2046.7000 1389.9200 ;
        RECT 2045.1000 1394.8800 2046.7000 1395.3600 ;
        RECT 2033.3400 1394.8800 2036.3400 1395.3600 ;
        RECT 2033.3400 1389.4400 2036.3400 1389.9200 ;
        RECT 2033.3400 1400.3200 2036.3400 1400.8000 ;
        RECT 2045.1000 1400.3200 2046.7000 1400.8000 ;
        RECT 2135.1000 1373.1200 2136.7000 1373.6000 ;
        RECT 2135.1000 1378.5600 2136.7000 1379.0400 ;
        RECT 2135.1000 1384.0000 2136.7000 1384.4800 ;
        RECT 2135.1000 1362.2400 2136.7000 1362.7200 ;
        RECT 2135.1000 1367.6800 2136.7000 1368.1600 ;
        RECT 2090.1000 1373.1200 2091.7000 1373.6000 ;
        RECT 2090.1000 1378.5600 2091.7000 1379.0400 ;
        RECT 2090.1000 1384.0000 2091.7000 1384.4800 ;
        RECT 2090.1000 1362.2400 2091.7000 1362.7200 ;
        RECT 2090.1000 1367.6800 2091.7000 1368.1600 ;
        RECT 2135.1000 1345.9200 2136.7000 1346.4000 ;
        RECT 2135.1000 1351.3600 2136.7000 1351.8400 ;
        RECT 2135.1000 1356.8000 2136.7000 1357.2800 ;
        RECT 2135.1000 1335.0400 2136.7000 1335.5200 ;
        RECT 2135.1000 1340.4800 2136.7000 1340.9600 ;
        RECT 2090.1000 1345.9200 2091.7000 1346.4000 ;
        RECT 2090.1000 1351.3600 2091.7000 1351.8400 ;
        RECT 2090.1000 1356.8000 2091.7000 1357.2800 ;
        RECT 2090.1000 1335.0400 2091.7000 1335.5200 ;
        RECT 2090.1000 1340.4800 2091.7000 1340.9600 ;
        RECT 2045.1000 1373.1200 2046.7000 1373.6000 ;
        RECT 2045.1000 1378.5600 2046.7000 1379.0400 ;
        RECT 2045.1000 1384.0000 2046.7000 1384.4800 ;
        RECT 2033.3400 1373.1200 2036.3400 1373.6000 ;
        RECT 2033.3400 1378.5600 2036.3400 1379.0400 ;
        RECT 2033.3400 1384.0000 2036.3400 1384.4800 ;
        RECT 2045.1000 1362.2400 2046.7000 1362.7200 ;
        RECT 2045.1000 1367.6800 2046.7000 1368.1600 ;
        RECT 2033.3400 1362.2400 2036.3400 1362.7200 ;
        RECT 2033.3400 1367.6800 2036.3400 1368.1600 ;
        RECT 2045.1000 1345.9200 2046.7000 1346.4000 ;
        RECT 2045.1000 1351.3600 2046.7000 1351.8400 ;
        RECT 2045.1000 1356.8000 2046.7000 1357.2800 ;
        RECT 2033.3400 1345.9200 2036.3400 1346.4000 ;
        RECT 2033.3400 1351.3600 2036.3400 1351.8400 ;
        RECT 2033.3400 1356.8000 2036.3400 1357.2800 ;
        RECT 2045.1000 1335.0400 2046.7000 1335.5200 ;
        RECT 2045.1000 1340.4800 2046.7000 1340.9600 ;
        RECT 2033.3400 1335.0400 2036.3400 1335.5200 ;
        RECT 2033.3400 1340.4800 2036.3400 1340.9600 ;
        RECT 2237.4400 1318.7200 2240.4400 1319.2000 ;
        RECT 2237.4400 1324.1600 2240.4400 1324.6400 ;
        RECT 2237.4400 1329.6000 2240.4400 1330.0800 ;
        RECT 2225.1000 1318.7200 2226.7000 1319.2000 ;
        RECT 2225.1000 1324.1600 2226.7000 1324.6400 ;
        RECT 2225.1000 1329.6000 2226.7000 1330.0800 ;
        RECT 2237.4400 1307.8400 2240.4400 1308.3200 ;
        RECT 2237.4400 1313.2800 2240.4400 1313.7600 ;
        RECT 2225.1000 1307.8400 2226.7000 1308.3200 ;
        RECT 2225.1000 1313.2800 2226.7000 1313.7600 ;
        RECT 2237.4400 1291.5200 2240.4400 1292.0000 ;
        RECT 2237.4400 1296.9600 2240.4400 1297.4400 ;
        RECT 2237.4400 1302.4000 2240.4400 1302.8800 ;
        RECT 2225.1000 1291.5200 2226.7000 1292.0000 ;
        RECT 2225.1000 1296.9600 2226.7000 1297.4400 ;
        RECT 2225.1000 1302.4000 2226.7000 1302.8800 ;
        RECT 2237.4400 1280.6400 2240.4400 1281.1200 ;
        RECT 2237.4400 1286.0800 2240.4400 1286.5600 ;
        RECT 2225.1000 1280.6400 2226.7000 1281.1200 ;
        RECT 2225.1000 1286.0800 2226.7000 1286.5600 ;
        RECT 2180.1000 1318.7200 2181.7000 1319.2000 ;
        RECT 2180.1000 1324.1600 2181.7000 1324.6400 ;
        RECT 2180.1000 1329.6000 2181.7000 1330.0800 ;
        RECT 2180.1000 1307.8400 2181.7000 1308.3200 ;
        RECT 2180.1000 1313.2800 2181.7000 1313.7600 ;
        RECT 2180.1000 1291.5200 2181.7000 1292.0000 ;
        RECT 2180.1000 1296.9600 2181.7000 1297.4400 ;
        RECT 2180.1000 1302.4000 2181.7000 1302.8800 ;
        RECT 2180.1000 1280.6400 2181.7000 1281.1200 ;
        RECT 2180.1000 1286.0800 2181.7000 1286.5600 ;
        RECT 2237.4400 1264.3200 2240.4400 1264.8000 ;
        RECT 2237.4400 1269.7600 2240.4400 1270.2400 ;
        RECT 2237.4400 1275.2000 2240.4400 1275.6800 ;
        RECT 2225.1000 1264.3200 2226.7000 1264.8000 ;
        RECT 2225.1000 1269.7600 2226.7000 1270.2400 ;
        RECT 2225.1000 1275.2000 2226.7000 1275.6800 ;
        RECT 2237.4400 1253.4400 2240.4400 1253.9200 ;
        RECT 2237.4400 1258.8800 2240.4400 1259.3600 ;
        RECT 2225.1000 1253.4400 2226.7000 1253.9200 ;
        RECT 2225.1000 1258.8800 2226.7000 1259.3600 ;
        RECT 2237.4400 1237.1200 2240.4400 1237.6000 ;
        RECT 2237.4400 1242.5600 2240.4400 1243.0400 ;
        RECT 2237.4400 1248.0000 2240.4400 1248.4800 ;
        RECT 2225.1000 1237.1200 2226.7000 1237.6000 ;
        RECT 2225.1000 1242.5600 2226.7000 1243.0400 ;
        RECT 2225.1000 1248.0000 2226.7000 1248.4800 ;
        RECT 2237.4400 1231.6800 2240.4400 1232.1600 ;
        RECT 2225.1000 1231.6800 2226.7000 1232.1600 ;
        RECT 2180.1000 1264.3200 2181.7000 1264.8000 ;
        RECT 2180.1000 1269.7600 2181.7000 1270.2400 ;
        RECT 2180.1000 1275.2000 2181.7000 1275.6800 ;
        RECT 2180.1000 1253.4400 2181.7000 1253.9200 ;
        RECT 2180.1000 1258.8800 2181.7000 1259.3600 ;
        RECT 2180.1000 1237.1200 2181.7000 1237.6000 ;
        RECT 2180.1000 1242.5600 2181.7000 1243.0400 ;
        RECT 2180.1000 1248.0000 2181.7000 1248.4800 ;
        RECT 2180.1000 1231.6800 2181.7000 1232.1600 ;
        RECT 2135.1000 1318.7200 2136.7000 1319.2000 ;
        RECT 2135.1000 1324.1600 2136.7000 1324.6400 ;
        RECT 2135.1000 1329.6000 2136.7000 1330.0800 ;
        RECT 2135.1000 1307.8400 2136.7000 1308.3200 ;
        RECT 2135.1000 1313.2800 2136.7000 1313.7600 ;
        RECT 2090.1000 1318.7200 2091.7000 1319.2000 ;
        RECT 2090.1000 1324.1600 2091.7000 1324.6400 ;
        RECT 2090.1000 1329.6000 2091.7000 1330.0800 ;
        RECT 2090.1000 1307.8400 2091.7000 1308.3200 ;
        RECT 2090.1000 1313.2800 2091.7000 1313.7600 ;
        RECT 2135.1000 1291.5200 2136.7000 1292.0000 ;
        RECT 2135.1000 1296.9600 2136.7000 1297.4400 ;
        RECT 2135.1000 1302.4000 2136.7000 1302.8800 ;
        RECT 2135.1000 1280.6400 2136.7000 1281.1200 ;
        RECT 2135.1000 1286.0800 2136.7000 1286.5600 ;
        RECT 2090.1000 1291.5200 2091.7000 1292.0000 ;
        RECT 2090.1000 1296.9600 2091.7000 1297.4400 ;
        RECT 2090.1000 1302.4000 2091.7000 1302.8800 ;
        RECT 2090.1000 1280.6400 2091.7000 1281.1200 ;
        RECT 2090.1000 1286.0800 2091.7000 1286.5600 ;
        RECT 2045.1000 1318.7200 2046.7000 1319.2000 ;
        RECT 2045.1000 1324.1600 2046.7000 1324.6400 ;
        RECT 2045.1000 1329.6000 2046.7000 1330.0800 ;
        RECT 2033.3400 1318.7200 2036.3400 1319.2000 ;
        RECT 2033.3400 1324.1600 2036.3400 1324.6400 ;
        RECT 2033.3400 1329.6000 2036.3400 1330.0800 ;
        RECT 2045.1000 1307.8400 2046.7000 1308.3200 ;
        RECT 2045.1000 1313.2800 2046.7000 1313.7600 ;
        RECT 2033.3400 1307.8400 2036.3400 1308.3200 ;
        RECT 2033.3400 1313.2800 2036.3400 1313.7600 ;
        RECT 2045.1000 1291.5200 2046.7000 1292.0000 ;
        RECT 2045.1000 1296.9600 2046.7000 1297.4400 ;
        RECT 2045.1000 1302.4000 2046.7000 1302.8800 ;
        RECT 2033.3400 1291.5200 2036.3400 1292.0000 ;
        RECT 2033.3400 1296.9600 2036.3400 1297.4400 ;
        RECT 2033.3400 1302.4000 2036.3400 1302.8800 ;
        RECT 2045.1000 1280.6400 2046.7000 1281.1200 ;
        RECT 2045.1000 1286.0800 2046.7000 1286.5600 ;
        RECT 2033.3400 1280.6400 2036.3400 1281.1200 ;
        RECT 2033.3400 1286.0800 2036.3400 1286.5600 ;
        RECT 2135.1000 1264.3200 2136.7000 1264.8000 ;
        RECT 2135.1000 1269.7600 2136.7000 1270.2400 ;
        RECT 2135.1000 1275.2000 2136.7000 1275.6800 ;
        RECT 2135.1000 1253.4400 2136.7000 1253.9200 ;
        RECT 2135.1000 1258.8800 2136.7000 1259.3600 ;
        RECT 2090.1000 1264.3200 2091.7000 1264.8000 ;
        RECT 2090.1000 1269.7600 2091.7000 1270.2400 ;
        RECT 2090.1000 1275.2000 2091.7000 1275.6800 ;
        RECT 2090.1000 1253.4400 2091.7000 1253.9200 ;
        RECT 2090.1000 1258.8800 2091.7000 1259.3600 ;
        RECT 2135.1000 1237.1200 2136.7000 1237.6000 ;
        RECT 2135.1000 1242.5600 2136.7000 1243.0400 ;
        RECT 2135.1000 1248.0000 2136.7000 1248.4800 ;
        RECT 2135.1000 1231.6800 2136.7000 1232.1600 ;
        RECT 2090.1000 1237.1200 2091.7000 1237.6000 ;
        RECT 2090.1000 1242.5600 2091.7000 1243.0400 ;
        RECT 2090.1000 1248.0000 2091.7000 1248.4800 ;
        RECT 2090.1000 1231.6800 2091.7000 1232.1600 ;
        RECT 2045.1000 1264.3200 2046.7000 1264.8000 ;
        RECT 2045.1000 1269.7600 2046.7000 1270.2400 ;
        RECT 2045.1000 1275.2000 2046.7000 1275.6800 ;
        RECT 2033.3400 1264.3200 2036.3400 1264.8000 ;
        RECT 2033.3400 1269.7600 2036.3400 1270.2400 ;
        RECT 2033.3400 1275.2000 2036.3400 1275.6800 ;
        RECT 2045.1000 1253.4400 2046.7000 1253.9200 ;
        RECT 2045.1000 1258.8800 2046.7000 1259.3600 ;
        RECT 2033.3400 1253.4400 2036.3400 1253.9200 ;
        RECT 2033.3400 1258.8800 2036.3400 1259.3600 ;
        RECT 2045.1000 1237.1200 2046.7000 1237.6000 ;
        RECT 2045.1000 1242.5600 2046.7000 1243.0400 ;
        RECT 2045.1000 1248.0000 2046.7000 1248.4800 ;
        RECT 2033.3400 1237.1200 2036.3400 1237.6000 ;
        RECT 2033.3400 1242.5600 2036.3400 1243.0400 ;
        RECT 2033.3400 1248.0000 2036.3400 1248.4800 ;
        RECT 2033.3400 1231.6800 2036.3400 1232.1600 ;
        RECT 2045.1000 1231.6800 2046.7000 1232.1600 ;
        RECT 2033.3400 1436.5900 2240.4400 1439.5900 ;
        RECT 2033.3400 1223.4900 2240.4400 1226.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 993.8500 2226.7000 1209.9500 ;
        RECT 2180.1000 993.8500 2181.7000 1209.9500 ;
        RECT 2135.1000 993.8500 2136.7000 1209.9500 ;
        RECT 2090.1000 993.8500 2091.7000 1209.9500 ;
        RECT 2045.1000 993.8500 2046.7000 1209.9500 ;
        RECT 2237.4400 993.8500 2240.4400 1209.9500 ;
        RECT 2033.3400 993.8500 2036.3400 1209.9500 ;
      LAYER met3 ;
        RECT 2237.4400 1187.0000 2240.4400 1187.4800 ;
        RECT 2237.4400 1192.4400 2240.4400 1192.9200 ;
        RECT 2225.1000 1187.0000 2226.7000 1187.4800 ;
        RECT 2225.1000 1192.4400 2226.7000 1192.9200 ;
        RECT 2237.4400 1197.8800 2240.4400 1198.3600 ;
        RECT 2225.1000 1197.8800 2226.7000 1198.3600 ;
        RECT 2237.4400 1176.1200 2240.4400 1176.6000 ;
        RECT 2237.4400 1181.5600 2240.4400 1182.0400 ;
        RECT 2225.1000 1176.1200 2226.7000 1176.6000 ;
        RECT 2225.1000 1181.5600 2226.7000 1182.0400 ;
        RECT 2237.4400 1159.8000 2240.4400 1160.2800 ;
        RECT 2237.4400 1165.2400 2240.4400 1165.7200 ;
        RECT 2225.1000 1159.8000 2226.7000 1160.2800 ;
        RECT 2225.1000 1165.2400 2226.7000 1165.7200 ;
        RECT 2237.4400 1170.6800 2240.4400 1171.1600 ;
        RECT 2225.1000 1170.6800 2226.7000 1171.1600 ;
        RECT 2180.1000 1187.0000 2181.7000 1187.4800 ;
        RECT 2180.1000 1192.4400 2181.7000 1192.9200 ;
        RECT 2180.1000 1197.8800 2181.7000 1198.3600 ;
        RECT 2180.1000 1176.1200 2181.7000 1176.6000 ;
        RECT 2180.1000 1181.5600 2181.7000 1182.0400 ;
        RECT 2180.1000 1159.8000 2181.7000 1160.2800 ;
        RECT 2180.1000 1165.2400 2181.7000 1165.7200 ;
        RECT 2180.1000 1170.6800 2181.7000 1171.1600 ;
        RECT 2237.4400 1143.4800 2240.4400 1143.9600 ;
        RECT 2237.4400 1148.9200 2240.4400 1149.4000 ;
        RECT 2237.4400 1154.3600 2240.4400 1154.8400 ;
        RECT 2225.1000 1143.4800 2226.7000 1143.9600 ;
        RECT 2225.1000 1148.9200 2226.7000 1149.4000 ;
        RECT 2225.1000 1154.3600 2226.7000 1154.8400 ;
        RECT 2237.4400 1132.6000 2240.4400 1133.0800 ;
        RECT 2237.4400 1138.0400 2240.4400 1138.5200 ;
        RECT 2225.1000 1132.6000 2226.7000 1133.0800 ;
        RECT 2225.1000 1138.0400 2226.7000 1138.5200 ;
        RECT 2237.4400 1116.2800 2240.4400 1116.7600 ;
        RECT 2237.4400 1121.7200 2240.4400 1122.2000 ;
        RECT 2237.4400 1127.1600 2240.4400 1127.6400 ;
        RECT 2225.1000 1116.2800 2226.7000 1116.7600 ;
        RECT 2225.1000 1121.7200 2226.7000 1122.2000 ;
        RECT 2225.1000 1127.1600 2226.7000 1127.6400 ;
        RECT 2237.4400 1105.4000 2240.4400 1105.8800 ;
        RECT 2237.4400 1110.8400 2240.4400 1111.3200 ;
        RECT 2225.1000 1105.4000 2226.7000 1105.8800 ;
        RECT 2225.1000 1110.8400 2226.7000 1111.3200 ;
        RECT 2180.1000 1143.4800 2181.7000 1143.9600 ;
        RECT 2180.1000 1148.9200 2181.7000 1149.4000 ;
        RECT 2180.1000 1154.3600 2181.7000 1154.8400 ;
        RECT 2180.1000 1132.6000 2181.7000 1133.0800 ;
        RECT 2180.1000 1138.0400 2181.7000 1138.5200 ;
        RECT 2180.1000 1116.2800 2181.7000 1116.7600 ;
        RECT 2180.1000 1121.7200 2181.7000 1122.2000 ;
        RECT 2180.1000 1127.1600 2181.7000 1127.6400 ;
        RECT 2180.1000 1105.4000 2181.7000 1105.8800 ;
        RECT 2180.1000 1110.8400 2181.7000 1111.3200 ;
        RECT 2135.1000 1187.0000 2136.7000 1187.4800 ;
        RECT 2135.1000 1192.4400 2136.7000 1192.9200 ;
        RECT 2135.1000 1197.8800 2136.7000 1198.3600 ;
        RECT 2090.1000 1187.0000 2091.7000 1187.4800 ;
        RECT 2090.1000 1192.4400 2091.7000 1192.9200 ;
        RECT 2090.1000 1197.8800 2091.7000 1198.3600 ;
        RECT 2135.1000 1176.1200 2136.7000 1176.6000 ;
        RECT 2135.1000 1181.5600 2136.7000 1182.0400 ;
        RECT 2135.1000 1159.8000 2136.7000 1160.2800 ;
        RECT 2135.1000 1165.2400 2136.7000 1165.7200 ;
        RECT 2135.1000 1170.6800 2136.7000 1171.1600 ;
        RECT 2090.1000 1176.1200 2091.7000 1176.6000 ;
        RECT 2090.1000 1181.5600 2091.7000 1182.0400 ;
        RECT 2090.1000 1159.8000 2091.7000 1160.2800 ;
        RECT 2090.1000 1165.2400 2091.7000 1165.7200 ;
        RECT 2090.1000 1170.6800 2091.7000 1171.1600 ;
        RECT 2045.1000 1187.0000 2046.7000 1187.4800 ;
        RECT 2045.1000 1192.4400 2046.7000 1192.9200 ;
        RECT 2033.3400 1192.4400 2036.3400 1192.9200 ;
        RECT 2033.3400 1187.0000 2036.3400 1187.4800 ;
        RECT 2033.3400 1197.8800 2036.3400 1198.3600 ;
        RECT 2045.1000 1197.8800 2046.7000 1198.3600 ;
        RECT 2045.1000 1176.1200 2046.7000 1176.6000 ;
        RECT 2045.1000 1181.5600 2046.7000 1182.0400 ;
        RECT 2033.3400 1181.5600 2036.3400 1182.0400 ;
        RECT 2033.3400 1176.1200 2036.3400 1176.6000 ;
        RECT 2045.1000 1159.8000 2046.7000 1160.2800 ;
        RECT 2045.1000 1165.2400 2046.7000 1165.7200 ;
        RECT 2033.3400 1165.2400 2036.3400 1165.7200 ;
        RECT 2033.3400 1159.8000 2036.3400 1160.2800 ;
        RECT 2033.3400 1170.6800 2036.3400 1171.1600 ;
        RECT 2045.1000 1170.6800 2046.7000 1171.1600 ;
        RECT 2135.1000 1143.4800 2136.7000 1143.9600 ;
        RECT 2135.1000 1148.9200 2136.7000 1149.4000 ;
        RECT 2135.1000 1154.3600 2136.7000 1154.8400 ;
        RECT 2135.1000 1132.6000 2136.7000 1133.0800 ;
        RECT 2135.1000 1138.0400 2136.7000 1138.5200 ;
        RECT 2090.1000 1143.4800 2091.7000 1143.9600 ;
        RECT 2090.1000 1148.9200 2091.7000 1149.4000 ;
        RECT 2090.1000 1154.3600 2091.7000 1154.8400 ;
        RECT 2090.1000 1132.6000 2091.7000 1133.0800 ;
        RECT 2090.1000 1138.0400 2091.7000 1138.5200 ;
        RECT 2135.1000 1116.2800 2136.7000 1116.7600 ;
        RECT 2135.1000 1121.7200 2136.7000 1122.2000 ;
        RECT 2135.1000 1127.1600 2136.7000 1127.6400 ;
        RECT 2135.1000 1105.4000 2136.7000 1105.8800 ;
        RECT 2135.1000 1110.8400 2136.7000 1111.3200 ;
        RECT 2090.1000 1116.2800 2091.7000 1116.7600 ;
        RECT 2090.1000 1121.7200 2091.7000 1122.2000 ;
        RECT 2090.1000 1127.1600 2091.7000 1127.6400 ;
        RECT 2090.1000 1105.4000 2091.7000 1105.8800 ;
        RECT 2090.1000 1110.8400 2091.7000 1111.3200 ;
        RECT 2045.1000 1143.4800 2046.7000 1143.9600 ;
        RECT 2045.1000 1148.9200 2046.7000 1149.4000 ;
        RECT 2045.1000 1154.3600 2046.7000 1154.8400 ;
        RECT 2033.3400 1143.4800 2036.3400 1143.9600 ;
        RECT 2033.3400 1148.9200 2036.3400 1149.4000 ;
        RECT 2033.3400 1154.3600 2036.3400 1154.8400 ;
        RECT 2045.1000 1132.6000 2046.7000 1133.0800 ;
        RECT 2045.1000 1138.0400 2046.7000 1138.5200 ;
        RECT 2033.3400 1132.6000 2036.3400 1133.0800 ;
        RECT 2033.3400 1138.0400 2036.3400 1138.5200 ;
        RECT 2045.1000 1116.2800 2046.7000 1116.7600 ;
        RECT 2045.1000 1121.7200 2046.7000 1122.2000 ;
        RECT 2045.1000 1127.1600 2046.7000 1127.6400 ;
        RECT 2033.3400 1116.2800 2036.3400 1116.7600 ;
        RECT 2033.3400 1121.7200 2036.3400 1122.2000 ;
        RECT 2033.3400 1127.1600 2036.3400 1127.6400 ;
        RECT 2045.1000 1105.4000 2046.7000 1105.8800 ;
        RECT 2045.1000 1110.8400 2046.7000 1111.3200 ;
        RECT 2033.3400 1105.4000 2036.3400 1105.8800 ;
        RECT 2033.3400 1110.8400 2036.3400 1111.3200 ;
        RECT 2237.4400 1089.0800 2240.4400 1089.5600 ;
        RECT 2237.4400 1094.5200 2240.4400 1095.0000 ;
        RECT 2237.4400 1099.9600 2240.4400 1100.4400 ;
        RECT 2225.1000 1089.0800 2226.7000 1089.5600 ;
        RECT 2225.1000 1094.5200 2226.7000 1095.0000 ;
        RECT 2225.1000 1099.9600 2226.7000 1100.4400 ;
        RECT 2237.4400 1078.2000 2240.4400 1078.6800 ;
        RECT 2237.4400 1083.6400 2240.4400 1084.1200 ;
        RECT 2225.1000 1078.2000 2226.7000 1078.6800 ;
        RECT 2225.1000 1083.6400 2226.7000 1084.1200 ;
        RECT 2237.4400 1061.8800 2240.4400 1062.3600 ;
        RECT 2237.4400 1067.3200 2240.4400 1067.8000 ;
        RECT 2237.4400 1072.7600 2240.4400 1073.2400 ;
        RECT 2225.1000 1061.8800 2226.7000 1062.3600 ;
        RECT 2225.1000 1067.3200 2226.7000 1067.8000 ;
        RECT 2225.1000 1072.7600 2226.7000 1073.2400 ;
        RECT 2237.4400 1051.0000 2240.4400 1051.4800 ;
        RECT 2237.4400 1056.4400 2240.4400 1056.9200 ;
        RECT 2225.1000 1051.0000 2226.7000 1051.4800 ;
        RECT 2225.1000 1056.4400 2226.7000 1056.9200 ;
        RECT 2180.1000 1089.0800 2181.7000 1089.5600 ;
        RECT 2180.1000 1094.5200 2181.7000 1095.0000 ;
        RECT 2180.1000 1099.9600 2181.7000 1100.4400 ;
        RECT 2180.1000 1078.2000 2181.7000 1078.6800 ;
        RECT 2180.1000 1083.6400 2181.7000 1084.1200 ;
        RECT 2180.1000 1061.8800 2181.7000 1062.3600 ;
        RECT 2180.1000 1067.3200 2181.7000 1067.8000 ;
        RECT 2180.1000 1072.7600 2181.7000 1073.2400 ;
        RECT 2180.1000 1051.0000 2181.7000 1051.4800 ;
        RECT 2180.1000 1056.4400 2181.7000 1056.9200 ;
        RECT 2237.4400 1034.6800 2240.4400 1035.1600 ;
        RECT 2237.4400 1040.1200 2240.4400 1040.6000 ;
        RECT 2237.4400 1045.5600 2240.4400 1046.0400 ;
        RECT 2225.1000 1034.6800 2226.7000 1035.1600 ;
        RECT 2225.1000 1040.1200 2226.7000 1040.6000 ;
        RECT 2225.1000 1045.5600 2226.7000 1046.0400 ;
        RECT 2237.4400 1023.8000 2240.4400 1024.2800 ;
        RECT 2237.4400 1029.2400 2240.4400 1029.7200 ;
        RECT 2225.1000 1023.8000 2226.7000 1024.2800 ;
        RECT 2225.1000 1029.2400 2226.7000 1029.7200 ;
        RECT 2237.4400 1007.4800 2240.4400 1007.9600 ;
        RECT 2237.4400 1012.9200 2240.4400 1013.4000 ;
        RECT 2237.4400 1018.3600 2240.4400 1018.8400 ;
        RECT 2225.1000 1007.4800 2226.7000 1007.9600 ;
        RECT 2225.1000 1012.9200 2226.7000 1013.4000 ;
        RECT 2225.1000 1018.3600 2226.7000 1018.8400 ;
        RECT 2237.4400 1002.0400 2240.4400 1002.5200 ;
        RECT 2225.1000 1002.0400 2226.7000 1002.5200 ;
        RECT 2180.1000 1034.6800 2181.7000 1035.1600 ;
        RECT 2180.1000 1040.1200 2181.7000 1040.6000 ;
        RECT 2180.1000 1045.5600 2181.7000 1046.0400 ;
        RECT 2180.1000 1023.8000 2181.7000 1024.2800 ;
        RECT 2180.1000 1029.2400 2181.7000 1029.7200 ;
        RECT 2180.1000 1007.4800 2181.7000 1007.9600 ;
        RECT 2180.1000 1012.9200 2181.7000 1013.4000 ;
        RECT 2180.1000 1018.3600 2181.7000 1018.8400 ;
        RECT 2180.1000 1002.0400 2181.7000 1002.5200 ;
        RECT 2135.1000 1089.0800 2136.7000 1089.5600 ;
        RECT 2135.1000 1094.5200 2136.7000 1095.0000 ;
        RECT 2135.1000 1099.9600 2136.7000 1100.4400 ;
        RECT 2135.1000 1078.2000 2136.7000 1078.6800 ;
        RECT 2135.1000 1083.6400 2136.7000 1084.1200 ;
        RECT 2090.1000 1089.0800 2091.7000 1089.5600 ;
        RECT 2090.1000 1094.5200 2091.7000 1095.0000 ;
        RECT 2090.1000 1099.9600 2091.7000 1100.4400 ;
        RECT 2090.1000 1078.2000 2091.7000 1078.6800 ;
        RECT 2090.1000 1083.6400 2091.7000 1084.1200 ;
        RECT 2135.1000 1061.8800 2136.7000 1062.3600 ;
        RECT 2135.1000 1067.3200 2136.7000 1067.8000 ;
        RECT 2135.1000 1072.7600 2136.7000 1073.2400 ;
        RECT 2135.1000 1051.0000 2136.7000 1051.4800 ;
        RECT 2135.1000 1056.4400 2136.7000 1056.9200 ;
        RECT 2090.1000 1061.8800 2091.7000 1062.3600 ;
        RECT 2090.1000 1067.3200 2091.7000 1067.8000 ;
        RECT 2090.1000 1072.7600 2091.7000 1073.2400 ;
        RECT 2090.1000 1051.0000 2091.7000 1051.4800 ;
        RECT 2090.1000 1056.4400 2091.7000 1056.9200 ;
        RECT 2045.1000 1089.0800 2046.7000 1089.5600 ;
        RECT 2045.1000 1094.5200 2046.7000 1095.0000 ;
        RECT 2045.1000 1099.9600 2046.7000 1100.4400 ;
        RECT 2033.3400 1089.0800 2036.3400 1089.5600 ;
        RECT 2033.3400 1094.5200 2036.3400 1095.0000 ;
        RECT 2033.3400 1099.9600 2036.3400 1100.4400 ;
        RECT 2045.1000 1078.2000 2046.7000 1078.6800 ;
        RECT 2045.1000 1083.6400 2046.7000 1084.1200 ;
        RECT 2033.3400 1078.2000 2036.3400 1078.6800 ;
        RECT 2033.3400 1083.6400 2036.3400 1084.1200 ;
        RECT 2045.1000 1061.8800 2046.7000 1062.3600 ;
        RECT 2045.1000 1067.3200 2046.7000 1067.8000 ;
        RECT 2045.1000 1072.7600 2046.7000 1073.2400 ;
        RECT 2033.3400 1061.8800 2036.3400 1062.3600 ;
        RECT 2033.3400 1067.3200 2036.3400 1067.8000 ;
        RECT 2033.3400 1072.7600 2036.3400 1073.2400 ;
        RECT 2045.1000 1051.0000 2046.7000 1051.4800 ;
        RECT 2045.1000 1056.4400 2046.7000 1056.9200 ;
        RECT 2033.3400 1051.0000 2036.3400 1051.4800 ;
        RECT 2033.3400 1056.4400 2036.3400 1056.9200 ;
        RECT 2135.1000 1034.6800 2136.7000 1035.1600 ;
        RECT 2135.1000 1040.1200 2136.7000 1040.6000 ;
        RECT 2135.1000 1045.5600 2136.7000 1046.0400 ;
        RECT 2135.1000 1023.8000 2136.7000 1024.2800 ;
        RECT 2135.1000 1029.2400 2136.7000 1029.7200 ;
        RECT 2090.1000 1034.6800 2091.7000 1035.1600 ;
        RECT 2090.1000 1040.1200 2091.7000 1040.6000 ;
        RECT 2090.1000 1045.5600 2091.7000 1046.0400 ;
        RECT 2090.1000 1023.8000 2091.7000 1024.2800 ;
        RECT 2090.1000 1029.2400 2091.7000 1029.7200 ;
        RECT 2135.1000 1007.4800 2136.7000 1007.9600 ;
        RECT 2135.1000 1012.9200 2136.7000 1013.4000 ;
        RECT 2135.1000 1018.3600 2136.7000 1018.8400 ;
        RECT 2135.1000 1002.0400 2136.7000 1002.5200 ;
        RECT 2090.1000 1007.4800 2091.7000 1007.9600 ;
        RECT 2090.1000 1012.9200 2091.7000 1013.4000 ;
        RECT 2090.1000 1018.3600 2091.7000 1018.8400 ;
        RECT 2090.1000 1002.0400 2091.7000 1002.5200 ;
        RECT 2045.1000 1034.6800 2046.7000 1035.1600 ;
        RECT 2045.1000 1040.1200 2046.7000 1040.6000 ;
        RECT 2045.1000 1045.5600 2046.7000 1046.0400 ;
        RECT 2033.3400 1034.6800 2036.3400 1035.1600 ;
        RECT 2033.3400 1040.1200 2036.3400 1040.6000 ;
        RECT 2033.3400 1045.5600 2036.3400 1046.0400 ;
        RECT 2045.1000 1023.8000 2046.7000 1024.2800 ;
        RECT 2045.1000 1029.2400 2046.7000 1029.7200 ;
        RECT 2033.3400 1023.8000 2036.3400 1024.2800 ;
        RECT 2033.3400 1029.2400 2036.3400 1029.7200 ;
        RECT 2045.1000 1007.4800 2046.7000 1007.9600 ;
        RECT 2045.1000 1012.9200 2046.7000 1013.4000 ;
        RECT 2045.1000 1018.3600 2046.7000 1018.8400 ;
        RECT 2033.3400 1007.4800 2036.3400 1007.9600 ;
        RECT 2033.3400 1012.9200 2036.3400 1013.4000 ;
        RECT 2033.3400 1018.3600 2036.3400 1018.8400 ;
        RECT 2033.3400 1002.0400 2036.3400 1002.5200 ;
        RECT 2045.1000 1002.0400 2046.7000 1002.5200 ;
        RECT 2033.3400 1206.9500 2240.4400 1209.9500 ;
        RECT 2033.3400 993.8500 2240.4400 996.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2225.1000 764.2100 2226.7000 980.3100 ;
        RECT 2180.1000 764.2100 2181.7000 980.3100 ;
        RECT 2135.1000 764.2100 2136.7000 980.3100 ;
        RECT 2090.1000 764.2100 2091.7000 980.3100 ;
        RECT 2045.1000 764.2100 2046.7000 980.3100 ;
        RECT 2237.4400 764.2100 2240.4400 980.3100 ;
        RECT 2033.3400 764.2100 2036.3400 980.3100 ;
      LAYER met3 ;
        RECT 2237.4400 957.3600 2240.4400 957.8400 ;
        RECT 2237.4400 962.8000 2240.4400 963.2800 ;
        RECT 2225.1000 957.3600 2226.7000 957.8400 ;
        RECT 2225.1000 962.8000 2226.7000 963.2800 ;
        RECT 2237.4400 968.2400 2240.4400 968.7200 ;
        RECT 2225.1000 968.2400 2226.7000 968.7200 ;
        RECT 2237.4400 946.4800 2240.4400 946.9600 ;
        RECT 2237.4400 951.9200 2240.4400 952.4000 ;
        RECT 2225.1000 946.4800 2226.7000 946.9600 ;
        RECT 2225.1000 951.9200 2226.7000 952.4000 ;
        RECT 2237.4400 930.1600 2240.4400 930.6400 ;
        RECT 2237.4400 935.6000 2240.4400 936.0800 ;
        RECT 2225.1000 930.1600 2226.7000 930.6400 ;
        RECT 2225.1000 935.6000 2226.7000 936.0800 ;
        RECT 2237.4400 941.0400 2240.4400 941.5200 ;
        RECT 2225.1000 941.0400 2226.7000 941.5200 ;
        RECT 2180.1000 957.3600 2181.7000 957.8400 ;
        RECT 2180.1000 962.8000 2181.7000 963.2800 ;
        RECT 2180.1000 968.2400 2181.7000 968.7200 ;
        RECT 2180.1000 946.4800 2181.7000 946.9600 ;
        RECT 2180.1000 951.9200 2181.7000 952.4000 ;
        RECT 2180.1000 930.1600 2181.7000 930.6400 ;
        RECT 2180.1000 935.6000 2181.7000 936.0800 ;
        RECT 2180.1000 941.0400 2181.7000 941.5200 ;
        RECT 2237.4400 913.8400 2240.4400 914.3200 ;
        RECT 2237.4400 919.2800 2240.4400 919.7600 ;
        RECT 2237.4400 924.7200 2240.4400 925.2000 ;
        RECT 2225.1000 913.8400 2226.7000 914.3200 ;
        RECT 2225.1000 919.2800 2226.7000 919.7600 ;
        RECT 2225.1000 924.7200 2226.7000 925.2000 ;
        RECT 2237.4400 902.9600 2240.4400 903.4400 ;
        RECT 2237.4400 908.4000 2240.4400 908.8800 ;
        RECT 2225.1000 902.9600 2226.7000 903.4400 ;
        RECT 2225.1000 908.4000 2226.7000 908.8800 ;
        RECT 2237.4400 886.6400 2240.4400 887.1200 ;
        RECT 2237.4400 892.0800 2240.4400 892.5600 ;
        RECT 2237.4400 897.5200 2240.4400 898.0000 ;
        RECT 2225.1000 886.6400 2226.7000 887.1200 ;
        RECT 2225.1000 892.0800 2226.7000 892.5600 ;
        RECT 2225.1000 897.5200 2226.7000 898.0000 ;
        RECT 2237.4400 875.7600 2240.4400 876.2400 ;
        RECT 2237.4400 881.2000 2240.4400 881.6800 ;
        RECT 2225.1000 875.7600 2226.7000 876.2400 ;
        RECT 2225.1000 881.2000 2226.7000 881.6800 ;
        RECT 2180.1000 913.8400 2181.7000 914.3200 ;
        RECT 2180.1000 919.2800 2181.7000 919.7600 ;
        RECT 2180.1000 924.7200 2181.7000 925.2000 ;
        RECT 2180.1000 902.9600 2181.7000 903.4400 ;
        RECT 2180.1000 908.4000 2181.7000 908.8800 ;
        RECT 2180.1000 886.6400 2181.7000 887.1200 ;
        RECT 2180.1000 892.0800 2181.7000 892.5600 ;
        RECT 2180.1000 897.5200 2181.7000 898.0000 ;
        RECT 2180.1000 875.7600 2181.7000 876.2400 ;
        RECT 2180.1000 881.2000 2181.7000 881.6800 ;
        RECT 2135.1000 957.3600 2136.7000 957.8400 ;
        RECT 2135.1000 962.8000 2136.7000 963.2800 ;
        RECT 2135.1000 968.2400 2136.7000 968.7200 ;
        RECT 2090.1000 957.3600 2091.7000 957.8400 ;
        RECT 2090.1000 962.8000 2091.7000 963.2800 ;
        RECT 2090.1000 968.2400 2091.7000 968.7200 ;
        RECT 2135.1000 946.4800 2136.7000 946.9600 ;
        RECT 2135.1000 951.9200 2136.7000 952.4000 ;
        RECT 2135.1000 930.1600 2136.7000 930.6400 ;
        RECT 2135.1000 935.6000 2136.7000 936.0800 ;
        RECT 2135.1000 941.0400 2136.7000 941.5200 ;
        RECT 2090.1000 946.4800 2091.7000 946.9600 ;
        RECT 2090.1000 951.9200 2091.7000 952.4000 ;
        RECT 2090.1000 930.1600 2091.7000 930.6400 ;
        RECT 2090.1000 935.6000 2091.7000 936.0800 ;
        RECT 2090.1000 941.0400 2091.7000 941.5200 ;
        RECT 2045.1000 957.3600 2046.7000 957.8400 ;
        RECT 2045.1000 962.8000 2046.7000 963.2800 ;
        RECT 2033.3400 962.8000 2036.3400 963.2800 ;
        RECT 2033.3400 957.3600 2036.3400 957.8400 ;
        RECT 2033.3400 968.2400 2036.3400 968.7200 ;
        RECT 2045.1000 968.2400 2046.7000 968.7200 ;
        RECT 2045.1000 946.4800 2046.7000 946.9600 ;
        RECT 2045.1000 951.9200 2046.7000 952.4000 ;
        RECT 2033.3400 951.9200 2036.3400 952.4000 ;
        RECT 2033.3400 946.4800 2036.3400 946.9600 ;
        RECT 2045.1000 930.1600 2046.7000 930.6400 ;
        RECT 2045.1000 935.6000 2046.7000 936.0800 ;
        RECT 2033.3400 935.6000 2036.3400 936.0800 ;
        RECT 2033.3400 930.1600 2036.3400 930.6400 ;
        RECT 2033.3400 941.0400 2036.3400 941.5200 ;
        RECT 2045.1000 941.0400 2046.7000 941.5200 ;
        RECT 2135.1000 913.8400 2136.7000 914.3200 ;
        RECT 2135.1000 919.2800 2136.7000 919.7600 ;
        RECT 2135.1000 924.7200 2136.7000 925.2000 ;
        RECT 2135.1000 902.9600 2136.7000 903.4400 ;
        RECT 2135.1000 908.4000 2136.7000 908.8800 ;
        RECT 2090.1000 913.8400 2091.7000 914.3200 ;
        RECT 2090.1000 919.2800 2091.7000 919.7600 ;
        RECT 2090.1000 924.7200 2091.7000 925.2000 ;
        RECT 2090.1000 902.9600 2091.7000 903.4400 ;
        RECT 2090.1000 908.4000 2091.7000 908.8800 ;
        RECT 2135.1000 886.6400 2136.7000 887.1200 ;
        RECT 2135.1000 892.0800 2136.7000 892.5600 ;
        RECT 2135.1000 897.5200 2136.7000 898.0000 ;
        RECT 2135.1000 875.7600 2136.7000 876.2400 ;
        RECT 2135.1000 881.2000 2136.7000 881.6800 ;
        RECT 2090.1000 886.6400 2091.7000 887.1200 ;
        RECT 2090.1000 892.0800 2091.7000 892.5600 ;
        RECT 2090.1000 897.5200 2091.7000 898.0000 ;
        RECT 2090.1000 875.7600 2091.7000 876.2400 ;
        RECT 2090.1000 881.2000 2091.7000 881.6800 ;
        RECT 2045.1000 913.8400 2046.7000 914.3200 ;
        RECT 2045.1000 919.2800 2046.7000 919.7600 ;
        RECT 2045.1000 924.7200 2046.7000 925.2000 ;
        RECT 2033.3400 913.8400 2036.3400 914.3200 ;
        RECT 2033.3400 919.2800 2036.3400 919.7600 ;
        RECT 2033.3400 924.7200 2036.3400 925.2000 ;
        RECT 2045.1000 902.9600 2046.7000 903.4400 ;
        RECT 2045.1000 908.4000 2046.7000 908.8800 ;
        RECT 2033.3400 902.9600 2036.3400 903.4400 ;
        RECT 2033.3400 908.4000 2036.3400 908.8800 ;
        RECT 2045.1000 886.6400 2046.7000 887.1200 ;
        RECT 2045.1000 892.0800 2046.7000 892.5600 ;
        RECT 2045.1000 897.5200 2046.7000 898.0000 ;
        RECT 2033.3400 886.6400 2036.3400 887.1200 ;
        RECT 2033.3400 892.0800 2036.3400 892.5600 ;
        RECT 2033.3400 897.5200 2036.3400 898.0000 ;
        RECT 2045.1000 875.7600 2046.7000 876.2400 ;
        RECT 2045.1000 881.2000 2046.7000 881.6800 ;
        RECT 2033.3400 875.7600 2036.3400 876.2400 ;
        RECT 2033.3400 881.2000 2036.3400 881.6800 ;
        RECT 2237.4400 859.4400 2240.4400 859.9200 ;
        RECT 2237.4400 864.8800 2240.4400 865.3600 ;
        RECT 2237.4400 870.3200 2240.4400 870.8000 ;
        RECT 2225.1000 859.4400 2226.7000 859.9200 ;
        RECT 2225.1000 864.8800 2226.7000 865.3600 ;
        RECT 2225.1000 870.3200 2226.7000 870.8000 ;
        RECT 2237.4400 848.5600 2240.4400 849.0400 ;
        RECT 2237.4400 854.0000 2240.4400 854.4800 ;
        RECT 2225.1000 848.5600 2226.7000 849.0400 ;
        RECT 2225.1000 854.0000 2226.7000 854.4800 ;
        RECT 2237.4400 832.2400 2240.4400 832.7200 ;
        RECT 2237.4400 837.6800 2240.4400 838.1600 ;
        RECT 2237.4400 843.1200 2240.4400 843.6000 ;
        RECT 2225.1000 832.2400 2226.7000 832.7200 ;
        RECT 2225.1000 837.6800 2226.7000 838.1600 ;
        RECT 2225.1000 843.1200 2226.7000 843.6000 ;
        RECT 2237.4400 821.3600 2240.4400 821.8400 ;
        RECT 2237.4400 826.8000 2240.4400 827.2800 ;
        RECT 2225.1000 821.3600 2226.7000 821.8400 ;
        RECT 2225.1000 826.8000 2226.7000 827.2800 ;
        RECT 2180.1000 859.4400 2181.7000 859.9200 ;
        RECT 2180.1000 864.8800 2181.7000 865.3600 ;
        RECT 2180.1000 870.3200 2181.7000 870.8000 ;
        RECT 2180.1000 848.5600 2181.7000 849.0400 ;
        RECT 2180.1000 854.0000 2181.7000 854.4800 ;
        RECT 2180.1000 832.2400 2181.7000 832.7200 ;
        RECT 2180.1000 837.6800 2181.7000 838.1600 ;
        RECT 2180.1000 843.1200 2181.7000 843.6000 ;
        RECT 2180.1000 821.3600 2181.7000 821.8400 ;
        RECT 2180.1000 826.8000 2181.7000 827.2800 ;
        RECT 2237.4400 805.0400 2240.4400 805.5200 ;
        RECT 2237.4400 810.4800 2240.4400 810.9600 ;
        RECT 2237.4400 815.9200 2240.4400 816.4000 ;
        RECT 2225.1000 805.0400 2226.7000 805.5200 ;
        RECT 2225.1000 810.4800 2226.7000 810.9600 ;
        RECT 2225.1000 815.9200 2226.7000 816.4000 ;
        RECT 2237.4400 794.1600 2240.4400 794.6400 ;
        RECT 2237.4400 799.6000 2240.4400 800.0800 ;
        RECT 2225.1000 794.1600 2226.7000 794.6400 ;
        RECT 2225.1000 799.6000 2226.7000 800.0800 ;
        RECT 2237.4400 777.8400 2240.4400 778.3200 ;
        RECT 2237.4400 783.2800 2240.4400 783.7600 ;
        RECT 2237.4400 788.7200 2240.4400 789.2000 ;
        RECT 2225.1000 777.8400 2226.7000 778.3200 ;
        RECT 2225.1000 783.2800 2226.7000 783.7600 ;
        RECT 2225.1000 788.7200 2226.7000 789.2000 ;
        RECT 2237.4400 772.4000 2240.4400 772.8800 ;
        RECT 2225.1000 772.4000 2226.7000 772.8800 ;
        RECT 2180.1000 805.0400 2181.7000 805.5200 ;
        RECT 2180.1000 810.4800 2181.7000 810.9600 ;
        RECT 2180.1000 815.9200 2181.7000 816.4000 ;
        RECT 2180.1000 794.1600 2181.7000 794.6400 ;
        RECT 2180.1000 799.6000 2181.7000 800.0800 ;
        RECT 2180.1000 777.8400 2181.7000 778.3200 ;
        RECT 2180.1000 783.2800 2181.7000 783.7600 ;
        RECT 2180.1000 788.7200 2181.7000 789.2000 ;
        RECT 2180.1000 772.4000 2181.7000 772.8800 ;
        RECT 2135.1000 859.4400 2136.7000 859.9200 ;
        RECT 2135.1000 864.8800 2136.7000 865.3600 ;
        RECT 2135.1000 870.3200 2136.7000 870.8000 ;
        RECT 2135.1000 848.5600 2136.7000 849.0400 ;
        RECT 2135.1000 854.0000 2136.7000 854.4800 ;
        RECT 2090.1000 859.4400 2091.7000 859.9200 ;
        RECT 2090.1000 864.8800 2091.7000 865.3600 ;
        RECT 2090.1000 870.3200 2091.7000 870.8000 ;
        RECT 2090.1000 848.5600 2091.7000 849.0400 ;
        RECT 2090.1000 854.0000 2091.7000 854.4800 ;
        RECT 2135.1000 832.2400 2136.7000 832.7200 ;
        RECT 2135.1000 837.6800 2136.7000 838.1600 ;
        RECT 2135.1000 843.1200 2136.7000 843.6000 ;
        RECT 2135.1000 821.3600 2136.7000 821.8400 ;
        RECT 2135.1000 826.8000 2136.7000 827.2800 ;
        RECT 2090.1000 832.2400 2091.7000 832.7200 ;
        RECT 2090.1000 837.6800 2091.7000 838.1600 ;
        RECT 2090.1000 843.1200 2091.7000 843.6000 ;
        RECT 2090.1000 821.3600 2091.7000 821.8400 ;
        RECT 2090.1000 826.8000 2091.7000 827.2800 ;
        RECT 2045.1000 859.4400 2046.7000 859.9200 ;
        RECT 2045.1000 864.8800 2046.7000 865.3600 ;
        RECT 2045.1000 870.3200 2046.7000 870.8000 ;
        RECT 2033.3400 859.4400 2036.3400 859.9200 ;
        RECT 2033.3400 864.8800 2036.3400 865.3600 ;
        RECT 2033.3400 870.3200 2036.3400 870.8000 ;
        RECT 2045.1000 848.5600 2046.7000 849.0400 ;
        RECT 2045.1000 854.0000 2046.7000 854.4800 ;
        RECT 2033.3400 848.5600 2036.3400 849.0400 ;
        RECT 2033.3400 854.0000 2036.3400 854.4800 ;
        RECT 2045.1000 832.2400 2046.7000 832.7200 ;
        RECT 2045.1000 837.6800 2046.7000 838.1600 ;
        RECT 2045.1000 843.1200 2046.7000 843.6000 ;
        RECT 2033.3400 832.2400 2036.3400 832.7200 ;
        RECT 2033.3400 837.6800 2036.3400 838.1600 ;
        RECT 2033.3400 843.1200 2036.3400 843.6000 ;
        RECT 2045.1000 821.3600 2046.7000 821.8400 ;
        RECT 2045.1000 826.8000 2046.7000 827.2800 ;
        RECT 2033.3400 821.3600 2036.3400 821.8400 ;
        RECT 2033.3400 826.8000 2036.3400 827.2800 ;
        RECT 2135.1000 805.0400 2136.7000 805.5200 ;
        RECT 2135.1000 810.4800 2136.7000 810.9600 ;
        RECT 2135.1000 815.9200 2136.7000 816.4000 ;
        RECT 2135.1000 794.1600 2136.7000 794.6400 ;
        RECT 2135.1000 799.6000 2136.7000 800.0800 ;
        RECT 2090.1000 805.0400 2091.7000 805.5200 ;
        RECT 2090.1000 810.4800 2091.7000 810.9600 ;
        RECT 2090.1000 815.9200 2091.7000 816.4000 ;
        RECT 2090.1000 794.1600 2091.7000 794.6400 ;
        RECT 2090.1000 799.6000 2091.7000 800.0800 ;
        RECT 2135.1000 777.8400 2136.7000 778.3200 ;
        RECT 2135.1000 783.2800 2136.7000 783.7600 ;
        RECT 2135.1000 788.7200 2136.7000 789.2000 ;
        RECT 2135.1000 772.4000 2136.7000 772.8800 ;
        RECT 2090.1000 777.8400 2091.7000 778.3200 ;
        RECT 2090.1000 783.2800 2091.7000 783.7600 ;
        RECT 2090.1000 788.7200 2091.7000 789.2000 ;
        RECT 2090.1000 772.4000 2091.7000 772.8800 ;
        RECT 2045.1000 805.0400 2046.7000 805.5200 ;
        RECT 2045.1000 810.4800 2046.7000 810.9600 ;
        RECT 2045.1000 815.9200 2046.7000 816.4000 ;
        RECT 2033.3400 805.0400 2036.3400 805.5200 ;
        RECT 2033.3400 810.4800 2036.3400 810.9600 ;
        RECT 2033.3400 815.9200 2036.3400 816.4000 ;
        RECT 2045.1000 794.1600 2046.7000 794.6400 ;
        RECT 2045.1000 799.6000 2046.7000 800.0800 ;
        RECT 2033.3400 794.1600 2036.3400 794.6400 ;
        RECT 2033.3400 799.6000 2036.3400 800.0800 ;
        RECT 2045.1000 777.8400 2046.7000 778.3200 ;
        RECT 2045.1000 783.2800 2046.7000 783.7600 ;
        RECT 2045.1000 788.7200 2046.7000 789.2000 ;
        RECT 2033.3400 777.8400 2036.3400 778.3200 ;
        RECT 2033.3400 783.2800 2036.3400 783.7600 ;
        RECT 2033.3400 788.7200 2036.3400 789.2000 ;
        RECT 2033.3400 772.4000 2036.3400 772.8800 ;
        RECT 2045.1000 772.4000 2046.7000 772.8800 ;
        RECT 2033.3400 977.3100 2240.4400 980.3100 ;
        RECT 2033.3400 764.2100 2240.4400 767.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 3390.2000 2889.6600 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 3390.2000 2889.6600 ;
    LAYER met2 ;
      RECT 3300.0200 2889.0350 3390.2000 2889.6600 ;
      RECT 3140.4000 2889.0350 3299.6000 2889.6600 ;
      RECT 2980.3200 2889.0350 3139.9800 2889.6600 ;
      RECT 2820.2400 2889.0350 2979.9000 2889.6600 ;
      RECT 2660.1600 2889.0350 2819.8200 2889.6600 ;
      RECT 2500.0800 2889.0350 2659.7400 2889.6600 ;
      RECT 2340.4600 2889.0350 2499.6600 2889.6600 ;
      RECT 2180.3800 2889.0350 2340.0400 2889.6600 ;
      RECT 2020.3000 2889.0350 2179.9600 2889.6600 ;
      RECT 1860.2200 2889.0350 2019.8800 2889.6600 ;
      RECT 1700.1400 2889.0350 1859.8000 2889.6600 ;
      RECT 1540.5200 2889.0350 1699.7200 2889.6600 ;
      RECT 1380.4400 2889.0350 1540.1000 2889.6600 ;
      RECT 1220.3600 2889.0350 1380.0200 2889.6600 ;
      RECT 1060.2800 2889.0350 1219.9400 2889.6600 ;
      RECT 900.2000 2889.0350 1059.8600 2889.6600 ;
      RECT 740.5800 2889.0350 899.7800 2889.6600 ;
      RECT 580.5000 2889.0350 740.1600 2889.6600 ;
      RECT 420.4200 2889.0350 580.0800 2889.6600 ;
      RECT 260.3400 2889.0350 420.0000 2889.6600 ;
      RECT 100.2600 2889.0350 259.9200 2889.6600 ;
      RECT 0.0000 2889.0350 99.8400 2889.6600 ;
      RECT 0.0000 0.6250 3390.2000 2889.0350 ;
      RECT 3300.0200 0.0000 3390.2000 0.6250 ;
      RECT 3227.3400 0.0000 3299.6000 0.6250 ;
      RECT 3154.6600 0.0000 3226.9200 0.6250 ;
      RECT 3081.9800 0.0000 3154.2400 0.6250 ;
      RECT 3009.3000 0.0000 3081.5600 0.6250 ;
      RECT 2936.6200 0.0000 3008.8800 0.6250 ;
      RECT 2863.9400 0.0000 2936.2000 0.6250 ;
      RECT 2791.2600 0.0000 2863.5200 0.6250 ;
      RECT 2718.5800 0.0000 2790.8400 0.6250 ;
      RECT 2645.9000 0.0000 2718.1600 0.6250 ;
      RECT 2573.2200 0.0000 2645.4800 0.6250 ;
      RECT 2500.5400 0.0000 2572.8000 0.6250 ;
      RECT 2427.4000 0.0000 2500.1200 0.6250 ;
      RECT 2354.7200 0.0000 2426.9800 0.6250 ;
      RECT 2282.0400 0.0000 2354.3000 0.6250 ;
      RECT 2209.3600 0.0000 2281.6200 0.6250 ;
      RECT 2136.6800 0.0000 2208.9400 0.6250 ;
      RECT 2064.0000 0.0000 2136.2600 0.6250 ;
      RECT 1991.3200 0.0000 2063.5800 0.6250 ;
      RECT 1918.6400 0.0000 1990.9000 0.6250 ;
      RECT 1845.9600 0.0000 1918.2200 0.6250 ;
      RECT 1773.2800 0.0000 1845.5400 0.6250 ;
      RECT 1700.6000 0.0000 1772.8600 0.6250 ;
      RECT 1627.4600 0.0000 1700.1800 0.6250 ;
      RECT 1554.7800 0.0000 1627.0400 0.6250 ;
      RECT 1482.1000 0.0000 1554.3600 0.6250 ;
      RECT 1409.4200 0.0000 1481.6800 0.6250 ;
      RECT 1336.7400 0.0000 1409.0000 0.6250 ;
      RECT 1264.0600 0.0000 1336.3200 0.6250 ;
      RECT 1191.3800 0.0000 1263.6400 0.6250 ;
      RECT 1118.7000 0.0000 1190.9600 0.6250 ;
      RECT 1046.0200 0.0000 1118.2800 0.6250 ;
      RECT 973.3400 0.0000 1045.6000 0.6250 ;
      RECT 900.6600 0.0000 972.9200 0.6250 ;
      RECT 827.5200 0.0000 900.2400 0.6250 ;
      RECT 754.8400 0.0000 827.1000 0.6250 ;
      RECT 682.1600 0.0000 754.4200 0.6250 ;
      RECT 609.4800 0.0000 681.7400 0.6250 ;
      RECT 536.8000 0.0000 609.0600 0.6250 ;
      RECT 464.1200 0.0000 536.3800 0.6250 ;
      RECT 391.4400 0.0000 463.7000 0.6250 ;
      RECT 318.7600 0.0000 391.0200 0.6250 ;
      RECT 246.0800 0.0000 318.3400 0.6250 ;
      RECT 173.4000 0.0000 245.6600 0.6250 ;
      RECT 100.7200 0.0000 172.9800 0.6250 ;
      RECT 0.0000 0.0000 100.3000 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 2887.9600 3390.2000 2889.6600 ;
      RECT 3388.5000 2884.3600 3390.2000 2887.9600 ;
      RECT 0.0000 2884.3600 1.7000 2887.9600 ;
      RECT 0.0000 2883.9600 3390.2000 2884.3600 ;
      RECT 3384.5000 2880.3600 3390.2000 2883.9600 ;
      RECT 0.0000 2880.3600 5.7000 2883.9600 ;
      RECT 0.0000 2880.0000 3390.2000 2880.3600 ;
      RECT 3388.5000 2878.9200 3390.2000 2880.0000 ;
      RECT 5.3000 2878.9200 3384.9000 2880.0000 ;
      RECT 0.0000 2878.9200 1.7000 2880.0000 ;
      RECT 0.0000 2877.2800 3390.2000 2878.9200 ;
      RECT 3384.5000 2876.2000 3390.2000 2877.2800 ;
      RECT 9.3000 2876.2000 3380.9000 2877.2800 ;
      RECT 0.0000 2876.2000 5.7000 2877.2800 ;
      RECT 0.0000 2874.5600 3390.2000 2876.2000 ;
      RECT 3388.5000 2873.4800 3390.2000 2874.5600 ;
      RECT 5.3000 2873.4800 3384.9000 2874.5600 ;
      RECT 0.0000 2873.4800 1.7000 2874.5600 ;
      RECT 0.0000 2871.8400 3390.2000 2873.4800 ;
      RECT 3384.5000 2870.7600 3390.2000 2871.8400 ;
      RECT 9.3000 2870.7600 3380.9000 2871.8400 ;
      RECT 0.0000 2870.7600 5.7000 2871.8400 ;
      RECT 0.0000 2869.1200 3390.2000 2870.7600 ;
      RECT 3388.5000 2868.0400 3390.2000 2869.1200 ;
      RECT 5.3000 2868.0400 3384.9000 2869.1200 ;
      RECT 0.0000 2868.0400 1.7000 2869.1200 ;
      RECT 0.0000 2866.4000 3390.2000 2868.0400 ;
      RECT 3384.5000 2865.3200 3390.2000 2866.4000 ;
      RECT 9.3000 2865.3200 3380.9000 2866.4000 ;
      RECT 0.0000 2865.3200 5.7000 2866.4000 ;
      RECT 0.0000 2863.6800 3390.2000 2865.3200 ;
      RECT 3388.5000 2862.6000 3390.2000 2863.6800 ;
      RECT 5.3000 2862.6000 3384.9000 2863.6800 ;
      RECT 0.0000 2862.6000 1.7000 2863.6800 ;
      RECT 0.0000 2860.9600 3390.2000 2862.6000 ;
      RECT 3384.5000 2859.8800 3390.2000 2860.9600 ;
      RECT 9.3000 2859.8800 3380.9000 2860.9600 ;
      RECT 0.0000 2859.8800 5.7000 2860.9600 ;
      RECT 0.0000 2858.2400 3390.2000 2859.8800 ;
      RECT 3388.5000 2857.1600 3390.2000 2858.2400 ;
      RECT 5.3000 2857.1600 3384.9000 2858.2400 ;
      RECT 0.0000 2857.1600 1.7000 2858.2400 ;
      RECT 0.0000 2855.5200 3390.2000 2857.1600 ;
      RECT 3384.5000 2854.4400 3390.2000 2855.5200 ;
      RECT 9.3000 2854.4400 3380.9000 2855.5200 ;
      RECT 0.0000 2854.4400 5.7000 2855.5200 ;
      RECT 0.0000 2852.8000 3390.2000 2854.4400 ;
      RECT 3388.5000 2851.7200 3390.2000 2852.8000 ;
      RECT 5.3000 2851.7200 3384.9000 2852.8000 ;
      RECT 0.0000 2851.7200 1.7000 2852.8000 ;
      RECT 0.0000 2850.0800 3390.2000 2851.7200 ;
      RECT 3384.5000 2849.0000 3390.2000 2850.0800 ;
      RECT 9.3000 2849.0000 3380.9000 2850.0800 ;
      RECT 0.0000 2849.0000 5.7000 2850.0800 ;
      RECT 0.0000 2847.3600 3390.2000 2849.0000 ;
      RECT 3388.5000 2846.2800 3390.2000 2847.3600 ;
      RECT 5.3000 2846.2800 3384.9000 2847.3600 ;
      RECT 0.0000 2846.2800 1.7000 2847.3600 ;
      RECT 0.0000 2844.6400 3390.2000 2846.2800 ;
      RECT 3384.5000 2843.5600 3390.2000 2844.6400 ;
      RECT 9.3000 2843.5600 3380.9000 2844.6400 ;
      RECT 0.0000 2843.5600 5.7000 2844.6400 ;
      RECT 0.0000 2841.9200 3390.2000 2843.5600 ;
      RECT 3388.5000 2840.8400 3390.2000 2841.9200 ;
      RECT 5.3000 2840.8400 3384.9000 2841.9200 ;
      RECT 0.0000 2840.8400 1.7000 2841.9200 ;
      RECT 0.0000 2839.2000 3390.2000 2840.8400 ;
      RECT 3384.5000 2838.1200 3390.2000 2839.2000 ;
      RECT 9.3000 2838.1200 3380.9000 2839.2000 ;
      RECT 0.0000 2838.1200 5.7000 2839.2000 ;
      RECT 0.0000 2836.4800 3390.2000 2838.1200 ;
      RECT 3388.5000 2835.4000 3390.2000 2836.4800 ;
      RECT 5.3000 2835.4000 3384.9000 2836.4800 ;
      RECT 0.0000 2835.4000 1.7000 2836.4800 ;
      RECT 0.0000 2833.7600 3390.2000 2835.4000 ;
      RECT 3384.5000 2832.6800 3390.2000 2833.7600 ;
      RECT 9.3000 2832.6800 3380.9000 2833.7600 ;
      RECT 0.0000 2832.6800 5.7000 2833.7600 ;
      RECT 0.0000 2831.0400 3390.2000 2832.6800 ;
      RECT 3388.5000 2829.9600 3390.2000 2831.0400 ;
      RECT 5.3000 2829.9600 3384.9000 2831.0400 ;
      RECT 0.0000 2829.9600 1.7000 2831.0400 ;
      RECT 0.0000 2828.3200 3390.2000 2829.9600 ;
      RECT 3384.5000 2827.2400 3390.2000 2828.3200 ;
      RECT 9.3000 2827.2400 3380.9000 2828.3200 ;
      RECT 0.0000 2827.2400 5.7000 2828.3200 ;
      RECT 0.0000 2825.6000 3390.2000 2827.2400 ;
      RECT 3388.5000 2824.5200 3390.2000 2825.6000 ;
      RECT 5.3000 2824.5200 3384.9000 2825.6000 ;
      RECT 0.0000 2824.5200 1.7000 2825.6000 ;
      RECT 0.0000 2822.8800 3390.2000 2824.5200 ;
      RECT 3384.5000 2821.8000 3390.2000 2822.8800 ;
      RECT 9.3000 2821.8000 3380.9000 2822.8800 ;
      RECT 0.0000 2821.8000 5.7000 2822.8800 ;
      RECT 0.0000 2820.1600 3390.2000 2821.8000 ;
      RECT 3388.5000 2819.0800 3390.2000 2820.1600 ;
      RECT 5.3000 2819.0800 3384.9000 2820.1600 ;
      RECT 0.0000 2819.0800 1.7000 2820.1600 ;
      RECT 0.0000 2817.4400 3390.2000 2819.0800 ;
      RECT 3384.5000 2816.3600 3390.2000 2817.4400 ;
      RECT 9.3000 2816.3600 3380.9000 2817.4400 ;
      RECT 0.0000 2816.3600 5.7000 2817.4400 ;
      RECT 0.0000 2814.7200 3390.2000 2816.3600 ;
      RECT 3388.5000 2813.6400 3390.2000 2814.7200 ;
      RECT 5.3000 2813.6400 3384.9000 2814.7200 ;
      RECT 0.0000 2813.6400 1.7000 2814.7200 ;
      RECT 0.0000 2812.0000 3390.2000 2813.6400 ;
      RECT 3384.5000 2810.9200 3390.2000 2812.0000 ;
      RECT 9.3000 2810.9200 3380.9000 2812.0000 ;
      RECT 0.0000 2810.9200 5.7000 2812.0000 ;
      RECT 0.0000 2809.2800 3390.2000 2810.9200 ;
      RECT 3388.5000 2808.2000 3390.2000 2809.2800 ;
      RECT 5.3000 2808.2000 3384.9000 2809.2800 ;
      RECT 0.0000 2808.2000 1.7000 2809.2800 ;
      RECT 0.0000 2806.5600 3390.2000 2808.2000 ;
      RECT 3384.5000 2805.4800 3390.2000 2806.5600 ;
      RECT 9.3000 2805.4800 3380.9000 2806.5600 ;
      RECT 0.0000 2805.4800 5.7000 2806.5600 ;
      RECT 0.0000 2803.8400 3390.2000 2805.4800 ;
      RECT 3388.5000 2802.7600 3390.2000 2803.8400 ;
      RECT 5.3000 2802.7600 3384.9000 2803.8400 ;
      RECT 0.0000 2802.7600 1.7000 2803.8400 ;
      RECT 0.0000 2801.1200 3390.2000 2802.7600 ;
      RECT 3384.5000 2800.0400 3390.2000 2801.1200 ;
      RECT 9.3000 2800.0400 3380.9000 2801.1200 ;
      RECT 0.0000 2800.0400 5.7000 2801.1200 ;
      RECT 0.0000 2800.0100 3390.2000 2800.0400 ;
      RECT 1.1000 2799.1100 3389.1000 2800.0100 ;
      RECT 0.0000 2798.4000 3390.2000 2799.1100 ;
      RECT 3388.5000 2797.3200 3390.2000 2798.4000 ;
      RECT 5.3000 2797.3200 3384.9000 2798.4000 ;
      RECT 0.0000 2797.3200 1.7000 2798.4000 ;
      RECT 0.0000 2795.6800 3390.2000 2797.3200 ;
      RECT 3384.5000 2794.6000 3390.2000 2795.6800 ;
      RECT 9.3000 2794.6000 3380.9000 2795.6800 ;
      RECT 0.0000 2794.6000 5.7000 2795.6800 ;
      RECT 0.0000 2792.9600 3390.2000 2794.6000 ;
      RECT 3388.5000 2791.8800 3390.2000 2792.9600 ;
      RECT 5.3000 2791.8800 3384.9000 2792.9600 ;
      RECT 0.0000 2791.8800 1.7000 2792.9600 ;
      RECT 0.0000 2790.2400 3390.2000 2791.8800 ;
      RECT 3384.5000 2789.1600 3390.2000 2790.2400 ;
      RECT 9.3000 2789.1600 3380.9000 2790.2400 ;
      RECT 0.0000 2789.1600 5.7000 2790.2400 ;
      RECT 0.0000 2787.5200 3390.2000 2789.1600 ;
      RECT 3388.5000 2786.4400 3390.2000 2787.5200 ;
      RECT 5.3000 2786.4400 3384.9000 2787.5200 ;
      RECT 0.0000 2786.4400 1.7000 2787.5200 ;
      RECT 0.0000 2784.8000 3390.2000 2786.4400 ;
      RECT 3384.5000 2783.7200 3390.2000 2784.8000 ;
      RECT 9.3000 2783.7200 3380.9000 2784.8000 ;
      RECT 0.0000 2783.7200 5.7000 2784.8000 ;
      RECT 0.0000 2782.0800 3390.2000 2783.7200 ;
      RECT 3388.5000 2781.0000 3390.2000 2782.0800 ;
      RECT 5.3000 2781.0000 3384.9000 2782.0800 ;
      RECT 0.0000 2781.0000 1.7000 2782.0800 ;
      RECT 0.0000 2779.3600 3390.2000 2781.0000 ;
      RECT 3384.5000 2778.2800 3390.2000 2779.3600 ;
      RECT 9.3000 2778.2800 3380.9000 2779.3600 ;
      RECT 0.0000 2778.2800 5.7000 2779.3600 ;
      RECT 0.0000 2776.6400 3390.2000 2778.2800 ;
      RECT 3388.5000 2775.5600 3390.2000 2776.6400 ;
      RECT 5.3000 2775.5600 3384.9000 2776.6400 ;
      RECT 0.0000 2775.5600 1.7000 2776.6400 ;
      RECT 0.0000 2775.0000 3390.2000 2775.5600 ;
      RECT 1.1000 2774.1000 3390.2000 2775.0000 ;
      RECT 0.0000 2773.9200 3390.2000 2774.1000 ;
      RECT 3384.5000 2772.8400 3390.2000 2773.9200 ;
      RECT 9.3000 2772.8400 3380.9000 2773.9200 ;
      RECT 0.0000 2772.8400 5.7000 2773.9200 ;
      RECT 0.0000 2771.2000 3390.2000 2772.8400 ;
      RECT 3388.5000 2770.1200 3390.2000 2771.2000 ;
      RECT 5.3000 2770.1200 3384.9000 2771.2000 ;
      RECT 0.0000 2770.1200 1.7000 2771.2000 ;
      RECT 0.0000 2768.4800 3390.2000 2770.1200 ;
      RECT 3384.5000 2767.4000 3390.2000 2768.4800 ;
      RECT 9.3000 2767.4000 3380.9000 2768.4800 ;
      RECT 0.0000 2767.4000 5.7000 2768.4800 ;
      RECT 0.0000 2765.7600 3390.2000 2767.4000 ;
      RECT 3388.5000 2764.6800 3390.2000 2765.7600 ;
      RECT 5.3000 2764.6800 3384.9000 2765.7600 ;
      RECT 0.0000 2764.6800 1.7000 2765.7600 ;
      RECT 0.0000 2763.0400 3390.2000 2764.6800 ;
      RECT 3384.5000 2761.9600 3390.2000 2763.0400 ;
      RECT 9.3000 2761.9600 3380.9000 2763.0400 ;
      RECT 0.0000 2761.9600 5.7000 2763.0400 ;
      RECT 0.0000 2760.3200 3390.2000 2761.9600 ;
      RECT 3388.5000 2759.2400 3390.2000 2760.3200 ;
      RECT 5.3000 2759.2400 3384.9000 2760.3200 ;
      RECT 0.0000 2759.2400 1.7000 2760.3200 ;
      RECT 0.0000 2757.6000 3390.2000 2759.2400 ;
      RECT 3384.5000 2756.5200 3390.2000 2757.6000 ;
      RECT 9.3000 2756.5200 3380.9000 2757.6000 ;
      RECT 0.0000 2756.5200 5.7000 2757.6000 ;
      RECT 0.0000 2754.8800 3390.2000 2756.5200 ;
      RECT 3388.5000 2753.8000 3390.2000 2754.8800 ;
      RECT 5.3000 2753.8000 3384.9000 2754.8800 ;
      RECT 0.0000 2753.8000 1.7000 2754.8800 ;
      RECT 0.0000 2752.1600 3390.2000 2753.8000 ;
      RECT 3384.5000 2751.0800 3390.2000 2752.1600 ;
      RECT 9.3000 2751.0800 3380.9000 2752.1600 ;
      RECT 0.0000 2751.0800 5.7000 2752.1600 ;
      RECT 0.0000 2749.9900 3390.2000 2751.0800 ;
      RECT 1.1000 2749.4400 3390.2000 2749.9900 ;
      RECT 1.1000 2749.0900 1.7000 2749.4400 ;
      RECT 3388.5000 2748.3600 3390.2000 2749.4400 ;
      RECT 5.3000 2748.3600 3384.9000 2749.4400 ;
      RECT 0.0000 2748.3600 1.7000 2749.0900 ;
      RECT 0.0000 2746.7200 3390.2000 2748.3600 ;
      RECT 3384.5000 2745.6400 3390.2000 2746.7200 ;
      RECT 9.3000 2745.6400 3380.9000 2746.7200 ;
      RECT 0.0000 2745.6400 5.7000 2746.7200 ;
      RECT 0.0000 2744.0000 3390.2000 2745.6400 ;
      RECT 3388.5000 2742.9200 3390.2000 2744.0000 ;
      RECT 5.3000 2742.9200 3384.9000 2744.0000 ;
      RECT 0.0000 2742.9200 1.7000 2744.0000 ;
      RECT 0.0000 2741.2800 3390.2000 2742.9200 ;
      RECT 3384.5000 2740.2000 3390.2000 2741.2800 ;
      RECT 9.3000 2740.2000 3380.9000 2741.2800 ;
      RECT 0.0000 2740.2000 5.7000 2741.2800 ;
      RECT 0.0000 2738.5600 3390.2000 2740.2000 ;
      RECT 3388.5000 2737.4800 3390.2000 2738.5600 ;
      RECT 5.3000 2737.4800 3384.9000 2738.5600 ;
      RECT 0.0000 2737.4800 1.7000 2738.5600 ;
      RECT 0.0000 2735.8400 3390.2000 2737.4800 ;
      RECT 3384.5000 2734.7600 3390.2000 2735.8400 ;
      RECT 9.3000 2734.7600 3380.9000 2735.8400 ;
      RECT 0.0000 2734.7600 5.7000 2735.8400 ;
      RECT 0.0000 2733.1200 3390.2000 2734.7600 ;
      RECT 3388.5000 2732.0400 3390.2000 2733.1200 ;
      RECT 5.3000 2732.0400 3384.9000 2733.1200 ;
      RECT 0.0000 2732.0400 1.7000 2733.1200 ;
      RECT 0.0000 2730.4000 3390.2000 2732.0400 ;
      RECT 3384.5000 2729.3200 3390.2000 2730.4000 ;
      RECT 9.3000 2729.3200 3380.9000 2730.4000 ;
      RECT 0.0000 2729.3200 5.7000 2730.4000 ;
      RECT 0.0000 2727.6800 3390.2000 2729.3200 ;
      RECT 3388.5000 2726.6000 3390.2000 2727.6800 ;
      RECT 5.3000 2726.6000 3384.9000 2727.6800 ;
      RECT 0.0000 2726.6000 1.7000 2727.6800 ;
      RECT 0.0000 2724.9600 3390.2000 2726.6000 ;
      RECT 0.0000 2724.3700 5.7000 2724.9600 ;
      RECT 3384.5000 2723.8800 3390.2000 2724.9600 ;
      RECT 9.3000 2723.8800 3380.9000 2724.9600 ;
      RECT 1.1000 2723.8800 5.7000 2724.3700 ;
      RECT 1.1000 2723.4700 3390.2000 2723.8800 ;
      RECT 0.0000 2722.2400 3390.2000 2723.4700 ;
      RECT 3388.5000 2721.1600 3390.2000 2722.2400 ;
      RECT 5.3000 2721.1600 3384.9000 2722.2400 ;
      RECT 0.0000 2721.1600 1.7000 2722.2400 ;
      RECT 0.0000 2719.5200 3390.2000 2721.1600 ;
      RECT 3384.5000 2718.4400 3390.2000 2719.5200 ;
      RECT 9.3000 2718.4400 3380.9000 2719.5200 ;
      RECT 0.0000 2718.4400 5.7000 2719.5200 ;
      RECT 0.0000 2716.8000 3390.2000 2718.4400 ;
      RECT 3388.5000 2715.7200 3390.2000 2716.8000 ;
      RECT 5.3000 2715.7200 3384.9000 2716.8000 ;
      RECT 0.0000 2715.7200 1.7000 2716.8000 ;
      RECT 0.0000 2714.0800 3390.2000 2715.7200 ;
      RECT 3384.5000 2713.0000 3390.2000 2714.0800 ;
      RECT 9.3000 2713.0000 3380.9000 2714.0800 ;
      RECT 0.0000 2713.0000 5.7000 2714.0800 ;
      RECT 0.0000 2711.3600 3390.2000 2713.0000 ;
      RECT 3388.5000 2710.2800 3390.2000 2711.3600 ;
      RECT 5.3000 2710.2800 3384.9000 2711.3600 ;
      RECT 0.0000 2710.2800 1.7000 2711.3600 ;
      RECT 0.0000 2708.6400 3390.2000 2710.2800 ;
      RECT 3384.5000 2707.5600 3390.2000 2708.6400 ;
      RECT 9.3000 2707.5600 3380.9000 2708.6400 ;
      RECT 0.0000 2707.5600 5.7000 2708.6400 ;
      RECT 0.0000 2705.9200 3390.2000 2707.5600 ;
      RECT 3388.5000 2704.8400 3390.2000 2705.9200 ;
      RECT 5.3000 2704.8400 3384.9000 2705.9200 ;
      RECT 0.0000 2704.8400 1.7000 2705.9200 ;
      RECT 0.0000 2703.2000 3390.2000 2704.8400 ;
      RECT 3384.5000 2702.1200 3390.2000 2703.2000 ;
      RECT 9.3000 2702.1200 3380.9000 2703.2000 ;
      RECT 0.0000 2702.1200 5.7000 2703.2000 ;
      RECT 0.0000 2700.4800 3390.2000 2702.1200 ;
      RECT 3388.5000 2699.4000 3390.2000 2700.4800 ;
      RECT 5.3000 2699.4000 3384.9000 2700.4800 ;
      RECT 0.0000 2699.4000 1.7000 2700.4800 ;
      RECT 0.0000 2699.3600 3390.2000 2699.4000 ;
      RECT 1.1000 2698.4600 3390.2000 2699.3600 ;
      RECT 0.0000 2697.7600 3390.2000 2698.4600 ;
      RECT 3384.5000 2696.6800 3390.2000 2697.7600 ;
      RECT 9.3000 2696.6800 3380.9000 2697.7600 ;
      RECT 0.0000 2696.6800 5.7000 2697.7600 ;
      RECT 0.0000 2696.3100 3390.2000 2696.6800 ;
      RECT 0.0000 2695.4100 3389.1000 2696.3100 ;
      RECT 0.0000 2695.0400 3390.2000 2695.4100 ;
      RECT 3388.5000 2693.9600 3390.2000 2695.0400 ;
      RECT 5.3000 2693.9600 3384.9000 2695.0400 ;
      RECT 0.0000 2693.9600 1.7000 2695.0400 ;
      RECT 0.0000 2692.3200 3390.2000 2693.9600 ;
      RECT 3384.5000 2691.2400 3390.2000 2692.3200 ;
      RECT 9.3000 2691.2400 3380.9000 2692.3200 ;
      RECT 0.0000 2691.2400 5.7000 2692.3200 ;
      RECT 0.0000 2689.6000 3390.2000 2691.2400 ;
      RECT 3388.5000 2688.5200 3390.2000 2689.6000 ;
      RECT 5.3000 2688.5200 3384.9000 2689.6000 ;
      RECT 0.0000 2688.5200 1.7000 2689.6000 ;
      RECT 0.0000 2686.8800 3390.2000 2688.5200 ;
      RECT 3384.5000 2685.8000 3390.2000 2686.8800 ;
      RECT 9.3000 2685.8000 3380.9000 2686.8800 ;
      RECT 0.0000 2685.8000 5.7000 2686.8800 ;
      RECT 0.0000 2684.1600 3390.2000 2685.8000 ;
      RECT 3388.5000 2683.0800 3390.2000 2684.1600 ;
      RECT 5.3000 2683.0800 3384.9000 2684.1600 ;
      RECT 0.0000 2683.0800 1.7000 2684.1600 ;
      RECT 0.0000 2681.4400 3390.2000 2683.0800 ;
      RECT 3384.5000 2680.3600 3390.2000 2681.4400 ;
      RECT 9.3000 2680.3600 3380.9000 2681.4400 ;
      RECT 0.0000 2680.3600 5.7000 2681.4400 ;
      RECT 0.0000 2678.7200 3390.2000 2680.3600 ;
      RECT 3388.5000 2677.6400 3390.2000 2678.7200 ;
      RECT 5.3000 2677.6400 3384.9000 2678.7200 ;
      RECT 0.0000 2677.6400 1.7000 2678.7200 ;
      RECT 0.0000 2676.0000 3390.2000 2677.6400 ;
      RECT 3384.5000 2674.9200 3390.2000 2676.0000 ;
      RECT 9.3000 2674.9200 3380.9000 2676.0000 ;
      RECT 0.0000 2674.9200 5.7000 2676.0000 ;
      RECT 0.0000 2674.3500 3390.2000 2674.9200 ;
      RECT 1.1000 2673.4500 3390.2000 2674.3500 ;
      RECT 0.0000 2673.2800 3390.2000 2673.4500 ;
      RECT 3388.5000 2672.2000 3390.2000 2673.2800 ;
      RECT 5.3000 2672.2000 3384.9000 2673.2800 ;
      RECT 0.0000 2672.2000 1.7000 2673.2800 ;
      RECT 0.0000 2670.5600 3390.2000 2672.2000 ;
      RECT 3384.5000 2669.4800 3390.2000 2670.5600 ;
      RECT 9.3000 2669.4800 3380.9000 2670.5600 ;
      RECT 0.0000 2669.4800 5.7000 2670.5600 ;
      RECT 0.0000 2667.8400 3390.2000 2669.4800 ;
      RECT 3388.5000 2666.7600 3390.2000 2667.8400 ;
      RECT 5.3000 2666.7600 3384.9000 2667.8400 ;
      RECT 0.0000 2666.7600 1.7000 2667.8400 ;
      RECT 0.0000 2665.1200 3390.2000 2666.7600 ;
      RECT 3384.5000 2664.0400 3390.2000 2665.1200 ;
      RECT 9.3000 2664.0400 3380.9000 2665.1200 ;
      RECT 0.0000 2664.0400 5.7000 2665.1200 ;
      RECT 0.0000 2662.4000 3390.2000 2664.0400 ;
      RECT 3388.5000 2661.3200 3390.2000 2662.4000 ;
      RECT 5.3000 2661.3200 3384.9000 2662.4000 ;
      RECT 0.0000 2661.3200 1.7000 2662.4000 ;
      RECT 0.0000 2659.6800 3390.2000 2661.3200 ;
      RECT 3384.5000 2658.6000 3390.2000 2659.6800 ;
      RECT 9.3000 2658.6000 3380.9000 2659.6800 ;
      RECT 0.0000 2658.6000 5.7000 2659.6800 ;
      RECT 0.0000 2656.9600 3390.2000 2658.6000 ;
      RECT 3388.5000 2655.8800 3390.2000 2656.9600 ;
      RECT 5.3000 2655.8800 3384.9000 2656.9600 ;
      RECT 0.0000 2655.8800 1.7000 2656.9600 ;
      RECT 0.0000 2654.2400 3390.2000 2655.8800 ;
      RECT 3384.5000 2653.1600 3390.2000 2654.2400 ;
      RECT 9.3000 2653.1600 3380.9000 2654.2400 ;
      RECT 0.0000 2653.1600 5.7000 2654.2400 ;
      RECT 0.0000 2651.5200 3390.2000 2653.1600 ;
      RECT 3388.5000 2650.4400 3390.2000 2651.5200 ;
      RECT 5.3000 2650.4400 3384.9000 2651.5200 ;
      RECT 0.0000 2650.4400 1.7000 2651.5200 ;
      RECT 0.0000 2648.8000 3390.2000 2650.4400 ;
      RECT 0.0000 2648.7300 5.7000 2648.8000 ;
      RECT 1.1000 2647.8300 5.7000 2648.7300 ;
      RECT 3384.5000 2647.7200 3390.2000 2648.8000 ;
      RECT 9.3000 2647.7200 3380.9000 2648.8000 ;
      RECT 0.0000 2647.7200 5.7000 2647.8300 ;
      RECT 0.0000 2646.0800 3390.2000 2647.7200 ;
      RECT 3388.5000 2645.0000 3390.2000 2646.0800 ;
      RECT 5.3000 2645.0000 3384.9000 2646.0800 ;
      RECT 0.0000 2645.0000 1.7000 2646.0800 ;
      RECT 0.0000 2643.3600 3390.2000 2645.0000 ;
      RECT 3384.5000 2642.2800 3390.2000 2643.3600 ;
      RECT 9.3000 2642.2800 3380.9000 2643.3600 ;
      RECT 0.0000 2642.2800 5.7000 2643.3600 ;
      RECT 0.0000 2640.6400 3390.2000 2642.2800 ;
      RECT 3388.5000 2639.5600 3390.2000 2640.6400 ;
      RECT 5.3000 2639.5600 3384.9000 2640.6400 ;
      RECT 0.0000 2639.5600 1.7000 2640.6400 ;
      RECT 0.0000 2637.9200 3390.2000 2639.5600 ;
      RECT 3384.5000 2636.8400 3390.2000 2637.9200 ;
      RECT 9.3000 2636.8400 3380.9000 2637.9200 ;
      RECT 0.0000 2636.8400 5.7000 2637.9200 ;
      RECT 0.0000 2635.2000 3390.2000 2636.8400 ;
      RECT 3388.5000 2634.1200 3390.2000 2635.2000 ;
      RECT 5.3000 2634.1200 3384.9000 2635.2000 ;
      RECT 0.0000 2634.1200 1.7000 2635.2000 ;
      RECT 0.0000 2632.4800 3390.2000 2634.1200 ;
      RECT 3384.5000 2631.4000 3390.2000 2632.4800 ;
      RECT 9.3000 2631.4000 3380.9000 2632.4800 ;
      RECT 0.0000 2631.4000 5.7000 2632.4800 ;
      RECT 0.0000 2629.7600 3390.2000 2631.4000 ;
      RECT 3388.5000 2628.6800 3390.2000 2629.7600 ;
      RECT 5.3000 2628.6800 3384.9000 2629.7600 ;
      RECT 0.0000 2628.6800 1.7000 2629.7600 ;
      RECT 0.0000 2627.0400 3390.2000 2628.6800 ;
      RECT 3384.5000 2625.9600 3390.2000 2627.0400 ;
      RECT 9.3000 2625.9600 3380.9000 2627.0400 ;
      RECT 0.0000 2625.9600 5.7000 2627.0400 ;
      RECT 0.0000 2624.3200 3390.2000 2625.9600 ;
      RECT 0.0000 2623.7200 1.7000 2624.3200 ;
      RECT 3388.5000 2623.2400 3390.2000 2624.3200 ;
      RECT 5.3000 2623.2400 3384.9000 2624.3200 ;
      RECT 1.1000 2623.2400 1.7000 2623.7200 ;
      RECT 1.1000 2622.8200 3390.2000 2623.2400 ;
      RECT 0.0000 2621.6000 3390.2000 2622.8200 ;
      RECT 3384.5000 2620.5200 3390.2000 2621.6000 ;
      RECT 9.3000 2620.5200 3380.9000 2621.6000 ;
      RECT 0.0000 2620.5200 5.7000 2621.6000 ;
      RECT 0.0000 2618.8800 3390.2000 2620.5200 ;
      RECT 3388.5000 2617.8000 3390.2000 2618.8800 ;
      RECT 5.3000 2617.8000 3384.9000 2618.8800 ;
      RECT 0.0000 2617.8000 1.7000 2618.8800 ;
      RECT 0.0000 2616.1600 3390.2000 2617.8000 ;
      RECT 3384.5000 2615.0800 3390.2000 2616.1600 ;
      RECT 9.3000 2615.0800 3380.9000 2616.1600 ;
      RECT 0.0000 2615.0800 5.7000 2616.1600 ;
      RECT 0.0000 2613.4400 3390.2000 2615.0800 ;
      RECT 3388.5000 2612.3600 3390.2000 2613.4400 ;
      RECT 5.3000 2612.3600 3384.9000 2613.4400 ;
      RECT 0.0000 2612.3600 1.7000 2613.4400 ;
      RECT 0.0000 2610.7200 3390.2000 2612.3600 ;
      RECT 3384.5000 2609.6400 3390.2000 2610.7200 ;
      RECT 9.3000 2609.6400 3380.9000 2610.7200 ;
      RECT 0.0000 2609.6400 5.7000 2610.7200 ;
      RECT 0.0000 2608.0000 3390.2000 2609.6400 ;
      RECT 3388.5000 2606.9200 3390.2000 2608.0000 ;
      RECT 5.3000 2606.9200 3384.9000 2608.0000 ;
      RECT 0.0000 2606.9200 1.7000 2608.0000 ;
      RECT 0.0000 2605.2800 3390.2000 2606.9200 ;
      RECT 3384.5000 2604.2000 3390.2000 2605.2800 ;
      RECT 9.3000 2604.2000 3380.9000 2605.2800 ;
      RECT 0.0000 2604.2000 5.7000 2605.2800 ;
      RECT 0.0000 2602.5600 3390.2000 2604.2000 ;
      RECT 3388.5000 2601.4800 3390.2000 2602.5600 ;
      RECT 5.3000 2601.4800 3384.9000 2602.5600 ;
      RECT 0.0000 2601.4800 1.7000 2602.5600 ;
      RECT 0.0000 2599.8400 3390.2000 2601.4800 ;
      RECT 3384.5000 2598.7600 3390.2000 2599.8400 ;
      RECT 9.3000 2598.7600 3380.9000 2599.8400 ;
      RECT 0.0000 2598.7600 5.7000 2599.8400 ;
      RECT 0.0000 2598.7100 3390.2000 2598.7600 ;
      RECT 1.1000 2597.8100 3390.2000 2598.7100 ;
      RECT 0.0000 2597.1200 3390.2000 2597.8100 ;
      RECT 3388.5000 2596.0400 3390.2000 2597.1200 ;
      RECT 5.3000 2596.0400 3384.9000 2597.1200 ;
      RECT 0.0000 2596.0400 1.7000 2597.1200 ;
      RECT 0.0000 2594.4000 3390.2000 2596.0400 ;
      RECT 3384.5000 2593.3200 3390.2000 2594.4000 ;
      RECT 9.3000 2593.3200 3380.9000 2594.4000 ;
      RECT 0.0000 2593.3200 5.7000 2594.4000 ;
      RECT 0.0000 2592.6100 3390.2000 2593.3200 ;
      RECT 0.0000 2591.7100 3389.1000 2592.6100 ;
      RECT 0.0000 2591.6800 3390.2000 2591.7100 ;
      RECT 3388.5000 2590.6000 3390.2000 2591.6800 ;
      RECT 5.3000 2590.6000 3384.9000 2591.6800 ;
      RECT 0.0000 2590.6000 1.7000 2591.6800 ;
      RECT 0.0000 2588.9600 3390.2000 2590.6000 ;
      RECT 3384.5000 2587.8800 3390.2000 2588.9600 ;
      RECT 9.3000 2587.8800 3380.9000 2588.9600 ;
      RECT 0.0000 2587.8800 5.7000 2588.9600 ;
      RECT 0.0000 2586.2400 3390.2000 2587.8800 ;
      RECT 3388.5000 2585.1600 3390.2000 2586.2400 ;
      RECT 5.3000 2585.1600 3384.9000 2586.2400 ;
      RECT 0.0000 2585.1600 1.7000 2586.2400 ;
      RECT 0.0000 2583.5200 3390.2000 2585.1600 ;
      RECT 3384.5000 2582.4400 3390.2000 2583.5200 ;
      RECT 9.3000 2582.4400 3380.9000 2583.5200 ;
      RECT 0.0000 2582.4400 5.7000 2583.5200 ;
      RECT 0.0000 2580.8000 3390.2000 2582.4400 ;
      RECT 3388.5000 2579.7200 3390.2000 2580.8000 ;
      RECT 5.3000 2579.7200 3384.9000 2580.8000 ;
      RECT 0.0000 2579.7200 1.7000 2580.8000 ;
      RECT 0.0000 2578.0800 3390.2000 2579.7200 ;
      RECT 3384.5000 2577.0000 3390.2000 2578.0800 ;
      RECT 9.3000 2577.0000 3380.9000 2578.0800 ;
      RECT 0.0000 2577.0000 5.7000 2578.0800 ;
      RECT 0.0000 2575.3600 3390.2000 2577.0000 ;
      RECT 3388.5000 2574.2800 3390.2000 2575.3600 ;
      RECT 5.3000 2574.2800 3384.9000 2575.3600 ;
      RECT 0.0000 2574.2800 1.7000 2575.3600 ;
      RECT 0.0000 2573.0900 3390.2000 2574.2800 ;
      RECT 1.1000 2572.6400 3390.2000 2573.0900 ;
      RECT 1.1000 2572.1900 5.7000 2572.6400 ;
      RECT 3384.5000 2571.5600 3390.2000 2572.6400 ;
      RECT 9.3000 2571.5600 3380.9000 2572.6400 ;
      RECT 0.0000 2571.5600 5.7000 2572.1900 ;
      RECT 0.0000 2569.9200 3390.2000 2571.5600 ;
      RECT 3388.5000 2568.8400 3390.2000 2569.9200 ;
      RECT 5.3000 2568.8400 3384.9000 2569.9200 ;
      RECT 0.0000 2568.8400 1.7000 2569.9200 ;
      RECT 0.0000 2567.2000 3390.2000 2568.8400 ;
      RECT 3384.5000 2566.1200 3390.2000 2567.2000 ;
      RECT 9.3000 2566.1200 3380.9000 2567.2000 ;
      RECT 0.0000 2566.1200 5.7000 2567.2000 ;
      RECT 0.0000 2564.4800 3390.2000 2566.1200 ;
      RECT 3388.5000 2563.4000 3390.2000 2564.4800 ;
      RECT 5.3000 2563.4000 3384.9000 2564.4800 ;
      RECT 0.0000 2563.4000 1.7000 2564.4800 ;
      RECT 0.0000 2561.7600 3390.2000 2563.4000 ;
      RECT 3384.5000 2560.6800 3390.2000 2561.7600 ;
      RECT 9.3000 2560.6800 3380.9000 2561.7600 ;
      RECT 0.0000 2560.6800 5.7000 2561.7600 ;
      RECT 0.0000 2559.0400 3390.2000 2560.6800 ;
      RECT 3388.5000 2557.9600 3390.2000 2559.0400 ;
      RECT 5.3000 2557.9600 3384.9000 2559.0400 ;
      RECT 0.0000 2557.9600 1.7000 2559.0400 ;
      RECT 0.0000 2556.3200 3390.2000 2557.9600 ;
      RECT 3384.5000 2555.2400 3390.2000 2556.3200 ;
      RECT 9.3000 2555.2400 3380.9000 2556.3200 ;
      RECT 0.0000 2555.2400 5.7000 2556.3200 ;
      RECT 0.0000 2553.6000 3390.2000 2555.2400 ;
      RECT 3388.5000 2552.5200 3390.2000 2553.6000 ;
      RECT 5.3000 2552.5200 3384.9000 2553.6000 ;
      RECT 0.0000 2552.5200 1.7000 2553.6000 ;
      RECT 0.0000 2550.8800 3390.2000 2552.5200 ;
      RECT 3384.5000 2549.8000 3390.2000 2550.8800 ;
      RECT 9.3000 2549.8000 3380.9000 2550.8800 ;
      RECT 0.0000 2549.8000 5.7000 2550.8800 ;
      RECT 0.0000 2548.1600 3390.2000 2549.8000 ;
      RECT 0.0000 2548.0800 1.7000 2548.1600 ;
      RECT 1.1000 2547.1800 1.7000 2548.0800 ;
      RECT 3388.5000 2547.0800 3390.2000 2548.1600 ;
      RECT 5.3000 2547.0800 3384.9000 2548.1600 ;
      RECT 0.0000 2547.0800 1.7000 2547.1800 ;
      RECT 0.0000 2545.4400 3390.2000 2547.0800 ;
      RECT 3384.5000 2544.3600 3390.2000 2545.4400 ;
      RECT 9.3000 2544.3600 3380.9000 2545.4400 ;
      RECT 0.0000 2544.3600 5.7000 2545.4400 ;
      RECT 0.0000 2542.7200 3390.2000 2544.3600 ;
      RECT 3388.5000 2541.6400 3390.2000 2542.7200 ;
      RECT 5.3000 2541.6400 3384.9000 2542.7200 ;
      RECT 0.0000 2541.6400 1.7000 2542.7200 ;
      RECT 0.0000 2540.0000 3390.2000 2541.6400 ;
      RECT 3384.5000 2538.9200 3390.2000 2540.0000 ;
      RECT 9.3000 2538.9200 3380.9000 2540.0000 ;
      RECT 0.0000 2538.9200 5.7000 2540.0000 ;
      RECT 0.0000 2537.2800 3390.2000 2538.9200 ;
      RECT 3388.5000 2536.2000 3390.2000 2537.2800 ;
      RECT 5.3000 2536.2000 3384.9000 2537.2800 ;
      RECT 0.0000 2536.2000 1.7000 2537.2800 ;
      RECT 0.0000 2534.5600 3390.2000 2536.2000 ;
      RECT 3384.5000 2533.4800 3390.2000 2534.5600 ;
      RECT 9.3000 2533.4800 3380.9000 2534.5600 ;
      RECT 0.0000 2533.4800 5.7000 2534.5600 ;
      RECT 0.0000 2531.8400 3390.2000 2533.4800 ;
      RECT 3388.5000 2530.7600 3390.2000 2531.8400 ;
      RECT 5.3000 2530.7600 3384.9000 2531.8400 ;
      RECT 0.0000 2530.7600 1.7000 2531.8400 ;
      RECT 0.0000 2529.1200 3390.2000 2530.7600 ;
      RECT 3384.5000 2528.0400 3390.2000 2529.1200 ;
      RECT 9.3000 2528.0400 3380.9000 2529.1200 ;
      RECT 0.0000 2528.0400 5.7000 2529.1200 ;
      RECT 0.0000 2526.4000 3390.2000 2528.0400 ;
      RECT 3388.5000 2525.3200 3390.2000 2526.4000 ;
      RECT 5.3000 2525.3200 3384.9000 2526.4000 ;
      RECT 0.0000 2525.3200 1.7000 2526.4000 ;
      RECT 0.0000 2523.6800 3390.2000 2525.3200 ;
      RECT 0.0000 2523.0700 5.7000 2523.6800 ;
      RECT 3384.5000 2522.6000 3390.2000 2523.6800 ;
      RECT 9.3000 2522.6000 3380.9000 2523.6800 ;
      RECT 1.1000 2522.6000 5.7000 2523.0700 ;
      RECT 1.1000 2522.1700 3390.2000 2522.6000 ;
      RECT 0.0000 2520.9600 3390.2000 2522.1700 ;
      RECT 3388.5000 2519.8800 3390.2000 2520.9600 ;
      RECT 5.3000 2519.8800 3384.9000 2520.9600 ;
      RECT 0.0000 2519.8800 1.7000 2520.9600 ;
      RECT 0.0000 2518.2400 3390.2000 2519.8800 ;
      RECT 3384.5000 2517.1600 3390.2000 2518.2400 ;
      RECT 9.3000 2517.1600 3380.9000 2518.2400 ;
      RECT 0.0000 2517.1600 5.7000 2518.2400 ;
      RECT 0.0000 2515.5200 3390.2000 2517.1600 ;
      RECT 3388.5000 2514.4400 3390.2000 2515.5200 ;
      RECT 5.3000 2514.4400 3384.9000 2515.5200 ;
      RECT 0.0000 2514.4400 1.7000 2515.5200 ;
      RECT 0.0000 2512.8000 3390.2000 2514.4400 ;
      RECT 3384.5000 2511.7200 3390.2000 2512.8000 ;
      RECT 9.3000 2511.7200 3380.9000 2512.8000 ;
      RECT 0.0000 2511.7200 5.7000 2512.8000 ;
      RECT 0.0000 2510.0800 3390.2000 2511.7200 ;
      RECT 3388.5000 2509.0000 3390.2000 2510.0800 ;
      RECT 5.3000 2509.0000 3384.9000 2510.0800 ;
      RECT 0.0000 2509.0000 1.7000 2510.0800 ;
      RECT 0.0000 2507.3600 3390.2000 2509.0000 ;
      RECT 3384.5000 2506.2800 3390.2000 2507.3600 ;
      RECT 9.3000 2506.2800 3380.9000 2507.3600 ;
      RECT 0.0000 2506.2800 5.7000 2507.3600 ;
      RECT 0.0000 2504.6400 3390.2000 2506.2800 ;
      RECT 3388.5000 2503.5600 3390.2000 2504.6400 ;
      RECT 5.3000 2503.5600 3384.9000 2504.6400 ;
      RECT 0.0000 2503.5600 1.7000 2504.6400 ;
      RECT 0.0000 2501.9200 3390.2000 2503.5600 ;
      RECT 3384.5000 2500.8400 3390.2000 2501.9200 ;
      RECT 9.3000 2500.8400 3380.9000 2501.9200 ;
      RECT 0.0000 2500.8400 5.7000 2501.9200 ;
      RECT 0.0000 2499.2000 3390.2000 2500.8400 ;
      RECT 3388.5000 2498.1200 3390.2000 2499.2000 ;
      RECT 5.3000 2498.1200 3384.9000 2499.2000 ;
      RECT 0.0000 2498.1200 1.7000 2499.2000 ;
      RECT 0.0000 2497.4500 3390.2000 2498.1200 ;
      RECT 1.1000 2496.5500 3390.2000 2497.4500 ;
      RECT 0.0000 2496.4800 3390.2000 2496.5500 ;
      RECT 3384.5000 2495.4000 3390.2000 2496.4800 ;
      RECT 9.3000 2495.4000 3380.9000 2496.4800 ;
      RECT 0.0000 2495.4000 5.7000 2496.4800 ;
      RECT 0.0000 2493.7600 3390.2000 2495.4000 ;
      RECT 3388.5000 2492.6800 3390.2000 2493.7600 ;
      RECT 5.3000 2492.6800 3384.9000 2493.7600 ;
      RECT 0.0000 2492.6800 1.7000 2493.7600 ;
      RECT 0.0000 2491.0400 3390.2000 2492.6800 ;
      RECT 3384.5000 2489.9600 3390.2000 2491.0400 ;
      RECT 9.3000 2489.9600 3380.9000 2491.0400 ;
      RECT 0.0000 2489.9600 5.7000 2491.0400 ;
      RECT 0.0000 2488.9100 3390.2000 2489.9600 ;
      RECT 0.0000 2488.3200 3389.1000 2488.9100 ;
      RECT 3388.5000 2488.0100 3389.1000 2488.3200 ;
      RECT 3388.5000 2487.2400 3390.2000 2488.0100 ;
      RECT 5.3000 2487.2400 3384.9000 2488.3200 ;
      RECT 0.0000 2487.2400 1.7000 2488.3200 ;
      RECT 0.0000 2485.6000 3390.2000 2487.2400 ;
      RECT 3384.5000 2484.5200 3390.2000 2485.6000 ;
      RECT 9.3000 2484.5200 3380.9000 2485.6000 ;
      RECT 0.0000 2484.5200 5.7000 2485.6000 ;
      RECT 0.0000 2482.8800 3390.2000 2484.5200 ;
      RECT 3388.5000 2481.8000 3390.2000 2482.8800 ;
      RECT 5.3000 2481.8000 3384.9000 2482.8800 ;
      RECT 0.0000 2481.8000 1.7000 2482.8800 ;
      RECT 0.0000 2480.1600 3390.2000 2481.8000 ;
      RECT 3384.5000 2479.0800 3390.2000 2480.1600 ;
      RECT 9.3000 2479.0800 3380.9000 2480.1600 ;
      RECT 0.0000 2479.0800 5.7000 2480.1600 ;
      RECT 0.0000 2477.4400 3390.2000 2479.0800 ;
      RECT 3388.5000 2476.3600 3390.2000 2477.4400 ;
      RECT 5.3000 2476.3600 3384.9000 2477.4400 ;
      RECT 0.0000 2476.3600 1.7000 2477.4400 ;
      RECT 0.0000 2474.7200 3390.2000 2476.3600 ;
      RECT 3384.5000 2473.6400 3390.2000 2474.7200 ;
      RECT 9.3000 2473.6400 3380.9000 2474.7200 ;
      RECT 0.0000 2473.6400 5.7000 2474.7200 ;
      RECT 0.0000 2472.4400 3390.2000 2473.6400 ;
      RECT 1.1000 2472.0000 3390.2000 2472.4400 ;
      RECT 1.1000 2471.5400 1.7000 2472.0000 ;
      RECT 3388.5000 2470.9200 3390.2000 2472.0000 ;
      RECT 5.3000 2470.9200 3384.9000 2472.0000 ;
      RECT 0.0000 2470.9200 1.7000 2471.5400 ;
      RECT 0.0000 2469.2800 3390.2000 2470.9200 ;
      RECT 3384.5000 2468.2000 3390.2000 2469.2800 ;
      RECT 9.3000 2468.2000 3380.9000 2469.2800 ;
      RECT 0.0000 2468.2000 5.7000 2469.2800 ;
      RECT 0.0000 2466.5600 3390.2000 2468.2000 ;
      RECT 3388.5000 2465.4800 3390.2000 2466.5600 ;
      RECT 5.3000 2465.4800 3384.9000 2466.5600 ;
      RECT 0.0000 2465.4800 1.7000 2466.5600 ;
      RECT 0.0000 2463.8400 3390.2000 2465.4800 ;
      RECT 3384.5000 2462.7600 3390.2000 2463.8400 ;
      RECT 9.3000 2462.7600 3380.9000 2463.8400 ;
      RECT 0.0000 2462.7600 5.7000 2463.8400 ;
      RECT 0.0000 2461.1200 3390.2000 2462.7600 ;
      RECT 3388.5000 2460.0400 3390.2000 2461.1200 ;
      RECT 5.3000 2460.0400 3384.9000 2461.1200 ;
      RECT 0.0000 2460.0400 1.7000 2461.1200 ;
      RECT 0.0000 2458.4000 3390.2000 2460.0400 ;
      RECT 3384.5000 2457.3200 3390.2000 2458.4000 ;
      RECT 9.3000 2457.3200 3380.9000 2458.4000 ;
      RECT 0.0000 2457.3200 5.7000 2458.4000 ;
      RECT 0.0000 2455.6800 3390.2000 2457.3200 ;
      RECT 3388.5000 2454.6000 3390.2000 2455.6800 ;
      RECT 5.3000 2454.6000 3384.9000 2455.6800 ;
      RECT 0.0000 2454.6000 1.7000 2455.6800 ;
      RECT 0.0000 2452.9600 3390.2000 2454.6000 ;
      RECT 3384.5000 2451.8800 3390.2000 2452.9600 ;
      RECT 9.3000 2451.8800 3380.9000 2452.9600 ;
      RECT 0.0000 2451.8800 5.7000 2452.9600 ;
      RECT 0.0000 2450.2400 3390.2000 2451.8800 ;
      RECT 3388.5000 2449.1600 3390.2000 2450.2400 ;
      RECT 5.3000 2449.1600 3384.9000 2450.2400 ;
      RECT 0.0000 2449.1600 1.7000 2450.2400 ;
      RECT 0.0000 2447.5200 3390.2000 2449.1600 ;
      RECT 0.0000 2447.4300 5.7000 2447.5200 ;
      RECT 1.1000 2446.5300 5.7000 2447.4300 ;
      RECT 3384.5000 2446.4400 3390.2000 2447.5200 ;
      RECT 9.3000 2446.4400 3380.9000 2447.5200 ;
      RECT 0.0000 2446.4400 5.7000 2446.5300 ;
      RECT 0.0000 2444.8000 3390.2000 2446.4400 ;
      RECT 3388.5000 2443.7200 3390.2000 2444.8000 ;
      RECT 5.3000 2443.7200 3384.9000 2444.8000 ;
      RECT 0.0000 2443.7200 1.7000 2444.8000 ;
      RECT 0.0000 2442.0800 3390.2000 2443.7200 ;
      RECT 3384.5000 2441.0000 3390.2000 2442.0800 ;
      RECT 9.3000 2441.0000 3380.9000 2442.0800 ;
      RECT 0.0000 2441.0000 5.7000 2442.0800 ;
      RECT 0.0000 2439.3600 3390.2000 2441.0000 ;
      RECT 3388.5000 2438.2800 3390.2000 2439.3600 ;
      RECT 5.3000 2438.2800 3384.9000 2439.3600 ;
      RECT 0.0000 2438.2800 1.7000 2439.3600 ;
      RECT 0.0000 2436.6400 3390.2000 2438.2800 ;
      RECT 3384.5000 2435.5600 3390.2000 2436.6400 ;
      RECT 9.3000 2435.5600 3380.9000 2436.6400 ;
      RECT 0.0000 2435.5600 5.7000 2436.6400 ;
      RECT 0.0000 2433.9200 3390.2000 2435.5600 ;
      RECT 3388.5000 2432.8400 3390.2000 2433.9200 ;
      RECT 5.3000 2432.8400 3384.9000 2433.9200 ;
      RECT 0.0000 2432.8400 1.7000 2433.9200 ;
      RECT 0.0000 2431.2000 3390.2000 2432.8400 ;
      RECT 3384.5000 2430.1200 3390.2000 2431.2000 ;
      RECT 9.3000 2430.1200 3380.9000 2431.2000 ;
      RECT 0.0000 2430.1200 5.7000 2431.2000 ;
      RECT 0.0000 2428.4800 3390.2000 2430.1200 ;
      RECT 3388.5000 2427.4000 3390.2000 2428.4800 ;
      RECT 5.3000 2427.4000 3384.9000 2428.4800 ;
      RECT 0.0000 2427.4000 1.7000 2428.4800 ;
      RECT 0.0000 2425.7600 3390.2000 2427.4000 ;
      RECT 3384.5000 2424.6800 3390.2000 2425.7600 ;
      RECT 9.3000 2424.6800 3380.9000 2425.7600 ;
      RECT 0.0000 2424.6800 5.7000 2425.7600 ;
      RECT 0.0000 2423.0400 3390.2000 2424.6800 ;
      RECT 3388.5000 2421.9600 3390.2000 2423.0400 ;
      RECT 5.3000 2421.9600 3384.9000 2423.0400 ;
      RECT 0.0000 2421.9600 1.7000 2423.0400 ;
      RECT 0.0000 2421.8100 3390.2000 2421.9600 ;
      RECT 1.1000 2420.9100 3390.2000 2421.8100 ;
      RECT 0.0000 2420.3200 3390.2000 2420.9100 ;
      RECT 3384.5000 2419.2400 3390.2000 2420.3200 ;
      RECT 9.3000 2419.2400 3380.9000 2420.3200 ;
      RECT 0.0000 2419.2400 5.7000 2420.3200 ;
      RECT 0.0000 2417.6000 3390.2000 2419.2400 ;
      RECT 3388.5000 2416.5200 3390.2000 2417.6000 ;
      RECT 5.3000 2416.5200 3384.9000 2417.6000 ;
      RECT 0.0000 2416.5200 1.7000 2417.6000 ;
      RECT 0.0000 2414.8800 3390.2000 2416.5200 ;
      RECT 3384.5000 2413.8000 3390.2000 2414.8800 ;
      RECT 9.3000 2413.8000 3380.9000 2414.8800 ;
      RECT 0.0000 2413.8000 5.7000 2414.8800 ;
      RECT 0.0000 2412.1600 3390.2000 2413.8000 ;
      RECT 3388.5000 2411.0800 3390.2000 2412.1600 ;
      RECT 5.3000 2411.0800 3384.9000 2412.1600 ;
      RECT 0.0000 2411.0800 1.7000 2412.1600 ;
      RECT 0.0000 2409.4400 3390.2000 2411.0800 ;
      RECT 3384.5000 2408.3600 3390.2000 2409.4400 ;
      RECT 9.3000 2408.3600 3380.9000 2409.4400 ;
      RECT 0.0000 2408.3600 5.7000 2409.4400 ;
      RECT 0.0000 2406.7200 3390.2000 2408.3600 ;
      RECT 3388.5000 2405.6400 3390.2000 2406.7200 ;
      RECT 5.3000 2405.6400 3384.9000 2406.7200 ;
      RECT 0.0000 2405.6400 1.7000 2406.7200 ;
      RECT 0.0000 2404.0000 3390.2000 2405.6400 ;
      RECT 3384.5000 2402.9200 3390.2000 2404.0000 ;
      RECT 9.3000 2402.9200 3380.9000 2404.0000 ;
      RECT 0.0000 2402.9200 5.7000 2404.0000 ;
      RECT 0.0000 2401.2800 3390.2000 2402.9200 ;
      RECT 3388.5000 2400.2000 3390.2000 2401.2800 ;
      RECT 5.3000 2400.2000 3384.9000 2401.2800 ;
      RECT 0.0000 2400.2000 1.7000 2401.2800 ;
      RECT 0.0000 2398.5600 3390.2000 2400.2000 ;
      RECT 3384.5000 2397.4800 3390.2000 2398.5600 ;
      RECT 9.3000 2397.4800 3380.9000 2398.5600 ;
      RECT 0.0000 2397.4800 5.7000 2398.5600 ;
      RECT 0.0000 2396.8000 3390.2000 2397.4800 ;
      RECT 1.1000 2395.9000 3390.2000 2396.8000 ;
      RECT 0.0000 2395.8400 3390.2000 2395.9000 ;
      RECT 3388.5000 2394.7600 3390.2000 2395.8400 ;
      RECT 5.3000 2394.7600 3384.9000 2395.8400 ;
      RECT 0.0000 2394.7600 1.7000 2395.8400 ;
      RECT 0.0000 2393.1200 3390.2000 2394.7600 ;
      RECT 3384.5000 2392.0400 3390.2000 2393.1200 ;
      RECT 9.3000 2392.0400 3380.9000 2393.1200 ;
      RECT 0.0000 2392.0400 5.7000 2393.1200 ;
      RECT 0.0000 2390.4000 3390.2000 2392.0400 ;
      RECT 3388.5000 2389.3200 3390.2000 2390.4000 ;
      RECT 5.3000 2389.3200 3384.9000 2390.4000 ;
      RECT 0.0000 2389.3200 1.7000 2390.4000 ;
      RECT 0.0000 2387.6800 3390.2000 2389.3200 ;
      RECT 3384.5000 2386.6000 3390.2000 2387.6800 ;
      RECT 9.3000 2386.6000 3380.9000 2387.6800 ;
      RECT 0.0000 2386.6000 5.7000 2387.6800 ;
      RECT 0.0000 2385.2100 3390.2000 2386.6000 ;
      RECT 0.0000 2384.9600 3389.1000 2385.2100 ;
      RECT 3388.5000 2384.3100 3389.1000 2384.9600 ;
      RECT 3388.5000 2383.8800 3390.2000 2384.3100 ;
      RECT 5.3000 2383.8800 3384.9000 2384.9600 ;
      RECT 0.0000 2383.8800 1.7000 2384.9600 ;
      RECT 0.0000 2382.2400 3390.2000 2383.8800 ;
      RECT 3384.5000 2381.1600 3390.2000 2382.2400 ;
      RECT 9.3000 2381.1600 3380.9000 2382.2400 ;
      RECT 0.0000 2381.1600 5.7000 2382.2400 ;
      RECT 0.0000 2379.5200 3390.2000 2381.1600 ;
      RECT 3388.5000 2378.4400 3390.2000 2379.5200 ;
      RECT 5.3000 2378.4400 3384.9000 2379.5200 ;
      RECT 0.0000 2378.4400 1.7000 2379.5200 ;
      RECT 0.0000 2376.8000 3390.2000 2378.4400 ;
      RECT 3384.5000 2375.7200 3390.2000 2376.8000 ;
      RECT 9.3000 2375.7200 3380.9000 2376.8000 ;
      RECT 0.0000 2375.7200 5.7000 2376.8000 ;
      RECT 0.0000 2374.0800 3390.2000 2375.7200 ;
      RECT 3388.5000 2373.0000 3390.2000 2374.0800 ;
      RECT 5.3000 2373.0000 3384.9000 2374.0800 ;
      RECT 0.0000 2373.0000 1.7000 2374.0800 ;
      RECT 0.0000 2371.3600 3390.2000 2373.0000 ;
      RECT 0.0000 2371.1800 5.7000 2371.3600 ;
      RECT 3384.5000 2370.2800 3390.2000 2371.3600 ;
      RECT 9.3000 2370.2800 3380.9000 2371.3600 ;
      RECT 1.1000 2370.2800 5.7000 2371.1800 ;
      RECT 0.0000 2368.6400 3390.2000 2370.2800 ;
      RECT 3388.5000 2367.5600 3390.2000 2368.6400 ;
      RECT 5.3000 2367.5600 3384.9000 2368.6400 ;
      RECT 0.0000 2367.5600 1.7000 2368.6400 ;
      RECT 0.0000 2365.9200 3390.2000 2367.5600 ;
      RECT 3384.5000 2364.8400 3390.2000 2365.9200 ;
      RECT 9.3000 2364.8400 3380.9000 2365.9200 ;
      RECT 0.0000 2364.8400 5.7000 2365.9200 ;
      RECT 0.0000 2363.2000 3390.2000 2364.8400 ;
      RECT 3388.5000 2362.1200 3390.2000 2363.2000 ;
      RECT 5.3000 2362.1200 3384.9000 2363.2000 ;
      RECT 0.0000 2362.1200 1.7000 2363.2000 ;
      RECT 0.0000 2360.4800 3390.2000 2362.1200 ;
      RECT 3384.5000 2359.4000 3390.2000 2360.4800 ;
      RECT 9.3000 2359.4000 3380.9000 2360.4800 ;
      RECT 0.0000 2359.4000 5.7000 2360.4800 ;
      RECT 0.0000 2357.7600 3390.2000 2359.4000 ;
      RECT 3388.5000 2356.6800 3390.2000 2357.7600 ;
      RECT 5.3000 2356.6800 3384.9000 2357.7600 ;
      RECT 0.0000 2356.6800 1.7000 2357.7600 ;
      RECT 0.0000 2355.0400 3390.2000 2356.6800 ;
      RECT 3384.5000 2353.9600 3390.2000 2355.0400 ;
      RECT 9.3000 2353.9600 3380.9000 2355.0400 ;
      RECT 0.0000 2353.9600 5.7000 2355.0400 ;
      RECT 0.0000 2352.3200 3390.2000 2353.9600 ;
      RECT 3388.5000 2351.2400 3390.2000 2352.3200 ;
      RECT 5.3000 2351.2400 3384.9000 2352.3200 ;
      RECT 0.0000 2351.2400 1.7000 2352.3200 ;
      RECT 0.0000 2349.6000 3390.2000 2351.2400 ;
      RECT 3384.5000 2348.5200 3390.2000 2349.6000 ;
      RECT 9.3000 2348.5200 3380.9000 2349.6000 ;
      RECT 0.0000 2348.5200 5.7000 2349.6000 ;
      RECT 0.0000 2346.8800 3390.2000 2348.5200 ;
      RECT 0.0000 2346.1700 1.7000 2346.8800 ;
      RECT 3388.5000 2345.8000 3390.2000 2346.8800 ;
      RECT 5.3000 2345.8000 3384.9000 2346.8800 ;
      RECT 1.1000 2345.8000 1.7000 2346.1700 ;
      RECT 1.1000 2345.2700 3390.2000 2345.8000 ;
      RECT 0.0000 2344.1600 3390.2000 2345.2700 ;
      RECT 3384.5000 2343.0800 3390.2000 2344.1600 ;
      RECT 9.3000 2343.0800 3380.9000 2344.1600 ;
      RECT 0.0000 2343.0800 5.7000 2344.1600 ;
      RECT 0.0000 2341.4400 3390.2000 2343.0800 ;
      RECT 3388.5000 2340.3600 3390.2000 2341.4400 ;
      RECT 5.3000 2340.3600 3384.9000 2341.4400 ;
      RECT 0.0000 2340.3600 1.7000 2341.4400 ;
      RECT 0.0000 2338.7200 3390.2000 2340.3600 ;
      RECT 3384.5000 2337.6400 3390.2000 2338.7200 ;
      RECT 9.3000 2337.6400 3380.9000 2338.7200 ;
      RECT 0.0000 2337.6400 5.7000 2338.7200 ;
      RECT 0.0000 2336.0000 3390.2000 2337.6400 ;
      RECT 3388.5000 2334.9200 3390.2000 2336.0000 ;
      RECT 5.3000 2334.9200 3384.9000 2336.0000 ;
      RECT 0.0000 2334.9200 1.7000 2336.0000 ;
      RECT 0.0000 2333.2800 3390.2000 2334.9200 ;
      RECT 3384.5000 2332.2000 3390.2000 2333.2800 ;
      RECT 9.3000 2332.2000 3380.9000 2333.2800 ;
      RECT 0.0000 2332.2000 5.7000 2333.2800 ;
      RECT 0.0000 2330.5600 3390.2000 2332.2000 ;
      RECT 3388.5000 2329.4800 3390.2000 2330.5600 ;
      RECT 5.3000 2329.4800 3384.9000 2330.5600 ;
      RECT 0.0000 2329.4800 1.7000 2330.5600 ;
      RECT 0.0000 2327.8400 3390.2000 2329.4800 ;
      RECT 3384.5000 2326.7600 3390.2000 2327.8400 ;
      RECT 9.3000 2326.7600 3380.9000 2327.8400 ;
      RECT 0.0000 2326.7600 5.7000 2327.8400 ;
      RECT 0.0000 2325.1200 3390.2000 2326.7600 ;
      RECT 3388.5000 2324.0400 3390.2000 2325.1200 ;
      RECT 5.3000 2324.0400 3384.9000 2325.1200 ;
      RECT 0.0000 2324.0400 1.7000 2325.1200 ;
      RECT 0.0000 2322.4000 3390.2000 2324.0400 ;
      RECT 3384.5000 2321.3200 3390.2000 2322.4000 ;
      RECT 9.3000 2321.3200 3380.9000 2322.4000 ;
      RECT 0.0000 2321.3200 5.7000 2322.4000 ;
      RECT 0.0000 2321.1600 3390.2000 2321.3200 ;
      RECT 1.1000 2320.2600 3390.2000 2321.1600 ;
      RECT 0.0000 2319.6800 3390.2000 2320.2600 ;
      RECT 3388.5000 2318.6000 3390.2000 2319.6800 ;
      RECT 5.3000 2318.6000 3384.9000 2319.6800 ;
      RECT 0.0000 2318.6000 1.7000 2319.6800 ;
      RECT 0.0000 2316.9600 3390.2000 2318.6000 ;
      RECT 3384.5000 2315.8800 3390.2000 2316.9600 ;
      RECT 9.3000 2315.8800 3380.9000 2316.9600 ;
      RECT 0.0000 2315.8800 5.7000 2316.9600 ;
      RECT 0.0000 2314.2400 3390.2000 2315.8800 ;
      RECT 3388.5000 2313.1600 3390.2000 2314.2400 ;
      RECT 5.3000 2313.1600 3384.9000 2314.2400 ;
      RECT 0.0000 2313.1600 1.7000 2314.2400 ;
      RECT 0.0000 2311.5200 3390.2000 2313.1600 ;
      RECT 3384.5000 2310.4400 3390.2000 2311.5200 ;
      RECT 9.3000 2310.4400 3380.9000 2311.5200 ;
      RECT 0.0000 2310.4400 5.7000 2311.5200 ;
      RECT 0.0000 2308.8000 3390.2000 2310.4400 ;
      RECT 3388.5000 2307.7200 3390.2000 2308.8000 ;
      RECT 5.3000 2307.7200 3384.9000 2308.8000 ;
      RECT 0.0000 2307.7200 1.7000 2308.8000 ;
      RECT 0.0000 2306.0800 3390.2000 2307.7200 ;
      RECT 3384.5000 2305.0000 3390.2000 2306.0800 ;
      RECT 9.3000 2305.0000 3380.9000 2306.0800 ;
      RECT 0.0000 2305.0000 5.7000 2306.0800 ;
      RECT 0.0000 2303.3600 3390.2000 2305.0000 ;
      RECT 3388.5000 2302.2800 3390.2000 2303.3600 ;
      RECT 5.3000 2302.2800 3384.9000 2303.3600 ;
      RECT 0.0000 2302.2800 1.7000 2303.3600 ;
      RECT 0.0000 2300.6400 3390.2000 2302.2800 ;
      RECT 3384.5000 2299.5600 3390.2000 2300.6400 ;
      RECT 9.3000 2299.5600 3380.9000 2300.6400 ;
      RECT 0.0000 2299.5600 5.7000 2300.6400 ;
      RECT 0.0000 2297.9200 3390.2000 2299.5600 ;
      RECT 3388.5000 2296.8400 3390.2000 2297.9200 ;
      RECT 5.3000 2296.8400 3384.9000 2297.9200 ;
      RECT 0.0000 2296.8400 1.7000 2297.9200 ;
      RECT 0.0000 2295.5400 3390.2000 2296.8400 ;
      RECT 1.1000 2295.2000 3390.2000 2295.5400 ;
      RECT 1.1000 2294.6400 5.7000 2295.2000 ;
      RECT 3384.5000 2294.1200 3390.2000 2295.2000 ;
      RECT 9.3000 2294.1200 3380.9000 2295.2000 ;
      RECT 0.0000 2294.1200 5.7000 2294.6400 ;
      RECT 0.0000 2292.4800 3390.2000 2294.1200 ;
      RECT 3388.5000 2291.4000 3390.2000 2292.4800 ;
      RECT 5.3000 2291.4000 3384.9000 2292.4800 ;
      RECT 0.0000 2291.4000 1.7000 2292.4800 ;
      RECT 0.0000 2289.7600 3390.2000 2291.4000 ;
      RECT 3384.5000 2288.6800 3390.2000 2289.7600 ;
      RECT 9.3000 2288.6800 3380.9000 2289.7600 ;
      RECT 0.0000 2288.6800 5.7000 2289.7600 ;
      RECT 0.0000 2287.0400 3390.2000 2288.6800 ;
      RECT 3388.5000 2285.9600 3390.2000 2287.0400 ;
      RECT 5.3000 2285.9600 3384.9000 2287.0400 ;
      RECT 0.0000 2285.9600 1.7000 2287.0400 ;
      RECT 0.0000 2284.3200 3390.2000 2285.9600 ;
      RECT 3384.5000 2283.2400 3390.2000 2284.3200 ;
      RECT 9.3000 2283.2400 3380.9000 2284.3200 ;
      RECT 0.0000 2283.2400 5.7000 2284.3200 ;
      RECT 0.0000 2281.6000 3390.2000 2283.2400 ;
      RECT 3388.5000 2281.5100 3390.2000 2281.6000 ;
      RECT 3388.5000 2280.6100 3389.1000 2281.5100 ;
      RECT 3388.5000 2280.5200 3390.2000 2280.6100 ;
      RECT 5.3000 2280.5200 3384.9000 2281.6000 ;
      RECT 0.0000 2280.5200 1.7000 2281.6000 ;
      RECT 0.0000 2278.8800 3390.2000 2280.5200 ;
      RECT 3384.5000 2277.8000 3390.2000 2278.8800 ;
      RECT 9.3000 2277.8000 3380.9000 2278.8800 ;
      RECT 0.0000 2277.8000 5.7000 2278.8800 ;
      RECT 0.0000 2276.1600 3390.2000 2277.8000 ;
      RECT 3388.5000 2275.0800 3390.2000 2276.1600 ;
      RECT 5.3000 2275.0800 3384.9000 2276.1600 ;
      RECT 0.0000 2275.0800 1.7000 2276.1600 ;
      RECT 0.0000 2273.4400 3390.2000 2275.0800 ;
      RECT 3384.5000 2272.3600 3390.2000 2273.4400 ;
      RECT 9.3000 2272.3600 3380.9000 2273.4400 ;
      RECT 0.0000 2272.3600 5.7000 2273.4400 ;
      RECT 0.0000 2270.7200 3390.2000 2272.3600 ;
      RECT 0.0000 2270.5300 1.7000 2270.7200 ;
      RECT 3388.5000 2269.6400 3390.2000 2270.7200 ;
      RECT 5.3000 2269.6400 3384.9000 2270.7200 ;
      RECT 1.1000 2269.6400 1.7000 2270.5300 ;
      RECT 1.1000 2269.6300 3390.2000 2269.6400 ;
      RECT 0.0000 2268.0000 3390.2000 2269.6300 ;
      RECT 3384.5000 2266.9200 3390.2000 2268.0000 ;
      RECT 9.3000 2266.9200 3380.9000 2268.0000 ;
      RECT 0.0000 2266.9200 5.7000 2268.0000 ;
      RECT 0.0000 2265.2800 3390.2000 2266.9200 ;
      RECT 3388.5000 2264.2000 3390.2000 2265.2800 ;
      RECT 5.3000 2264.2000 3384.9000 2265.2800 ;
      RECT 0.0000 2264.2000 1.7000 2265.2800 ;
      RECT 0.0000 2262.5600 3390.2000 2264.2000 ;
      RECT 3384.5000 2261.4800 3390.2000 2262.5600 ;
      RECT 9.3000 2261.4800 3380.9000 2262.5600 ;
      RECT 0.0000 2261.4800 5.7000 2262.5600 ;
      RECT 0.0000 2259.8400 3390.2000 2261.4800 ;
      RECT 3388.5000 2258.7600 3390.2000 2259.8400 ;
      RECT 5.3000 2258.7600 3384.9000 2259.8400 ;
      RECT 0.0000 2258.7600 1.7000 2259.8400 ;
      RECT 0.0000 2257.1200 3390.2000 2258.7600 ;
      RECT 3384.5000 2256.0400 3390.2000 2257.1200 ;
      RECT 9.3000 2256.0400 3380.9000 2257.1200 ;
      RECT 0.0000 2256.0400 5.7000 2257.1200 ;
      RECT 0.0000 2254.4000 3390.2000 2256.0400 ;
      RECT 3388.5000 2253.3200 3390.2000 2254.4000 ;
      RECT 5.3000 2253.3200 3384.9000 2254.4000 ;
      RECT 0.0000 2253.3200 1.7000 2254.4000 ;
      RECT 0.0000 2251.6800 3390.2000 2253.3200 ;
      RECT 3384.5000 2250.6000 3390.2000 2251.6800 ;
      RECT 9.3000 2250.6000 3380.9000 2251.6800 ;
      RECT 0.0000 2250.6000 5.7000 2251.6800 ;
      RECT 0.0000 2248.9600 3390.2000 2250.6000 ;
      RECT 3388.5000 2247.8800 3390.2000 2248.9600 ;
      RECT 5.3000 2247.8800 3384.9000 2248.9600 ;
      RECT 0.0000 2247.8800 1.7000 2248.9600 ;
      RECT 0.0000 2246.2400 3390.2000 2247.8800 ;
      RECT 0.0000 2245.5200 5.7000 2246.2400 ;
      RECT 3384.5000 2245.1600 3390.2000 2246.2400 ;
      RECT 9.3000 2245.1600 3380.9000 2246.2400 ;
      RECT 1.1000 2245.1600 5.7000 2245.5200 ;
      RECT 1.1000 2244.6200 3390.2000 2245.1600 ;
      RECT 0.0000 2243.5200 3390.2000 2244.6200 ;
      RECT 3388.5000 2242.4400 3390.2000 2243.5200 ;
      RECT 5.3000 2242.4400 3384.9000 2243.5200 ;
      RECT 0.0000 2242.4400 1.7000 2243.5200 ;
      RECT 0.0000 2240.8000 3390.2000 2242.4400 ;
      RECT 3384.5000 2239.7200 3390.2000 2240.8000 ;
      RECT 9.3000 2239.7200 3380.9000 2240.8000 ;
      RECT 0.0000 2239.7200 5.7000 2240.8000 ;
      RECT 0.0000 2238.0800 3390.2000 2239.7200 ;
      RECT 3388.5000 2237.0000 3390.2000 2238.0800 ;
      RECT 5.3000 2237.0000 3384.9000 2238.0800 ;
      RECT 0.0000 2237.0000 1.7000 2238.0800 ;
      RECT 0.0000 2235.3600 3390.2000 2237.0000 ;
      RECT 3384.5000 2234.2800 3390.2000 2235.3600 ;
      RECT 9.3000 2234.2800 3380.9000 2235.3600 ;
      RECT 0.0000 2234.2800 5.7000 2235.3600 ;
      RECT 0.0000 2232.6400 3390.2000 2234.2800 ;
      RECT 3388.5000 2231.5600 3390.2000 2232.6400 ;
      RECT 5.3000 2231.5600 3384.9000 2232.6400 ;
      RECT 0.0000 2231.5600 1.7000 2232.6400 ;
      RECT 0.0000 2229.9200 3390.2000 2231.5600 ;
      RECT 3384.5000 2228.8400 3390.2000 2229.9200 ;
      RECT 9.3000 2228.8400 3380.9000 2229.9200 ;
      RECT 0.0000 2228.8400 5.7000 2229.9200 ;
      RECT 0.0000 2227.2000 3390.2000 2228.8400 ;
      RECT 3388.5000 2226.1200 3390.2000 2227.2000 ;
      RECT 5.3000 2226.1200 3384.9000 2227.2000 ;
      RECT 0.0000 2226.1200 1.7000 2227.2000 ;
      RECT 0.0000 2224.4800 3390.2000 2226.1200 ;
      RECT 3384.5000 2223.4000 3390.2000 2224.4800 ;
      RECT 9.3000 2223.4000 3380.9000 2224.4800 ;
      RECT 0.0000 2223.4000 5.7000 2224.4800 ;
      RECT 0.0000 2221.7600 3390.2000 2223.4000 ;
      RECT 3388.5000 2220.6800 3390.2000 2221.7600 ;
      RECT 5.3000 2220.6800 3384.9000 2221.7600 ;
      RECT 0.0000 2220.6800 1.7000 2221.7600 ;
      RECT 0.0000 2219.9000 3390.2000 2220.6800 ;
      RECT 1.1000 2219.0400 3390.2000 2219.9000 ;
      RECT 1.1000 2219.0000 5.7000 2219.0400 ;
      RECT 3384.5000 2217.9600 3390.2000 2219.0400 ;
      RECT 9.3000 2217.9600 3380.9000 2219.0400 ;
      RECT 0.0000 2217.9600 5.7000 2219.0000 ;
      RECT 0.0000 2216.3200 3390.2000 2217.9600 ;
      RECT 3388.5000 2215.2400 3390.2000 2216.3200 ;
      RECT 5.3000 2215.2400 3384.9000 2216.3200 ;
      RECT 0.0000 2215.2400 1.7000 2216.3200 ;
      RECT 0.0000 2213.6000 3390.2000 2215.2400 ;
      RECT 3384.5000 2212.5200 3390.2000 2213.6000 ;
      RECT 9.3000 2212.5200 3380.9000 2213.6000 ;
      RECT 0.0000 2212.5200 5.7000 2213.6000 ;
      RECT 0.0000 2210.8800 3390.2000 2212.5200 ;
      RECT 3388.5000 2209.8000 3390.2000 2210.8800 ;
      RECT 5.3000 2209.8000 3384.9000 2210.8800 ;
      RECT 0.0000 2209.8000 1.7000 2210.8800 ;
      RECT 0.0000 2208.1600 3390.2000 2209.8000 ;
      RECT 3384.5000 2207.0800 3390.2000 2208.1600 ;
      RECT 9.3000 2207.0800 3380.9000 2208.1600 ;
      RECT 0.0000 2207.0800 5.7000 2208.1600 ;
      RECT 0.0000 2205.4400 3390.2000 2207.0800 ;
      RECT 3388.5000 2204.3600 3390.2000 2205.4400 ;
      RECT 5.3000 2204.3600 3384.9000 2205.4400 ;
      RECT 0.0000 2204.3600 1.7000 2205.4400 ;
      RECT 0.0000 2202.7200 3390.2000 2204.3600 ;
      RECT 3384.5000 2201.6400 3390.2000 2202.7200 ;
      RECT 9.3000 2201.6400 3380.9000 2202.7200 ;
      RECT 0.0000 2201.6400 5.7000 2202.7200 ;
      RECT 0.0000 2200.0000 3390.2000 2201.6400 ;
      RECT 3388.5000 2198.9200 3390.2000 2200.0000 ;
      RECT 5.3000 2198.9200 3384.9000 2200.0000 ;
      RECT 0.0000 2198.9200 1.7000 2200.0000 ;
      RECT 0.0000 2197.2800 3390.2000 2198.9200 ;
      RECT 3384.5000 2196.2000 3390.2000 2197.2800 ;
      RECT 9.3000 2196.2000 3380.9000 2197.2800 ;
      RECT 0.0000 2196.2000 5.7000 2197.2800 ;
      RECT 0.0000 2194.8900 3390.2000 2196.2000 ;
      RECT 1.1000 2194.5600 3390.2000 2194.8900 ;
      RECT 1.1000 2193.9900 1.7000 2194.5600 ;
      RECT 3388.5000 2193.4800 3390.2000 2194.5600 ;
      RECT 5.3000 2193.4800 3384.9000 2194.5600 ;
      RECT 0.0000 2193.4800 1.7000 2193.9900 ;
      RECT 0.0000 2191.8400 3390.2000 2193.4800 ;
      RECT 3384.5000 2190.7600 3390.2000 2191.8400 ;
      RECT 9.3000 2190.7600 3380.9000 2191.8400 ;
      RECT 0.0000 2190.7600 5.7000 2191.8400 ;
      RECT 0.0000 2189.1200 3390.2000 2190.7600 ;
      RECT 3388.5000 2188.0400 3390.2000 2189.1200 ;
      RECT 5.3000 2188.0400 3384.9000 2189.1200 ;
      RECT 0.0000 2188.0400 1.7000 2189.1200 ;
      RECT 0.0000 2186.4000 3390.2000 2188.0400 ;
      RECT 3384.5000 2185.3200 3390.2000 2186.4000 ;
      RECT 9.3000 2185.3200 3380.9000 2186.4000 ;
      RECT 0.0000 2185.3200 5.7000 2186.4000 ;
      RECT 0.0000 2183.6800 3390.2000 2185.3200 ;
      RECT 3388.5000 2182.6000 3390.2000 2183.6800 ;
      RECT 5.3000 2182.6000 3384.9000 2183.6800 ;
      RECT 0.0000 2182.6000 1.7000 2183.6800 ;
      RECT 0.0000 2180.9600 3390.2000 2182.6000 ;
      RECT 3384.5000 2179.8800 3390.2000 2180.9600 ;
      RECT 9.3000 2179.8800 3380.9000 2180.9600 ;
      RECT 0.0000 2179.8800 5.7000 2180.9600 ;
      RECT 0.0000 2178.2400 3390.2000 2179.8800 ;
      RECT 3388.5000 2177.2000 3390.2000 2178.2400 ;
      RECT 3388.5000 2177.1600 3389.1000 2177.2000 ;
      RECT 5.3000 2177.1600 3384.9000 2178.2400 ;
      RECT 0.0000 2177.1600 1.7000 2178.2400 ;
      RECT 0.0000 2176.3000 3389.1000 2177.1600 ;
      RECT 0.0000 2175.5200 3390.2000 2176.3000 ;
      RECT 3384.5000 2174.4400 3390.2000 2175.5200 ;
      RECT 9.3000 2174.4400 3380.9000 2175.5200 ;
      RECT 0.0000 2174.4400 5.7000 2175.5200 ;
      RECT 0.0000 2172.8000 3390.2000 2174.4400 ;
      RECT 3388.5000 2171.7200 3390.2000 2172.8000 ;
      RECT 5.3000 2171.7200 3384.9000 2172.8000 ;
      RECT 0.0000 2171.7200 1.7000 2172.8000 ;
      RECT 0.0000 2170.0800 3390.2000 2171.7200 ;
      RECT 0.0000 2169.8800 5.7000 2170.0800 ;
      RECT 3384.5000 2169.0000 3390.2000 2170.0800 ;
      RECT 9.3000 2169.0000 3380.9000 2170.0800 ;
      RECT 1.1000 2169.0000 5.7000 2169.8800 ;
      RECT 1.1000 2168.9800 3390.2000 2169.0000 ;
      RECT 0.0000 2167.3600 3390.2000 2168.9800 ;
      RECT 3388.5000 2166.2800 3390.2000 2167.3600 ;
      RECT 5.3000 2166.2800 3384.9000 2167.3600 ;
      RECT 0.0000 2166.2800 1.7000 2167.3600 ;
      RECT 0.0000 2164.6400 3390.2000 2166.2800 ;
      RECT 3384.5000 2163.5600 3390.2000 2164.6400 ;
      RECT 9.3000 2163.5600 3380.9000 2164.6400 ;
      RECT 0.0000 2163.5600 5.7000 2164.6400 ;
      RECT 0.0000 2161.9200 3390.2000 2163.5600 ;
      RECT 3388.5000 2160.8400 3390.2000 2161.9200 ;
      RECT 5.3000 2160.8400 3384.9000 2161.9200 ;
      RECT 0.0000 2160.8400 1.7000 2161.9200 ;
      RECT 0.0000 2159.2000 3390.2000 2160.8400 ;
      RECT 3384.5000 2158.1200 3390.2000 2159.2000 ;
      RECT 9.3000 2158.1200 3380.9000 2159.2000 ;
      RECT 0.0000 2158.1200 5.7000 2159.2000 ;
      RECT 0.0000 2156.4800 3390.2000 2158.1200 ;
      RECT 3388.5000 2155.4000 3390.2000 2156.4800 ;
      RECT 5.3000 2155.4000 3384.9000 2156.4800 ;
      RECT 0.0000 2155.4000 1.7000 2156.4800 ;
      RECT 0.0000 2153.7600 3390.2000 2155.4000 ;
      RECT 3384.5000 2152.6800 3390.2000 2153.7600 ;
      RECT 9.3000 2152.6800 3380.9000 2153.7600 ;
      RECT 0.0000 2152.6800 5.7000 2153.7600 ;
      RECT 0.0000 2151.0400 3390.2000 2152.6800 ;
      RECT 3388.5000 2149.9600 3390.2000 2151.0400 ;
      RECT 5.3000 2149.9600 3384.9000 2151.0400 ;
      RECT 0.0000 2149.9600 1.7000 2151.0400 ;
      RECT 0.0000 2148.3200 3390.2000 2149.9600 ;
      RECT 3384.5000 2147.2400 3390.2000 2148.3200 ;
      RECT 9.3000 2147.2400 3380.9000 2148.3200 ;
      RECT 0.0000 2147.2400 5.7000 2148.3200 ;
      RECT 0.0000 2145.6000 3390.2000 2147.2400 ;
      RECT 3388.5000 2144.5200 3390.2000 2145.6000 ;
      RECT 5.3000 2144.5200 3384.9000 2145.6000 ;
      RECT 0.0000 2144.5200 1.7000 2145.6000 ;
      RECT 0.0000 2144.2600 3390.2000 2144.5200 ;
      RECT 1.1000 2143.3600 3390.2000 2144.2600 ;
      RECT 0.0000 2142.8800 3390.2000 2143.3600 ;
      RECT 3384.5000 2141.8000 3390.2000 2142.8800 ;
      RECT 9.3000 2141.8000 3380.9000 2142.8800 ;
      RECT 0.0000 2141.8000 5.7000 2142.8800 ;
      RECT 0.0000 2140.1600 3390.2000 2141.8000 ;
      RECT 3388.5000 2139.0800 3390.2000 2140.1600 ;
      RECT 5.3000 2139.0800 3384.9000 2140.1600 ;
      RECT 0.0000 2139.0800 1.7000 2140.1600 ;
      RECT 0.0000 2137.4400 3390.2000 2139.0800 ;
      RECT 3384.5000 2136.3600 3390.2000 2137.4400 ;
      RECT 9.3000 2136.3600 3380.9000 2137.4400 ;
      RECT 0.0000 2136.3600 5.7000 2137.4400 ;
      RECT 0.0000 2134.7200 3390.2000 2136.3600 ;
      RECT 3388.5000 2133.6400 3390.2000 2134.7200 ;
      RECT 5.3000 2133.6400 3384.9000 2134.7200 ;
      RECT 0.0000 2133.6400 1.7000 2134.7200 ;
      RECT 0.0000 2132.0000 3390.2000 2133.6400 ;
      RECT 3384.5000 2130.9200 3390.2000 2132.0000 ;
      RECT 9.3000 2130.9200 3380.9000 2132.0000 ;
      RECT 0.0000 2130.9200 5.7000 2132.0000 ;
      RECT 0.0000 2129.2800 3390.2000 2130.9200 ;
      RECT 3388.5000 2128.2000 3390.2000 2129.2800 ;
      RECT 5.3000 2128.2000 3384.9000 2129.2800 ;
      RECT 0.0000 2128.2000 1.7000 2129.2800 ;
      RECT 0.0000 2126.5600 3390.2000 2128.2000 ;
      RECT 3384.5000 2125.4800 3390.2000 2126.5600 ;
      RECT 9.3000 2125.4800 3380.9000 2126.5600 ;
      RECT 0.0000 2125.4800 5.7000 2126.5600 ;
      RECT 0.0000 2123.8400 3390.2000 2125.4800 ;
      RECT 3388.5000 2122.7600 3390.2000 2123.8400 ;
      RECT 5.3000 2122.7600 3384.9000 2123.8400 ;
      RECT 0.0000 2122.7600 1.7000 2123.8400 ;
      RECT 0.0000 2121.1200 3390.2000 2122.7600 ;
      RECT 3384.5000 2120.0400 3390.2000 2121.1200 ;
      RECT 9.3000 2120.0400 3380.9000 2121.1200 ;
      RECT 0.0000 2120.0400 5.7000 2121.1200 ;
      RECT 0.0000 2119.2500 3390.2000 2120.0400 ;
      RECT 1.1000 2118.4000 3390.2000 2119.2500 ;
      RECT 1.1000 2118.3500 1.7000 2118.4000 ;
      RECT 3388.5000 2117.3200 3390.2000 2118.4000 ;
      RECT 5.3000 2117.3200 3384.9000 2118.4000 ;
      RECT 0.0000 2117.3200 1.7000 2118.3500 ;
      RECT 0.0000 2115.6800 3390.2000 2117.3200 ;
      RECT 3384.5000 2114.6000 3390.2000 2115.6800 ;
      RECT 9.3000 2114.6000 3380.9000 2115.6800 ;
      RECT 0.0000 2114.6000 5.7000 2115.6800 ;
      RECT 0.0000 2112.9600 3390.2000 2114.6000 ;
      RECT 3388.5000 2111.8800 3390.2000 2112.9600 ;
      RECT 5.3000 2111.8800 3384.9000 2112.9600 ;
      RECT 0.0000 2111.8800 1.7000 2112.9600 ;
      RECT 0.0000 2110.2400 3390.2000 2111.8800 ;
      RECT 3384.5000 2109.1600 3390.2000 2110.2400 ;
      RECT 9.3000 2109.1600 3380.9000 2110.2400 ;
      RECT 0.0000 2109.1600 5.7000 2110.2400 ;
      RECT 0.0000 2107.5200 3390.2000 2109.1600 ;
      RECT 3388.5000 2106.4400 3390.2000 2107.5200 ;
      RECT 5.3000 2106.4400 3384.9000 2107.5200 ;
      RECT 0.0000 2106.4400 1.7000 2107.5200 ;
      RECT 0.0000 2104.8000 3390.2000 2106.4400 ;
      RECT 3384.5000 2103.7200 3390.2000 2104.8000 ;
      RECT 9.3000 2103.7200 3380.9000 2104.8000 ;
      RECT 0.0000 2103.7200 5.7000 2104.8000 ;
      RECT 0.0000 2102.0800 3390.2000 2103.7200 ;
      RECT 3388.5000 2101.0000 3390.2000 2102.0800 ;
      RECT 5.3000 2101.0000 3384.9000 2102.0800 ;
      RECT 0.0000 2101.0000 1.7000 2102.0800 ;
      RECT 0.0000 2099.3600 3390.2000 2101.0000 ;
      RECT 3384.5000 2098.2800 3390.2000 2099.3600 ;
      RECT 9.3000 2098.2800 3380.9000 2099.3600 ;
      RECT 0.0000 2098.2800 5.7000 2099.3600 ;
      RECT 0.0000 2096.6400 3390.2000 2098.2800 ;
      RECT 3388.5000 2095.5600 3390.2000 2096.6400 ;
      RECT 5.3000 2095.5600 3384.9000 2096.6400 ;
      RECT 0.0000 2095.5600 1.7000 2096.6400 ;
      RECT 0.0000 2094.2400 3390.2000 2095.5600 ;
      RECT 1.1000 2093.9200 3390.2000 2094.2400 ;
      RECT 1.1000 2093.3400 5.7000 2093.9200 ;
      RECT 3384.5000 2092.8400 3390.2000 2093.9200 ;
      RECT 9.3000 2092.8400 3380.9000 2093.9200 ;
      RECT 0.0000 2092.8400 5.7000 2093.3400 ;
      RECT 0.0000 2091.2000 3390.2000 2092.8400 ;
      RECT 3388.5000 2090.1200 3390.2000 2091.2000 ;
      RECT 5.3000 2090.1200 3384.9000 2091.2000 ;
      RECT 0.0000 2090.1200 1.7000 2091.2000 ;
      RECT 0.0000 2088.4800 3390.2000 2090.1200 ;
      RECT 3384.5000 2087.4000 3390.2000 2088.4800 ;
      RECT 9.3000 2087.4000 3380.9000 2088.4800 ;
      RECT 0.0000 2087.4000 5.7000 2088.4800 ;
      RECT 0.0000 2085.7600 3390.2000 2087.4000 ;
      RECT 3388.5000 2084.6800 3390.2000 2085.7600 ;
      RECT 5.3000 2084.6800 3384.9000 2085.7600 ;
      RECT 0.0000 2084.6800 1.7000 2085.7600 ;
      RECT 0.0000 2083.0400 3390.2000 2084.6800 ;
      RECT 3384.5000 2081.9600 3390.2000 2083.0400 ;
      RECT 9.3000 2081.9600 3380.9000 2083.0400 ;
      RECT 0.0000 2081.9600 5.7000 2083.0400 ;
      RECT 0.0000 2080.3200 3390.2000 2081.9600 ;
      RECT 3388.5000 2079.2400 3390.2000 2080.3200 ;
      RECT 5.3000 2079.2400 3384.9000 2080.3200 ;
      RECT 0.0000 2079.2400 1.7000 2080.3200 ;
      RECT 0.0000 2077.6000 3390.2000 2079.2400 ;
      RECT 3384.5000 2076.5200 3390.2000 2077.6000 ;
      RECT 9.3000 2076.5200 3380.9000 2077.6000 ;
      RECT 0.0000 2076.5200 5.7000 2077.6000 ;
      RECT 0.0000 2074.8800 3390.2000 2076.5200 ;
      RECT 3388.5000 2073.8000 3390.2000 2074.8800 ;
      RECT 5.3000 2073.8000 3384.9000 2074.8800 ;
      RECT 0.0000 2073.8000 1.7000 2074.8800 ;
      RECT 0.0000 2073.5000 3390.2000 2073.8000 ;
      RECT 0.0000 2072.6000 3389.1000 2073.5000 ;
      RECT 0.0000 2072.1600 3390.2000 2072.6000 ;
      RECT 3384.5000 2071.0800 3390.2000 2072.1600 ;
      RECT 9.3000 2071.0800 3380.9000 2072.1600 ;
      RECT 0.0000 2071.0800 5.7000 2072.1600 ;
      RECT 0.0000 2069.4400 3390.2000 2071.0800 ;
      RECT 0.0000 2068.6200 1.7000 2069.4400 ;
      RECT 3388.5000 2068.3600 3390.2000 2069.4400 ;
      RECT 5.3000 2068.3600 3384.9000 2069.4400 ;
      RECT 1.1000 2068.3600 1.7000 2068.6200 ;
      RECT 1.1000 2067.7200 3390.2000 2068.3600 ;
      RECT 0.0000 2066.7200 3390.2000 2067.7200 ;
      RECT 3384.5000 2065.6400 3390.2000 2066.7200 ;
      RECT 9.3000 2065.6400 3380.9000 2066.7200 ;
      RECT 0.0000 2065.6400 5.7000 2066.7200 ;
      RECT 0.0000 2064.0000 3390.2000 2065.6400 ;
      RECT 3388.5000 2062.9200 3390.2000 2064.0000 ;
      RECT 5.3000 2062.9200 3384.9000 2064.0000 ;
      RECT 0.0000 2062.9200 1.7000 2064.0000 ;
      RECT 0.0000 2061.2800 3390.2000 2062.9200 ;
      RECT 3384.5000 2060.2000 3390.2000 2061.2800 ;
      RECT 9.3000 2060.2000 3380.9000 2061.2800 ;
      RECT 0.0000 2060.2000 5.7000 2061.2800 ;
      RECT 0.0000 2058.5600 3390.2000 2060.2000 ;
      RECT 3388.5000 2057.4800 3390.2000 2058.5600 ;
      RECT 5.3000 2057.4800 3384.9000 2058.5600 ;
      RECT 0.0000 2057.4800 1.7000 2058.5600 ;
      RECT 0.0000 2055.8400 3390.2000 2057.4800 ;
      RECT 3384.5000 2054.7600 3390.2000 2055.8400 ;
      RECT 9.3000 2054.7600 3380.9000 2055.8400 ;
      RECT 0.0000 2054.7600 5.7000 2055.8400 ;
      RECT 0.0000 2053.1200 3390.2000 2054.7600 ;
      RECT 3388.5000 2052.0400 3390.2000 2053.1200 ;
      RECT 5.3000 2052.0400 3384.9000 2053.1200 ;
      RECT 0.0000 2052.0400 1.7000 2053.1200 ;
      RECT 0.0000 2050.4000 3390.2000 2052.0400 ;
      RECT 3384.5000 2049.3200 3390.2000 2050.4000 ;
      RECT 9.3000 2049.3200 3380.9000 2050.4000 ;
      RECT 0.0000 2049.3200 5.7000 2050.4000 ;
      RECT 0.0000 2047.6800 3390.2000 2049.3200 ;
      RECT 3388.5000 2046.6000 3390.2000 2047.6800 ;
      RECT 5.3000 2046.6000 3384.9000 2047.6800 ;
      RECT 0.0000 2046.6000 1.7000 2047.6800 ;
      RECT 0.0000 2044.9600 3390.2000 2046.6000 ;
      RECT 3384.5000 2043.8800 3390.2000 2044.9600 ;
      RECT 9.3000 2043.8800 3380.9000 2044.9600 ;
      RECT 0.0000 2043.8800 5.7000 2044.9600 ;
      RECT 0.0000 2043.6100 3390.2000 2043.8800 ;
      RECT 1.1000 2042.7100 3390.2000 2043.6100 ;
      RECT 0.0000 2042.2400 3390.2000 2042.7100 ;
      RECT 3388.5000 2041.1600 3390.2000 2042.2400 ;
      RECT 5.3000 2041.1600 3384.9000 2042.2400 ;
      RECT 0.0000 2041.1600 1.7000 2042.2400 ;
      RECT 0.0000 2039.5200 3390.2000 2041.1600 ;
      RECT 3384.5000 2038.4400 3390.2000 2039.5200 ;
      RECT 9.3000 2038.4400 3380.9000 2039.5200 ;
      RECT 0.0000 2038.4400 5.7000 2039.5200 ;
      RECT 0.0000 2036.8000 3390.2000 2038.4400 ;
      RECT 3388.5000 2035.7200 3390.2000 2036.8000 ;
      RECT 5.3000 2035.7200 3384.9000 2036.8000 ;
      RECT 0.0000 2035.7200 1.7000 2036.8000 ;
      RECT 0.0000 2034.0800 3390.2000 2035.7200 ;
      RECT 3384.5000 2033.0000 3390.2000 2034.0800 ;
      RECT 9.3000 2033.0000 3380.9000 2034.0800 ;
      RECT 0.0000 2033.0000 5.7000 2034.0800 ;
      RECT 0.0000 2031.3600 3390.2000 2033.0000 ;
      RECT 3388.5000 2030.2800 3390.2000 2031.3600 ;
      RECT 5.3000 2030.2800 3384.9000 2031.3600 ;
      RECT 0.0000 2030.2800 1.7000 2031.3600 ;
      RECT 0.0000 2028.6400 3390.2000 2030.2800 ;
      RECT 3384.5000 2027.5600 3390.2000 2028.6400 ;
      RECT 9.3000 2027.5600 3380.9000 2028.6400 ;
      RECT 0.0000 2027.5600 5.7000 2028.6400 ;
      RECT 0.0000 2025.9200 3390.2000 2027.5600 ;
      RECT 3388.5000 2024.8400 3390.2000 2025.9200 ;
      RECT 5.3000 2024.8400 3384.9000 2025.9200 ;
      RECT 0.0000 2024.8400 1.7000 2025.9200 ;
      RECT 0.0000 2023.2000 3390.2000 2024.8400 ;
      RECT 3384.5000 2022.1200 3390.2000 2023.2000 ;
      RECT 9.3000 2022.1200 3380.9000 2023.2000 ;
      RECT 0.0000 2022.1200 5.7000 2023.2000 ;
      RECT 0.0000 2020.4800 3390.2000 2022.1200 ;
      RECT 3388.5000 2019.4000 3390.2000 2020.4800 ;
      RECT 5.3000 2019.4000 3384.9000 2020.4800 ;
      RECT 0.0000 2019.4000 1.7000 2020.4800 ;
      RECT 0.0000 2017.9900 3390.2000 2019.4000 ;
      RECT 1.1000 2017.7600 3390.2000 2017.9900 ;
      RECT 1.1000 2017.0900 5.7000 2017.7600 ;
      RECT 3384.5000 2016.6800 3390.2000 2017.7600 ;
      RECT 9.3000 2016.6800 3380.9000 2017.7600 ;
      RECT 0.0000 2016.6800 5.7000 2017.0900 ;
      RECT 0.0000 2015.0400 3390.2000 2016.6800 ;
      RECT 3388.5000 2013.9600 3390.2000 2015.0400 ;
      RECT 5.3000 2013.9600 3384.9000 2015.0400 ;
      RECT 0.0000 2013.9600 1.7000 2015.0400 ;
      RECT 0.0000 2012.3200 3390.2000 2013.9600 ;
      RECT 3384.5000 2011.2400 3390.2000 2012.3200 ;
      RECT 9.3000 2011.2400 3380.9000 2012.3200 ;
      RECT 0.0000 2011.2400 5.7000 2012.3200 ;
      RECT 0.0000 2009.6000 3390.2000 2011.2400 ;
      RECT 3388.5000 2008.5200 3390.2000 2009.6000 ;
      RECT 5.3000 2008.5200 3384.9000 2009.6000 ;
      RECT 0.0000 2008.5200 1.7000 2009.6000 ;
      RECT 0.0000 2006.8800 3390.2000 2008.5200 ;
      RECT 3384.5000 2005.8000 3390.2000 2006.8800 ;
      RECT 9.3000 2005.8000 3380.9000 2006.8800 ;
      RECT 0.0000 2005.8000 5.7000 2006.8800 ;
      RECT 0.0000 2004.1600 3390.2000 2005.8000 ;
      RECT 3388.5000 2003.0800 3390.2000 2004.1600 ;
      RECT 5.3000 2003.0800 3384.9000 2004.1600 ;
      RECT 0.0000 2003.0800 1.7000 2004.1600 ;
      RECT 0.0000 2001.4400 3390.2000 2003.0800 ;
      RECT 3384.5000 2000.3600 3390.2000 2001.4400 ;
      RECT 9.3000 2000.3600 3380.9000 2001.4400 ;
      RECT 0.0000 2000.3600 5.7000 2001.4400 ;
      RECT 0.0000 1998.7200 3390.2000 2000.3600 ;
      RECT 3388.5000 1997.6400 3390.2000 1998.7200 ;
      RECT 5.3000 1997.6400 3384.9000 1998.7200 ;
      RECT 0.0000 1997.6400 1.7000 1998.7200 ;
      RECT 0.0000 1996.0000 3390.2000 1997.6400 ;
      RECT 3384.5000 1994.9200 3390.2000 1996.0000 ;
      RECT 9.3000 1994.9200 3380.9000 1996.0000 ;
      RECT 0.0000 1994.9200 5.7000 1996.0000 ;
      RECT 0.0000 1993.2800 3390.2000 1994.9200 ;
      RECT 0.0000 1992.9800 1.7000 1993.2800 ;
      RECT 3388.5000 1992.2000 3390.2000 1993.2800 ;
      RECT 5.3000 1992.2000 3384.9000 1993.2800 ;
      RECT 1.1000 1992.2000 1.7000 1992.9800 ;
      RECT 1.1000 1992.0800 3390.2000 1992.2000 ;
      RECT 0.0000 1990.5600 3390.2000 1992.0800 ;
      RECT 3384.5000 1989.4800 3390.2000 1990.5600 ;
      RECT 9.3000 1989.4800 3380.9000 1990.5600 ;
      RECT 0.0000 1989.4800 5.7000 1990.5600 ;
      RECT 0.0000 1987.8400 3390.2000 1989.4800 ;
      RECT 3388.5000 1986.7600 3390.2000 1987.8400 ;
      RECT 5.3000 1986.7600 3384.9000 1987.8400 ;
      RECT 0.0000 1986.7600 1.7000 1987.8400 ;
      RECT 0.0000 1985.1200 3390.2000 1986.7600 ;
      RECT 3384.5000 1984.0400 3390.2000 1985.1200 ;
      RECT 9.3000 1984.0400 3380.9000 1985.1200 ;
      RECT 0.0000 1984.0400 5.7000 1985.1200 ;
      RECT 0.0000 1982.4000 3390.2000 1984.0400 ;
      RECT 3388.5000 1981.3200 3390.2000 1982.4000 ;
      RECT 5.3000 1981.3200 3384.9000 1982.4000 ;
      RECT 0.0000 1981.3200 1.7000 1982.4000 ;
      RECT 0.0000 1979.6800 3390.2000 1981.3200 ;
      RECT 3384.5000 1978.6000 3390.2000 1979.6800 ;
      RECT 9.3000 1978.6000 3380.9000 1979.6800 ;
      RECT 0.0000 1978.6000 5.7000 1979.6800 ;
      RECT 0.0000 1976.9600 3390.2000 1978.6000 ;
      RECT 3388.5000 1975.8800 3390.2000 1976.9600 ;
      RECT 5.3000 1975.8800 3384.9000 1976.9600 ;
      RECT 0.0000 1975.8800 1.7000 1976.9600 ;
      RECT 0.0000 1974.2400 3390.2000 1975.8800 ;
      RECT 3384.5000 1973.1600 3390.2000 1974.2400 ;
      RECT 9.3000 1973.1600 3380.9000 1974.2400 ;
      RECT 0.0000 1973.1600 5.7000 1974.2400 ;
      RECT 0.0000 1971.5200 3390.2000 1973.1600 ;
      RECT 3388.5000 1970.4400 3390.2000 1971.5200 ;
      RECT 5.3000 1970.4400 3384.9000 1971.5200 ;
      RECT 0.0000 1970.4400 1.7000 1971.5200 ;
      RECT 0.0000 1969.8000 3390.2000 1970.4400 ;
      RECT 0.0000 1968.9000 3389.1000 1969.8000 ;
      RECT 0.0000 1968.8000 3390.2000 1968.9000 ;
      RECT 0.0000 1967.9700 5.7000 1968.8000 ;
      RECT 3384.5000 1967.7200 3390.2000 1968.8000 ;
      RECT 9.3000 1967.7200 3380.9000 1968.8000 ;
      RECT 1.1000 1967.7200 5.7000 1967.9700 ;
      RECT 1.1000 1967.0700 3390.2000 1967.7200 ;
      RECT 0.0000 1966.0800 3390.2000 1967.0700 ;
      RECT 3388.5000 1965.0000 3390.2000 1966.0800 ;
      RECT 5.3000 1965.0000 3384.9000 1966.0800 ;
      RECT 0.0000 1965.0000 1.7000 1966.0800 ;
      RECT 0.0000 1963.3600 3390.2000 1965.0000 ;
      RECT 3384.5000 1962.2800 3390.2000 1963.3600 ;
      RECT 9.3000 1962.2800 3380.9000 1963.3600 ;
      RECT 0.0000 1962.2800 5.7000 1963.3600 ;
      RECT 0.0000 1960.6400 3390.2000 1962.2800 ;
      RECT 3388.5000 1959.5600 3390.2000 1960.6400 ;
      RECT 5.3000 1959.5600 3384.9000 1960.6400 ;
      RECT 0.0000 1959.5600 1.7000 1960.6400 ;
      RECT 0.0000 1957.9200 3390.2000 1959.5600 ;
      RECT 3384.5000 1956.8400 3390.2000 1957.9200 ;
      RECT 9.3000 1956.8400 3380.9000 1957.9200 ;
      RECT 0.0000 1956.8400 5.7000 1957.9200 ;
      RECT 0.0000 1955.2000 3390.2000 1956.8400 ;
      RECT 3388.5000 1954.1200 3390.2000 1955.2000 ;
      RECT 5.3000 1954.1200 3384.9000 1955.2000 ;
      RECT 0.0000 1954.1200 1.7000 1955.2000 ;
      RECT 0.0000 1952.4800 3390.2000 1954.1200 ;
      RECT 3384.5000 1951.4000 3390.2000 1952.4800 ;
      RECT 9.3000 1951.4000 3380.9000 1952.4800 ;
      RECT 0.0000 1951.4000 5.7000 1952.4800 ;
      RECT 0.0000 1949.7600 3390.2000 1951.4000 ;
      RECT 3388.5000 1948.6800 3390.2000 1949.7600 ;
      RECT 5.3000 1948.6800 3384.9000 1949.7600 ;
      RECT 0.0000 1948.6800 1.7000 1949.7600 ;
      RECT 0.0000 1947.0400 3390.2000 1948.6800 ;
      RECT 3384.5000 1945.9600 3390.2000 1947.0400 ;
      RECT 9.3000 1945.9600 3380.9000 1947.0400 ;
      RECT 0.0000 1945.9600 5.7000 1947.0400 ;
      RECT 0.0000 1944.3200 3390.2000 1945.9600 ;
      RECT 3388.5000 1943.2400 3390.2000 1944.3200 ;
      RECT 5.3000 1943.2400 3384.9000 1944.3200 ;
      RECT 0.0000 1943.2400 1.7000 1944.3200 ;
      RECT 0.0000 1942.3500 3390.2000 1943.2400 ;
      RECT 1.1000 1941.6000 3390.2000 1942.3500 ;
      RECT 1.1000 1941.4500 5.7000 1941.6000 ;
      RECT 3384.5000 1940.5200 3390.2000 1941.6000 ;
      RECT 9.3000 1940.5200 3380.9000 1941.6000 ;
      RECT 0.0000 1940.5200 5.7000 1941.4500 ;
      RECT 0.0000 1938.8800 3390.2000 1940.5200 ;
      RECT 3388.5000 1937.8000 3390.2000 1938.8800 ;
      RECT 5.3000 1937.8000 3384.9000 1938.8800 ;
      RECT 0.0000 1937.8000 1.7000 1938.8800 ;
      RECT 0.0000 1936.1600 3390.2000 1937.8000 ;
      RECT 3384.5000 1935.0800 3390.2000 1936.1600 ;
      RECT 9.3000 1935.0800 3380.9000 1936.1600 ;
      RECT 0.0000 1935.0800 5.7000 1936.1600 ;
      RECT 0.0000 1933.4400 3390.2000 1935.0800 ;
      RECT 3388.5000 1932.3600 3390.2000 1933.4400 ;
      RECT 5.3000 1932.3600 3384.9000 1933.4400 ;
      RECT 0.0000 1932.3600 1.7000 1933.4400 ;
      RECT 0.0000 1930.7200 3390.2000 1932.3600 ;
      RECT 3384.5000 1929.6400 3390.2000 1930.7200 ;
      RECT 9.3000 1929.6400 3380.9000 1930.7200 ;
      RECT 0.0000 1929.6400 5.7000 1930.7200 ;
      RECT 0.0000 1928.0000 3390.2000 1929.6400 ;
      RECT 3388.5000 1926.9200 3390.2000 1928.0000 ;
      RECT 5.3000 1926.9200 3384.9000 1928.0000 ;
      RECT 0.0000 1926.9200 1.7000 1928.0000 ;
      RECT 0.0000 1925.2800 3390.2000 1926.9200 ;
      RECT 3384.5000 1924.2000 3390.2000 1925.2800 ;
      RECT 9.3000 1924.2000 3380.9000 1925.2800 ;
      RECT 0.0000 1924.2000 5.7000 1925.2800 ;
      RECT 0.0000 1922.5600 3390.2000 1924.2000 ;
      RECT 3388.5000 1921.4800 3390.2000 1922.5600 ;
      RECT 5.3000 1921.4800 3384.9000 1922.5600 ;
      RECT 0.0000 1921.4800 1.7000 1922.5600 ;
      RECT 0.0000 1919.8400 3390.2000 1921.4800 ;
      RECT 3384.5000 1918.7600 3390.2000 1919.8400 ;
      RECT 9.3000 1918.7600 3380.9000 1919.8400 ;
      RECT 0.0000 1918.7600 5.7000 1919.8400 ;
      RECT 0.0000 1917.3400 3390.2000 1918.7600 ;
      RECT 1.1000 1917.1200 3390.2000 1917.3400 ;
      RECT 1.1000 1916.4400 1.7000 1917.1200 ;
      RECT 3388.5000 1916.0400 3390.2000 1917.1200 ;
      RECT 5.3000 1916.0400 3384.9000 1917.1200 ;
      RECT 0.0000 1916.0400 1.7000 1916.4400 ;
      RECT 0.0000 1914.4000 3390.2000 1916.0400 ;
      RECT 3384.5000 1913.3200 3390.2000 1914.4000 ;
      RECT 9.3000 1913.3200 3380.9000 1914.4000 ;
      RECT 0.0000 1913.3200 5.7000 1914.4000 ;
      RECT 0.0000 1911.6800 3390.2000 1913.3200 ;
      RECT 3388.5000 1910.6000 3390.2000 1911.6800 ;
      RECT 5.3000 1910.6000 3384.9000 1911.6800 ;
      RECT 0.0000 1910.6000 1.7000 1911.6800 ;
      RECT 0.0000 1908.9600 3390.2000 1910.6000 ;
      RECT 3384.5000 1907.8800 3390.2000 1908.9600 ;
      RECT 9.3000 1907.8800 3380.9000 1908.9600 ;
      RECT 0.0000 1907.8800 5.7000 1908.9600 ;
      RECT 0.0000 1906.2400 3390.2000 1907.8800 ;
      RECT 3388.5000 1905.1600 3390.2000 1906.2400 ;
      RECT 5.3000 1905.1600 3384.9000 1906.2400 ;
      RECT 0.0000 1905.1600 1.7000 1906.2400 ;
      RECT 0.0000 1903.5200 3390.2000 1905.1600 ;
      RECT 3384.5000 1902.4400 3390.2000 1903.5200 ;
      RECT 9.3000 1902.4400 3380.9000 1903.5200 ;
      RECT 0.0000 1902.4400 5.7000 1903.5200 ;
      RECT 0.0000 1900.8000 3390.2000 1902.4400 ;
      RECT 3388.5000 1899.7200 3390.2000 1900.8000 ;
      RECT 5.3000 1899.7200 3384.9000 1900.8000 ;
      RECT 0.0000 1899.7200 1.7000 1900.8000 ;
      RECT 0.0000 1898.0800 3390.2000 1899.7200 ;
      RECT 3384.5000 1897.0000 3390.2000 1898.0800 ;
      RECT 9.3000 1897.0000 3380.9000 1898.0800 ;
      RECT 0.0000 1897.0000 5.7000 1898.0800 ;
      RECT 0.0000 1895.3600 3390.2000 1897.0000 ;
      RECT 3388.5000 1894.2800 3390.2000 1895.3600 ;
      RECT 5.3000 1894.2800 3384.9000 1895.3600 ;
      RECT 0.0000 1894.2800 1.7000 1895.3600 ;
      RECT 0.0000 1892.6400 3390.2000 1894.2800 ;
      RECT 0.0000 1892.3300 5.7000 1892.6400 ;
      RECT 3384.5000 1891.5600 3390.2000 1892.6400 ;
      RECT 9.3000 1891.5600 3380.9000 1892.6400 ;
      RECT 1.1000 1891.5600 5.7000 1892.3300 ;
      RECT 1.1000 1891.4300 3390.2000 1891.5600 ;
      RECT 0.0000 1889.9200 3390.2000 1891.4300 ;
      RECT 3388.5000 1888.8400 3390.2000 1889.9200 ;
      RECT 5.3000 1888.8400 3384.9000 1889.9200 ;
      RECT 0.0000 1888.8400 1.7000 1889.9200 ;
      RECT 0.0000 1887.2000 3390.2000 1888.8400 ;
      RECT 3384.5000 1886.1200 3390.2000 1887.2000 ;
      RECT 9.3000 1886.1200 3380.9000 1887.2000 ;
      RECT 0.0000 1886.1200 5.7000 1887.2000 ;
      RECT 0.0000 1884.4800 3390.2000 1886.1200 ;
      RECT 3388.5000 1883.4000 3390.2000 1884.4800 ;
      RECT 5.3000 1883.4000 3384.9000 1884.4800 ;
      RECT 0.0000 1883.4000 1.7000 1884.4800 ;
      RECT 0.0000 1881.7600 3390.2000 1883.4000 ;
      RECT 3384.5000 1880.6800 3390.2000 1881.7600 ;
      RECT 9.3000 1880.6800 3380.9000 1881.7600 ;
      RECT 0.0000 1880.6800 5.7000 1881.7600 ;
      RECT 0.0000 1879.0400 3390.2000 1880.6800 ;
      RECT 3388.5000 1877.9600 3390.2000 1879.0400 ;
      RECT 5.3000 1877.9600 3384.9000 1879.0400 ;
      RECT 0.0000 1877.9600 1.7000 1879.0400 ;
      RECT 0.0000 1876.3200 3390.2000 1877.9600 ;
      RECT 3384.5000 1875.2400 3390.2000 1876.3200 ;
      RECT 9.3000 1875.2400 3380.9000 1876.3200 ;
      RECT 0.0000 1875.2400 5.7000 1876.3200 ;
      RECT 0.0000 1873.6000 3390.2000 1875.2400 ;
      RECT 3388.5000 1872.5200 3390.2000 1873.6000 ;
      RECT 5.3000 1872.5200 3384.9000 1873.6000 ;
      RECT 0.0000 1872.5200 1.7000 1873.6000 ;
      RECT 0.0000 1870.8800 3390.2000 1872.5200 ;
      RECT 3384.5000 1869.8000 3390.2000 1870.8800 ;
      RECT 9.3000 1869.8000 3380.9000 1870.8800 ;
      RECT 0.0000 1869.8000 5.7000 1870.8800 ;
      RECT 0.0000 1868.1600 3390.2000 1869.8000 ;
      RECT 3388.5000 1867.0800 3390.2000 1868.1600 ;
      RECT 5.3000 1867.0800 3384.9000 1868.1600 ;
      RECT 0.0000 1867.0800 1.7000 1868.1600 ;
      RECT 0.0000 1866.7100 3390.2000 1867.0800 ;
      RECT 1.1000 1866.1000 3390.2000 1866.7100 ;
      RECT 1.1000 1865.8100 3389.1000 1866.1000 ;
      RECT 0.0000 1865.4400 3389.1000 1865.8100 ;
      RECT 3384.5000 1865.2000 3389.1000 1865.4400 ;
      RECT 3384.5000 1864.3600 3390.2000 1865.2000 ;
      RECT 9.3000 1864.3600 3380.9000 1865.4400 ;
      RECT 0.0000 1864.3600 5.7000 1865.4400 ;
      RECT 0.0000 1862.7200 3390.2000 1864.3600 ;
      RECT 3388.5000 1861.6400 3390.2000 1862.7200 ;
      RECT 5.3000 1861.6400 3384.9000 1862.7200 ;
      RECT 0.0000 1861.6400 1.7000 1862.7200 ;
      RECT 0.0000 1860.0000 3390.2000 1861.6400 ;
      RECT 3384.5000 1858.9200 3390.2000 1860.0000 ;
      RECT 9.3000 1858.9200 3380.9000 1860.0000 ;
      RECT 0.0000 1858.9200 5.7000 1860.0000 ;
      RECT 0.0000 1857.2800 3390.2000 1858.9200 ;
      RECT 3388.5000 1856.2000 3390.2000 1857.2800 ;
      RECT 5.3000 1856.2000 3384.9000 1857.2800 ;
      RECT 0.0000 1856.2000 1.7000 1857.2800 ;
      RECT 0.0000 1854.5600 3390.2000 1856.2000 ;
      RECT 3384.5000 1853.4800 3390.2000 1854.5600 ;
      RECT 9.3000 1853.4800 3380.9000 1854.5600 ;
      RECT 0.0000 1853.4800 5.7000 1854.5600 ;
      RECT 0.0000 1851.8400 3390.2000 1853.4800 ;
      RECT 3388.5000 1850.7600 3390.2000 1851.8400 ;
      RECT 5.3000 1850.7600 3384.9000 1851.8400 ;
      RECT 0.0000 1850.7600 1.7000 1851.8400 ;
      RECT 0.0000 1849.1200 3390.2000 1850.7600 ;
      RECT 3384.5000 1848.0400 3390.2000 1849.1200 ;
      RECT 9.3000 1848.0400 3380.9000 1849.1200 ;
      RECT 0.0000 1848.0400 5.7000 1849.1200 ;
      RECT 0.0000 1846.4000 3390.2000 1848.0400 ;
      RECT 3388.5000 1845.3200 3390.2000 1846.4000 ;
      RECT 5.3000 1845.3200 3384.9000 1846.4000 ;
      RECT 0.0000 1845.3200 1.7000 1846.4000 ;
      RECT 0.0000 1843.6800 3390.2000 1845.3200 ;
      RECT 3384.5000 1842.6000 3390.2000 1843.6800 ;
      RECT 9.3000 1842.6000 3380.9000 1843.6800 ;
      RECT 0.0000 1842.6000 5.7000 1843.6800 ;
      RECT 0.0000 1841.7000 3390.2000 1842.6000 ;
      RECT 1.1000 1840.9600 3390.2000 1841.7000 ;
      RECT 1.1000 1840.8000 1.7000 1840.9600 ;
      RECT 3388.5000 1839.8800 3390.2000 1840.9600 ;
      RECT 5.3000 1839.8800 3384.9000 1840.9600 ;
      RECT 0.0000 1839.8800 1.7000 1840.8000 ;
      RECT 0.0000 1838.2400 3390.2000 1839.8800 ;
      RECT 3384.5000 1837.1600 3390.2000 1838.2400 ;
      RECT 9.3000 1837.1600 3380.9000 1838.2400 ;
      RECT 0.0000 1837.1600 5.7000 1838.2400 ;
      RECT 0.0000 1835.5200 3390.2000 1837.1600 ;
      RECT 3388.5000 1834.4400 3390.2000 1835.5200 ;
      RECT 5.3000 1834.4400 3384.9000 1835.5200 ;
      RECT 0.0000 1834.4400 1.7000 1835.5200 ;
      RECT 0.0000 1832.8000 3390.2000 1834.4400 ;
      RECT 3384.5000 1831.7200 3390.2000 1832.8000 ;
      RECT 9.3000 1831.7200 3380.9000 1832.8000 ;
      RECT 0.0000 1831.7200 5.7000 1832.8000 ;
      RECT 0.0000 1830.0800 3390.2000 1831.7200 ;
      RECT 3388.5000 1829.0000 3390.2000 1830.0800 ;
      RECT 5.3000 1829.0000 3384.9000 1830.0800 ;
      RECT 0.0000 1829.0000 1.7000 1830.0800 ;
      RECT 0.0000 1827.3600 3390.2000 1829.0000 ;
      RECT 3384.5000 1826.2800 3390.2000 1827.3600 ;
      RECT 9.3000 1826.2800 3380.9000 1827.3600 ;
      RECT 0.0000 1826.2800 5.7000 1827.3600 ;
      RECT 0.0000 1824.6400 3390.2000 1826.2800 ;
      RECT 3388.5000 1823.5600 3390.2000 1824.6400 ;
      RECT 5.3000 1823.5600 3384.9000 1824.6400 ;
      RECT 0.0000 1823.5600 1.7000 1824.6400 ;
      RECT 0.0000 1821.9200 3390.2000 1823.5600 ;
      RECT 3384.5000 1820.8400 3390.2000 1821.9200 ;
      RECT 9.3000 1820.8400 3380.9000 1821.9200 ;
      RECT 0.0000 1820.8400 5.7000 1821.9200 ;
      RECT 0.0000 1819.2000 3390.2000 1820.8400 ;
      RECT 3388.5000 1818.1200 3390.2000 1819.2000 ;
      RECT 5.3000 1818.1200 3384.9000 1819.2000 ;
      RECT 0.0000 1818.1200 1.7000 1819.2000 ;
      RECT 0.0000 1816.6900 3390.2000 1818.1200 ;
      RECT 1.1000 1816.4800 3390.2000 1816.6900 ;
      RECT 1.1000 1815.7900 5.7000 1816.4800 ;
      RECT 3384.5000 1815.4000 3390.2000 1816.4800 ;
      RECT 9.3000 1815.4000 3380.9000 1816.4800 ;
      RECT 0.0000 1815.4000 5.7000 1815.7900 ;
      RECT 0.0000 1813.7600 3390.2000 1815.4000 ;
      RECT 3388.5000 1812.6800 3390.2000 1813.7600 ;
      RECT 5.3000 1812.6800 3384.9000 1813.7600 ;
      RECT 0.0000 1812.6800 1.7000 1813.7600 ;
      RECT 0.0000 1811.0400 3390.2000 1812.6800 ;
      RECT 3384.5000 1809.9600 3390.2000 1811.0400 ;
      RECT 9.3000 1809.9600 3380.9000 1811.0400 ;
      RECT 0.0000 1809.9600 5.7000 1811.0400 ;
      RECT 0.0000 1808.3200 3390.2000 1809.9600 ;
      RECT 3388.5000 1807.2400 3390.2000 1808.3200 ;
      RECT 5.3000 1807.2400 3384.9000 1808.3200 ;
      RECT 0.0000 1807.2400 1.7000 1808.3200 ;
      RECT 0.0000 1805.6000 3390.2000 1807.2400 ;
      RECT 3384.5000 1804.5200 3390.2000 1805.6000 ;
      RECT 9.3000 1804.5200 3380.9000 1805.6000 ;
      RECT 0.0000 1804.5200 5.7000 1805.6000 ;
      RECT 0.0000 1802.8800 3390.2000 1804.5200 ;
      RECT 3388.5000 1801.8000 3390.2000 1802.8800 ;
      RECT 5.3000 1801.8000 3384.9000 1802.8800 ;
      RECT 0.0000 1801.8000 1.7000 1802.8800 ;
      RECT 0.0000 1800.1600 3390.2000 1801.8000 ;
      RECT 3384.5000 1799.0800 3390.2000 1800.1600 ;
      RECT 9.3000 1799.0800 3380.9000 1800.1600 ;
      RECT 0.0000 1799.0800 5.7000 1800.1600 ;
      RECT 0.0000 1797.4400 3390.2000 1799.0800 ;
      RECT 3388.5000 1796.3600 3390.2000 1797.4400 ;
      RECT 5.3000 1796.3600 3384.9000 1797.4400 ;
      RECT 0.0000 1796.3600 1.7000 1797.4400 ;
      RECT 0.0000 1794.7200 3390.2000 1796.3600 ;
      RECT 3384.5000 1793.6400 3390.2000 1794.7200 ;
      RECT 9.3000 1793.6400 3380.9000 1794.7200 ;
      RECT 0.0000 1793.6400 5.7000 1794.7200 ;
      RECT 0.0000 1792.0000 3390.2000 1793.6400 ;
      RECT 0.0000 1791.0700 1.7000 1792.0000 ;
      RECT 3388.5000 1790.9200 3390.2000 1792.0000 ;
      RECT 5.3000 1790.9200 3384.9000 1792.0000 ;
      RECT 1.1000 1790.9200 1.7000 1791.0700 ;
      RECT 1.1000 1790.1700 3390.2000 1790.9200 ;
      RECT 0.0000 1789.2800 3390.2000 1790.1700 ;
      RECT 3384.5000 1788.2000 3390.2000 1789.2800 ;
      RECT 9.3000 1788.2000 3380.9000 1789.2800 ;
      RECT 0.0000 1788.2000 5.7000 1789.2800 ;
      RECT 0.0000 1786.5600 3390.2000 1788.2000 ;
      RECT 3388.5000 1785.4800 3390.2000 1786.5600 ;
      RECT 5.3000 1785.4800 3384.9000 1786.5600 ;
      RECT 0.0000 1785.4800 1.7000 1786.5600 ;
      RECT 0.0000 1783.8400 3390.2000 1785.4800 ;
      RECT 3384.5000 1782.7600 3390.2000 1783.8400 ;
      RECT 9.3000 1782.7600 3380.9000 1783.8400 ;
      RECT 0.0000 1782.7600 5.7000 1783.8400 ;
      RECT 0.0000 1781.1200 3390.2000 1782.7600 ;
      RECT 3388.5000 1780.0400 3390.2000 1781.1200 ;
      RECT 5.3000 1780.0400 3384.9000 1781.1200 ;
      RECT 0.0000 1780.0400 1.7000 1781.1200 ;
      RECT 0.0000 1778.4000 3390.2000 1780.0400 ;
      RECT 3384.5000 1777.3200 3390.2000 1778.4000 ;
      RECT 9.3000 1777.3200 3380.9000 1778.4000 ;
      RECT 0.0000 1777.3200 5.7000 1778.4000 ;
      RECT 0.0000 1775.6800 3390.2000 1777.3200 ;
      RECT 3388.5000 1774.6000 3390.2000 1775.6800 ;
      RECT 5.3000 1774.6000 3384.9000 1775.6800 ;
      RECT 0.0000 1774.6000 1.7000 1775.6800 ;
      RECT 0.0000 1772.9600 3390.2000 1774.6000 ;
      RECT 3384.5000 1771.8800 3390.2000 1772.9600 ;
      RECT 9.3000 1771.8800 3380.9000 1772.9600 ;
      RECT 0.0000 1771.8800 5.7000 1772.9600 ;
      RECT 0.0000 1770.2400 3390.2000 1771.8800 ;
      RECT 3388.5000 1769.1600 3390.2000 1770.2400 ;
      RECT 5.3000 1769.1600 3384.9000 1770.2400 ;
      RECT 0.0000 1769.1600 1.7000 1770.2400 ;
      RECT 0.0000 1767.5200 3390.2000 1769.1600 ;
      RECT 3384.5000 1766.4400 3390.2000 1767.5200 ;
      RECT 9.3000 1766.4400 3380.9000 1767.5200 ;
      RECT 0.0000 1766.4400 5.7000 1767.5200 ;
      RECT 0.0000 1766.0600 3390.2000 1766.4400 ;
      RECT 1.1000 1765.1600 3390.2000 1766.0600 ;
      RECT 0.0000 1764.8000 3390.2000 1765.1600 ;
      RECT 3388.5000 1763.7200 3390.2000 1764.8000 ;
      RECT 5.3000 1763.7200 3384.9000 1764.8000 ;
      RECT 0.0000 1763.7200 1.7000 1764.8000 ;
      RECT 0.0000 1762.4000 3390.2000 1763.7200 ;
      RECT 0.0000 1762.0800 3389.1000 1762.4000 ;
      RECT 3384.5000 1761.5000 3389.1000 1762.0800 ;
      RECT 3384.5000 1761.0000 3390.2000 1761.5000 ;
      RECT 9.3000 1761.0000 3380.9000 1762.0800 ;
      RECT 0.0000 1761.0000 5.7000 1762.0800 ;
      RECT 0.0000 1759.3600 3390.2000 1761.0000 ;
      RECT 3388.5000 1758.2800 3390.2000 1759.3600 ;
      RECT 5.3000 1758.2800 3384.9000 1759.3600 ;
      RECT 0.0000 1758.2800 1.7000 1759.3600 ;
      RECT 0.0000 1756.6400 3390.2000 1758.2800 ;
      RECT 3384.5000 1755.5600 3390.2000 1756.6400 ;
      RECT 9.3000 1755.5600 3380.9000 1756.6400 ;
      RECT 0.0000 1755.5600 5.7000 1756.6400 ;
      RECT 0.0000 1753.9200 3390.2000 1755.5600 ;
      RECT 3388.5000 1752.8400 3390.2000 1753.9200 ;
      RECT 5.3000 1752.8400 3384.9000 1753.9200 ;
      RECT 0.0000 1752.8400 1.7000 1753.9200 ;
      RECT 0.0000 1751.2000 3390.2000 1752.8400 ;
      RECT 3384.5000 1750.1200 3390.2000 1751.2000 ;
      RECT 9.3000 1750.1200 3380.9000 1751.2000 ;
      RECT 0.0000 1750.1200 5.7000 1751.2000 ;
      RECT 0.0000 1748.4800 3390.2000 1750.1200 ;
      RECT 3388.5000 1747.4000 3390.2000 1748.4800 ;
      RECT 5.3000 1747.4000 3384.9000 1748.4800 ;
      RECT 0.0000 1747.4000 1.7000 1748.4800 ;
      RECT 0.0000 1745.7600 3390.2000 1747.4000 ;
      RECT 3384.5000 1744.6800 3390.2000 1745.7600 ;
      RECT 9.3000 1744.6800 3380.9000 1745.7600 ;
      RECT 0.0000 1744.6800 5.7000 1745.7600 ;
      RECT 0.0000 1743.0400 3390.2000 1744.6800 ;
      RECT 3388.5000 1741.9600 3390.2000 1743.0400 ;
      RECT 5.3000 1741.9600 3384.9000 1743.0400 ;
      RECT 0.0000 1741.9600 1.7000 1743.0400 ;
      RECT 0.0000 1741.0500 3390.2000 1741.9600 ;
      RECT 1.1000 1740.3200 3390.2000 1741.0500 ;
      RECT 1.1000 1740.1500 5.7000 1740.3200 ;
      RECT 3384.5000 1739.2400 3390.2000 1740.3200 ;
      RECT 9.3000 1739.2400 3380.9000 1740.3200 ;
      RECT 0.0000 1739.2400 5.7000 1740.1500 ;
      RECT 0.0000 1737.6000 3390.2000 1739.2400 ;
      RECT 3388.5000 1736.5200 3390.2000 1737.6000 ;
      RECT 5.3000 1736.5200 3384.9000 1737.6000 ;
      RECT 0.0000 1736.5200 1.7000 1737.6000 ;
      RECT 0.0000 1734.8800 3390.2000 1736.5200 ;
      RECT 3384.5000 1733.8000 3390.2000 1734.8800 ;
      RECT 9.3000 1733.8000 3380.9000 1734.8800 ;
      RECT 0.0000 1733.8000 5.7000 1734.8800 ;
      RECT 0.0000 1732.1600 3390.2000 1733.8000 ;
      RECT 3388.5000 1731.0800 3390.2000 1732.1600 ;
      RECT 5.3000 1731.0800 3384.9000 1732.1600 ;
      RECT 0.0000 1731.0800 1.7000 1732.1600 ;
      RECT 0.0000 1729.4400 3390.2000 1731.0800 ;
      RECT 3384.5000 1728.3600 3390.2000 1729.4400 ;
      RECT 9.3000 1728.3600 3380.9000 1729.4400 ;
      RECT 0.0000 1728.3600 5.7000 1729.4400 ;
      RECT 0.0000 1726.7200 3390.2000 1728.3600 ;
      RECT 3388.5000 1725.6400 3390.2000 1726.7200 ;
      RECT 5.3000 1725.6400 3384.9000 1726.7200 ;
      RECT 0.0000 1725.6400 1.7000 1726.7200 ;
      RECT 0.0000 1724.0000 3390.2000 1725.6400 ;
      RECT 3384.5000 1722.9200 3390.2000 1724.0000 ;
      RECT 9.3000 1722.9200 3380.9000 1724.0000 ;
      RECT 0.0000 1722.9200 5.7000 1724.0000 ;
      RECT 0.0000 1721.2800 3390.2000 1722.9200 ;
      RECT 3388.5000 1720.2000 3390.2000 1721.2800 ;
      RECT 5.3000 1720.2000 3384.9000 1721.2800 ;
      RECT 0.0000 1720.2000 1.7000 1721.2800 ;
      RECT 0.0000 1718.5600 3390.2000 1720.2000 ;
      RECT 3384.5000 1717.4800 3390.2000 1718.5600 ;
      RECT 9.3000 1717.4800 3380.9000 1718.5600 ;
      RECT 0.0000 1717.4800 5.7000 1718.5600 ;
      RECT 0.0000 1715.8400 3390.2000 1717.4800 ;
      RECT 0.0000 1715.4300 1.7000 1715.8400 ;
      RECT 3388.5000 1714.7600 3390.2000 1715.8400 ;
      RECT 5.3000 1714.7600 3384.9000 1715.8400 ;
      RECT 1.1000 1714.7600 1.7000 1715.4300 ;
      RECT 1.1000 1714.5300 3390.2000 1714.7600 ;
      RECT 0.0000 1713.1200 3390.2000 1714.5300 ;
      RECT 3384.5000 1712.0400 3390.2000 1713.1200 ;
      RECT 9.3000 1712.0400 3380.9000 1713.1200 ;
      RECT 0.0000 1712.0400 5.7000 1713.1200 ;
      RECT 0.0000 1710.4000 3390.2000 1712.0400 ;
      RECT 3388.5000 1709.3200 3390.2000 1710.4000 ;
      RECT 5.3000 1709.3200 3384.9000 1710.4000 ;
      RECT 0.0000 1709.3200 1.7000 1710.4000 ;
      RECT 0.0000 1707.6800 3390.2000 1709.3200 ;
      RECT 3384.5000 1706.6000 3390.2000 1707.6800 ;
      RECT 9.3000 1706.6000 3380.9000 1707.6800 ;
      RECT 0.0000 1706.6000 5.7000 1707.6800 ;
      RECT 0.0000 1704.9600 3390.2000 1706.6000 ;
      RECT 3388.5000 1703.8800 3390.2000 1704.9600 ;
      RECT 5.3000 1703.8800 3384.9000 1704.9600 ;
      RECT 0.0000 1703.8800 1.7000 1704.9600 ;
      RECT 0.0000 1702.2400 3390.2000 1703.8800 ;
      RECT 3384.5000 1701.1600 3390.2000 1702.2400 ;
      RECT 9.3000 1701.1600 3380.9000 1702.2400 ;
      RECT 0.0000 1701.1600 5.7000 1702.2400 ;
      RECT 0.0000 1699.5200 3390.2000 1701.1600 ;
      RECT 3388.5000 1698.4400 3390.2000 1699.5200 ;
      RECT 5.3000 1698.4400 3384.9000 1699.5200 ;
      RECT 0.0000 1698.4400 1.7000 1699.5200 ;
      RECT 0.0000 1696.8000 3390.2000 1698.4400 ;
      RECT 3384.5000 1695.7200 3390.2000 1696.8000 ;
      RECT 9.3000 1695.7200 3380.9000 1696.8000 ;
      RECT 0.0000 1695.7200 5.7000 1696.8000 ;
      RECT 0.0000 1694.0800 3390.2000 1695.7200 ;
      RECT 3388.5000 1693.0000 3390.2000 1694.0800 ;
      RECT 5.3000 1693.0000 3384.9000 1694.0800 ;
      RECT 0.0000 1693.0000 1.7000 1694.0800 ;
      RECT 0.0000 1691.3600 3390.2000 1693.0000 ;
      RECT 0.0000 1690.4200 5.7000 1691.3600 ;
      RECT 3384.5000 1690.2800 3390.2000 1691.3600 ;
      RECT 9.3000 1690.2800 3380.9000 1691.3600 ;
      RECT 1.1000 1690.2800 5.7000 1690.4200 ;
      RECT 1.1000 1689.5200 3390.2000 1690.2800 ;
      RECT 0.0000 1688.6400 3390.2000 1689.5200 ;
      RECT 3388.5000 1687.5600 3390.2000 1688.6400 ;
      RECT 5.3000 1687.5600 3384.9000 1688.6400 ;
      RECT 0.0000 1687.5600 1.7000 1688.6400 ;
      RECT 0.0000 1685.9200 3390.2000 1687.5600 ;
      RECT 3384.5000 1684.8400 3390.2000 1685.9200 ;
      RECT 9.3000 1684.8400 3380.9000 1685.9200 ;
      RECT 0.0000 1684.8400 5.7000 1685.9200 ;
      RECT 0.0000 1683.2000 3390.2000 1684.8400 ;
      RECT 3388.5000 1682.1200 3390.2000 1683.2000 ;
      RECT 5.3000 1682.1200 3384.9000 1683.2000 ;
      RECT 0.0000 1682.1200 1.7000 1683.2000 ;
      RECT 0.0000 1680.4800 3390.2000 1682.1200 ;
      RECT 3384.5000 1679.4000 3390.2000 1680.4800 ;
      RECT 9.3000 1679.4000 3380.9000 1680.4800 ;
      RECT 0.0000 1679.4000 5.7000 1680.4800 ;
      RECT 0.0000 1677.7600 3390.2000 1679.4000 ;
      RECT 3388.5000 1676.6800 3390.2000 1677.7600 ;
      RECT 5.3000 1676.6800 3384.9000 1677.7600 ;
      RECT 0.0000 1676.6800 1.7000 1677.7600 ;
      RECT 0.0000 1675.0400 3390.2000 1676.6800 ;
      RECT 3384.5000 1673.9600 3390.2000 1675.0400 ;
      RECT 9.3000 1673.9600 3380.9000 1675.0400 ;
      RECT 0.0000 1673.9600 5.7000 1675.0400 ;
      RECT 0.0000 1672.3200 3390.2000 1673.9600 ;
      RECT 3388.5000 1671.2400 3390.2000 1672.3200 ;
      RECT 5.3000 1671.2400 3384.9000 1672.3200 ;
      RECT 0.0000 1671.2400 1.7000 1672.3200 ;
      RECT 0.0000 1669.6000 3390.2000 1671.2400 ;
      RECT 3384.5000 1668.5200 3390.2000 1669.6000 ;
      RECT 9.3000 1668.5200 3380.9000 1669.6000 ;
      RECT 0.0000 1668.5200 5.7000 1669.6000 ;
      RECT 0.0000 1666.8800 3390.2000 1668.5200 ;
      RECT 3388.5000 1665.8000 3390.2000 1666.8800 ;
      RECT 5.3000 1665.8000 3384.9000 1666.8800 ;
      RECT 0.0000 1665.8000 1.7000 1666.8800 ;
      RECT 0.0000 1665.4100 3390.2000 1665.8000 ;
      RECT 1.1000 1664.5100 3390.2000 1665.4100 ;
      RECT 0.0000 1664.1600 3390.2000 1664.5100 ;
      RECT 3384.5000 1663.0800 3390.2000 1664.1600 ;
      RECT 9.3000 1663.0800 3380.9000 1664.1600 ;
      RECT 0.0000 1663.0800 5.7000 1664.1600 ;
      RECT 0.0000 1661.4400 3390.2000 1663.0800 ;
      RECT 3388.5000 1660.3600 3390.2000 1661.4400 ;
      RECT 5.3000 1660.3600 3384.9000 1661.4400 ;
      RECT 0.0000 1660.3600 1.7000 1661.4400 ;
      RECT 0.0000 1658.7200 3390.2000 1660.3600 ;
      RECT 3384.5000 1658.0900 3390.2000 1658.7200 ;
      RECT 3384.5000 1657.6400 3389.1000 1658.0900 ;
      RECT 9.3000 1657.6400 3380.9000 1658.7200 ;
      RECT 0.0000 1657.6400 5.7000 1658.7200 ;
      RECT 0.0000 1657.1900 3389.1000 1657.6400 ;
      RECT 0.0000 1656.0000 3390.2000 1657.1900 ;
      RECT 3388.5000 1654.9200 3390.2000 1656.0000 ;
      RECT 5.3000 1654.9200 3384.9000 1656.0000 ;
      RECT 0.0000 1654.9200 1.7000 1656.0000 ;
      RECT 0.0000 1653.2800 3390.2000 1654.9200 ;
      RECT 3384.5000 1652.2000 3390.2000 1653.2800 ;
      RECT 9.3000 1652.2000 3380.9000 1653.2800 ;
      RECT 0.0000 1652.2000 5.7000 1653.2800 ;
      RECT 0.0000 1650.5600 3390.2000 1652.2000 ;
      RECT 3388.5000 1649.4800 3390.2000 1650.5600 ;
      RECT 5.3000 1649.4800 3384.9000 1650.5600 ;
      RECT 0.0000 1649.4800 1.7000 1650.5600 ;
      RECT 0.0000 1647.8400 3390.2000 1649.4800 ;
      RECT 3384.5000 1646.7600 3390.2000 1647.8400 ;
      RECT 9.3000 1646.7600 3380.9000 1647.8400 ;
      RECT 0.0000 1646.7600 5.7000 1647.8400 ;
      RECT 0.0000 1645.1200 3390.2000 1646.7600 ;
      RECT 3388.5000 1644.0400 3390.2000 1645.1200 ;
      RECT 5.3000 1644.0400 3384.9000 1645.1200 ;
      RECT 0.0000 1644.0400 1.7000 1645.1200 ;
      RECT 0.0000 1642.4000 3390.2000 1644.0400 ;
      RECT 3384.5000 1641.3200 3390.2000 1642.4000 ;
      RECT 9.3000 1641.3200 3380.9000 1642.4000 ;
      RECT 0.0000 1641.3200 5.7000 1642.4000 ;
      RECT 0.0000 1639.7900 3390.2000 1641.3200 ;
      RECT 1.1000 1639.6800 3390.2000 1639.7900 ;
      RECT 1.1000 1638.8900 1.7000 1639.6800 ;
      RECT 3388.5000 1638.6000 3390.2000 1639.6800 ;
      RECT 5.3000 1638.6000 3384.9000 1639.6800 ;
      RECT 0.0000 1638.6000 1.7000 1638.8900 ;
      RECT 0.0000 1636.9600 3390.2000 1638.6000 ;
      RECT 3384.5000 1635.8800 3390.2000 1636.9600 ;
      RECT 9.3000 1635.8800 3380.9000 1636.9600 ;
      RECT 0.0000 1635.8800 5.7000 1636.9600 ;
      RECT 0.0000 1634.2400 3390.2000 1635.8800 ;
      RECT 3388.5000 1633.1600 3390.2000 1634.2400 ;
      RECT 5.3000 1633.1600 3384.9000 1634.2400 ;
      RECT 0.0000 1633.1600 1.7000 1634.2400 ;
      RECT 0.0000 1631.5200 3390.2000 1633.1600 ;
      RECT 3384.5000 1630.4400 3390.2000 1631.5200 ;
      RECT 9.3000 1630.4400 3380.9000 1631.5200 ;
      RECT 0.0000 1630.4400 5.7000 1631.5200 ;
      RECT 0.0000 1628.8000 3390.2000 1630.4400 ;
      RECT 3388.5000 1627.7200 3390.2000 1628.8000 ;
      RECT 5.3000 1627.7200 3384.9000 1628.8000 ;
      RECT 0.0000 1627.7200 1.7000 1628.8000 ;
      RECT 0.0000 1626.0800 3390.2000 1627.7200 ;
      RECT 3384.5000 1625.0000 3390.2000 1626.0800 ;
      RECT 9.3000 1625.0000 3380.9000 1626.0800 ;
      RECT 0.0000 1625.0000 5.7000 1626.0800 ;
      RECT 0.0000 1623.3600 3390.2000 1625.0000 ;
      RECT 3388.5000 1622.2800 3390.2000 1623.3600 ;
      RECT 5.3000 1622.2800 3384.9000 1623.3600 ;
      RECT 0.0000 1622.2800 1.7000 1623.3600 ;
      RECT 0.0000 1620.6400 3390.2000 1622.2800 ;
      RECT 3384.5000 1619.5600 3390.2000 1620.6400 ;
      RECT 9.3000 1619.5600 3380.9000 1620.6400 ;
      RECT 0.0000 1619.5600 5.7000 1620.6400 ;
      RECT 0.0000 1617.9200 3390.2000 1619.5600 ;
      RECT 3388.5000 1616.8400 3390.2000 1617.9200 ;
      RECT 5.3000 1616.8400 3384.9000 1617.9200 ;
      RECT 0.0000 1616.8400 1.7000 1617.9200 ;
      RECT 0.0000 1615.2000 3390.2000 1616.8400 ;
      RECT 0.0000 1614.7800 5.7000 1615.2000 ;
      RECT 3384.5000 1614.1200 3390.2000 1615.2000 ;
      RECT 9.3000 1614.1200 3380.9000 1615.2000 ;
      RECT 1.1000 1614.1200 5.7000 1614.7800 ;
      RECT 1.1000 1613.8800 3390.2000 1614.1200 ;
      RECT 0.0000 1612.4800 3390.2000 1613.8800 ;
      RECT 3388.5000 1611.4000 3390.2000 1612.4800 ;
      RECT 5.3000 1611.4000 3384.9000 1612.4800 ;
      RECT 0.0000 1611.4000 1.7000 1612.4800 ;
      RECT 0.0000 1609.7600 3390.2000 1611.4000 ;
      RECT 3384.5000 1608.6800 3390.2000 1609.7600 ;
      RECT 9.3000 1608.6800 3380.9000 1609.7600 ;
      RECT 0.0000 1608.6800 5.7000 1609.7600 ;
      RECT 0.0000 1607.0400 3390.2000 1608.6800 ;
      RECT 3388.5000 1605.9600 3390.2000 1607.0400 ;
      RECT 5.3000 1605.9600 3384.9000 1607.0400 ;
      RECT 0.0000 1605.9600 1.7000 1607.0400 ;
      RECT 0.0000 1604.3200 3390.2000 1605.9600 ;
      RECT 3384.5000 1603.2400 3390.2000 1604.3200 ;
      RECT 9.3000 1603.2400 3380.9000 1604.3200 ;
      RECT 0.0000 1603.2400 5.7000 1604.3200 ;
      RECT 0.0000 1601.6000 3390.2000 1603.2400 ;
      RECT 3388.5000 1600.5200 3390.2000 1601.6000 ;
      RECT 5.3000 1600.5200 3384.9000 1601.6000 ;
      RECT 0.0000 1600.5200 1.7000 1601.6000 ;
      RECT 0.0000 1598.8800 3390.2000 1600.5200 ;
      RECT 3384.5000 1597.8000 3390.2000 1598.8800 ;
      RECT 9.3000 1597.8000 3380.9000 1598.8800 ;
      RECT 0.0000 1597.8000 5.7000 1598.8800 ;
      RECT 0.0000 1596.1600 3390.2000 1597.8000 ;
      RECT 3388.5000 1595.0800 3390.2000 1596.1600 ;
      RECT 5.3000 1595.0800 3384.9000 1596.1600 ;
      RECT 0.0000 1595.0800 1.7000 1596.1600 ;
      RECT 0.0000 1593.4400 3390.2000 1595.0800 ;
      RECT 3384.5000 1592.3600 3390.2000 1593.4400 ;
      RECT 9.3000 1592.3600 3380.9000 1593.4400 ;
      RECT 0.0000 1592.3600 5.7000 1593.4400 ;
      RECT 0.0000 1590.7200 3390.2000 1592.3600 ;
      RECT 3388.5000 1589.6400 3390.2000 1590.7200 ;
      RECT 5.3000 1589.6400 3384.9000 1590.7200 ;
      RECT 0.0000 1589.6400 1.7000 1590.7200 ;
      RECT 0.0000 1589.1600 3390.2000 1589.6400 ;
      RECT 1.1000 1588.2600 3390.2000 1589.1600 ;
      RECT 0.0000 1588.0000 3390.2000 1588.2600 ;
      RECT 3384.5000 1586.9200 3390.2000 1588.0000 ;
      RECT 9.3000 1586.9200 3380.9000 1588.0000 ;
      RECT 0.0000 1586.9200 5.7000 1588.0000 ;
      RECT 0.0000 1585.2800 3390.2000 1586.9200 ;
      RECT 3388.5000 1584.2000 3390.2000 1585.2800 ;
      RECT 5.3000 1584.2000 3384.9000 1585.2800 ;
      RECT 0.0000 1584.2000 1.7000 1585.2800 ;
      RECT 0.0000 1582.5600 3390.2000 1584.2000 ;
      RECT 3384.5000 1581.4800 3390.2000 1582.5600 ;
      RECT 9.3000 1581.4800 3380.9000 1582.5600 ;
      RECT 0.0000 1581.4800 5.7000 1582.5600 ;
      RECT 0.0000 1579.8400 3390.2000 1581.4800 ;
      RECT 3388.5000 1578.7600 3390.2000 1579.8400 ;
      RECT 5.3000 1578.7600 3384.9000 1579.8400 ;
      RECT 0.0000 1578.7600 1.7000 1579.8400 ;
      RECT 0.0000 1577.1200 3390.2000 1578.7600 ;
      RECT 3384.5000 1576.0400 3390.2000 1577.1200 ;
      RECT 9.3000 1576.0400 3380.9000 1577.1200 ;
      RECT 0.0000 1576.0400 5.7000 1577.1200 ;
      RECT 0.0000 1574.4000 3390.2000 1576.0400 ;
      RECT 3388.5000 1573.3200 3390.2000 1574.4000 ;
      RECT 5.3000 1573.3200 3384.9000 1574.4000 ;
      RECT 0.0000 1573.3200 1.7000 1574.4000 ;
      RECT 0.0000 1571.6800 3390.2000 1573.3200 ;
      RECT 3384.5000 1570.6000 3390.2000 1571.6800 ;
      RECT 9.3000 1570.6000 3380.9000 1571.6800 ;
      RECT 0.0000 1570.6000 5.7000 1571.6800 ;
      RECT 0.0000 1568.9600 3390.2000 1570.6000 ;
      RECT 3388.5000 1567.8800 3390.2000 1568.9600 ;
      RECT 5.3000 1567.8800 3384.9000 1568.9600 ;
      RECT 0.0000 1567.8800 1.7000 1568.9600 ;
      RECT 0.0000 1566.2400 3390.2000 1567.8800 ;
      RECT 3384.5000 1565.1600 3390.2000 1566.2400 ;
      RECT 9.3000 1565.1600 3380.9000 1566.2400 ;
      RECT 0.0000 1565.1600 5.7000 1566.2400 ;
      RECT 0.0000 1564.1500 3390.2000 1565.1600 ;
      RECT 1.1000 1563.5200 3390.2000 1564.1500 ;
      RECT 1.1000 1563.2500 1.7000 1563.5200 ;
      RECT 3388.5000 1562.4400 3390.2000 1563.5200 ;
      RECT 5.3000 1562.4400 3384.9000 1563.5200 ;
      RECT 0.0000 1562.4400 1.7000 1563.2500 ;
      RECT 0.0000 1560.8000 3390.2000 1562.4400 ;
      RECT 3384.5000 1559.7200 3390.2000 1560.8000 ;
      RECT 9.3000 1559.7200 3380.9000 1560.8000 ;
      RECT 0.0000 1559.7200 5.7000 1560.8000 ;
      RECT 0.0000 1558.0800 3390.2000 1559.7200 ;
      RECT 3388.5000 1557.0000 3390.2000 1558.0800 ;
      RECT 5.3000 1557.0000 3384.9000 1558.0800 ;
      RECT 0.0000 1557.0000 1.7000 1558.0800 ;
      RECT 0.0000 1555.3600 3390.2000 1557.0000 ;
      RECT 3384.5000 1554.3900 3390.2000 1555.3600 ;
      RECT 3384.5000 1554.2800 3389.1000 1554.3900 ;
      RECT 9.3000 1554.2800 3380.9000 1555.3600 ;
      RECT 0.0000 1554.2800 5.7000 1555.3600 ;
      RECT 0.0000 1553.4900 3389.1000 1554.2800 ;
      RECT 0.0000 1552.6400 3390.2000 1553.4900 ;
      RECT 3388.5000 1551.5600 3390.2000 1552.6400 ;
      RECT 5.3000 1551.5600 3384.9000 1552.6400 ;
      RECT 0.0000 1551.5600 1.7000 1552.6400 ;
      RECT 0.0000 1549.9200 3390.2000 1551.5600 ;
      RECT 3384.5000 1548.8400 3390.2000 1549.9200 ;
      RECT 9.3000 1548.8400 3380.9000 1549.9200 ;
      RECT 0.0000 1548.8400 5.7000 1549.9200 ;
      RECT 0.0000 1547.2000 3390.2000 1548.8400 ;
      RECT 3388.5000 1546.1200 3390.2000 1547.2000 ;
      RECT 5.3000 1546.1200 3384.9000 1547.2000 ;
      RECT 0.0000 1546.1200 1.7000 1547.2000 ;
      RECT 0.0000 1544.4800 3390.2000 1546.1200 ;
      RECT 3384.5000 1543.4000 3390.2000 1544.4800 ;
      RECT 9.3000 1543.4000 3380.9000 1544.4800 ;
      RECT 0.0000 1543.4000 5.7000 1544.4800 ;
      RECT 0.0000 1541.7600 3390.2000 1543.4000 ;
      RECT 3388.5000 1540.6800 3390.2000 1541.7600 ;
      RECT 5.3000 1540.6800 3384.9000 1541.7600 ;
      RECT 0.0000 1540.6800 1.7000 1541.7600 ;
      RECT 0.0000 1539.1400 3390.2000 1540.6800 ;
      RECT 1.1000 1539.0400 3390.2000 1539.1400 ;
      RECT 1.1000 1538.2400 5.7000 1539.0400 ;
      RECT 3384.5000 1537.9600 3390.2000 1539.0400 ;
      RECT 9.3000 1537.9600 3380.9000 1539.0400 ;
      RECT 0.0000 1537.9600 5.7000 1538.2400 ;
      RECT 0.0000 1536.3200 3390.2000 1537.9600 ;
      RECT 3388.5000 1535.2400 3390.2000 1536.3200 ;
      RECT 5.3000 1535.2400 3384.9000 1536.3200 ;
      RECT 0.0000 1535.2400 1.7000 1536.3200 ;
      RECT 0.0000 1533.6000 3390.2000 1535.2400 ;
      RECT 3384.5000 1532.5200 3390.2000 1533.6000 ;
      RECT 9.3000 1532.5200 3380.9000 1533.6000 ;
      RECT 0.0000 1532.5200 5.7000 1533.6000 ;
      RECT 0.0000 1530.8800 3390.2000 1532.5200 ;
      RECT 3388.5000 1529.8000 3390.2000 1530.8800 ;
      RECT 5.3000 1529.8000 3384.9000 1530.8800 ;
      RECT 0.0000 1529.8000 1.7000 1530.8800 ;
      RECT 0.0000 1528.1600 3390.2000 1529.8000 ;
      RECT 3384.5000 1527.0800 3390.2000 1528.1600 ;
      RECT 9.3000 1527.0800 3380.9000 1528.1600 ;
      RECT 0.0000 1527.0800 5.7000 1528.1600 ;
      RECT 0.0000 1525.4400 3390.2000 1527.0800 ;
      RECT 3388.5000 1524.3600 3390.2000 1525.4400 ;
      RECT 5.3000 1524.3600 3384.9000 1525.4400 ;
      RECT 0.0000 1524.3600 1.7000 1525.4400 ;
      RECT 0.0000 1522.7200 3390.2000 1524.3600 ;
      RECT 3384.5000 1521.6400 3390.2000 1522.7200 ;
      RECT 9.3000 1521.6400 3380.9000 1522.7200 ;
      RECT 0.0000 1521.6400 5.7000 1522.7200 ;
      RECT 0.0000 1520.0000 3390.2000 1521.6400 ;
      RECT 3388.5000 1518.9200 3390.2000 1520.0000 ;
      RECT 5.3000 1518.9200 3384.9000 1520.0000 ;
      RECT 0.0000 1518.9200 1.7000 1520.0000 ;
      RECT 0.0000 1517.2800 3390.2000 1518.9200 ;
      RECT 3384.5000 1516.2000 3390.2000 1517.2800 ;
      RECT 9.3000 1516.2000 3380.9000 1517.2800 ;
      RECT 0.0000 1516.2000 5.7000 1517.2800 ;
      RECT 0.0000 1514.5600 3390.2000 1516.2000 ;
      RECT 0.0000 1513.5200 1.7000 1514.5600 ;
      RECT 3388.5000 1513.4800 3390.2000 1514.5600 ;
      RECT 5.3000 1513.4800 3384.9000 1514.5600 ;
      RECT 1.1000 1513.4800 1.7000 1513.5200 ;
      RECT 1.1000 1512.6200 3390.2000 1513.4800 ;
      RECT 0.0000 1511.8400 3390.2000 1512.6200 ;
      RECT 3384.5000 1510.7600 3390.2000 1511.8400 ;
      RECT 9.3000 1510.7600 3380.9000 1511.8400 ;
      RECT 0.0000 1510.7600 5.7000 1511.8400 ;
      RECT 0.0000 1509.1200 3390.2000 1510.7600 ;
      RECT 3388.5000 1508.0400 3390.2000 1509.1200 ;
      RECT 5.3000 1508.0400 3384.9000 1509.1200 ;
      RECT 0.0000 1508.0400 1.7000 1509.1200 ;
      RECT 0.0000 1506.4000 3390.2000 1508.0400 ;
      RECT 3384.5000 1505.3200 3390.2000 1506.4000 ;
      RECT 9.3000 1505.3200 3380.9000 1506.4000 ;
      RECT 0.0000 1505.3200 5.7000 1506.4000 ;
      RECT 0.0000 1503.6800 3390.2000 1505.3200 ;
      RECT 3388.5000 1502.6000 3390.2000 1503.6800 ;
      RECT 5.3000 1502.6000 3384.9000 1503.6800 ;
      RECT 0.0000 1502.6000 1.7000 1503.6800 ;
      RECT 0.0000 1500.9600 3390.2000 1502.6000 ;
      RECT 3384.5000 1499.8800 3390.2000 1500.9600 ;
      RECT 9.3000 1499.8800 3380.9000 1500.9600 ;
      RECT 0.0000 1499.8800 5.7000 1500.9600 ;
      RECT 0.0000 1498.2400 3390.2000 1499.8800 ;
      RECT 3388.5000 1497.1600 3390.2000 1498.2400 ;
      RECT 5.3000 1497.1600 3384.9000 1498.2400 ;
      RECT 0.0000 1497.1600 1.7000 1498.2400 ;
      RECT 0.0000 1495.5200 3390.2000 1497.1600 ;
      RECT 3384.5000 1494.4400 3390.2000 1495.5200 ;
      RECT 9.3000 1494.4400 3380.9000 1495.5200 ;
      RECT 0.0000 1494.4400 5.7000 1495.5200 ;
      RECT 0.0000 1492.8000 3390.2000 1494.4400 ;
      RECT 3388.5000 1491.7200 3390.2000 1492.8000 ;
      RECT 5.3000 1491.7200 3384.9000 1492.8000 ;
      RECT 0.0000 1491.7200 1.7000 1492.8000 ;
      RECT 0.0000 1490.0800 3390.2000 1491.7200 ;
      RECT 3384.5000 1489.0000 3390.2000 1490.0800 ;
      RECT 9.3000 1489.0000 3380.9000 1490.0800 ;
      RECT 0.0000 1489.0000 5.7000 1490.0800 ;
      RECT 0.0000 1488.5100 3390.2000 1489.0000 ;
      RECT 1.1000 1487.6100 3390.2000 1488.5100 ;
      RECT 0.0000 1487.3600 3390.2000 1487.6100 ;
      RECT 3388.5000 1486.2800 3390.2000 1487.3600 ;
      RECT 5.3000 1486.2800 3384.9000 1487.3600 ;
      RECT 0.0000 1486.2800 1.7000 1487.3600 ;
      RECT 0.0000 1484.6400 3390.2000 1486.2800 ;
      RECT 3384.5000 1483.5600 3390.2000 1484.6400 ;
      RECT 9.3000 1483.5600 3380.9000 1484.6400 ;
      RECT 0.0000 1483.5600 5.7000 1484.6400 ;
      RECT 0.0000 1481.9200 3390.2000 1483.5600 ;
      RECT 3388.5000 1480.8400 3390.2000 1481.9200 ;
      RECT 5.3000 1480.8400 3384.9000 1481.9200 ;
      RECT 0.0000 1480.8400 1.7000 1481.9200 ;
      RECT 0.0000 1479.2000 3390.2000 1480.8400 ;
      RECT 3384.5000 1478.1200 3390.2000 1479.2000 ;
      RECT 9.3000 1478.1200 3380.9000 1479.2000 ;
      RECT 0.0000 1478.1200 5.7000 1479.2000 ;
      RECT 0.0000 1476.4800 3390.2000 1478.1200 ;
      RECT 3388.5000 1475.4000 3390.2000 1476.4800 ;
      RECT 5.3000 1475.4000 3384.9000 1476.4800 ;
      RECT 0.0000 1475.4000 1.7000 1476.4800 ;
      RECT 0.0000 1473.7600 3390.2000 1475.4000 ;
      RECT 3384.5000 1472.6800 3390.2000 1473.7600 ;
      RECT 9.3000 1472.6800 3380.9000 1473.7600 ;
      RECT 0.0000 1472.6800 5.7000 1473.7600 ;
      RECT 0.0000 1471.0400 3390.2000 1472.6800 ;
      RECT 3388.5000 1469.9600 3390.2000 1471.0400 ;
      RECT 5.3000 1469.9600 3384.9000 1471.0400 ;
      RECT 0.0000 1469.9600 1.7000 1471.0400 ;
      RECT 0.0000 1468.3200 3390.2000 1469.9600 ;
      RECT 3384.5000 1467.2400 3390.2000 1468.3200 ;
      RECT 9.3000 1467.2400 3380.9000 1468.3200 ;
      RECT 0.0000 1467.2400 5.7000 1468.3200 ;
      RECT 0.0000 1465.6000 3390.2000 1467.2400 ;
      RECT 3388.5000 1464.5200 3390.2000 1465.6000 ;
      RECT 5.3000 1464.5200 3384.9000 1465.6000 ;
      RECT 0.0000 1464.5200 1.7000 1465.6000 ;
      RECT 0.0000 1463.5000 3390.2000 1464.5200 ;
      RECT 1.1000 1462.8800 3390.2000 1463.5000 ;
      RECT 1.1000 1462.6000 5.7000 1462.8800 ;
      RECT 3384.5000 1461.8000 3390.2000 1462.8800 ;
      RECT 9.3000 1461.8000 3380.9000 1462.8800 ;
      RECT 0.0000 1461.8000 5.7000 1462.6000 ;
      RECT 0.0000 1460.1600 3390.2000 1461.8000 ;
      RECT 3388.5000 1459.0800 3390.2000 1460.1600 ;
      RECT 5.3000 1459.0800 3384.9000 1460.1600 ;
      RECT 0.0000 1459.0800 1.7000 1460.1600 ;
      RECT 0.0000 1457.4400 3390.2000 1459.0800 ;
      RECT 3384.5000 1456.3600 3390.2000 1457.4400 ;
      RECT 9.3000 1456.3600 3380.9000 1457.4400 ;
      RECT 0.0000 1456.3600 5.7000 1457.4400 ;
      RECT 0.0000 1454.7200 3390.2000 1456.3600 ;
      RECT 3388.5000 1453.6400 3390.2000 1454.7200 ;
      RECT 5.3000 1453.6400 3384.9000 1454.7200 ;
      RECT 0.0000 1453.6400 1.7000 1454.7200 ;
      RECT 0.0000 1452.0000 3390.2000 1453.6400 ;
      RECT 3384.5000 1450.9200 3390.2000 1452.0000 ;
      RECT 9.3000 1450.9200 3380.9000 1452.0000 ;
      RECT 0.0000 1450.9200 5.7000 1452.0000 ;
      RECT 0.0000 1450.6900 3390.2000 1450.9200 ;
      RECT 0.0000 1449.7900 3389.1000 1450.6900 ;
      RECT 0.0000 1449.2800 3390.2000 1449.7900 ;
      RECT 3388.5000 1448.2000 3390.2000 1449.2800 ;
      RECT 5.3000 1448.2000 3384.9000 1449.2800 ;
      RECT 0.0000 1448.2000 1.7000 1449.2800 ;
      RECT 0.0000 1446.5600 3390.2000 1448.2000 ;
      RECT 3384.5000 1445.4800 3390.2000 1446.5600 ;
      RECT 9.3000 1445.4800 3380.9000 1446.5600 ;
      RECT 0.0000 1445.4800 5.7000 1446.5600 ;
      RECT 0.0000 1443.8400 3390.2000 1445.4800 ;
      RECT 3388.5000 1442.7600 3390.2000 1443.8400 ;
      RECT 5.3000 1442.7600 3384.9000 1443.8400 ;
      RECT 0.0000 1442.7600 1.7000 1443.8400 ;
      RECT 0.0000 1441.1200 3390.2000 1442.7600 ;
      RECT 3384.5000 1440.0400 3390.2000 1441.1200 ;
      RECT 9.3000 1440.0400 3380.9000 1441.1200 ;
      RECT 0.0000 1440.0400 5.7000 1441.1200 ;
      RECT 0.0000 1438.4000 3390.2000 1440.0400 ;
      RECT 0.0000 1437.8800 1.7000 1438.4000 ;
      RECT 3388.5000 1437.3200 3390.2000 1438.4000 ;
      RECT 5.3000 1437.3200 3384.9000 1438.4000 ;
      RECT 1.1000 1437.3200 1.7000 1437.8800 ;
      RECT 1.1000 1436.9800 3390.2000 1437.3200 ;
      RECT 0.0000 1435.6800 3390.2000 1436.9800 ;
      RECT 3384.5000 1434.6000 3390.2000 1435.6800 ;
      RECT 9.3000 1434.6000 3380.9000 1435.6800 ;
      RECT 0.0000 1434.6000 5.7000 1435.6800 ;
      RECT 0.0000 1432.9600 3390.2000 1434.6000 ;
      RECT 3388.5000 1431.8800 3390.2000 1432.9600 ;
      RECT 5.3000 1431.8800 3384.9000 1432.9600 ;
      RECT 0.0000 1431.8800 1.7000 1432.9600 ;
      RECT 0.0000 1430.2400 3390.2000 1431.8800 ;
      RECT 3384.5000 1429.1600 3390.2000 1430.2400 ;
      RECT 9.3000 1429.1600 3380.9000 1430.2400 ;
      RECT 0.0000 1429.1600 5.7000 1430.2400 ;
      RECT 0.0000 1427.5200 3390.2000 1429.1600 ;
      RECT 3388.5000 1426.4400 3390.2000 1427.5200 ;
      RECT 5.3000 1426.4400 3384.9000 1427.5200 ;
      RECT 0.0000 1426.4400 1.7000 1427.5200 ;
      RECT 0.0000 1424.8000 3390.2000 1426.4400 ;
      RECT 3384.5000 1423.7200 3390.2000 1424.8000 ;
      RECT 9.3000 1423.7200 3380.9000 1424.8000 ;
      RECT 0.0000 1423.7200 5.7000 1424.8000 ;
      RECT 0.0000 1422.0800 3390.2000 1423.7200 ;
      RECT 3388.5000 1421.0000 3390.2000 1422.0800 ;
      RECT 5.3000 1421.0000 3384.9000 1422.0800 ;
      RECT 0.0000 1421.0000 1.7000 1422.0800 ;
      RECT 0.0000 1419.3600 3390.2000 1421.0000 ;
      RECT 3384.5000 1418.2800 3390.2000 1419.3600 ;
      RECT 9.3000 1418.2800 3380.9000 1419.3600 ;
      RECT 0.0000 1418.2800 5.7000 1419.3600 ;
      RECT 0.0000 1416.6400 3390.2000 1418.2800 ;
      RECT 3388.5000 1415.5600 3390.2000 1416.6400 ;
      RECT 5.3000 1415.5600 3384.9000 1416.6400 ;
      RECT 0.0000 1415.5600 1.7000 1416.6400 ;
      RECT 0.0000 1413.9200 3390.2000 1415.5600 ;
      RECT 0.0000 1412.8700 5.7000 1413.9200 ;
      RECT 3384.5000 1412.8400 3390.2000 1413.9200 ;
      RECT 9.3000 1412.8400 3380.9000 1413.9200 ;
      RECT 1.1000 1412.8400 5.7000 1412.8700 ;
      RECT 1.1000 1411.9700 3390.2000 1412.8400 ;
      RECT 0.0000 1411.2000 3390.2000 1411.9700 ;
      RECT 3388.5000 1410.1200 3390.2000 1411.2000 ;
      RECT 5.3000 1410.1200 3384.9000 1411.2000 ;
      RECT 0.0000 1410.1200 1.7000 1411.2000 ;
      RECT 0.0000 1408.4800 3390.2000 1410.1200 ;
      RECT 3384.5000 1407.4000 3390.2000 1408.4800 ;
      RECT 9.3000 1407.4000 3380.9000 1408.4800 ;
      RECT 0.0000 1407.4000 5.7000 1408.4800 ;
      RECT 0.0000 1405.7600 3390.2000 1407.4000 ;
      RECT 3388.5000 1404.6800 3390.2000 1405.7600 ;
      RECT 5.3000 1404.6800 3384.9000 1405.7600 ;
      RECT 0.0000 1404.6800 1.7000 1405.7600 ;
      RECT 0.0000 1403.0400 3390.2000 1404.6800 ;
      RECT 3384.5000 1401.9600 3390.2000 1403.0400 ;
      RECT 9.3000 1401.9600 3380.9000 1403.0400 ;
      RECT 0.0000 1401.9600 5.7000 1403.0400 ;
      RECT 0.0000 1400.3200 3390.2000 1401.9600 ;
      RECT 3388.5000 1399.2400 3390.2000 1400.3200 ;
      RECT 5.3000 1399.2400 3384.9000 1400.3200 ;
      RECT 0.0000 1399.2400 1.7000 1400.3200 ;
      RECT 0.0000 1397.6000 3390.2000 1399.2400 ;
      RECT 3384.5000 1396.5200 3390.2000 1397.6000 ;
      RECT 9.3000 1396.5200 3380.9000 1397.6000 ;
      RECT 0.0000 1396.5200 5.7000 1397.6000 ;
      RECT 0.0000 1394.8800 3390.2000 1396.5200 ;
      RECT 3388.5000 1393.8000 3390.2000 1394.8800 ;
      RECT 5.3000 1393.8000 3384.9000 1394.8800 ;
      RECT 0.0000 1393.8000 1.7000 1394.8800 ;
      RECT 0.0000 1392.1600 3390.2000 1393.8000 ;
      RECT 3384.5000 1391.0800 3390.2000 1392.1600 ;
      RECT 9.3000 1391.0800 3380.9000 1392.1600 ;
      RECT 0.0000 1391.0800 5.7000 1392.1600 ;
      RECT 0.0000 1389.4400 3390.2000 1391.0800 ;
      RECT 3388.5000 1388.3600 3390.2000 1389.4400 ;
      RECT 5.3000 1388.3600 3384.9000 1389.4400 ;
      RECT 0.0000 1388.3600 1.7000 1389.4400 ;
      RECT 0.0000 1387.8600 3390.2000 1388.3600 ;
      RECT 1.1000 1386.9600 3390.2000 1387.8600 ;
      RECT 0.0000 1386.7200 3390.2000 1386.9600 ;
      RECT 3384.5000 1385.6400 3390.2000 1386.7200 ;
      RECT 9.3000 1385.6400 3380.9000 1386.7200 ;
      RECT 0.0000 1385.6400 5.7000 1386.7200 ;
      RECT 0.0000 1384.0000 3390.2000 1385.6400 ;
      RECT 3388.5000 1382.9200 3390.2000 1384.0000 ;
      RECT 5.3000 1382.9200 3384.9000 1384.0000 ;
      RECT 0.0000 1382.9200 1.7000 1384.0000 ;
      RECT 0.0000 1381.2800 3390.2000 1382.9200 ;
      RECT 3384.5000 1380.2000 3390.2000 1381.2800 ;
      RECT 9.3000 1380.2000 3380.9000 1381.2800 ;
      RECT 0.0000 1380.2000 5.7000 1381.2800 ;
      RECT 0.0000 1378.5600 3390.2000 1380.2000 ;
      RECT 3388.5000 1377.4800 3390.2000 1378.5600 ;
      RECT 5.3000 1377.4800 3384.9000 1378.5600 ;
      RECT 0.0000 1377.4800 1.7000 1378.5600 ;
      RECT 0.0000 1375.8400 3390.2000 1377.4800 ;
      RECT 3384.5000 1374.7600 3390.2000 1375.8400 ;
      RECT 9.3000 1374.7600 3380.9000 1375.8400 ;
      RECT 0.0000 1374.7600 5.7000 1375.8400 ;
      RECT 0.0000 1373.1200 3390.2000 1374.7600 ;
      RECT 3388.5000 1372.0400 3390.2000 1373.1200 ;
      RECT 5.3000 1372.0400 3384.9000 1373.1200 ;
      RECT 0.0000 1372.0400 1.7000 1373.1200 ;
      RECT 0.0000 1370.4000 3390.2000 1372.0400 ;
      RECT 3384.5000 1369.3200 3390.2000 1370.4000 ;
      RECT 9.3000 1369.3200 3380.9000 1370.4000 ;
      RECT 0.0000 1369.3200 5.7000 1370.4000 ;
      RECT 0.0000 1367.6800 3390.2000 1369.3200 ;
      RECT 3388.5000 1366.6000 3390.2000 1367.6800 ;
      RECT 5.3000 1366.6000 3384.9000 1367.6800 ;
      RECT 0.0000 1366.6000 1.7000 1367.6800 ;
      RECT 0.0000 1364.9600 3390.2000 1366.6000 ;
      RECT 3384.5000 1363.8800 3390.2000 1364.9600 ;
      RECT 9.3000 1363.8800 3380.9000 1364.9600 ;
      RECT 0.0000 1363.8800 5.7000 1364.9600 ;
      RECT 0.0000 1362.2400 3390.2000 1363.8800 ;
      RECT 1.1000 1361.3400 1.7000 1362.2400 ;
      RECT 3388.5000 1361.1600 3390.2000 1362.2400 ;
      RECT 5.3000 1361.1600 3384.9000 1362.2400 ;
      RECT 0.0000 1361.1600 1.7000 1361.3400 ;
      RECT 0.0000 1359.5200 3390.2000 1361.1600 ;
      RECT 3384.5000 1358.4400 3390.2000 1359.5200 ;
      RECT 9.3000 1358.4400 3380.9000 1359.5200 ;
      RECT 0.0000 1358.4400 5.7000 1359.5200 ;
      RECT 0.0000 1356.8000 3390.2000 1358.4400 ;
      RECT 3388.5000 1355.7200 3390.2000 1356.8000 ;
      RECT 5.3000 1355.7200 3384.9000 1356.8000 ;
      RECT 0.0000 1355.7200 1.7000 1356.8000 ;
      RECT 0.0000 1354.0800 3390.2000 1355.7200 ;
      RECT 3384.5000 1353.0000 3390.2000 1354.0800 ;
      RECT 9.3000 1353.0000 3380.9000 1354.0800 ;
      RECT 0.0000 1353.0000 5.7000 1354.0800 ;
      RECT 0.0000 1351.3600 3390.2000 1353.0000 ;
      RECT 3388.5000 1350.2800 3390.2000 1351.3600 ;
      RECT 5.3000 1350.2800 3384.9000 1351.3600 ;
      RECT 0.0000 1350.2800 1.7000 1351.3600 ;
      RECT 0.0000 1348.6400 3390.2000 1350.2800 ;
      RECT 3384.5000 1347.5600 3390.2000 1348.6400 ;
      RECT 9.3000 1347.5600 3380.9000 1348.6400 ;
      RECT 0.0000 1347.5600 5.7000 1348.6400 ;
      RECT 0.0000 1346.9900 3390.2000 1347.5600 ;
      RECT 0.0000 1346.0900 3389.1000 1346.9900 ;
      RECT 0.0000 1345.9200 3390.2000 1346.0900 ;
      RECT 3388.5000 1344.8400 3390.2000 1345.9200 ;
      RECT 5.3000 1344.8400 3384.9000 1345.9200 ;
      RECT 0.0000 1344.8400 1.7000 1345.9200 ;
      RECT 0.0000 1343.2000 3390.2000 1344.8400 ;
      RECT 3384.5000 1342.1200 3390.2000 1343.2000 ;
      RECT 9.3000 1342.1200 3380.9000 1343.2000 ;
      RECT 0.0000 1342.1200 5.7000 1343.2000 ;
      RECT 0.0000 1340.4800 3390.2000 1342.1200 ;
      RECT 3388.5000 1339.4000 3390.2000 1340.4800 ;
      RECT 5.3000 1339.4000 3384.9000 1340.4800 ;
      RECT 0.0000 1339.4000 1.7000 1340.4800 ;
      RECT 0.0000 1337.7600 3390.2000 1339.4000 ;
      RECT 0.0000 1337.2300 5.7000 1337.7600 ;
      RECT 3384.5000 1336.6800 3390.2000 1337.7600 ;
      RECT 9.3000 1336.6800 3380.9000 1337.7600 ;
      RECT 1.1000 1336.6800 5.7000 1337.2300 ;
      RECT 1.1000 1336.3300 3390.2000 1336.6800 ;
      RECT 0.0000 1335.0400 3390.2000 1336.3300 ;
      RECT 3388.5000 1333.9600 3390.2000 1335.0400 ;
      RECT 5.3000 1333.9600 3384.9000 1335.0400 ;
      RECT 0.0000 1333.9600 1.7000 1335.0400 ;
      RECT 0.0000 1332.3200 3390.2000 1333.9600 ;
      RECT 3384.5000 1331.2400 3390.2000 1332.3200 ;
      RECT 9.3000 1331.2400 3380.9000 1332.3200 ;
      RECT 0.0000 1331.2400 5.7000 1332.3200 ;
      RECT 0.0000 1329.6000 3390.2000 1331.2400 ;
      RECT 3388.5000 1328.5200 3390.2000 1329.6000 ;
      RECT 5.3000 1328.5200 3384.9000 1329.6000 ;
      RECT 0.0000 1328.5200 1.7000 1329.6000 ;
      RECT 0.0000 1326.8800 3390.2000 1328.5200 ;
      RECT 3384.5000 1325.8000 3390.2000 1326.8800 ;
      RECT 9.3000 1325.8000 3380.9000 1326.8800 ;
      RECT 0.0000 1325.8000 5.7000 1326.8800 ;
      RECT 0.0000 1324.1600 3390.2000 1325.8000 ;
      RECT 3388.5000 1323.0800 3390.2000 1324.1600 ;
      RECT 5.3000 1323.0800 3384.9000 1324.1600 ;
      RECT 0.0000 1323.0800 1.7000 1324.1600 ;
      RECT 0.0000 1321.4400 3390.2000 1323.0800 ;
      RECT 3384.5000 1320.3600 3390.2000 1321.4400 ;
      RECT 9.3000 1320.3600 3380.9000 1321.4400 ;
      RECT 0.0000 1320.3600 5.7000 1321.4400 ;
      RECT 0.0000 1318.7200 3390.2000 1320.3600 ;
      RECT 3388.5000 1317.6400 3390.2000 1318.7200 ;
      RECT 5.3000 1317.6400 3384.9000 1318.7200 ;
      RECT 0.0000 1317.6400 1.7000 1318.7200 ;
      RECT 0.0000 1316.0000 3390.2000 1317.6400 ;
      RECT 3384.5000 1314.9200 3390.2000 1316.0000 ;
      RECT 9.3000 1314.9200 3380.9000 1316.0000 ;
      RECT 0.0000 1314.9200 5.7000 1316.0000 ;
      RECT 0.0000 1313.2800 3390.2000 1314.9200 ;
      RECT 0.0000 1312.2200 1.7000 1313.2800 ;
      RECT 3388.5000 1312.2000 3390.2000 1313.2800 ;
      RECT 5.3000 1312.2000 3384.9000 1313.2800 ;
      RECT 1.1000 1312.2000 1.7000 1312.2200 ;
      RECT 1.1000 1311.3200 3390.2000 1312.2000 ;
      RECT 0.0000 1310.5600 3390.2000 1311.3200 ;
      RECT 3384.5000 1309.4800 3390.2000 1310.5600 ;
      RECT 9.3000 1309.4800 3380.9000 1310.5600 ;
      RECT 0.0000 1309.4800 5.7000 1310.5600 ;
      RECT 0.0000 1307.8400 3390.2000 1309.4800 ;
      RECT 3388.5000 1306.7600 3390.2000 1307.8400 ;
      RECT 5.3000 1306.7600 3384.9000 1307.8400 ;
      RECT 0.0000 1306.7600 1.7000 1307.8400 ;
      RECT 0.0000 1305.1200 3390.2000 1306.7600 ;
      RECT 3384.5000 1304.0400 3390.2000 1305.1200 ;
      RECT 9.3000 1304.0400 3380.9000 1305.1200 ;
      RECT 0.0000 1304.0400 5.7000 1305.1200 ;
      RECT 0.0000 1302.4000 3390.2000 1304.0400 ;
      RECT 3388.5000 1301.3200 3390.2000 1302.4000 ;
      RECT 5.3000 1301.3200 3384.9000 1302.4000 ;
      RECT 0.0000 1301.3200 1.7000 1302.4000 ;
      RECT 0.0000 1299.6800 3390.2000 1301.3200 ;
      RECT 3384.5000 1298.6000 3390.2000 1299.6800 ;
      RECT 9.3000 1298.6000 3380.9000 1299.6800 ;
      RECT 0.0000 1298.6000 5.7000 1299.6800 ;
      RECT 0.0000 1296.9600 3390.2000 1298.6000 ;
      RECT 3388.5000 1295.8800 3390.2000 1296.9600 ;
      RECT 5.3000 1295.8800 3384.9000 1296.9600 ;
      RECT 0.0000 1295.8800 1.7000 1296.9600 ;
      RECT 0.0000 1294.2400 3390.2000 1295.8800 ;
      RECT 3384.5000 1293.1600 3390.2000 1294.2400 ;
      RECT 9.3000 1293.1600 3380.9000 1294.2400 ;
      RECT 0.0000 1293.1600 5.7000 1294.2400 ;
      RECT 0.0000 1291.5200 3390.2000 1293.1600 ;
      RECT 3388.5000 1290.4400 3390.2000 1291.5200 ;
      RECT 5.3000 1290.4400 3384.9000 1291.5200 ;
      RECT 0.0000 1290.4400 1.7000 1291.5200 ;
      RECT 0.0000 1288.8000 3390.2000 1290.4400 ;
      RECT 3384.5000 1287.7200 3390.2000 1288.8000 ;
      RECT 9.3000 1287.7200 3380.9000 1288.8000 ;
      RECT 0.0000 1287.7200 5.7000 1288.8000 ;
      RECT 0.0000 1286.6000 3390.2000 1287.7200 ;
      RECT 1.1000 1286.0800 3390.2000 1286.6000 ;
      RECT 1.1000 1285.7000 1.7000 1286.0800 ;
      RECT 3388.5000 1285.0000 3390.2000 1286.0800 ;
      RECT 5.3000 1285.0000 3384.9000 1286.0800 ;
      RECT 0.0000 1285.0000 1.7000 1285.7000 ;
      RECT 0.0000 1283.3600 3390.2000 1285.0000 ;
      RECT 3384.5000 1282.2800 3390.2000 1283.3600 ;
      RECT 9.3000 1282.2800 3380.9000 1283.3600 ;
      RECT 0.0000 1282.2800 5.7000 1283.3600 ;
      RECT 0.0000 1280.6400 3390.2000 1282.2800 ;
      RECT 3388.5000 1279.5600 3390.2000 1280.6400 ;
      RECT 5.3000 1279.5600 3384.9000 1280.6400 ;
      RECT 0.0000 1279.5600 1.7000 1280.6400 ;
      RECT 0.0000 1277.9200 3390.2000 1279.5600 ;
      RECT 3384.5000 1276.8400 3390.2000 1277.9200 ;
      RECT 9.3000 1276.8400 3380.9000 1277.9200 ;
      RECT 0.0000 1276.8400 5.7000 1277.9200 ;
      RECT 0.0000 1275.2000 3390.2000 1276.8400 ;
      RECT 3388.5000 1274.1200 3390.2000 1275.2000 ;
      RECT 5.3000 1274.1200 3384.9000 1275.2000 ;
      RECT 0.0000 1274.1200 1.7000 1275.2000 ;
      RECT 0.0000 1272.4800 3390.2000 1274.1200 ;
      RECT 3384.5000 1271.4000 3390.2000 1272.4800 ;
      RECT 9.3000 1271.4000 3380.9000 1272.4800 ;
      RECT 0.0000 1271.4000 5.7000 1272.4800 ;
      RECT 0.0000 1269.7600 3390.2000 1271.4000 ;
      RECT 3388.5000 1268.6800 3390.2000 1269.7600 ;
      RECT 5.3000 1268.6800 3384.9000 1269.7600 ;
      RECT 0.0000 1268.6800 1.7000 1269.7600 ;
      RECT 0.0000 1267.0400 3390.2000 1268.6800 ;
      RECT 3384.5000 1265.9600 3390.2000 1267.0400 ;
      RECT 9.3000 1265.9600 3380.9000 1267.0400 ;
      RECT 0.0000 1265.9600 5.7000 1267.0400 ;
      RECT 0.0000 1264.3200 3390.2000 1265.9600 ;
      RECT 3388.5000 1263.2400 3390.2000 1264.3200 ;
      RECT 5.3000 1263.2400 3384.9000 1264.3200 ;
      RECT 0.0000 1263.2400 1.7000 1264.3200 ;
      RECT 0.0000 1261.6000 3390.2000 1263.2400 ;
      RECT 0.0000 1261.5900 5.7000 1261.6000 ;
      RECT 1.1000 1260.6900 5.7000 1261.5900 ;
      RECT 3384.5000 1260.5200 3390.2000 1261.6000 ;
      RECT 9.3000 1260.5200 3380.9000 1261.6000 ;
      RECT 0.0000 1260.5200 5.7000 1260.6900 ;
      RECT 0.0000 1258.8800 3390.2000 1260.5200 ;
      RECT 3388.5000 1257.8000 3390.2000 1258.8800 ;
      RECT 5.3000 1257.8000 3384.9000 1258.8800 ;
      RECT 0.0000 1257.8000 1.7000 1258.8800 ;
      RECT 0.0000 1256.1600 3390.2000 1257.8000 ;
      RECT 3384.5000 1255.0800 3390.2000 1256.1600 ;
      RECT 9.3000 1255.0800 3380.9000 1256.1600 ;
      RECT 0.0000 1255.0800 5.7000 1256.1600 ;
      RECT 0.0000 1253.4400 3390.2000 1255.0800 ;
      RECT 3388.5000 1252.3600 3390.2000 1253.4400 ;
      RECT 5.3000 1252.3600 3384.9000 1253.4400 ;
      RECT 0.0000 1252.3600 1.7000 1253.4400 ;
      RECT 0.0000 1250.7200 3390.2000 1252.3600 ;
      RECT 3384.5000 1249.6400 3390.2000 1250.7200 ;
      RECT 9.3000 1249.6400 3380.9000 1250.7200 ;
      RECT 0.0000 1249.6400 5.7000 1250.7200 ;
      RECT 0.0000 1248.0000 3390.2000 1249.6400 ;
      RECT 3388.5000 1246.9200 3390.2000 1248.0000 ;
      RECT 5.3000 1246.9200 3384.9000 1248.0000 ;
      RECT 0.0000 1246.9200 1.7000 1248.0000 ;
      RECT 0.0000 1245.2800 3390.2000 1246.9200 ;
      RECT 3384.5000 1244.2000 3390.2000 1245.2800 ;
      RECT 9.3000 1244.2000 3380.9000 1245.2800 ;
      RECT 0.0000 1244.2000 5.7000 1245.2800 ;
      RECT 0.0000 1243.2900 3390.2000 1244.2000 ;
      RECT 0.0000 1242.5600 3389.1000 1243.2900 ;
      RECT 3388.5000 1242.3900 3389.1000 1242.5600 ;
      RECT 3388.5000 1241.4800 3390.2000 1242.3900 ;
      RECT 5.3000 1241.4800 3384.9000 1242.5600 ;
      RECT 0.0000 1241.4800 1.7000 1242.5600 ;
      RECT 0.0000 1239.8400 3390.2000 1241.4800 ;
      RECT 3384.5000 1238.7600 3390.2000 1239.8400 ;
      RECT 9.3000 1238.7600 3380.9000 1239.8400 ;
      RECT 0.0000 1238.7600 5.7000 1239.8400 ;
      RECT 0.0000 1237.1200 3390.2000 1238.7600 ;
      RECT 3388.5000 1236.0400 3390.2000 1237.1200 ;
      RECT 5.3000 1236.0400 3384.9000 1237.1200 ;
      RECT 0.0000 1236.0400 1.7000 1237.1200 ;
      RECT 0.0000 1235.9700 3390.2000 1236.0400 ;
      RECT 1.1000 1235.0700 3390.2000 1235.9700 ;
      RECT 0.0000 1234.4000 3390.2000 1235.0700 ;
      RECT 3384.5000 1233.3200 3390.2000 1234.4000 ;
      RECT 9.3000 1233.3200 3380.9000 1234.4000 ;
      RECT 0.0000 1233.3200 5.7000 1234.4000 ;
      RECT 0.0000 1231.6800 3390.2000 1233.3200 ;
      RECT 3388.5000 1230.6000 3390.2000 1231.6800 ;
      RECT 5.3000 1230.6000 3384.9000 1231.6800 ;
      RECT 0.0000 1230.6000 1.7000 1231.6800 ;
      RECT 0.0000 1228.9600 3390.2000 1230.6000 ;
      RECT 3384.5000 1227.8800 3390.2000 1228.9600 ;
      RECT 9.3000 1227.8800 3380.9000 1228.9600 ;
      RECT 0.0000 1227.8800 5.7000 1228.9600 ;
      RECT 0.0000 1226.2400 3390.2000 1227.8800 ;
      RECT 3388.5000 1225.1600 3390.2000 1226.2400 ;
      RECT 5.3000 1225.1600 3384.9000 1226.2400 ;
      RECT 0.0000 1225.1600 1.7000 1226.2400 ;
      RECT 0.0000 1223.5200 3390.2000 1225.1600 ;
      RECT 3384.5000 1222.4400 3390.2000 1223.5200 ;
      RECT 9.3000 1222.4400 3380.9000 1223.5200 ;
      RECT 0.0000 1222.4400 5.7000 1223.5200 ;
      RECT 0.0000 1220.8000 3390.2000 1222.4400 ;
      RECT 3388.5000 1219.7200 3390.2000 1220.8000 ;
      RECT 5.3000 1219.7200 3384.9000 1220.8000 ;
      RECT 0.0000 1219.7200 1.7000 1220.8000 ;
      RECT 0.0000 1218.0800 3390.2000 1219.7200 ;
      RECT 3384.5000 1217.0000 3390.2000 1218.0800 ;
      RECT 9.3000 1217.0000 3380.9000 1218.0800 ;
      RECT 0.0000 1217.0000 5.7000 1218.0800 ;
      RECT 0.0000 1215.3600 3390.2000 1217.0000 ;
      RECT 3388.5000 1214.2800 3390.2000 1215.3600 ;
      RECT 5.3000 1214.2800 3384.9000 1215.3600 ;
      RECT 0.0000 1214.2800 1.7000 1215.3600 ;
      RECT 0.0000 1212.6400 3390.2000 1214.2800 ;
      RECT 3384.5000 1211.5600 3390.2000 1212.6400 ;
      RECT 9.3000 1211.5600 3380.9000 1212.6400 ;
      RECT 0.0000 1211.5600 5.7000 1212.6400 ;
      RECT 0.0000 1210.9600 3390.2000 1211.5600 ;
      RECT 1.1000 1210.0600 3390.2000 1210.9600 ;
      RECT 0.0000 1209.9200 3390.2000 1210.0600 ;
      RECT 3388.5000 1208.8400 3390.2000 1209.9200 ;
      RECT 5.3000 1208.8400 3384.9000 1209.9200 ;
      RECT 0.0000 1208.8400 1.7000 1209.9200 ;
      RECT 0.0000 1207.2000 3390.2000 1208.8400 ;
      RECT 3384.5000 1206.1200 3390.2000 1207.2000 ;
      RECT 9.3000 1206.1200 3380.9000 1207.2000 ;
      RECT 0.0000 1206.1200 5.7000 1207.2000 ;
      RECT 0.0000 1204.4800 3390.2000 1206.1200 ;
      RECT 3388.5000 1203.4000 3390.2000 1204.4800 ;
      RECT 5.3000 1203.4000 3384.9000 1204.4800 ;
      RECT 0.0000 1203.4000 1.7000 1204.4800 ;
      RECT 0.0000 1201.7600 3390.2000 1203.4000 ;
      RECT 3384.5000 1200.6800 3390.2000 1201.7600 ;
      RECT 9.3000 1200.6800 3380.9000 1201.7600 ;
      RECT 0.0000 1200.6800 5.7000 1201.7600 ;
      RECT 0.0000 1199.0400 3390.2000 1200.6800 ;
      RECT 3388.5000 1197.9600 3390.2000 1199.0400 ;
      RECT 5.3000 1197.9600 3384.9000 1199.0400 ;
      RECT 0.0000 1197.9600 1.7000 1199.0400 ;
      RECT 0.0000 1196.3200 3390.2000 1197.9600 ;
      RECT 3384.5000 1195.2400 3390.2000 1196.3200 ;
      RECT 9.3000 1195.2400 3380.9000 1196.3200 ;
      RECT 0.0000 1195.2400 5.7000 1196.3200 ;
      RECT 0.0000 1193.6000 3390.2000 1195.2400 ;
      RECT 3388.5000 1192.5200 3390.2000 1193.6000 ;
      RECT 5.3000 1192.5200 3384.9000 1193.6000 ;
      RECT 0.0000 1192.5200 1.7000 1193.6000 ;
      RECT 0.0000 1190.8800 3390.2000 1192.5200 ;
      RECT 3384.5000 1189.8000 3390.2000 1190.8800 ;
      RECT 9.3000 1189.8000 3380.9000 1190.8800 ;
      RECT 0.0000 1189.8000 5.7000 1190.8800 ;
      RECT 0.0000 1188.1600 3390.2000 1189.8000 ;
      RECT 3388.5000 1187.0800 3390.2000 1188.1600 ;
      RECT 5.3000 1187.0800 3384.9000 1188.1600 ;
      RECT 0.0000 1187.0800 1.7000 1188.1600 ;
      RECT 0.0000 1185.9500 3390.2000 1187.0800 ;
      RECT 1.1000 1185.4400 3390.2000 1185.9500 ;
      RECT 1.1000 1185.0500 5.7000 1185.4400 ;
      RECT 3384.5000 1184.3600 3390.2000 1185.4400 ;
      RECT 9.3000 1184.3600 3380.9000 1185.4400 ;
      RECT 0.0000 1184.3600 5.7000 1185.0500 ;
      RECT 0.0000 1182.7200 3390.2000 1184.3600 ;
      RECT 3388.5000 1181.6400 3390.2000 1182.7200 ;
      RECT 5.3000 1181.6400 3384.9000 1182.7200 ;
      RECT 0.0000 1181.6400 1.7000 1182.7200 ;
      RECT 0.0000 1180.0000 3390.2000 1181.6400 ;
      RECT 3384.5000 1178.9200 3390.2000 1180.0000 ;
      RECT 9.3000 1178.9200 3380.9000 1180.0000 ;
      RECT 0.0000 1178.9200 5.7000 1180.0000 ;
      RECT 0.0000 1177.2800 3390.2000 1178.9200 ;
      RECT 3388.5000 1176.2000 3390.2000 1177.2800 ;
      RECT 5.3000 1176.2000 3384.9000 1177.2800 ;
      RECT 0.0000 1176.2000 1.7000 1177.2800 ;
      RECT 0.0000 1174.5600 3390.2000 1176.2000 ;
      RECT 3384.5000 1173.4800 3390.2000 1174.5600 ;
      RECT 9.3000 1173.4800 3380.9000 1174.5600 ;
      RECT 0.0000 1173.4800 5.7000 1174.5600 ;
      RECT 0.0000 1171.8400 3390.2000 1173.4800 ;
      RECT 3388.5000 1170.7600 3390.2000 1171.8400 ;
      RECT 5.3000 1170.7600 3384.9000 1171.8400 ;
      RECT 0.0000 1170.7600 1.7000 1171.8400 ;
      RECT 0.0000 1169.1200 3390.2000 1170.7600 ;
      RECT 3384.5000 1168.0400 3390.2000 1169.1200 ;
      RECT 9.3000 1168.0400 3380.9000 1169.1200 ;
      RECT 0.0000 1168.0400 5.7000 1169.1200 ;
      RECT 0.0000 1166.4000 3390.2000 1168.0400 ;
      RECT 3388.5000 1165.3200 3390.2000 1166.4000 ;
      RECT 5.3000 1165.3200 3384.9000 1166.4000 ;
      RECT 0.0000 1165.3200 1.7000 1166.4000 ;
      RECT 0.0000 1163.6800 3390.2000 1165.3200 ;
      RECT 3384.5000 1162.6000 3390.2000 1163.6800 ;
      RECT 9.3000 1162.6000 3380.9000 1163.6800 ;
      RECT 0.0000 1162.6000 5.7000 1163.6800 ;
      RECT 0.0000 1160.9600 3390.2000 1162.6000 ;
      RECT 0.0000 1160.3300 1.7000 1160.9600 ;
      RECT 3388.5000 1159.8800 3390.2000 1160.9600 ;
      RECT 5.3000 1159.8800 3384.9000 1160.9600 ;
      RECT 1.1000 1159.8800 1.7000 1160.3300 ;
      RECT 1.1000 1159.4300 3390.2000 1159.8800 ;
      RECT 0.0000 1158.2400 3390.2000 1159.4300 ;
      RECT 3384.5000 1157.1600 3390.2000 1158.2400 ;
      RECT 9.3000 1157.1600 3380.9000 1158.2400 ;
      RECT 0.0000 1157.1600 5.7000 1158.2400 ;
      RECT 0.0000 1155.5200 3390.2000 1157.1600 ;
      RECT 3388.5000 1154.4400 3390.2000 1155.5200 ;
      RECT 5.3000 1154.4400 3384.9000 1155.5200 ;
      RECT 0.0000 1154.4400 1.7000 1155.5200 ;
      RECT 0.0000 1152.8000 3390.2000 1154.4400 ;
      RECT 3384.5000 1151.7200 3390.2000 1152.8000 ;
      RECT 9.3000 1151.7200 3380.9000 1152.8000 ;
      RECT 0.0000 1151.7200 5.7000 1152.8000 ;
      RECT 0.0000 1150.0800 3390.2000 1151.7200 ;
      RECT 3388.5000 1149.0000 3390.2000 1150.0800 ;
      RECT 5.3000 1149.0000 3384.9000 1150.0800 ;
      RECT 0.0000 1149.0000 1.7000 1150.0800 ;
      RECT 0.0000 1147.3600 3390.2000 1149.0000 ;
      RECT 3384.5000 1146.2800 3390.2000 1147.3600 ;
      RECT 9.3000 1146.2800 3380.9000 1147.3600 ;
      RECT 0.0000 1146.2800 5.7000 1147.3600 ;
      RECT 0.0000 1144.6400 3390.2000 1146.2800 ;
      RECT 3388.5000 1143.5600 3390.2000 1144.6400 ;
      RECT 5.3000 1143.5600 3384.9000 1144.6400 ;
      RECT 0.0000 1143.5600 1.7000 1144.6400 ;
      RECT 0.0000 1141.9200 3390.2000 1143.5600 ;
      RECT 3384.5000 1140.8400 3390.2000 1141.9200 ;
      RECT 9.3000 1140.8400 3380.9000 1141.9200 ;
      RECT 0.0000 1140.8400 5.7000 1141.9200 ;
      RECT 0.0000 1139.2000 3390.2000 1140.8400 ;
      RECT 3388.5000 1138.9800 3390.2000 1139.2000 ;
      RECT 3388.5000 1138.1200 3389.1000 1138.9800 ;
      RECT 5.3000 1138.1200 3384.9000 1139.2000 ;
      RECT 0.0000 1138.1200 1.7000 1139.2000 ;
      RECT 0.0000 1138.0800 3389.1000 1138.1200 ;
      RECT 0.0000 1136.4800 3390.2000 1138.0800 ;
      RECT 3384.5000 1135.4000 3390.2000 1136.4800 ;
      RECT 9.3000 1135.4000 3380.9000 1136.4800 ;
      RECT 0.0000 1135.4000 5.7000 1136.4800 ;
      RECT 0.0000 1135.3200 3390.2000 1135.4000 ;
      RECT 1.1000 1134.4200 3390.2000 1135.3200 ;
      RECT 0.0000 1133.7600 3390.2000 1134.4200 ;
      RECT 3388.5000 1132.6800 3390.2000 1133.7600 ;
      RECT 5.3000 1132.6800 3384.9000 1133.7600 ;
      RECT 0.0000 1132.6800 1.7000 1133.7600 ;
      RECT 0.0000 1131.0400 3390.2000 1132.6800 ;
      RECT 3384.5000 1129.9600 3390.2000 1131.0400 ;
      RECT 9.3000 1129.9600 3380.9000 1131.0400 ;
      RECT 0.0000 1129.9600 5.7000 1131.0400 ;
      RECT 0.0000 1128.3200 3390.2000 1129.9600 ;
      RECT 3388.5000 1127.2400 3390.2000 1128.3200 ;
      RECT 5.3000 1127.2400 3384.9000 1128.3200 ;
      RECT 0.0000 1127.2400 1.7000 1128.3200 ;
      RECT 0.0000 1125.6000 3390.2000 1127.2400 ;
      RECT 3384.5000 1124.5200 3390.2000 1125.6000 ;
      RECT 9.3000 1124.5200 3380.9000 1125.6000 ;
      RECT 0.0000 1124.5200 5.7000 1125.6000 ;
      RECT 0.0000 1122.8800 3390.2000 1124.5200 ;
      RECT 3388.5000 1121.8000 3390.2000 1122.8800 ;
      RECT 5.3000 1121.8000 3384.9000 1122.8800 ;
      RECT 0.0000 1121.8000 1.7000 1122.8800 ;
      RECT 0.0000 1120.1600 3390.2000 1121.8000 ;
      RECT 3384.5000 1119.0800 3390.2000 1120.1600 ;
      RECT 9.3000 1119.0800 3380.9000 1120.1600 ;
      RECT 0.0000 1119.0800 5.7000 1120.1600 ;
      RECT 0.0000 1117.4400 3390.2000 1119.0800 ;
      RECT 3388.5000 1116.3600 3390.2000 1117.4400 ;
      RECT 5.3000 1116.3600 3384.9000 1117.4400 ;
      RECT 0.0000 1116.3600 1.7000 1117.4400 ;
      RECT 0.0000 1114.7200 3390.2000 1116.3600 ;
      RECT 3384.5000 1113.6400 3390.2000 1114.7200 ;
      RECT 9.3000 1113.6400 3380.9000 1114.7200 ;
      RECT 0.0000 1113.6400 5.7000 1114.7200 ;
      RECT 0.0000 1112.0000 3390.2000 1113.6400 ;
      RECT 3388.5000 1110.9200 3390.2000 1112.0000 ;
      RECT 5.3000 1110.9200 3384.9000 1112.0000 ;
      RECT 0.0000 1110.9200 1.7000 1112.0000 ;
      RECT 0.0000 1110.3100 3390.2000 1110.9200 ;
      RECT 1.1000 1109.4100 3390.2000 1110.3100 ;
      RECT 0.0000 1109.2800 3390.2000 1109.4100 ;
      RECT 3384.5000 1108.2000 3390.2000 1109.2800 ;
      RECT 9.3000 1108.2000 3380.9000 1109.2800 ;
      RECT 0.0000 1108.2000 5.7000 1109.2800 ;
      RECT 0.0000 1106.5600 3390.2000 1108.2000 ;
      RECT 3388.5000 1105.4800 3390.2000 1106.5600 ;
      RECT 5.3000 1105.4800 3384.9000 1106.5600 ;
      RECT 0.0000 1105.4800 1.7000 1106.5600 ;
      RECT 0.0000 1103.8400 3390.2000 1105.4800 ;
      RECT 3384.5000 1102.7600 3390.2000 1103.8400 ;
      RECT 9.3000 1102.7600 3380.9000 1103.8400 ;
      RECT 0.0000 1102.7600 5.7000 1103.8400 ;
      RECT 0.0000 1101.1200 3390.2000 1102.7600 ;
      RECT 3388.5000 1100.0400 3390.2000 1101.1200 ;
      RECT 5.3000 1100.0400 3384.9000 1101.1200 ;
      RECT 0.0000 1100.0400 1.7000 1101.1200 ;
      RECT 0.0000 1098.4000 3390.2000 1100.0400 ;
      RECT 3384.5000 1097.3200 3390.2000 1098.4000 ;
      RECT 9.3000 1097.3200 3380.9000 1098.4000 ;
      RECT 0.0000 1097.3200 5.7000 1098.4000 ;
      RECT 0.0000 1095.6800 3390.2000 1097.3200 ;
      RECT 3388.5000 1094.6000 3390.2000 1095.6800 ;
      RECT 5.3000 1094.6000 3384.9000 1095.6800 ;
      RECT 0.0000 1094.6000 1.7000 1095.6800 ;
      RECT 0.0000 1092.9600 3390.2000 1094.6000 ;
      RECT 3384.5000 1091.8800 3390.2000 1092.9600 ;
      RECT 9.3000 1091.8800 3380.9000 1092.9600 ;
      RECT 0.0000 1091.8800 5.7000 1092.9600 ;
      RECT 0.0000 1090.2400 3390.2000 1091.8800 ;
      RECT 3388.5000 1089.1600 3390.2000 1090.2400 ;
      RECT 5.3000 1089.1600 3384.9000 1090.2400 ;
      RECT 0.0000 1089.1600 1.7000 1090.2400 ;
      RECT 0.0000 1087.5200 3390.2000 1089.1600 ;
      RECT 3384.5000 1086.4400 3390.2000 1087.5200 ;
      RECT 9.3000 1086.4400 3380.9000 1087.5200 ;
      RECT 0.0000 1086.4400 5.7000 1087.5200 ;
      RECT 0.0000 1084.8000 3390.2000 1086.4400 ;
      RECT 0.0000 1084.6900 1.7000 1084.8000 ;
      RECT 1.1000 1083.7900 1.7000 1084.6900 ;
      RECT 3388.5000 1083.7200 3390.2000 1084.8000 ;
      RECT 5.3000 1083.7200 3384.9000 1084.8000 ;
      RECT 0.0000 1083.7200 1.7000 1083.7900 ;
      RECT 0.0000 1082.0800 3390.2000 1083.7200 ;
      RECT 3384.5000 1081.0000 3390.2000 1082.0800 ;
      RECT 9.3000 1081.0000 3380.9000 1082.0800 ;
      RECT 0.0000 1081.0000 5.7000 1082.0800 ;
      RECT 0.0000 1079.3600 3390.2000 1081.0000 ;
      RECT 3388.5000 1078.2800 3390.2000 1079.3600 ;
      RECT 5.3000 1078.2800 3384.9000 1079.3600 ;
      RECT 0.0000 1078.2800 1.7000 1079.3600 ;
      RECT 0.0000 1076.6400 3390.2000 1078.2800 ;
      RECT 3384.5000 1075.5600 3390.2000 1076.6400 ;
      RECT 9.3000 1075.5600 3380.9000 1076.6400 ;
      RECT 0.0000 1075.5600 5.7000 1076.6400 ;
      RECT 0.0000 1073.9200 3390.2000 1075.5600 ;
      RECT 3388.5000 1072.8400 3390.2000 1073.9200 ;
      RECT 5.3000 1072.8400 3384.9000 1073.9200 ;
      RECT 0.0000 1072.8400 1.7000 1073.9200 ;
      RECT 0.0000 1071.2000 3390.2000 1072.8400 ;
      RECT 3384.5000 1070.1200 3390.2000 1071.2000 ;
      RECT 9.3000 1070.1200 3380.9000 1071.2000 ;
      RECT 0.0000 1070.1200 5.7000 1071.2000 ;
      RECT 0.0000 1068.4800 3390.2000 1070.1200 ;
      RECT 3388.5000 1067.4000 3390.2000 1068.4800 ;
      RECT 5.3000 1067.4000 3384.9000 1068.4800 ;
      RECT 0.0000 1067.4000 1.7000 1068.4800 ;
      RECT 0.0000 1065.7600 3390.2000 1067.4000 ;
      RECT 3384.5000 1064.6800 3390.2000 1065.7600 ;
      RECT 9.3000 1064.6800 3380.9000 1065.7600 ;
      RECT 0.0000 1064.6800 5.7000 1065.7600 ;
      RECT 0.0000 1063.0400 3390.2000 1064.6800 ;
      RECT 3388.5000 1061.9600 3390.2000 1063.0400 ;
      RECT 5.3000 1061.9600 3384.9000 1063.0400 ;
      RECT 0.0000 1061.9600 1.7000 1063.0400 ;
      RECT 0.0000 1060.3200 3390.2000 1061.9600 ;
      RECT 0.0000 1059.6800 5.7000 1060.3200 ;
      RECT 3384.5000 1059.2400 3390.2000 1060.3200 ;
      RECT 9.3000 1059.2400 3380.9000 1060.3200 ;
      RECT 1.1000 1059.2400 5.7000 1059.6800 ;
      RECT 1.1000 1058.7800 3390.2000 1059.2400 ;
      RECT 0.0000 1057.6000 3390.2000 1058.7800 ;
      RECT 3388.5000 1056.5200 3390.2000 1057.6000 ;
      RECT 5.3000 1056.5200 3384.9000 1057.6000 ;
      RECT 0.0000 1056.5200 1.7000 1057.6000 ;
      RECT 0.0000 1054.8800 3390.2000 1056.5200 ;
      RECT 3384.5000 1053.8000 3390.2000 1054.8800 ;
      RECT 9.3000 1053.8000 3380.9000 1054.8800 ;
      RECT 0.0000 1053.8000 5.7000 1054.8800 ;
      RECT 0.0000 1052.1600 3390.2000 1053.8000 ;
      RECT 3388.5000 1051.0800 3390.2000 1052.1600 ;
      RECT 5.3000 1051.0800 3384.9000 1052.1600 ;
      RECT 0.0000 1051.0800 1.7000 1052.1600 ;
      RECT 0.0000 1049.4400 3390.2000 1051.0800 ;
      RECT 3384.5000 1048.3600 3390.2000 1049.4400 ;
      RECT 9.3000 1048.3600 3380.9000 1049.4400 ;
      RECT 0.0000 1048.3600 5.7000 1049.4400 ;
      RECT 0.0000 1046.7200 3390.2000 1048.3600 ;
      RECT 3388.5000 1045.6400 3390.2000 1046.7200 ;
      RECT 5.3000 1045.6400 3384.9000 1046.7200 ;
      RECT 0.0000 1045.6400 1.7000 1046.7200 ;
      RECT 0.0000 1044.0000 3390.2000 1045.6400 ;
      RECT 3384.5000 1042.9200 3390.2000 1044.0000 ;
      RECT 9.3000 1042.9200 3380.9000 1044.0000 ;
      RECT 0.0000 1042.9200 5.7000 1044.0000 ;
      RECT 0.0000 1041.2800 3390.2000 1042.9200 ;
      RECT 3388.5000 1040.2000 3390.2000 1041.2800 ;
      RECT 5.3000 1040.2000 3384.9000 1041.2800 ;
      RECT 0.0000 1040.2000 1.7000 1041.2800 ;
      RECT 0.0000 1038.5600 3390.2000 1040.2000 ;
      RECT 3384.5000 1037.4800 3390.2000 1038.5600 ;
      RECT 9.3000 1037.4800 3380.9000 1038.5600 ;
      RECT 0.0000 1037.4800 5.7000 1038.5600 ;
      RECT 0.0000 1035.8400 3390.2000 1037.4800 ;
      RECT 3388.5000 1035.2800 3390.2000 1035.8400 ;
      RECT 3388.5000 1034.7600 3389.1000 1035.2800 ;
      RECT 5.3000 1034.7600 3384.9000 1035.8400 ;
      RECT 0.0000 1034.7600 1.7000 1035.8400 ;
      RECT 0.0000 1034.6700 3389.1000 1034.7600 ;
      RECT 1.1000 1034.3800 3389.1000 1034.6700 ;
      RECT 1.1000 1033.7700 3390.2000 1034.3800 ;
      RECT 0.0000 1033.1200 3390.2000 1033.7700 ;
      RECT 3384.5000 1032.0400 3390.2000 1033.1200 ;
      RECT 9.3000 1032.0400 3380.9000 1033.1200 ;
      RECT 0.0000 1032.0400 5.7000 1033.1200 ;
      RECT 0.0000 1030.4000 3390.2000 1032.0400 ;
      RECT 3388.5000 1029.3200 3390.2000 1030.4000 ;
      RECT 5.3000 1029.3200 3384.9000 1030.4000 ;
      RECT 0.0000 1029.3200 1.7000 1030.4000 ;
      RECT 0.0000 1027.6800 3390.2000 1029.3200 ;
      RECT 3384.5000 1026.6000 3390.2000 1027.6800 ;
      RECT 9.3000 1026.6000 3380.9000 1027.6800 ;
      RECT 0.0000 1026.6000 5.7000 1027.6800 ;
      RECT 0.0000 1024.9600 3390.2000 1026.6000 ;
      RECT 3388.5000 1023.8800 3390.2000 1024.9600 ;
      RECT 5.3000 1023.8800 3384.9000 1024.9600 ;
      RECT 0.0000 1023.8800 1.7000 1024.9600 ;
      RECT 0.0000 1022.2400 3390.2000 1023.8800 ;
      RECT 3384.5000 1021.1600 3390.2000 1022.2400 ;
      RECT 9.3000 1021.1600 3380.9000 1022.2400 ;
      RECT 0.0000 1021.1600 5.7000 1022.2400 ;
      RECT 0.0000 1019.5200 3390.2000 1021.1600 ;
      RECT 3388.5000 1018.4400 3390.2000 1019.5200 ;
      RECT 5.3000 1018.4400 3384.9000 1019.5200 ;
      RECT 0.0000 1018.4400 1.7000 1019.5200 ;
      RECT 0.0000 1016.8000 3390.2000 1018.4400 ;
      RECT 3384.5000 1015.7200 3390.2000 1016.8000 ;
      RECT 9.3000 1015.7200 3380.9000 1016.8000 ;
      RECT 0.0000 1015.7200 5.7000 1016.8000 ;
      RECT 0.0000 1014.0800 3390.2000 1015.7200 ;
      RECT 3388.5000 1013.0000 3390.2000 1014.0800 ;
      RECT 5.3000 1013.0000 3384.9000 1014.0800 ;
      RECT 0.0000 1013.0000 1.7000 1014.0800 ;
      RECT 0.0000 1011.3600 3390.2000 1013.0000 ;
      RECT 3384.5000 1010.2800 3390.2000 1011.3600 ;
      RECT 9.3000 1010.2800 3380.9000 1011.3600 ;
      RECT 0.0000 1010.2800 5.7000 1011.3600 ;
      RECT 0.0000 1009.0500 3390.2000 1010.2800 ;
      RECT 1.1000 1008.6400 3390.2000 1009.0500 ;
      RECT 1.1000 1008.1500 1.7000 1008.6400 ;
      RECT 3388.5000 1007.5600 3390.2000 1008.6400 ;
      RECT 5.3000 1007.5600 3384.9000 1008.6400 ;
      RECT 0.0000 1007.5600 1.7000 1008.1500 ;
      RECT 0.0000 1005.9200 3390.2000 1007.5600 ;
      RECT 3384.5000 1004.8400 3390.2000 1005.9200 ;
      RECT 9.3000 1004.8400 3380.9000 1005.9200 ;
      RECT 0.0000 1004.8400 5.7000 1005.9200 ;
      RECT 0.0000 1003.2000 3390.2000 1004.8400 ;
      RECT 3388.5000 1002.1200 3390.2000 1003.2000 ;
      RECT 5.3000 1002.1200 3384.9000 1003.2000 ;
      RECT 0.0000 1002.1200 1.7000 1003.2000 ;
      RECT 0.0000 1000.4800 3390.2000 1002.1200 ;
      RECT 3384.5000 999.4000 3390.2000 1000.4800 ;
      RECT 9.3000 999.4000 3380.9000 1000.4800 ;
      RECT 0.0000 999.4000 5.7000 1000.4800 ;
      RECT 0.0000 997.7600 3390.2000 999.4000 ;
      RECT 3388.5000 996.6800 3390.2000 997.7600 ;
      RECT 5.3000 996.6800 3384.9000 997.7600 ;
      RECT 0.0000 996.6800 1.7000 997.7600 ;
      RECT 0.0000 995.0400 3390.2000 996.6800 ;
      RECT 3384.5000 993.9600 3390.2000 995.0400 ;
      RECT 9.3000 993.9600 3380.9000 995.0400 ;
      RECT 0.0000 993.9600 5.7000 995.0400 ;
      RECT 0.0000 992.3200 3390.2000 993.9600 ;
      RECT 3388.5000 991.2400 3390.2000 992.3200 ;
      RECT 5.3000 991.2400 3384.9000 992.3200 ;
      RECT 0.0000 991.2400 1.7000 992.3200 ;
      RECT 0.0000 989.6000 3390.2000 991.2400 ;
      RECT 3384.5000 988.5200 3390.2000 989.6000 ;
      RECT 9.3000 988.5200 3380.9000 989.6000 ;
      RECT 0.0000 988.5200 5.7000 989.6000 ;
      RECT 0.0000 986.8800 3390.2000 988.5200 ;
      RECT 3388.5000 985.8000 3390.2000 986.8800 ;
      RECT 5.3000 985.8000 3384.9000 986.8800 ;
      RECT 0.0000 985.8000 1.7000 986.8800 ;
      RECT 0.0000 984.1600 3390.2000 985.8000 ;
      RECT 0.0000 984.0400 5.7000 984.1600 ;
      RECT 1.1000 983.1400 5.7000 984.0400 ;
      RECT 3384.5000 983.0800 3390.2000 984.1600 ;
      RECT 9.3000 983.0800 3380.9000 984.1600 ;
      RECT 0.0000 983.0800 5.7000 983.1400 ;
      RECT 0.0000 981.4400 3390.2000 983.0800 ;
      RECT 3388.5000 980.3600 3390.2000 981.4400 ;
      RECT 5.3000 980.3600 3384.9000 981.4400 ;
      RECT 0.0000 980.3600 1.7000 981.4400 ;
      RECT 0.0000 978.7200 3390.2000 980.3600 ;
      RECT 3384.5000 977.6400 3390.2000 978.7200 ;
      RECT 9.3000 977.6400 3380.9000 978.7200 ;
      RECT 0.0000 977.6400 5.7000 978.7200 ;
      RECT 0.0000 976.0000 3390.2000 977.6400 ;
      RECT 3388.5000 974.9200 3390.2000 976.0000 ;
      RECT 5.3000 974.9200 3384.9000 976.0000 ;
      RECT 0.0000 974.9200 1.7000 976.0000 ;
      RECT 0.0000 973.2800 3390.2000 974.9200 ;
      RECT 3384.5000 972.2000 3390.2000 973.2800 ;
      RECT 9.3000 972.2000 3380.9000 973.2800 ;
      RECT 0.0000 972.2000 5.7000 973.2800 ;
      RECT 0.0000 970.5600 3390.2000 972.2000 ;
      RECT 3388.5000 969.4800 3390.2000 970.5600 ;
      RECT 5.3000 969.4800 3384.9000 970.5600 ;
      RECT 0.0000 969.4800 1.7000 970.5600 ;
      RECT 0.0000 967.8400 3390.2000 969.4800 ;
      RECT 3384.5000 966.7600 3390.2000 967.8400 ;
      RECT 9.3000 966.7600 3380.9000 967.8400 ;
      RECT 0.0000 966.7600 5.7000 967.8400 ;
      RECT 0.0000 965.1200 3390.2000 966.7600 ;
      RECT 3388.5000 964.0400 3390.2000 965.1200 ;
      RECT 5.3000 964.0400 3384.9000 965.1200 ;
      RECT 0.0000 964.0400 1.7000 965.1200 ;
      RECT 0.0000 962.4000 3390.2000 964.0400 ;
      RECT 3384.5000 961.3200 3390.2000 962.4000 ;
      RECT 9.3000 961.3200 3380.9000 962.4000 ;
      RECT 0.0000 961.3200 5.7000 962.4000 ;
      RECT 0.0000 959.6800 3390.2000 961.3200 ;
      RECT 0.0000 959.0300 1.7000 959.6800 ;
      RECT 3388.5000 958.6000 3390.2000 959.6800 ;
      RECT 5.3000 958.6000 3384.9000 959.6800 ;
      RECT 1.1000 958.6000 1.7000 959.0300 ;
      RECT 1.1000 958.1300 3390.2000 958.6000 ;
      RECT 0.0000 956.9600 3390.2000 958.1300 ;
      RECT 3384.5000 955.8800 3390.2000 956.9600 ;
      RECT 9.3000 955.8800 3380.9000 956.9600 ;
      RECT 0.0000 955.8800 5.7000 956.9600 ;
      RECT 0.0000 954.2400 3390.2000 955.8800 ;
      RECT 3388.5000 953.1600 3390.2000 954.2400 ;
      RECT 5.3000 953.1600 3384.9000 954.2400 ;
      RECT 0.0000 953.1600 1.7000 954.2400 ;
      RECT 0.0000 951.5200 3390.2000 953.1600 ;
      RECT 3384.5000 950.4400 3390.2000 951.5200 ;
      RECT 9.3000 950.4400 3380.9000 951.5200 ;
      RECT 0.0000 950.4400 5.7000 951.5200 ;
      RECT 0.0000 948.8000 3390.2000 950.4400 ;
      RECT 3388.5000 947.7200 3390.2000 948.8000 ;
      RECT 5.3000 947.7200 3384.9000 948.8000 ;
      RECT 0.0000 947.7200 1.7000 948.8000 ;
      RECT 0.0000 946.0800 3390.2000 947.7200 ;
      RECT 3384.5000 945.0000 3390.2000 946.0800 ;
      RECT 9.3000 945.0000 3380.9000 946.0800 ;
      RECT 0.0000 945.0000 5.7000 946.0800 ;
      RECT 0.0000 943.3600 3390.2000 945.0000 ;
      RECT 3388.5000 942.2800 3390.2000 943.3600 ;
      RECT 5.3000 942.2800 3384.9000 943.3600 ;
      RECT 0.0000 942.2800 1.7000 943.3600 ;
      RECT 0.0000 940.6400 3390.2000 942.2800 ;
      RECT 3384.5000 939.5600 3390.2000 940.6400 ;
      RECT 9.3000 939.5600 3380.9000 940.6400 ;
      RECT 0.0000 939.5600 5.7000 940.6400 ;
      RECT 0.0000 937.9200 3390.2000 939.5600 ;
      RECT 3388.5000 936.8400 3390.2000 937.9200 ;
      RECT 5.3000 936.8400 3384.9000 937.9200 ;
      RECT 0.0000 936.8400 1.7000 937.9200 ;
      RECT 0.0000 935.2000 3390.2000 936.8400 ;
      RECT 3384.5000 934.1200 3390.2000 935.2000 ;
      RECT 9.3000 934.1200 3380.9000 935.2000 ;
      RECT 0.0000 934.1200 5.7000 935.2000 ;
      RECT 0.0000 933.4100 3390.2000 934.1200 ;
      RECT 1.1000 932.5100 3390.2000 933.4100 ;
      RECT 0.0000 932.4800 3390.2000 932.5100 ;
      RECT 3388.5000 931.5800 3390.2000 932.4800 ;
      RECT 3388.5000 931.4000 3389.1000 931.5800 ;
      RECT 5.3000 931.4000 3384.9000 932.4800 ;
      RECT 0.0000 931.4000 1.7000 932.4800 ;
      RECT 0.0000 930.6800 3389.1000 931.4000 ;
      RECT 0.0000 929.7600 3390.2000 930.6800 ;
      RECT 3384.5000 928.6800 3390.2000 929.7600 ;
      RECT 9.3000 928.6800 3380.9000 929.7600 ;
      RECT 0.0000 928.6800 5.7000 929.7600 ;
      RECT 0.0000 927.0400 3390.2000 928.6800 ;
      RECT 3388.5000 925.9600 3390.2000 927.0400 ;
      RECT 5.3000 925.9600 3384.9000 927.0400 ;
      RECT 0.0000 925.9600 1.7000 927.0400 ;
      RECT 0.0000 924.3200 3390.2000 925.9600 ;
      RECT 3384.5000 923.2400 3390.2000 924.3200 ;
      RECT 9.3000 923.2400 3380.9000 924.3200 ;
      RECT 0.0000 923.2400 5.7000 924.3200 ;
      RECT 0.0000 921.6000 3390.2000 923.2400 ;
      RECT 3388.5000 920.5200 3390.2000 921.6000 ;
      RECT 5.3000 920.5200 3384.9000 921.6000 ;
      RECT 0.0000 920.5200 1.7000 921.6000 ;
      RECT 0.0000 918.8800 3390.2000 920.5200 ;
      RECT 3384.5000 917.8000 3390.2000 918.8800 ;
      RECT 9.3000 917.8000 3380.9000 918.8800 ;
      RECT 0.0000 917.8000 5.7000 918.8800 ;
      RECT 0.0000 916.1600 3390.2000 917.8000 ;
      RECT 3388.5000 915.0800 3390.2000 916.1600 ;
      RECT 5.3000 915.0800 3384.9000 916.1600 ;
      RECT 0.0000 915.0800 1.7000 916.1600 ;
      RECT 0.0000 913.4400 3390.2000 915.0800 ;
      RECT 3384.5000 912.3600 3390.2000 913.4400 ;
      RECT 9.3000 912.3600 3380.9000 913.4400 ;
      RECT 0.0000 912.3600 5.7000 913.4400 ;
      RECT 0.0000 910.7200 3390.2000 912.3600 ;
      RECT 3388.5000 909.6400 3390.2000 910.7200 ;
      RECT 5.3000 909.6400 3384.9000 910.7200 ;
      RECT 0.0000 909.6400 1.7000 910.7200 ;
      RECT 0.0000 908.4000 3390.2000 909.6400 ;
      RECT 1.1000 908.0000 3390.2000 908.4000 ;
      RECT 1.1000 907.5000 5.7000 908.0000 ;
      RECT 3384.5000 906.9200 3390.2000 908.0000 ;
      RECT 9.3000 906.9200 3380.9000 908.0000 ;
      RECT 0.0000 906.9200 5.7000 907.5000 ;
      RECT 0.0000 905.2800 3390.2000 906.9200 ;
      RECT 3388.5000 904.2000 3390.2000 905.2800 ;
      RECT 5.3000 904.2000 3384.9000 905.2800 ;
      RECT 0.0000 904.2000 1.7000 905.2800 ;
      RECT 0.0000 902.5600 3390.2000 904.2000 ;
      RECT 3384.5000 901.4800 3390.2000 902.5600 ;
      RECT 9.3000 901.4800 3380.9000 902.5600 ;
      RECT 0.0000 901.4800 5.7000 902.5600 ;
      RECT 0.0000 899.8400 3390.2000 901.4800 ;
      RECT 3388.5000 898.7600 3390.2000 899.8400 ;
      RECT 5.3000 898.7600 3384.9000 899.8400 ;
      RECT 0.0000 898.7600 1.7000 899.8400 ;
      RECT 0.0000 897.1200 3390.2000 898.7600 ;
      RECT 3384.5000 896.0400 3390.2000 897.1200 ;
      RECT 9.3000 896.0400 3380.9000 897.1200 ;
      RECT 0.0000 896.0400 5.7000 897.1200 ;
      RECT 0.0000 894.4000 3390.2000 896.0400 ;
      RECT 3388.5000 893.3200 3390.2000 894.4000 ;
      RECT 5.3000 893.3200 3384.9000 894.4000 ;
      RECT 0.0000 893.3200 1.7000 894.4000 ;
      RECT 0.0000 891.6800 3390.2000 893.3200 ;
      RECT 3384.5000 890.6000 3390.2000 891.6800 ;
      RECT 9.3000 890.6000 3380.9000 891.6800 ;
      RECT 0.0000 890.6000 5.7000 891.6800 ;
      RECT 0.0000 888.9600 3390.2000 890.6000 ;
      RECT 3388.5000 887.8800 3390.2000 888.9600 ;
      RECT 5.3000 887.8800 3384.9000 888.9600 ;
      RECT 0.0000 887.8800 1.7000 888.9600 ;
      RECT 0.0000 886.2400 3390.2000 887.8800 ;
      RECT 3384.5000 885.1600 3390.2000 886.2400 ;
      RECT 9.3000 885.1600 3380.9000 886.2400 ;
      RECT 0.0000 885.1600 5.7000 886.2400 ;
      RECT 0.0000 883.5200 3390.2000 885.1600 ;
      RECT 0.0000 883.3900 1.7000 883.5200 ;
      RECT 1.1000 882.4900 1.7000 883.3900 ;
      RECT 3388.5000 882.4400 3390.2000 883.5200 ;
      RECT 5.3000 882.4400 3384.9000 883.5200 ;
      RECT 0.0000 882.4400 1.7000 882.4900 ;
      RECT 0.0000 880.8000 3390.2000 882.4400 ;
      RECT 3384.5000 879.7200 3390.2000 880.8000 ;
      RECT 9.3000 879.7200 3380.9000 880.8000 ;
      RECT 0.0000 879.7200 5.7000 880.8000 ;
      RECT 0.0000 878.0800 3390.2000 879.7200 ;
      RECT 3388.5000 877.0000 3390.2000 878.0800 ;
      RECT 5.3000 877.0000 3384.9000 878.0800 ;
      RECT 0.0000 877.0000 1.7000 878.0800 ;
      RECT 0.0000 875.3600 3390.2000 877.0000 ;
      RECT 3384.5000 874.2800 3390.2000 875.3600 ;
      RECT 9.3000 874.2800 3380.9000 875.3600 ;
      RECT 0.0000 874.2800 5.7000 875.3600 ;
      RECT 0.0000 872.6400 3390.2000 874.2800 ;
      RECT 3388.5000 871.5600 3390.2000 872.6400 ;
      RECT 5.3000 871.5600 3384.9000 872.6400 ;
      RECT 0.0000 871.5600 1.7000 872.6400 ;
      RECT 0.0000 869.9200 3390.2000 871.5600 ;
      RECT 3384.5000 868.8400 3390.2000 869.9200 ;
      RECT 9.3000 868.8400 3380.9000 869.9200 ;
      RECT 0.0000 868.8400 5.7000 869.9200 ;
      RECT 0.0000 867.2000 3390.2000 868.8400 ;
      RECT 3388.5000 866.1200 3390.2000 867.2000 ;
      RECT 5.3000 866.1200 3384.9000 867.2000 ;
      RECT 0.0000 866.1200 1.7000 867.2000 ;
      RECT 0.0000 864.4800 3390.2000 866.1200 ;
      RECT 3384.5000 863.4000 3390.2000 864.4800 ;
      RECT 9.3000 863.4000 3380.9000 864.4800 ;
      RECT 0.0000 863.4000 5.7000 864.4800 ;
      RECT 0.0000 861.7600 3390.2000 863.4000 ;
      RECT 3388.5000 860.6800 3390.2000 861.7600 ;
      RECT 5.3000 860.6800 3384.9000 861.7600 ;
      RECT 0.0000 860.6800 1.7000 861.7600 ;
      RECT 0.0000 859.0400 3390.2000 860.6800 ;
      RECT 3384.5000 857.9600 3390.2000 859.0400 ;
      RECT 9.3000 857.9600 3380.9000 859.0400 ;
      RECT 0.0000 857.9600 5.7000 859.0400 ;
      RECT 0.0000 857.7700 3390.2000 857.9600 ;
      RECT 1.1000 856.8700 3390.2000 857.7700 ;
      RECT 0.0000 856.3200 3390.2000 856.8700 ;
      RECT 3388.5000 855.2400 3390.2000 856.3200 ;
      RECT 5.3000 855.2400 3384.9000 856.3200 ;
      RECT 0.0000 855.2400 1.7000 856.3200 ;
      RECT 0.0000 853.6000 3390.2000 855.2400 ;
      RECT 3384.5000 852.5200 3390.2000 853.6000 ;
      RECT 9.3000 852.5200 3380.9000 853.6000 ;
      RECT 0.0000 852.5200 5.7000 853.6000 ;
      RECT 0.0000 850.8800 3390.2000 852.5200 ;
      RECT 3388.5000 849.8000 3390.2000 850.8800 ;
      RECT 5.3000 849.8000 3384.9000 850.8800 ;
      RECT 0.0000 849.8000 1.7000 850.8800 ;
      RECT 0.0000 848.1600 3390.2000 849.8000 ;
      RECT 3384.5000 847.0800 3390.2000 848.1600 ;
      RECT 9.3000 847.0800 3380.9000 848.1600 ;
      RECT 0.0000 847.0800 5.7000 848.1600 ;
      RECT 0.0000 845.4400 3390.2000 847.0800 ;
      RECT 3388.5000 844.3600 3390.2000 845.4400 ;
      RECT 5.3000 844.3600 3384.9000 845.4400 ;
      RECT 0.0000 844.3600 1.7000 845.4400 ;
      RECT 0.0000 842.7200 3390.2000 844.3600 ;
      RECT 3384.5000 841.6400 3390.2000 842.7200 ;
      RECT 9.3000 841.6400 3380.9000 842.7200 ;
      RECT 0.0000 841.6400 5.7000 842.7200 ;
      RECT 0.0000 840.0000 3390.2000 841.6400 ;
      RECT 3388.5000 838.9200 3390.2000 840.0000 ;
      RECT 5.3000 838.9200 3384.9000 840.0000 ;
      RECT 0.0000 838.9200 1.7000 840.0000 ;
      RECT 0.0000 837.2800 3390.2000 838.9200 ;
      RECT 3384.5000 836.2000 3390.2000 837.2800 ;
      RECT 9.3000 836.2000 3380.9000 837.2800 ;
      RECT 0.0000 836.2000 5.7000 837.2800 ;
      RECT 0.0000 834.5600 3390.2000 836.2000 ;
      RECT 3388.5000 833.4800 3390.2000 834.5600 ;
      RECT 5.3000 833.4800 3384.9000 834.5600 ;
      RECT 0.0000 833.4800 1.7000 834.5600 ;
      RECT 0.0000 832.7600 3390.2000 833.4800 ;
      RECT 1.1000 831.8600 3390.2000 832.7600 ;
      RECT 0.0000 831.8400 3390.2000 831.8600 ;
      RECT 3384.5000 830.7600 3390.2000 831.8400 ;
      RECT 9.3000 830.7600 3380.9000 831.8400 ;
      RECT 0.0000 830.7600 5.7000 831.8400 ;
      RECT 0.0000 829.1200 3390.2000 830.7600 ;
      RECT 3388.5000 828.0400 3390.2000 829.1200 ;
      RECT 5.3000 828.0400 3384.9000 829.1200 ;
      RECT 0.0000 828.0400 1.7000 829.1200 ;
      RECT 0.0000 827.8800 3390.2000 828.0400 ;
      RECT 0.0000 826.9800 3389.1000 827.8800 ;
      RECT 0.0000 826.4000 3390.2000 826.9800 ;
      RECT 3384.5000 825.3200 3390.2000 826.4000 ;
      RECT 9.3000 825.3200 3380.9000 826.4000 ;
      RECT 0.0000 825.3200 5.7000 826.4000 ;
      RECT 0.0000 823.6800 3390.2000 825.3200 ;
      RECT 3388.5000 822.6000 3390.2000 823.6800 ;
      RECT 5.3000 822.6000 3384.9000 823.6800 ;
      RECT 0.0000 822.6000 1.7000 823.6800 ;
      RECT 0.0000 820.9600 3390.2000 822.6000 ;
      RECT 3384.5000 819.8800 3390.2000 820.9600 ;
      RECT 9.3000 819.8800 3380.9000 820.9600 ;
      RECT 0.0000 819.8800 5.7000 820.9600 ;
      RECT 0.0000 818.2400 3390.2000 819.8800 ;
      RECT 3388.5000 817.1600 3390.2000 818.2400 ;
      RECT 5.3000 817.1600 3384.9000 818.2400 ;
      RECT 0.0000 817.1600 1.7000 818.2400 ;
      RECT 0.0000 815.5200 3390.2000 817.1600 ;
      RECT 3384.5000 814.4400 3390.2000 815.5200 ;
      RECT 9.3000 814.4400 3380.9000 815.5200 ;
      RECT 0.0000 814.4400 5.7000 815.5200 ;
      RECT 0.0000 812.8000 3390.2000 814.4400 ;
      RECT 3388.5000 811.7200 3390.2000 812.8000 ;
      RECT 5.3000 811.7200 3384.9000 812.8000 ;
      RECT 0.0000 811.7200 1.7000 812.8000 ;
      RECT 0.0000 810.0800 3390.2000 811.7200 ;
      RECT 3384.5000 809.0000 3390.2000 810.0800 ;
      RECT 9.3000 809.0000 3380.9000 810.0800 ;
      RECT 0.0000 809.0000 5.7000 810.0800 ;
      RECT 0.0000 807.3600 3390.2000 809.0000 ;
      RECT 0.0000 807.1400 1.7000 807.3600 ;
      RECT 3388.5000 806.2800 3390.2000 807.3600 ;
      RECT 5.3000 806.2800 3384.9000 807.3600 ;
      RECT 1.1000 806.2800 1.7000 807.1400 ;
      RECT 1.1000 806.2400 3390.2000 806.2800 ;
      RECT 0.0000 804.6400 3390.2000 806.2400 ;
      RECT 3384.5000 803.5600 3390.2000 804.6400 ;
      RECT 9.3000 803.5600 3380.9000 804.6400 ;
      RECT 0.0000 803.5600 5.7000 804.6400 ;
      RECT 0.0000 801.9200 3390.2000 803.5600 ;
      RECT 3388.5000 800.8400 3390.2000 801.9200 ;
      RECT 5.3000 800.8400 3384.9000 801.9200 ;
      RECT 0.0000 800.8400 1.7000 801.9200 ;
      RECT 0.0000 799.2000 3390.2000 800.8400 ;
      RECT 3384.5000 798.1200 3390.2000 799.2000 ;
      RECT 9.3000 798.1200 3380.9000 799.2000 ;
      RECT 0.0000 798.1200 5.7000 799.2000 ;
      RECT 0.0000 796.4800 3390.2000 798.1200 ;
      RECT 3388.5000 795.4000 3390.2000 796.4800 ;
      RECT 5.3000 795.4000 3384.9000 796.4800 ;
      RECT 0.0000 795.4000 1.7000 796.4800 ;
      RECT 0.0000 793.7600 3390.2000 795.4000 ;
      RECT 3384.5000 792.6800 3390.2000 793.7600 ;
      RECT 9.3000 792.6800 3380.9000 793.7600 ;
      RECT 0.0000 792.6800 5.7000 793.7600 ;
      RECT 0.0000 791.0400 3390.2000 792.6800 ;
      RECT 3388.5000 789.9600 3390.2000 791.0400 ;
      RECT 5.3000 789.9600 3384.9000 791.0400 ;
      RECT 0.0000 789.9600 1.7000 791.0400 ;
      RECT 0.0000 788.3200 3390.2000 789.9600 ;
      RECT 3384.5000 787.2400 3390.2000 788.3200 ;
      RECT 9.3000 787.2400 3380.9000 788.3200 ;
      RECT 0.0000 787.2400 5.7000 788.3200 ;
      RECT 0.0000 785.6000 3390.2000 787.2400 ;
      RECT 3388.5000 784.5200 3390.2000 785.6000 ;
      RECT 5.3000 784.5200 3384.9000 785.6000 ;
      RECT 0.0000 784.5200 1.7000 785.6000 ;
      RECT 0.0000 782.8800 3390.2000 784.5200 ;
      RECT 0.0000 782.1300 5.7000 782.8800 ;
      RECT 3384.5000 781.8000 3390.2000 782.8800 ;
      RECT 9.3000 781.8000 3380.9000 782.8800 ;
      RECT 1.1000 781.8000 5.7000 782.1300 ;
      RECT 1.1000 781.2300 3390.2000 781.8000 ;
      RECT 0.0000 780.1600 3390.2000 781.2300 ;
      RECT 3388.5000 779.0800 3390.2000 780.1600 ;
      RECT 5.3000 779.0800 3384.9000 780.1600 ;
      RECT 0.0000 779.0800 1.7000 780.1600 ;
      RECT 0.0000 777.4400 3390.2000 779.0800 ;
      RECT 3384.5000 776.3600 3390.2000 777.4400 ;
      RECT 9.3000 776.3600 3380.9000 777.4400 ;
      RECT 0.0000 776.3600 5.7000 777.4400 ;
      RECT 0.0000 774.7200 3390.2000 776.3600 ;
      RECT 3388.5000 773.6400 3390.2000 774.7200 ;
      RECT 5.3000 773.6400 3384.9000 774.7200 ;
      RECT 0.0000 773.6400 1.7000 774.7200 ;
      RECT 0.0000 772.0000 3390.2000 773.6400 ;
      RECT 3384.5000 770.9200 3390.2000 772.0000 ;
      RECT 9.3000 770.9200 3380.9000 772.0000 ;
      RECT 0.0000 770.9200 5.7000 772.0000 ;
      RECT 0.0000 769.2800 3390.2000 770.9200 ;
      RECT 3388.5000 768.2000 3390.2000 769.2800 ;
      RECT 5.3000 768.2000 3384.9000 769.2800 ;
      RECT 0.0000 768.2000 1.7000 769.2800 ;
      RECT 0.0000 766.5600 3390.2000 768.2000 ;
      RECT 3384.5000 765.4800 3390.2000 766.5600 ;
      RECT 9.3000 765.4800 3380.9000 766.5600 ;
      RECT 0.0000 765.4800 5.7000 766.5600 ;
      RECT 0.0000 763.8400 3390.2000 765.4800 ;
      RECT 3388.5000 762.7600 3390.2000 763.8400 ;
      RECT 5.3000 762.7600 3384.9000 763.8400 ;
      RECT 0.0000 762.7600 1.7000 763.8400 ;
      RECT 0.0000 761.1200 3390.2000 762.7600 ;
      RECT 3384.5000 760.0400 3390.2000 761.1200 ;
      RECT 9.3000 760.0400 3380.9000 761.1200 ;
      RECT 0.0000 760.0400 5.7000 761.1200 ;
      RECT 0.0000 758.4000 3390.2000 760.0400 ;
      RECT 3388.5000 757.3200 3390.2000 758.4000 ;
      RECT 5.3000 757.3200 3384.9000 758.4000 ;
      RECT 0.0000 757.3200 1.7000 758.4000 ;
      RECT 0.0000 757.1200 3390.2000 757.3200 ;
      RECT 1.1000 756.2200 3390.2000 757.1200 ;
      RECT 0.0000 755.6800 3390.2000 756.2200 ;
      RECT 3384.5000 754.6000 3390.2000 755.6800 ;
      RECT 9.3000 754.6000 3380.9000 755.6800 ;
      RECT 0.0000 754.6000 5.7000 755.6800 ;
      RECT 0.0000 752.9600 3390.2000 754.6000 ;
      RECT 3388.5000 751.8800 3390.2000 752.9600 ;
      RECT 5.3000 751.8800 3384.9000 752.9600 ;
      RECT 0.0000 751.8800 1.7000 752.9600 ;
      RECT 0.0000 750.2400 3390.2000 751.8800 ;
      RECT 3384.5000 749.1600 3390.2000 750.2400 ;
      RECT 9.3000 749.1600 3380.9000 750.2400 ;
      RECT 0.0000 749.1600 5.7000 750.2400 ;
      RECT 0.0000 747.5200 3390.2000 749.1600 ;
      RECT 3388.5000 746.4400 3390.2000 747.5200 ;
      RECT 5.3000 746.4400 3384.9000 747.5200 ;
      RECT 0.0000 746.4400 1.7000 747.5200 ;
      RECT 0.0000 744.8000 3390.2000 746.4400 ;
      RECT 3384.5000 743.7200 3390.2000 744.8000 ;
      RECT 9.3000 743.7200 3380.9000 744.8000 ;
      RECT 0.0000 743.7200 5.7000 744.8000 ;
      RECT 0.0000 742.0800 3390.2000 743.7200 ;
      RECT 3388.5000 741.0000 3390.2000 742.0800 ;
      RECT 5.3000 741.0000 3384.9000 742.0800 ;
      RECT 0.0000 741.0000 1.7000 742.0800 ;
      RECT 0.0000 739.3600 3390.2000 741.0000 ;
      RECT 3384.5000 738.2800 3390.2000 739.3600 ;
      RECT 9.3000 738.2800 3380.9000 739.3600 ;
      RECT 0.0000 738.2800 5.7000 739.3600 ;
      RECT 0.0000 736.6400 3390.2000 738.2800 ;
      RECT 3388.5000 735.5600 3390.2000 736.6400 ;
      RECT 5.3000 735.5600 3384.9000 736.6400 ;
      RECT 0.0000 735.5600 1.7000 736.6400 ;
      RECT 0.0000 733.9200 3390.2000 735.5600 ;
      RECT 3384.5000 732.8400 3390.2000 733.9200 ;
      RECT 9.3000 732.8400 3380.9000 733.9200 ;
      RECT 0.0000 732.8400 5.7000 733.9200 ;
      RECT 0.0000 731.5000 3390.2000 732.8400 ;
      RECT 1.1000 731.2000 3390.2000 731.5000 ;
      RECT 1.1000 730.6000 1.7000 731.2000 ;
      RECT 3388.5000 730.1200 3390.2000 731.2000 ;
      RECT 5.3000 730.1200 3384.9000 731.2000 ;
      RECT 0.0000 730.1200 1.7000 730.6000 ;
      RECT 0.0000 728.4800 3390.2000 730.1200 ;
      RECT 3384.5000 727.4000 3390.2000 728.4800 ;
      RECT 9.3000 727.4000 3380.9000 728.4800 ;
      RECT 0.0000 727.4000 5.7000 728.4800 ;
      RECT 0.0000 725.7600 3390.2000 727.4000 ;
      RECT 3388.5000 724.6800 3390.2000 725.7600 ;
      RECT 5.3000 724.6800 3384.9000 725.7600 ;
      RECT 0.0000 724.6800 1.7000 725.7600 ;
      RECT 0.0000 724.1800 3390.2000 724.6800 ;
      RECT 0.0000 723.2800 3389.1000 724.1800 ;
      RECT 0.0000 723.0400 3390.2000 723.2800 ;
      RECT 3384.5000 721.9600 3390.2000 723.0400 ;
      RECT 9.3000 721.9600 3380.9000 723.0400 ;
      RECT 0.0000 721.9600 5.7000 723.0400 ;
      RECT 0.0000 720.3200 3390.2000 721.9600 ;
      RECT 3388.5000 719.2400 3390.2000 720.3200 ;
      RECT 5.3000 719.2400 3384.9000 720.3200 ;
      RECT 0.0000 719.2400 1.7000 720.3200 ;
      RECT 0.0000 717.6000 3390.2000 719.2400 ;
      RECT 3384.5000 716.5200 3390.2000 717.6000 ;
      RECT 9.3000 716.5200 3380.9000 717.6000 ;
      RECT 0.0000 716.5200 5.7000 717.6000 ;
      RECT 0.0000 714.8800 3390.2000 716.5200 ;
      RECT 3388.5000 713.8000 3390.2000 714.8800 ;
      RECT 5.3000 713.8000 3384.9000 714.8800 ;
      RECT 0.0000 713.8000 1.7000 714.8800 ;
      RECT 0.0000 712.1600 3390.2000 713.8000 ;
      RECT 3384.5000 711.0800 3390.2000 712.1600 ;
      RECT 9.3000 711.0800 3380.9000 712.1600 ;
      RECT 0.0000 711.0800 5.7000 712.1600 ;
      RECT 0.0000 709.4400 3390.2000 711.0800 ;
      RECT 3388.5000 708.3600 3390.2000 709.4400 ;
      RECT 5.3000 708.3600 3384.9000 709.4400 ;
      RECT 0.0000 708.3600 1.7000 709.4400 ;
      RECT 0.0000 706.7200 3390.2000 708.3600 ;
      RECT 0.0000 706.4900 5.7000 706.7200 ;
      RECT 3384.5000 705.6400 3390.2000 706.7200 ;
      RECT 9.3000 705.6400 3380.9000 706.7200 ;
      RECT 1.1000 705.6400 5.7000 706.4900 ;
      RECT 1.1000 705.5900 3390.2000 705.6400 ;
      RECT 0.0000 704.0000 3390.2000 705.5900 ;
      RECT 3388.5000 702.9200 3390.2000 704.0000 ;
      RECT 5.3000 702.9200 3384.9000 704.0000 ;
      RECT 0.0000 702.9200 1.7000 704.0000 ;
      RECT 0.0000 701.2800 3390.2000 702.9200 ;
      RECT 3384.5000 700.2000 3390.2000 701.2800 ;
      RECT 9.3000 700.2000 3380.9000 701.2800 ;
      RECT 0.0000 700.2000 5.7000 701.2800 ;
      RECT 0.0000 698.5600 3390.2000 700.2000 ;
      RECT 3388.5000 697.4800 3390.2000 698.5600 ;
      RECT 5.3000 697.4800 3384.9000 698.5600 ;
      RECT 0.0000 697.4800 1.7000 698.5600 ;
      RECT 0.0000 695.8400 3390.2000 697.4800 ;
      RECT 3384.5000 694.7600 3390.2000 695.8400 ;
      RECT 9.3000 694.7600 3380.9000 695.8400 ;
      RECT 0.0000 694.7600 5.7000 695.8400 ;
      RECT 0.0000 693.1200 3390.2000 694.7600 ;
      RECT 3388.5000 692.0400 3390.2000 693.1200 ;
      RECT 5.3000 692.0400 3384.9000 693.1200 ;
      RECT 0.0000 692.0400 1.7000 693.1200 ;
      RECT 0.0000 690.4000 3390.2000 692.0400 ;
      RECT 3384.5000 689.3200 3390.2000 690.4000 ;
      RECT 9.3000 689.3200 3380.9000 690.4000 ;
      RECT 0.0000 689.3200 5.7000 690.4000 ;
      RECT 0.0000 687.6800 3390.2000 689.3200 ;
      RECT 3388.5000 686.6000 3390.2000 687.6800 ;
      RECT 5.3000 686.6000 3384.9000 687.6800 ;
      RECT 0.0000 686.6000 1.7000 687.6800 ;
      RECT 0.0000 684.9600 3390.2000 686.6000 ;
      RECT 3384.5000 683.8800 3390.2000 684.9600 ;
      RECT 9.3000 683.8800 3380.9000 684.9600 ;
      RECT 0.0000 683.8800 5.7000 684.9600 ;
      RECT 0.0000 682.2400 3390.2000 683.8800 ;
      RECT 0.0000 681.4800 1.7000 682.2400 ;
      RECT 3388.5000 681.1600 3390.2000 682.2400 ;
      RECT 5.3000 681.1600 3384.9000 682.2400 ;
      RECT 1.1000 681.1600 1.7000 681.4800 ;
      RECT 1.1000 680.5800 3390.2000 681.1600 ;
      RECT 0.0000 679.5200 3390.2000 680.5800 ;
      RECT 3384.5000 678.4400 3390.2000 679.5200 ;
      RECT 9.3000 678.4400 3380.9000 679.5200 ;
      RECT 0.0000 678.4400 5.7000 679.5200 ;
      RECT 0.0000 676.8000 3390.2000 678.4400 ;
      RECT 3388.5000 675.7200 3390.2000 676.8000 ;
      RECT 5.3000 675.7200 3384.9000 676.8000 ;
      RECT 0.0000 675.7200 1.7000 676.8000 ;
      RECT 0.0000 674.0800 3390.2000 675.7200 ;
      RECT 3384.5000 673.0000 3390.2000 674.0800 ;
      RECT 9.3000 673.0000 3380.9000 674.0800 ;
      RECT 0.0000 673.0000 5.7000 674.0800 ;
      RECT 0.0000 671.3600 3390.2000 673.0000 ;
      RECT 3388.5000 670.2800 3390.2000 671.3600 ;
      RECT 5.3000 670.2800 3384.9000 671.3600 ;
      RECT 0.0000 670.2800 1.7000 671.3600 ;
      RECT 0.0000 668.6400 3390.2000 670.2800 ;
      RECT 3384.5000 667.5600 3390.2000 668.6400 ;
      RECT 9.3000 667.5600 3380.9000 668.6400 ;
      RECT 0.0000 667.5600 5.7000 668.6400 ;
      RECT 0.0000 665.9200 3390.2000 667.5600 ;
      RECT 3388.5000 664.8400 3390.2000 665.9200 ;
      RECT 5.3000 664.8400 3384.9000 665.9200 ;
      RECT 0.0000 664.8400 1.7000 665.9200 ;
      RECT 0.0000 663.2000 3390.2000 664.8400 ;
      RECT 3384.5000 662.1200 3390.2000 663.2000 ;
      RECT 9.3000 662.1200 3380.9000 663.2000 ;
      RECT 0.0000 662.1200 5.7000 663.2000 ;
      RECT 0.0000 660.4800 3390.2000 662.1200 ;
      RECT 3388.5000 659.4000 3390.2000 660.4800 ;
      RECT 5.3000 659.4000 3384.9000 660.4800 ;
      RECT 0.0000 659.4000 1.7000 660.4800 ;
      RECT 0.0000 657.7600 3390.2000 659.4000 ;
      RECT 3384.5000 656.6800 3390.2000 657.7600 ;
      RECT 9.3000 656.6800 3380.9000 657.7600 ;
      RECT 0.0000 656.6800 5.7000 657.7600 ;
      RECT 0.0000 655.8600 3390.2000 656.6800 ;
      RECT 1.1000 655.0400 3390.2000 655.8600 ;
      RECT 1.1000 654.9600 1.7000 655.0400 ;
      RECT 3388.5000 653.9600 3390.2000 655.0400 ;
      RECT 5.3000 653.9600 3384.9000 655.0400 ;
      RECT 0.0000 653.9600 1.7000 654.9600 ;
      RECT 0.0000 652.3200 3390.2000 653.9600 ;
      RECT 3384.5000 651.2400 3390.2000 652.3200 ;
      RECT 9.3000 651.2400 3380.9000 652.3200 ;
      RECT 0.0000 651.2400 5.7000 652.3200 ;
      RECT 0.0000 649.6000 3390.2000 651.2400 ;
      RECT 3388.5000 648.5200 3390.2000 649.6000 ;
      RECT 5.3000 648.5200 3384.9000 649.6000 ;
      RECT 0.0000 648.5200 1.7000 649.6000 ;
      RECT 0.0000 646.8800 3390.2000 648.5200 ;
      RECT 3384.5000 645.8000 3390.2000 646.8800 ;
      RECT 9.3000 645.8000 3380.9000 646.8800 ;
      RECT 0.0000 645.8000 5.7000 646.8800 ;
      RECT 0.0000 644.1600 3390.2000 645.8000 ;
      RECT 3388.5000 643.0800 3390.2000 644.1600 ;
      RECT 5.3000 643.0800 3384.9000 644.1600 ;
      RECT 0.0000 643.0800 1.7000 644.1600 ;
      RECT 0.0000 641.4400 3390.2000 643.0800 ;
      RECT 3384.5000 640.3600 3390.2000 641.4400 ;
      RECT 9.3000 640.3600 3380.9000 641.4400 ;
      RECT 0.0000 640.3600 5.7000 641.4400 ;
      RECT 0.0000 638.7200 3390.2000 640.3600 ;
      RECT 3388.5000 637.6400 3390.2000 638.7200 ;
      RECT 5.3000 637.6400 3384.9000 638.7200 ;
      RECT 0.0000 637.6400 1.7000 638.7200 ;
      RECT 0.0000 636.0000 3390.2000 637.6400 ;
      RECT 3384.5000 634.9200 3390.2000 636.0000 ;
      RECT 9.3000 634.9200 3380.9000 636.0000 ;
      RECT 0.0000 634.9200 5.7000 636.0000 ;
      RECT 0.0000 633.2800 3390.2000 634.9200 ;
      RECT 3388.5000 632.2000 3390.2000 633.2800 ;
      RECT 5.3000 632.2000 3384.9000 633.2800 ;
      RECT 0.0000 632.2000 1.7000 633.2800 ;
      RECT 0.0000 630.8500 3390.2000 632.2000 ;
      RECT 1.1000 630.5600 3390.2000 630.8500 ;
      RECT 1.1000 629.9500 5.7000 630.5600 ;
      RECT 3384.5000 629.4800 3390.2000 630.5600 ;
      RECT 9.3000 629.4800 3380.9000 630.5600 ;
      RECT 0.0000 629.4800 5.7000 629.9500 ;
      RECT 0.0000 627.8400 3390.2000 629.4800 ;
      RECT 3388.5000 626.7600 3390.2000 627.8400 ;
      RECT 5.3000 626.7600 3384.9000 627.8400 ;
      RECT 0.0000 626.7600 1.7000 627.8400 ;
      RECT 0.0000 625.1200 3390.2000 626.7600 ;
      RECT 3384.5000 624.0400 3390.2000 625.1200 ;
      RECT 9.3000 624.0400 3380.9000 625.1200 ;
      RECT 0.0000 624.0400 5.7000 625.1200 ;
      RECT 0.0000 622.4000 3390.2000 624.0400 ;
      RECT 3388.5000 621.3200 3390.2000 622.4000 ;
      RECT 5.3000 621.3200 3384.9000 622.4000 ;
      RECT 0.0000 621.3200 1.7000 622.4000 ;
      RECT 0.0000 619.8700 3390.2000 621.3200 ;
      RECT 0.0000 619.6800 3389.1000 619.8700 ;
      RECT 3384.5000 618.9700 3389.1000 619.6800 ;
      RECT 3384.5000 618.6000 3390.2000 618.9700 ;
      RECT 9.3000 618.6000 3380.9000 619.6800 ;
      RECT 0.0000 618.6000 5.7000 619.6800 ;
      RECT 0.0000 616.9600 3390.2000 618.6000 ;
      RECT 3388.5000 615.8800 3390.2000 616.9600 ;
      RECT 5.3000 615.8800 3384.9000 616.9600 ;
      RECT 0.0000 615.8800 1.7000 616.9600 ;
      RECT 0.0000 614.2400 3390.2000 615.8800 ;
      RECT 3384.5000 613.1600 3390.2000 614.2400 ;
      RECT 9.3000 613.1600 3380.9000 614.2400 ;
      RECT 0.0000 613.1600 5.7000 614.2400 ;
      RECT 0.0000 611.5200 3390.2000 613.1600 ;
      RECT 3388.5000 610.4400 3390.2000 611.5200 ;
      RECT 5.3000 610.4400 3384.9000 611.5200 ;
      RECT 0.0000 610.4400 1.7000 611.5200 ;
      RECT 0.0000 608.8000 3390.2000 610.4400 ;
      RECT 3384.5000 607.7200 3390.2000 608.8000 ;
      RECT 9.3000 607.7200 3380.9000 608.8000 ;
      RECT 0.0000 607.7200 5.7000 608.8000 ;
      RECT 0.0000 606.0800 3390.2000 607.7200 ;
      RECT 0.0000 605.8400 1.7000 606.0800 ;
      RECT 3388.5000 605.0000 3390.2000 606.0800 ;
      RECT 5.3000 605.0000 3384.9000 606.0800 ;
      RECT 1.1000 605.0000 1.7000 605.8400 ;
      RECT 1.1000 604.9400 3390.2000 605.0000 ;
      RECT 0.0000 603.3600 3390.2000 604.9400 ;
      RECT 3384.5000 602.2800 3390.2000 603.3600 ;
      RECT 9.3000 602.2800 3380.9000 603.3600 ;
      RECT 0.0000 602.2800 5.7000 603.3600 ;
      RECT 0.0000 600.6400 3390.2000 602.2800 ;
      RECT 3388.5000 599.5600 3390.2000 600.6400 ;
      RECT 5.3000 599.5600 3384.9000 600.6400 ;
      RECT 0.0000 599.5600 1.7000 600.6400 ;
      RECT 0.0000 597.9200 3390.2000 599.5600 ;
      RECT 3384.5000 596.8400 3390.2000 597.9200 ;
      RECT 9.3000 596.8400 3380.9000 597.9200 ;
      RECT 0.0000 596.8400 5.7000 597.9200 ;
      RECT 0.0000 595.2000 3390.2000 596.8400 ;
      RECT 3388.5000 594.1200 3390.2000 595.2000 ;
      RECT 5.3000 594.1200 3384.9000 595.2000 ;
      RECT 0.0000 594.1200 1.7000 595.2000 ;
      RECT 0.0000 592.4800 3390.2000 594.1200 ;
      RECT 3384.5000 591.4000 3390.2000 592.4800 ;
      RECT 9.3000 591.4000 3380.9000 592.4800 ;
      RECT 0.0000 591.4000 5.7000 592.4800 ;
      RECT 0.0000 589.7600 3390.2000 591.4000 ;
      RECT 3388.5000 588.6800 3390.2000 589.7600 ;
      RECT 5.3000 588.6800 3384.9000 589.7600 ;
      RECT 0.0000 588.6800 1.7000 589.7600 ;
      RECT 0.0000 587.0400 3390.2000 588.6800 ;
      RECT 3384.5000 585.9600 3390.2000 587.0400 ;
      RECT 9.3000 585.9600 3380.9000 587.0400 ;
      RECT 0.0000 585.9600 5.7000 587.0400 ;
      RECT 0.0000 584.3200 3390.2000 585.9600 ;
      RECT 3388.5000 583.2400 3390.2000 584.3200 ;
      RECT 5.3000 583.2400 3384.9000 584.3200 ;
      RECT 0.0000 583.2400 1.7000 584.3200 ;
      RECT 0.0000 581.6000 3390.2000 583.2400 ;
      RECT 3384.5000 580.5200 3390.2000 581.6000 ;
      RECT 9.3000 580.5200 3380.9000 581.6000 ;
      RECT 0.0000 580.5200 5.7000 581.6000 ;
      RECT 0.0000 580.2200 3390.2000 580.5200 ;
      RECT 1.1000 579.3200 3390.2000 580.2200 ;
      RECT 0.0000 578.8800 3390.2000 579.3200 ;
      RECT 3388.5000 577.8000 3390.2000 578.8800 ;
      RECT 5.3000 577.8000 3384.9000 578.8800 ;
      RECT 0.0000 577.8000 1.7000 578.8800 ;
      RECT 0.0000 576.1600 3390.2000 577.8000 ;
      RECT 3384.5000 575.0800 3390.2000 576.1600 ;
      RECT 9.3000 575.0800 3380.9000 576.1600 ;
      RECT 0.0000 575.0800 5.7000 576.1600 ;
      RECT 0.0000 573.4400 3390.2000 575.0800 ;
      RECT 3388.5000 572.3600 3390.2000 573.4400 ;
      RECT 5.3000 572.3600 3384.9000 573.4400 ;
      RECT 0.0000 572.3600 1.7000 573.4400 ;
      RECT 0.0000 570.7200 3390.2000 572.3600 ;
      RECT 3384.5000 569.6400 3390.2000 570.7200 ;
      RECT 9.3000 569.6400 3380.9000 570.7200 ;
      RECT 0.0000 569.6400 5.7000 570.7200 ;
      RECT 0.0000 568.0000 3390.2000 569.6400 ;
      RECT 3388.5000 566.9200 3390.2000 568.0000 ;
      RECT 5.3000 566.9200 3384.9000 568.0000 ;
      RECT 0.0000 566.9200 1.7000 568.0000 ;
      RECT 0.0000 565.2800 3390.2000 566.9200 ;
      RECT 3384.5000 564.2000 3390.2000 565.2800 ;
      RECT 9.3000 564.2000 3380.9000 565.2800 ;
      RECT 0.0000 564.2000 5.7000 565.2800 ;
      RECT 0.0000 562.5600 3390.2000 564.2000 ;
      RECT 3388.5000 561.4800 3390.2000 562.5600 ;
      RECT 5.3000 561.4800 3384.9000 562.5600 ;
      RECT 0.0000 561.4800 1.7000 562.5600 ;
      RECT 0.0000 559.8400 3390.2000 561.4800 ;
      RECT 3384.5000 558.7600 3390.2000 559.8400 ;
      RECT 9.3000 558.7600 3380.9000 559.8400 ;
      RECT 0.0000 558.7600 5.7000 559.8400 ;
      RECT 0.0000 557.1200 3390.2000 558.7600 ;
      RECT 3388.5000 556.0400 3390.2000 557.1200 ;
      RECT 5.3000 556.0400 3384.9000 557.1200 ;
      RECT 0.0000 556.0400 1.7000 557.1200 ;
      RECT 0.0000 555.2100 3390.2000 556.0400 ;
      RECT 1.1000 554.4000 3390.2000 555.2100 ;
      RECT 1.1000 554.3100 5.7000 554.4000 ;
      RECT 3384.5000 553.3200 3390.2000 554.4000 ;
      RECT 9.3000 553.3200 3380.9000 554.4000 ;
      RECT 0.0000 553.3200 5.7000 554.3100 ;
      RECT 0.0000 551.6800 3390.2000 553.3200 ;
      RECT 3388.5000 550.6000 3390.2000 551.6800 ;
      RECT 5.3000 550.6000 3384.9000 551.6800 ;
      RECT 0.0000 550.6000 1.7000 551.6800 ;
      RECT 0.0000 548.9600 3390.2000 550.6000 ;
      RECT 3384.5000 547.8800 3390.2000 548.9600 ;
      RECT 9.3000 547.8800 3380.9000 548.9600 ;
      RECT 0.0000 547.8800 5.7000 548.9600 ;
      RECT 0.0000 546.2400 3390.2000 547.8800 ;
      RECT 3388.5000 545.1600 3390.2000 546.2400 ;
      RECT 5.3000 545.1600 3384.9000 546.2400 ;
      RECT 0.0000 545.1600 1.7000 546.2400 ;
      RECT 0.0000 543.5200 3390.2000 545.1600 ;
      RECT 3384.5000 542.4400 3390.2000 543.5200 ;
      RECT 9.3000 542.4400 3380.9000 543.5200 ;
      RECT 0.0000 542.4400 5.7000 543.5200 ;
      RECT 0.0000 540.8000 3390.2000 542.4400 ;
      RECT 3388.5000 539.7200 3390.2000 540.8000 ;
      RECT 5.3000 539.7200 3384.9000 540.8000 ;
      RECT 0.0000 539.7200 1.7000 540.8000 ;
      RECT 0.0000 538.0800 3390.2000 539.7200 ;
      RECT 3384.5000 537.0000 3390.2000 538.0800 ;
      RECT 9.3000 537.0000 3380.9000 538.0800 ;
      RECT 0.0000 537.0000 5.7000 538.0800 ;
      RECT 0.0000 535.3600 3390.2000 537.0000 ;
      RECT 3388.5000 534.2800 3390.2000 535.3600 ;
      RECT 5.3000 534.2800 3384.9000 535.3600 ;
      RECT 0.0000 534.2800 1.7000 535.3600 ;
      RECT 0.0000 532.6400 3390.2000 534.2800 ;
      RECT 3384.5000 531.5600 3390.2000 532.6400 ;
      RECT 9.3000 531.5600 3380.9000 532.6400 ;
      RECT 0.0000 531.5600 5.7000 532.6400 ;
      RECT 0.0000 530.2000 3390.2000 531.5600 ;
      RECT 1.1000 529.9200 3390.2000 530.2000 ;
      RECT 1.1000 529.3000 1.7000 529.9200 ;
      RECT 3388.5000 528.8400 3390.2000 529.9200 ;
      RECT 5.3000 528.8400 3384.9000 529.9200 ;
      RECT 0.0000 528.8400 1.7000 529.3000 ;
      RECT 0.0000 527.2000 3390.2000 528.8400 ;
      RECT 3384.5000 526.1200 3390.2000 527.2000 ;
      RECT 9.3000 526.1200 3380.9000 527.2000 ;
      RECT 0.0000 526.1200 5.7000 527.2000 ;
      RECT 0.0000 524.4800 3390.2000 526.1200 ;
      RECT 3388.5000 523.4000 3390.2000 524.4800 ;
      RECT 5.3000 523.4000 3384.9000 524.4800 ;
      RECT 0.0000 523.4000 1.7000 524.4800 ;
      RECT 0.0000 521.7600 3390.2000 523.4000 ;
      RECT 3384.5000 520.6800 3390.2000 521.7600 ;
      RECT 9.3000 520.6800 3380.9000 521.7600 ;
      RECT 0.0000 520.6800 5.7000 521.7600 ;
      RECT 0.0000 519.0400 3390.2000 520.6800 ;
      RECT 3388.5000 517.9600 3390.2000 519.0400 ;
      RECT 5.3000 517.9600 3384.9000 519.0400 ;
      RECT 0.0000 517.9600 1.7000 519.0400 ;
      RECT 0.0000 516.3200 3390.2000 517.9600 ;
      RECT 3384.5000 516.1700 3390.2000 516.3200 ;
      RECT 3384.5000 515.2700 3389.1000 516.1700 ;
      RECT 3384.5000 515.2400 3390.2000 515.2700 ;
      RECT 9.3000 515.2400 3380.9000 516.3200 ;
      RECT 0.0000 515.2400 5.7000 516.3200 ;
      RECT 0.0000 513.6000 3390.2000 515.2400 ;
      RECT 3388.5000 512.5200 3390.2000 513.6000 ;
      RECT 5.3000 512.5200 3384.9000 513.6000 ;
      RECT 0.0000 512.5200 1.7000 513.6000 ;
      RECT 0.0000 510.8800 3390.2000 512.5200 ;
      RECT 3384.5000 509.8000 3390.2000 510.8800 ;
      RECT 9.3000 509.8000 3380.9000 510.8800 ;
      RECT 0.0000 509.8000 5.7000 510.8800 ;
      RECT 0.0000 508.1600 3390.2000 509.8000 ;
      RECT 3388.5000 507.0800 3390.2000 508.1600 ;
      RECT 5.3000 507.0800 3384.9000 508.1600 ;
      RECT 0.0000 507.0800 1.7000 508.1600 ;
      RECT 0.0000 505.4400 3390.2000 507.0800 ;
      RECT 0.0000 504.5800 5.7000 505.4400 ;
      RECT 3384.5000 504.3600 3390.2000 505.4400 ;
      RECT 9.3000 504.3600 3380.9000 505.4400 ;
      RECT 1.1000 504.3600 5.7000 504.5800 ;
      RECT 1.1000 503.6800 3390.2000 504.3600 ;
      RECT 0.0000 502.7200 3390.2000 503.6800 ;
      RECT 3388.5000 501.6400 3390.2000 502.7200 ;
      RECT 5.3000 501.6400 3384.9000 502.7200 ;
      RECT 0.0000 501.6400 1.7000 502.7200 ;
      RECT 0.0000 500.0000 3390.2000 501.6400 ;
      RECT 3384.5000 498.9200 3390.2000 500.0000 ;
      RECT 9.3000 498.9200 3380.9000 500.0000 ;
      RECT 0.0000 498.9200 5.7000 500.0000 ;
      RECT 0.0000 497.2800 3390.2000 498.9200 ;
      RECT 3388.5000 496.2000 3390.2000 497.2800 ;
      RECT 5.3000 496.2000 3384.9000 497.2800 ;
      RECT 0.0000 496.2000 1.7000 497.2800 ;
      RECT 0.0000 494.5600 3390.2000 496.2000 ;
      RECT 3384.5000 493.4800 3390.2000 494.5600 ;
      RECT 9.3000 493.4800 3380.9000 494.5600 ;
      RECT 0.0000 493.4800 5.7000 494.5600 ;
      RECT 0.0000 491.8400 3390.2000 493.4800 ;
      RECT 3388.5000 490.7600 3390.2000 491.8400 ;
      RECT 5.3000 490.7600 3384.9000 491.8400 ;
      RECT 0.0000 490.7600 1.7000 491.8400 ;
      RECT 0.0000 489.1200 3390.2000 490.7600 ;
      RECT 3384.5000 488.0400 3390.2000 489.1200 ;
      RECT 9.3000 488.0400 3380.9000 489.1200 ;
      RECT 0.0000 488.0400 5.7000 489.1200 ;
      RECT 0.0000 486.4000 3390.2000 488.0400 ;
      RECT 3388.5000 485.3200 3390.2000 486.4000 ;
      RECT 5.3000 485.3200 3384.9000 486.4000 ;
      RECT 0.0000 485.3200 1.7000 486.4000 ;
      RECT 0.0000 483.6800 3390.2000 485.3200 ;
      RECT 3384.5000 482.6000 3390.2000 483.6800 ;
      RECT 9.3000 482.6000 3380.9000 483.6800 ;
      RECT 0.0000 482.6000 5.7000 483.6800 ;
      RECT 0.0000 480.9600 3390.2000 482.6000 ;
      RECT 3388.5000 479.8800 3390.2000 480.9600 ;
      RECT 5.3000 479.8800 3384.9000 480.9600 ;
      RECT 0.0000 479.8800 1.7000 480.9600 ;
      RECT 0.0000 479.5700 3390.2000 479.8800 ;
      RECT 1.1000 478.6700 3390.2000 479.5700 ;
      RECT 0.0000 478.2400 3390.2000 478.6700 ;
      RECT 3384.5000 477.1600 3390.2000 478.2400 ;
      RECT 9.3000 477.1600 3380.9000 478.2400 ;
      RECT 0.0000 477.1600 5.7000 478.2400 ;
      RECT 0.0000 475.5200 3390.2000 477.1600 ;
      RECT 3388.5000 474.4400 3390.2000 475.5200 ;
      RECT 5.3000 474.4400 3384.9000 475.5200 ;
      RECT 0.0000 474.4400 1.7000 475.5200 ;
      RECT 0.0000 472.8000 3390.2000 474.4400 ;
      RECT 3384.5000 471.7200 3390.2000 472.8000 ;
      RECT 9.3000 471.7200 3380.9000 472.8000 ;
      RECT 0.0000 471.7200 5.7000 472.8000 ;
      RECT 0.0000 470.0800 3390.2000 471.7200 ;
      RECT 3388.5000 469.0000 3390.2000 470.0800 ;
      RECT 5.3000 469.0000 3384.9000 470.0800 ;
      RECT 0.0000 469.0000 1.7000 470.0800 ;
      RECT 0.0000 467.3600 3390.2000 469.0000 ;
      RECT 3384.5000 466.2800 3390.2000 467.3600 ;
      RECT 9.3000 466.2800 3380.9000 467.3600 ;
      RECT 0.0000 466.2800 5.7000 467.3600 ;
      RECT 0.0000 464.6400 3390.2000 466.2800 ;
      RECT 3388.5000 463.5600 3390.2000 464.6400 ;
      RECT 5.3000 463.5600 3384.9000 464.6400 ;
      RECT 0.0000 463.5600 1.7000 464.6400 ;
      RECT 0.0000 461.9200 3390.2000 463.5600 ;
      RECT 3384.5000 460.8400 3390.2000 461.9200 ;
      RECT 9.3000 460.8400 3380.9000 461.9200 ;
      RECT 0.0000 460.8400 5.7000 461.9200 ;
      RECT 0.0000 459.2000 3390.2000 460.8400 ;
      RECT 3388.5000 458.1200 3390.2000 459.2000 ;
      RECT 5.3000 458.1200 3384.9000 459.2000 ;
      RECT 0.0000 458.1200 1.7000 459.2000 ;
      RECT 0.0000 456.4800 3390.2000 458.1200 ;
      RECT 3384.5000 455.4000 3390.2000 456.4800 ;
      RECT 9.3000 455.4000 3380.9000 456.4800 ;
      RECT 0.0000 455.4000 5.7000 456.4800 ;
      RECT 0.0000 453.9500 3390.2000 455.4000 ;
      RECT 1.1000 453.7600 3390.2000 453.9500 ;
      RECT 1.1000 453.0500 1.7000 453.7600 ;
      RECT 3388.5000 452.6800 3390.2000 453.7600 ;
      RECT 5.3000 452.6800 3384.9000 453.7600 ;
      RECT 0.0000 452.6800 1.7000 453.0500 ;
      RECT 0.0000 451.0400 3390.2000 452.6800 ;
      RECT 3384.5000 449.9600 3390.2000 451.0400 ;
      RECT 9.3000 449.9600 3380.9000 451.0400 ;
      RECT 0.0000 449.9600 5.7000 451.0400 ;
      RECT 0.0000 448.3200 3390.2000 449.9600 ;
      RECT 3388.5000 447.2400 3390.2000 448.3200 ;
      RECT 5.3000 447.2400 3384.9000 448.3200 ;
      RECT 0.0000 447.2400 1.7000 448.3200 ;
      RECT 0.0000 445.6000 3390.2000 447.2400 ;
      RECT 3384.5000 444.5200 3390.2000 445.6000 ;
      RECT 9.3000 444.5200 3380.9000 445.6000 ;
      RECT 0.0000 444.5200 5.7000 445.6000 ;
      RECT 0.0000 442.8800 3390.2000 444.5200 ;
      RECT 3388.5000 441.8000 3390.2000 442.8800 ;
      RECT 5.3000 441.8000 3384.9000 442.8800 ;
      RECT 0.0000 441.8000 1.7000 442.8800 ;
      RECT 0.0000 440.1600 3390.2000 441.8000 ;
      RECT 3384.5000 439.0800 3390.2000 440.1600 ;
      RECT 9.3000 439.0800 3380.9000 440.1600 ;
      RECT 0.0000 439.0800 5.7000 440.1600 ;
      RECT 0.0000 437.4400 3390.2000 439.0800 ;
      RECT 3388.5000 436.3600 3390.2000 437.4400 ;
      RECT 5.3000 436.3600 3384.9000 437.4400 ;
      RECT 0.0000 436.3600 1.7000 437.4400 ;
      RECT 0.0000 434.7200 3390.2000 436.3600 ;
      RECT 3384.5000 433.6400 3390.2000 434.7200 ;
      RECT 9.3000 433.6400 3380.9000 434.7200 ;
      RECT 0.0000 433.6400 5.7000 434.7200 ;
      RECT 0.0000 432.0000 3390.2000 433.6400 ;
      RECT 3388.5000 430.9200 3390.2000 432.0000 ;
      RECT 5.3000 430.9200 3384.9000 432.0000 ;
      RECT 0.0000 430.9200 1.7000 432.0000 ;
      RECT 0.0000 429.2800 3390.2000 430.9200 ;
      RECT 0.0000 428.9400 5.7000 429.2800 ;
      RECT 3384.5000 428.2000 3390.2000 429.2800 ;
      RECT 9.3000 428.2000 3380.9000 429.2800 ;
      RECT 1.1000 428.2000 5.7000 428.9400 ;
      RECT 1.1000 428.0400 3390.2000 428.2000 ;
      RECT 0.0000 426.5600 3390.2000 428.0400 ;
      RECT 3388.5000 425.4800 3390.2000 426.5600 ;
      RECT 5.3000 425.4800 3384.9000 426.5600 ;
      RECT 0.0000 425.4800 1.7000 426.5600 ;
      RECT 0.0000 423.8400 3390.2000 425.4800 ;
      RECT 3384.5000 422.7600 3390.2000 423.8400 ;
      RECT 9.3000 422.7600 3380.9000 423.8400 ;
      RECT 0.0000 422.7600 5.7000 423.8400 ;
      RECT 0.0000 421.1200 3390.2000 422.7600 ;
      RECT 3388.5000 420.0400 3390.2000 421.1200 ;
      RECT 5.3000 420.0400 3384.9000 421.1200 ;
      RECT 0.0000 420.0400 1.7000 421.1200 ;
      RECT 0.0000 418.4000 3390.2000 420.0400 ;
      RECT 3384.5000 417.3200 3390.2000 418.4000 ;
      RECT 9.3000 417.3200 3380.9000 418.4000 ;
      RECT 0.0000 417.3200 5.7000 418.4000 ;
      RECT 0.0000 415.6800 3390.2000 417.3200 ;
      RECT 3388.5000 414.6000 3390.2000 415.6800 ;
      RECT 5.3000 414.6000 3384.9000 415.6800 ;
      RECT 0.0000 414.6000 1.7000 415.6800 ;
      RECT 0.0000 412.9600 3390.2000 414.6000 ;
      RECT 3384.5000 412.4700 3390.2000 412.9600 ;
      RECT 3384.5000 411.8800 3389.1000 412.4700 ;
      RECT 9.3000 411.8800 3380.9000 412.9600 ;
      RECT 0.0000 411.8800 5.7000 412.9600 ;
      RECT 0.0000 411.5700 3389.1000 411.8800 ;
      RECT 0.0000 410.2400 3390.2000 411.5700 ;
      RECT 3388.5000 409.1600 3390.2000 410.2400 ;
      RECT 5.3000 409.1600 3384.9000 410.2400 ;
      RECT 0.0000 409.1600 1.7000 410.2400 ;
      RECT 0.0000 407.5200 3390.2000 409.1600 ;
      RECT 3384.5000 406.4400 3390.2000 407.5200 ;
      RECT 9.3000 406.4400 3380.9000 407.5200 ;
      RECT 0.0000 406.4400 5.7000 407.5200 ;
      RECT 0.0000 404.8000 3390.2000 406.4400 ;
      RECT 0.0000 403.9300 1.7000 404.8000 ;
      RECT 3388.5000 403.7200 3390.2000 404.8000 ;
      RECT 5.3000 403.7200 3384.9000 404.8000 ;
      RECT 1.1000 403.7200 1.7000 403.9300 ;
      RECT 1.1000 403.0300 3390.2000 403.7200 ;
      RECT 0.0000 402.0800 3390.2000 403.0300 ;
      RECT 3384.5000 401.0000 3390.2000 402.0800 ;
      RECT 9.3000 401.0000 3380.9000 402.0800 ;
      RECT 0.0000 401.0000 5.7000 402.0800 ;
      RECT 0.0000 399.3600 3390.2000 401.0000 ;
      RECT 3388.5000 398.2800 3390.2000 399.3600 ;
      RECT 5.3000 398.2800 3384.9000 399.3600 ;
      RECT 0.0000 398.2800 1.7000 399.3600 ;
      RECT 0.0000 396.6400 3390.2000 398.2800 ;
      RECT 3384.5000 395.5600 3390.2000 396.6400 ;
      RECT 9.3000 395.5600 3380.9000 396.6400 ;
      RECT 0.0000 395.5600 5.7000 396.6400 ;
      RECT 0.0000 393.9200 3390.2000 395.5600 ;
      RECT 3388.5000 392.8400 3390.2000 393.9200 ;
      RECT 5.3000 392.8400 3384.9000 393.9200 ;
      RECT 0.0000 392.8400 1.7000 393.9200 ;
      RECT 0.0000 391.2000 3390.2000 392.8400 ;
      RECT 3384.5000 390.1200 3390.2000 391.2000 ;
      RECT 9.3000 390.1200 3380.9000 391.2000 ;
      RECT 0.0000 390.1200 5.7000 391.2000 ;
      RECT 0.0000 388.4800 3390.2000 390.1200 ;
      RECT 3388.5000 387.4000 3390.2000 388.4800 ;
      RECT 5.3000 387.4000 3384.9000 388.4800 ;
      RECT 0.0000 387.4000 1.7000 388.4800 ;
      RECT 0.0000 385.7600 3390.2000 387.4000 ;
      RECT 3384.5000 384.6800 3390.2000 385.7600 ;
      RECT 9.3000 384.6800 3380.9000 385.7600 ;
      RECT 0.0000 384.6800 5.7000 385.7600 ;
      RECT 0.0000 383.0400 3390.2000 384.6800 ;
      RECT 3388.5000 381.9600 3390.2000 383.0400 ;
      RECT 5.3000 381.9600 3384.9000 383.0400 ;
      RECT 0.0000 381.9600 1.7000 383.0400 ;
      RECT 0.0000 380.3200 3390.2000 381.9600 ;
      RECT 3384.5000 379.2400 3390.2000 380.3200 ;
      RECT 9.3000 379.2400 3380.9000 380.3200 ;
      RECT 0.0000 379.2400 5.7000 380.3200 ;
      RECT 0.0000 378.3100 3390.2000 379.2400 ;
      RECT 1.1000 377.6000 3390.2000 378.3100 ;
      RECT 1.1000 377.4100 1.7000 377.6000 ;
      RECT 3388.5000 376.5200 3390.2000 377.6000 ;
      RECT 5.3000 376.5200 3384.9000 377.6000 ;
      RECT 0.0000 376.5200 1.7000 377.4100 ;
      RECT 0.0000 374.8800 3390.2000 376.5200 ;
      RECT 3384.5000 373.8000 3390.2000 374.8800 ;
      RECT 9.3000 373.8000 3380.9000 374.8800 ;
      RECT 0.0000 373.8000 5.7000 374.8800 ;
      RECT 0.0000 372.1600 3390.2000 373.8000 ;
      RECT 3388.5000 371.0800 3390.2000 372.1600 ;
      RECT 5.3000 371.0800 3384.9000 372.1600 ;
      RECT 0.0000 371.0800 1.7000 372.1600 ;
      RECT 0.0000 369.4400 3390.2000 371.0800 ;
      RECT 3384.5000 368.3600 3390.2000 369.4400 ;
      RECT 9.3000 368.3600 3380.9000 369.4400 ;
      RECT 0.0000 368.3600 5.7000 369.4400 ;
      RECT 0.0000 366.7200 3390.2000 368.3600 ;
      RECT 3388.5000 365.6400 3390.2000 366.7200 ;
      RECT 5.3000 365.6400 3384.9000 366.7200 ;
      RECT 0.0000 365.6400 1.7000 366.7200 ;
      RECT 0.0000 364.0000 3390.2000 365.6400 ;
      RECT 3384.5000 362.9200 3390.2000 364.0000 ;
      RECT 9.3000 362.9200 3380.9000 364.0000 ;
      RECT 0.0000 362.9200 5.7000 364.0000 ;
      RECT 0.0000 361.2800 3390.2000 362.9200 ;
      RECT 3388.5000 360.2000 3390.2000 361.2800 ;
      RECT 5.3000 360.2000 3384.9000 361.2800 ;
      RECT 0.0000 360.2000 1.7000 361.2800 ;
      RECT 0.0000 358.5600 3390.2000 360.2000 ;
      RECT 3384.5000 357.4800 3390.2000 358.5600 ;
      RECT 9.3000 357.4800 3380.9000 358.5600 ;
      RECT 0.0000 357.4800 5.7000 358.5600 ;
      RECT 0.0000 355.8400 3390.2000 357.4800 ;
      RECT 3388.5000 354.7600 3390.2000 355.8400 ;
      RECT 5.3000 354.7600 3384.9000 355.8400 ;
      RECT 0.0000 354.7600 1.7000 355.8400 ;
      RECT 0.0000 353.3000 3390.2000 354.7600 ;
      RECT 1.1000 353.1200 3390.2000 353.3000 ;
      RECT 1.1000 352.4000 5.7000 353.1200 ;
      RECT 3384.5000 352.0400 3390.2000 353.1200 ;
      RECT 9.3000 352.0400 3380.9000 353.1200 ;
      RECT 0.0000 352.0400 5.7000 352.4000 ;
      RECT 0.0000 350.4000 3390.2000 352.0400 ;
      RECT 3388.5000 349.3200 3390.2000 350.4000 ;
      RECT 5.3000 349.3200 3384.9000 350.4000 ;
      RECT 0.0000 349.3200 1.7000 350.4000 ;
      RECT 0.0000 347.6800 3390.2000 349.3200 ;
      RECT 3384.5000 346.6000 3390.2000 347.6800 ;
      RECT 9.3000 346.6000 3380.9000 347.6800 ;
      RECT 0.0000 346.6000 5.7000 347.6800 ;
      RECT 0.0000 344.9600 3390.2000 346.6000 ;
      RECT 3388.5000 343.8800 3390.2000 344.9600 ;
      RECT 5.3000 343.8800 3384.9000 344.9600 ;
      RECT 0.0000 343.8800 1.7000 344.9600 ;
      RECT 0.0000 342.2400 3390.2000 343.8800 ;
      RECT 3384.5000 341.1600 3390.2000 342.2400 ;
      RECT 9.3000 341.1600 3380.9000 342.2400 ;
      RECT 0.0000 341.1600 5.7000 342.2400 ;
      RECT 0.0000 339.5200 3390.2000 341.1600 ;
      RECT 3388.5000 338.4400 3390.2000 339.5200 ;
      RECT 5.3000 338.4400 3384.9000 339.5200 ;
      RECT 0.0000 338.4400 1.7000 339.5200 ;
      RECT 0.0000 336.8000 3390.2000 338.4400 ;
      RECT 3384.5000 335.7200 3390.2000 336.8000 ;
      RECT 9.3000 335.7200 3380.9000 336.8000 ;
      RECT 0.0000 335.7200 5.7000 336.8000 ;
      RECT 0.0000 334.0800 3390.2000 335.7200 ;
      RECT 3388.5000 333.0000 3390.2000 334.0800 ;
      RECT 5.3000 333.0000 3384.9000 334.0800 ;
      RECT 0.0000 333.0000 1.7000 334.0800 ;
      RECT 0.0000 331.3600 3390.2000 333.0000 ;
      RECT 3384.5000 330.2800 3390.2000 331.3600 ;
      RECT 9.3000 330.2800 3380.9000 331.3600 ;
      RECT 0.0000 330.2800 5.7000 331.3600 ;
      RECT 0.0000 328.6400 3390.2000 330.2800 ;
      RECT 0.0000 328.2900 1.7000 328.6400 ;
      RECT 3388.5000 327.5600 3390.2000 328.6400 ;
      RECT 5.3000 327.5600 3384.9000 328.6400 ;
      RECT 1.1000 327.5600 1.7000 328.2900 ;
      RECT 1.1000 327.3900 3390.2000 327.5600 ;
      RECT 0.0000 325.9200 3390.2000 327.3900 ;
      RECT 3384.5000 324.8400 3390.2000 325.9200 ;
      RECT 9.3000 324.8400 3380.9000 325.9200 ;
      RECT 0.0000 324.8400 5.7000 325.9200 ;
      RECT 0.0000 323.2000 3390.2000 324.8400 ;
      RECT 3388.5000 322.1200 3390.2000 323.2000 ;
      RECT 5.3000 322.1200 3384.9000 323.2000 ;
      RECT 0.0000 322.1200 1.7000 323.2000 ;
      RECT 0.0000 320.4800 3390.2000 322.1200 ;
      RECT 3384.5000 319.4000 3390.2000 320.4800 ;
      RECT 9.3000 319.4000 3380.9000 320.4800 ;
      RECT 0.0000 319.4000 5.7000 320.4800 ;
      RECT 0.0000 317.7600 3390.2000 319.4000 ;
      RECT 3388.5000 316.6800 3390.2000 317.7600 ;
      RECT 5.3000 316.6800 3384.9000 317.7600 ;
      RECT 0.0000 316.6800 1.7000 317.7600 ;
      RECT 0.0000 315.0400 3390.2000 316.6800 ;
      RECT 3384.5000 313.9600 3390.2000 315.0400 ;
      RECT 9.3000 313.9600 3380.9000 315.0400 ;
      RECT 0.0000 313.9600 5.7000 315.0400 ;
      RECT 0.0000 312.3200 3390.2000 313.9600 ;
      RECT 3388.5000 311.2400 3390.2000 312.3200 ;
      RECT 5.3000 311.2400 3384.9000 312.3200 ;
      RECT 0.0000 311.2400 1.7000 312.3200 ;
      RECT 0.0000 309.6000 3390.2000 311.2400 ;
      RECT 3384.5000 308.7700 3390.2000 309.6000 ;
      RECT 3384.5000 308.5200 3389.1000 308.7700 ;
      RECT 9.3000 308.5200 3380.9000 309.6000 ;
      RECT 0.0000 308.5200 5.7000 309.6000 ;
      RECT 0.0000 307.8700 3389.1000 308.5200 ;
      RECT 0.0000 306.8800 3390.2000 307.8700 ;
      RECT 3388.5000 305.8000 3390.2000 306.8800 ;
      RECT 5.3000 305.8000 3384.9000 306.8800 ;
      RECT 0.0000 305.8000 1.7000 306.8800 ;
      RECT 0.0000 304.1600 3390.2000 305.8000 ;
      RECT 3384.5000 303.0800 3390.2000 304.1600 ;
      RECT 9.3000 303.0800 3380.9000 304.1600 ;
      RECT 0.0000 303.0800 5.7000 304.1600 ;
      RECT 0.0000 302.6700 3390.2000 303.0800 ;
      RECT 1.1000 301.7700 3390.2000 302.6700 ;
      RECT 0.0000 301.4400 3390.2000 301.7700 ;
      RECT 3388.5000 300.3600 3390.2000 301.4400 ;
      RECT 5.3000 300.3600 3384.9000 301.4400 ;
      RECT 0.0000 300.3600 1.7000 301.4400 ;
      RECT 0.0000 298.7200 3390.2000 300.3600 ;
      RECT 3384.5000 297.6400 3390.2000 298.7200 ;
      RECT 9.3000 297.6400 3380.9000 298.7200 ;
      RECT 0.0000 297.6400 5.7000 298.7200 ;
      RECT 0.0000 296.0000 3390.2000 297.6400 ;
      RECT 3388.5000 294.9200 3390.2000 296.0000 ;
      RECT 5.3000 294.9200 3384.9000 296.0000 ;
      RECT 0.0000 294.9200 1.7000 296.0000 ;
      RECT 0.0000 293.2800 3390.2000 294.9200 ;
      RECT 3384.5000 292.2000 3390.2000 293.2800 ;
      RECT 9.3000 292.2000 3380.9000 293.2800 ;
      RECT 0.0000 292.2000 5.7000 293.2800 ;
      RECT 0.0000 290.5600 3390.2000 292.2000 ;
      RECT 3388.5000 289.4800 3390.2000 290.5600 ;
      RECT 5.3000 289.4800 3384.9000 290.5600 ;
      RECT 0.0000 289.4800 1.7000 290.5600 ;
      RECT 0.0000 287.8400 3390.2000 289.4800 ;
      RECT 3384.5000 286.7600 3390.2000 287.8400 ;
      RECT 9.3000 286.7600 3380.9000 287.8400 ;
      RECT 0.0000 286.7600 5.7000 287.8400 ;
      RECT 0.0000 285.1200 3390.2000 286.7600 ;
      RECT 3388.5000 284.0400 3390.2000 285.1200 ;
      RECT 5.3000 284.0400 3384.9000 285.1200 ;
      RECT 0.0000 284.0400 1.7000 285.1200 ;
      RECT 0.0000 282.4000 3390.2000 284.0400 ;
      RECT 3384.5000 281.3200 3390.2000 282.4000 ;
      RECT 9.3000 281.3200 3380.9000 282.4000 ;
      RECT 0.0000 281.3200 5.7000 282.4000 ;
      RECT 0.0000 279.6800 3390.2000 281.3200 ;
      RECT 3388.5000 278.6000 3390.2000 279.6800 ;
      RECT 5.3000 278.6000 3384.9000 279.6800 ;
      RECT 0.0000 278.6000 1.7000 279.6800 ;
      RECT 0.0000 277.6600 3390.2000 278.6000 ;
      RECT 1.1000 276.9600 3390.2000 277.6600 ;
      RECT 1.1000 276.7600 5.7000 276.9600 ;
      RECT 3384.5000 275.8800 3390.2000 276.9600 ;
      RECT 9.3000 275.8800 3380.9000 276.9600 ;
      RECT 0.0000 275.8800 5.7000 276.7600 ;
      RECT 0.0000 274.2400 3390.2000 275.8800 ;
      RECT 3388.5000 273.1600 3390.2000 274.2400 ;
      RECT 5.3000 273.1600 3384.9000 274.2400 ;
      RECT 0.0000 273.1600 1.7000 274.2400 ;
      RECT 0.0000 271.5200 3390.2000 273.1600 ;
      RECT 3384.5000 270.4400 3390.2000 271.5200 ;
      RECT 9.3000 270.4400 3380.9000 271.5200 ;
      RECT 0.0000 270.4400 5.7000 271.5200 ;
      RECT 0.0000 268.8000 3390.2000 270.4400 ;
      RECT 3388.5000 267.7200 3390.2000 268.8000 ;
      RECT 5.3000 267.7200 3384.9000 268.8000 ;
      RECT 0.0000 267.7200 1.7000 268.8000 ;
      RECT 0.0000 266.0800 3390.2000 267.7200 ;
      RECT 3384.5000 265.0000 3390.2000 266.0800 ;
      RECT 9.3000 265.0000 3380.9000 266.0800 ;
      RECT 0.0000 265.0000 5.7000 266.0800 ;
      RECT 0.0000 263.3600 3390.2000 265.0000 ;
      RECT 3388.5000 262.2800 3390.2000 263.3600 ;
      RECT 5.3000 262.2800 3384.9000 263.3600 ;
      RECT 0.0000 262.2800 1.7000 263.3600 ;
      RECT 0.0000 260.6400 3390.2000 262.2800 ;
      RECT 3384.5000 259.5600 3390.2000 260.6400 ;
      RECT 9.3000 259.5600 3380.9000 260.6400 ;
      RECT 0.0000 259.5600 5.7000 260.6400 ;
      RECT 0.0000 257.9200 3390.2000 259.5600 ;
      RECT 3388.5000 256.8400 3390.2000 257.9200 ;
      RECT 5.3000 256.8400 3384.9000 257.9200 ;
      RECT 0.0000 256.8400 1.7000 257.9200 ;
      RECT 0.0000 255.2000 3390.2000 256.8400 ;
      RECT 3384.5000 254.1200 3390.2000 255.2000 ;
      RECT 9.3000 254.1200 3380.9000 255.2000 ;
      RECT 0.0000 254.1200 5.7000 255.2000 ;
      RECT 0.0000 252.6500 3390.2000 254.1200 ;
      RECT 1.1000 252.4800 3390.2000 252.6500 ;
      RECT 1.1000 251.7500 1.7000 252.4800 ;
      RECT 3388.5000 251.4000 3390.2000 252.4800 ;
      RECT 5.3000 251.4000 3384.9000 252.4800 ;
      RECT 0.0000 251.4000 1.7000 251.7500 ;
      RECT 0.0000 249.7600 3390.2000 251.4000 ;
      RECT 3384.5000 248.6800 3390.2000 249.7600 ;
      RECT 9.3000 248.6800 3380.9000 249.7600 ;
      RECT 0.0000 248.6800 5.7000 249.7600 ;
      RECT 0.0000 247.0400 3390.2000 248.6800 ;
      RECT 3388.5000 245.9600 3390.2000 247.0400 ;
      RECT 5.3000 245.9600 3384.9000 247.0400 ;
      RECT 0.0000 245.9600 1.7000 247.0400 ;
      RECT 0.0000 244.3200 3390.2000 245.9600 ;
      RECT 3384.5000 243.2400 3390.2000 244.3200 ;
      RECT 9.3000 243.2400 3380.9000 244.3200 ;
      RECT 0.0000 243.2400 5.7000 244.3200 ;
      RECT 0.0000 241.6000 3390.2000 243.2400 ;
      RECT 3388.5000 240.5200 3390.2000 241.6000 ;
      RECT 5.3000 240.5200 3384.9000 241.6000 ;
      RECT 0.0000 240.5200 1.7000 241.6000 ;
      RECT 0.0000 238.8800 3390.2000 240.5200 ;
      RECT 3384.5000 237.8000 3390.2000 238.8800 ;
      RECT 9.3000 237.8000 3380.9000 238.8800 ;
      RECT 0.0000 237.8000 5.7000 238.8800 ;
      RECT 0.0000 236.1600 3390.2000 237.8000 ;
      RECT 3388.5000 235.0800 3390.2000 236.1600 ;
      RECT 5.3000 235.0800 3384.9000 236.1600 ;
      RECT 0.0000 235.0800 1.7000 236.1600 ;
      RECT 0.0000 233.4400 3390.2000 235.0800 ;
      RECT 3384.5000 232.3600 3390.2000 233.4400 ;
      RECT 9.3000 232.3600 3380.9000 233.4400 ;
      RECT 0.0000 232.3600 5.7000 233.4400 ;
      RECT 0.0000 230.7200 3390.2000 232.3600 ;
      RECT 3388.5000 229.6400 3390.2000 230.7200 ;
      RECT 5.3000 229.6400 3384.9000 230.7200 ;
      RECT 0.0000 229.6400 1.7000 230.7200 ;
      RECT 0.0000 228.0000 3390.2000 229.6400 ;
      RECT 0.0000 227.0300 5.7000 228.0000 ;
      RECT 3384.5000 226.9200 3390.2000 228.0000 ;
      RECT 9.3000 226.9200 3380.9000 228.0000 ;
      RECT 1.1000 226.9200 5.7000 227.0300 ;
      RECT 1.1000 226.1300 3390.2000 226.9200 ;
      RECT 0.0000 225.2800 3390.2000 226.1300 ;
      RECT 3388.5000 224.2000 3390.2000 225.2800 ;
      RECT 5.3000 224.2000 3384.9000 225.2800 ;
      RECT 0.0000 224.2000 1.7000 225.2800 ;
      RECT 0.0000 222.5600 3390.2000 224.2000 ;
      RECT 3384.5000 221.4800 3390.2000 222.5600 ;
      RECT 9.3000 221.4800 3380.9000 222.5600 ;
      RECT 0.0000 221.4800 5.7000 222.5600 ;
      RECT 0.0000 219.8400 3390.2000 221.4800 ;
      RECT 3388.5000 218.7600 3390.2000 219.8400 ;
      RECT 5.3000 218.7600 3384.9000 219.8400 ;
      RECT 0.0000 218.7600 1.7000 219.8400 ;
      RECT 0.0000 217.1200 3390.2000 218.7600 ;
      RECT 3384.5000 216.0400 3390.2000 217.1200 ;
      RECT 9.3000 216.0400 3380.9000 217.1200 ;
      RECT 0.0000 216.0400 5.7000 217.1200 ;
      RECT 0.0000 214.4000 3390.2000 216.0400 ;
      RECT 3388.5000 213.3200 3390.2000 214.4000 ;
      RECT 5.3000 213.3200 3384.9000 214.4000 ;
      RECT 0.0000 213.3200 1.7000 214.4000 ;
      RECT 0.0000 211.6800 3390.2000 213.3200 ;
      RECT 3384.5000 210.6000 3390.2000 211.6800 ;
      RECT 9.3000 210.6000 3380.9000 211.6800 ;
      RECT 0.0000 210.6000 5.7000 211.6800 ;
      RECT 0.0000 208.9600 3390.2000 210.6000 ;
      RECT 3388.5000 207.8800 3390.2000 208.9600 ;
      RECT 5.3000 207.8800 3384.9000 208.9600 ;
      RECT 0.0000 207.8800 1.7000 208.9600 ;
      RECT 0.0000 206.2400 3390.2000 207.8800 ;
      RECT 3384.5000 205.1600 3390.2000 206.2400 ;
      RECT 9.3000 205.1600 3380.9000 206.2400 ;
      RECT 0.0000 205.1600 5.7000 206.2400 ;
      RECT 0.0000 205.0700 3390.2000 205.1600 ;
      RECT 0.0000 204.1700 3389.1000 205.0700 ;
      RECT 0.0000 203.5200 3390.2000 204.1700 ;
      RECT 3388.5000 202.4400 3390.2000 203.5200 ;
      RECT 5.3000 202.4400 3384.9000 203.5200 ;
      RECT 0.0000 202.4400 1.7000 203.5200 ;
      RECT 0.0000 202.0200 3390.2000 202.4400 ;
      RECT 1.1000 201.1200 3390.2000 202.0200 ;
      RECT 0.0000 200.8000 3390.2000 201.1200 ;
      RECT 3384.5000 199.7200 3390.2000 200.8000 ;
      RECT 9.3000 199.7200 3380.9000 200.8000 ;
      RECT 0.0000 199.7200 5.7000 200.8000 ;
      RECT 0.0000 198.0800 3390.2000 199.7200 ;
      RECT 3388.5000 197.0000 3390.2000 198.0800 ;
      RECT 5.3000 197.0000 3384.9000 198.0800 ;
      RECT 0.0000 197.0000 1.7000 198.0800 ;
      RECT 0.0000 195.3600 3390.2000 197.0000 ;
      RECT 3384.5000 194.2800 3390.2000 195.3600 ;
      RECT 9.3000 194.2800 3380.9000 195.3600 ;
      RECT 0.0000 194.2800 5.7000 195.3600 ;
      RECT 0.0000 192.6400 3390.2000 194.2800 ;
      RECT 3388.5000 191.5600 3390.2000 192.6400 ;
      RECT 5.3000 191.5600 3384.9000 192.6400 ;
      RECT 0.0000 191.5600 1.7000 192.6400 ;
      RECT 0.0000 189.9200 3390.2000 191.5600 ;
      RECT 3384.5000 188.8400 3390.2000 189.9200 ;
      RECT 9.3000 188.8400 3380.9000 189.9200 ;
      RECT 0.0000 188.8400 5.7000 189.9200 ;
      RECT 0.0000 187.2000 3390.2000 188.8400 ;
      RECT 3388.5000 186.1200 3390.2000 187.2000 ;
      RECT 5.3000 186.1200 3384.9000 187.2000 ;
      RECT 0.0000 186.1200 1.7000 187.2000 ;
      RECT 0.0000 184.4800 3390.2000 186.1200 ;
      RECT 3384.5000 183.4000 3390.2000 184.4800 ;
      RECT 9.3000 183.4000 3380.9000 184.4800 ;
      RECT 0.0000 183.4000 5.7000 184.4800 ;
      RECT 0.0000 181.7600 3390.2000 183.4000 ;
      RECT 3388.5000 180.6800 3390.2000 181.7600 ;
      RECT 5.3000 180.6800 3384.9000 181.7600 ;
      RECT 0.0000 180.6800 1.7000 181.7600 ;
      RECT 0.0000 179.0400 3390.2000 180.6800 ;
      RECT 3384.5000 177.9600 3390.2000 179.0400 ;
      RECT 9.3000 177.9600 3380.9000 179.0400 ;
      RECT 0.0000 177.9600 5.7000 179.0400 ;
      RECT 0.0000 177.0100 3390.2000 177.9600 ;
      RECT 1.1000 176.3200 3390.2000 177.0100 ;
      RECT 1.1000 176.1100 1.7000 176.3200 ;
      RECT 3388.5000 175.2400 3390.2000 176.3200 ;
      RECT 5.3000 175.2400 3384.9000 176.3200 ;
      RECT 0.0000 175.2400 1.7000 176.1100 ;
      RECT 0.0000 173.6000 3390.2000 175.2400 ;
      RECT 3384.5000 172.5200 3390.2000 173.6000 ;
      RECT 9.3000 172.5200 3380.9000 173.6000 ;
      RECT 0.0000 172.5200 5.7000 173.6000 ;
      RECT 0.0000 170.8800 3390.2000 172.5200 ;
      RECT 3388.5000 169.8000 3390.2000 170.8800 ;
      RECT 5.3000 169.8000 3384.9000 170.8800 ;
      RECT 0.0000 169.8000 1.7000 170.8800 ;
      RECT 0.0000 168.1600 3390.2000 169.8000 ;
      RECT 3384.5000 167.0800 3390.2000 168.1600 ;
      RECT 9.3000 167.0800 3380.9000 168.1600 ;
      RECT 0.0000 167.0800 5.7000 168.1600 ;
      RECT 0.0000 165.4400 3390.2000 167.0800 ;
      RECT 3388.5000 164.3600 3390.2000 165.4400 ;
      RECT 5.3000 164.3600 3384.9000 165.4400 ;
      RECT 0.0000 164.3600 1.7000 165.4400 ;
      RECT 0.0000 162.7200 3390.2000 164.3600 ;
      RECT 3384.5000 161.6400 3390.2000 162.7200 ;
      RECT 9.3000 161.6400 3380.9000 162.7200 ;
      RECT 0.0000 161.6400 5.7000 162.7200 ;
      RECT 0.0000 160.0000 3390.2000 161.6400 ;
      RECT 3388.5000 158.9200 3390.2000 160.0000 ;
      RECT 5.3000 158.9200 3384.9000 160.0000 ;
      RECT 0.0000 158.9200 1.7000 160.0000 ;
      RECT 0.0000 157.2800 3390.2000 158.9200 ;
      RECT 3384.5000 156.2000 3390.2000 157.2800 ;
      RECT 9.3000 156.2000 3380.9000 157.2800 ;
      RECT 0.0000 156.2000 5.7000 157.2800 ;
      RECT 0.0000 154.5600 3390.2000 156.2000 ;
      RECT 3388.5000 153.4800 3390.2000 154.5600 ;
      RECT 5.3000 153.4800 3384.9000 154.5600 ;
      RECT 0.0000 153.4800 1.7000 154.5600 ;
      RECT 0.0000 151.8400 3390.2000 153.4800 ;
      RECT 0.0000 151.3900 5.7000 151.8400 ;
      RECT 3384.5000 150.7600 3390.2000 151.8400 ;
      RECT 9.3000 150.7600 3380.9000 151.8400 ;
      RECT 1.1000 150.7600 5.7000 151.3900 ;
      RECT 1.1000 150.4900 3390.2000 150.7600 ;
      RECT 0.0000 149.1200 3390.2000 150.4900 ;
      RECT 3388.5000 148.0400 3390.2000 149.1200 ;
      RECT 5.3000 148.0400 3384.9000 149.1200 ;
      RECT 0.0000 148.0400 1.7000 149.1200 ;
      RECT 0.0000 146.4000 3390.2000 148.0400 ;
      RECT 3384.5000 145.3200 3390.2000 146.4000 ;
      RECT 9.3000 145.3200 3380.9000 146.4000 ;
      RECT 0.0000 145.3200 5.7000 146.4000 ;
      RECT 0.0000 143.6800 3390.2000 145.3200 ;
      RECT 3388.5000 142.6000 3390.2000 143.6800 ;
      RECT 5.3000 142.6000 3384.9000 143.6800 ;
      RECT 0.0000 142.6000 1.7000 143.6800 ;
      RECT 0.0000 140.9600 3390.2000 142.6000 ;
      RECT 3384.5000 139.8800 3390.2000 140.9600 ;
      RECT 9.3000 139.8800 3380.9000 140.9600 ;
      RECT 0.0000 139.8800 5.7000 140.9600 ;
      RECT 0.0000 138.2400 3390.2000 139.8800 ;
      RECT 3388.5000 137.1600 3390.2000 138.2400 ;
      RECT 5.3000 137.1600 3384.9000 138.2400 ;
      RECT 0.0000 137.1600 1.7000 138.2400 ;
      RECT 0.0000 135.5200 3390.2000 137.1600 ;
      RECT 3384.5000 134.4400 3390.2000 135.5200 ;
      RECT 9.3000 134.4400 3380.9000 135.5200 ;
      RECT 0.0000 134.4400 5.7000 135.5200 ;
      RECT 0.0000 132.8000 3390.2000 134.4400 ;
      RECT 3388.5000 131.7200 3390.2000 132.8000 ;
      RECT 5.3000 131.7200 3384.9000 132.8000 ;
      RECT 0.0000 131.7200 1.7000 132.8000 ;
      RECT 0.0000 130.0800 3390.2000 131.7200 ;
      RECT 3384.5000 129.0000 3390.2000 130.0800 ;
      RECT 9.3000 129.0000 3380.9000 130.0800 ;
      RECT 0.0000 129.0000 5.7000 130.0800 ;
      RECT 0.0000 127.3600 3390.2000 129.0000 ;
      RECT 0.0000 126.3800 1.7000 127.3600 ;
      RECT 3388.5000 126.2800 3390.2000 127.3600 ;
      RECT 5.3000 126.2800 3384.9000 127.3600 ;
      RECT 1.1000 126.2800 1.7000 126.3800 ;
      RECT 1.1000 125.4800 3390.2000 126.2800 ;
      RECT 0.0000 124.6400 3390.2000 125.4800 ;
      RECT 3384.5000 123.5600 3390.2000 124.6400 ;
      RECT 9.3000 123.5600 3380.9000 124.6400 ;
      RECT 0.0000 123.5600 5.7000 124.6400 ;
      RECT 0.0000 121.9200 3390.2000 123.5600 ;
      RECT 3388.5000 120.8400 3390.2000 121.9200 ;
      RECT 5.3000 120.8400 3384.9000 121.9200 ;
      RECT 0.0000 120.8400 1.7000 121.9200 ;
      RECT 0.0000 119.2000 3390.2000 120.8400 ;
      RECT 3384.5000 118.1200 3390.2000 119.2000 ;
      RECT 9.3000 118.1200 3380.9000 119.2000 ;
      RECT 0.0000 118.1200 5.7000 119.2000 ;
      RECT 0.0000 116.4800 3390.2000 118.1200 ;
      RECT 3388.5000 115.4000 3390.2000 116.4800 ;
      RECT 5.3000 115.4000 3384.9000 116.4800 ;
      RECT 0.0000 115.4000 1.7000 116.4800 ;
      RECT 0.0000 113.7600 3390.2000 115.4000 ;
      RECT 3384.5000 112.6800 3390.2000 113.7600 ;
      RECT 9.3000 112.6800 3380.9000 113.7600 ;
      RECT 0.0000 112.6800 5.7000 113.7600 ;
      RECT 0.0000 111.0400 3390.2000 112.6800 ;
      RECT 3388.5000 109.9600 3390.2000 111.0400 ;
      RECT 5.3000 109.9600 3384.9000 111.0400 ;
      RECT 0.0000 109.9600 1.7000 111.0400 ;
      RECT 0.0000 108.3200 3390.2000 109.9600 ;
      RECT 3384.5000 107.2400 3390.2000 108.3200 ;
      RECT 9.3000 107.2400 3380.9000 108.3200 ;
      RECT 0.0000 107.2400 5.7000 108.3200 ;
      RECT 0.0000 105.6000 3390.2000 107.2400 ;
      RECT 3388.5000 104.5200 3390.2000 105.6000 ;
      RECT 5.3000 104.5200 3384.9000 105.6000 ;
      RECT 0.0000 104.5200 1.7000 105.6000 ;
      RECT 0.0000 102.8800 3390.2000 104.5200 ;
      RECT 3384.5000 101.8000 3390.2000 102.8800 ;
      RECT 9.3000 101.8000 3380.9000 102.8800 ;
      RECT 0.0000 101.8000 5.7000 102.8800 ;
      RECT 0.0000 101.3700 3390.2000 101.8000 ;
      RECT 1.1000 100.4700 3389.1000 101.3700 ;
      RECT 0.0000 100.1600 3390.2000 100.4700 ;
      RECT 3388.5000 99.0800 3390.2000 100.1600 ;
      RECT 5.3000 99.0800 3384.9000 100.1600 ;
      RECT 0.0000 99.0800 1.7000 100.1600 ;
      RECT 0.0000 97.4400 3390.2000 99.0800 ;
      RECT 3384.5000 96.3600 3390.2000 97.4400 ;
      RECT 9.3000 96.3600 3380.9000 97.4400 ;
      RECT 0.0000 96.3600 5.7000 97.4400 ;
      RECT 0.0000 94.7200 3390.2000 96.3600 ;
      RECT 3388.5000 93.6400 3390.2000 94.7200 ;
      RECT 5.3000 93.6400 3384.9000 94.7200 ;
      RECT 0.0000 93.6400 1.7000 94.7200 ;
      RECT 0.0000 92.0000 3390.2000 93.6400 ;
      RECT 3384.5000 90.9200 3390.2000 92.0000 ;
      RECT 9.3000 90.9200 3380.9000 92.0000 ;
      RECT 0.0000 90.9200 5.7000 92.0000 ;
      RECT 0.0000 89.2800 3390.2000 90.9200 ;
      RECT 3388.5000 88.2000 3390.2000 89.2800 ;
      RECT 5.3000 88.2000 3384.9000 89.2800 ;
      RECT 0.0000 88.2000 1.7000 89.2800 ;
      RECT 0.0000 86.5600 3390.2000 88.2000 ;
      RECT 3384.5000 85.4800 3390.2000 86.5600 ;
      RECT 9.3000 85.4800 3380.9000 86.5600 ;
      RECT 0.0000 85.4800 5.7000 86.5600 ;
      RECT 0.0000 83.8400 3390.2000 85.4800 ;
      RECT 3388.5000 82.7600 3390.2000 83.8400 ;
      RECT 5.3000 82.7600 3384.9000 83.8400 ;
      RECT 0.0000 82.7600 1.7000 83.8400 ;
      RECT 0.0000 81.1200 3390.2000 82.7600 ;
      RECT 3384.5000 80.0400 3390.2000 81.1200 ;
      RECT 9.3000 80.0400 3380.9000 81.1200 ;
      RECT 0.0000 80.0400 5.7000 81.1200 ;
      RECT 0.0000 78.4000 3390.2000 80.0400 ;
      RECT 3388.5000 77.3200 3390.2000 78.4000 ;
      RECT 5.3000 77.3200 3384.9000 78.4000 ;
      RECT 0.0000 77.3200 1.7000 78.4000 ;
      RECT 0.0000 75.6800 3390.2000 77.3200 ;
      RECT 3384.5000 74.6000 3390.2000 75.6800 ;
      RECT 9.3000 74.6000 3380.9000 75.6800 ;
      RECT 0.0000 74.6000 5.7000 75.6800 ;
      RECT 0.0000 72.9600 3390.2000 74.6000 ;
      RECT 3388.5000 71.8800 3390.2000 72.9600 ;
      RECT 5.3000 71.8800 3384.9000 72.9600 ;
      RECT 0.0000 71.8800 1.7000 72.9600 ;
      RECT 0.0000 70.2400 3390.2000 71.8800 ;
      RECT 3384.5000 69.1600 3390.2000 70.2400 ;
      RECT 9.3000 69.1600 3380.9000 70.2400 ;
      RECT 0.0000 69.1600 5.7000 70.2400 ;
      RECT 0.0000 67.5200 3390.2000 69.1600 ;
      RECT 3388.5000 66.4400 3390.2000 67.5200 ;
      RECT 5.3000 66.4400 3384.9000 67.5200 ;
      RECT 0.0000 66.4400 1.7000 67.5200 ;
      RECT 0.0000 64.8000 3390.2000 66.4400 ;
      RECT 3384.5000 63.7200 3390.2000 64.8000 ;
      RECT 9.3000 63.7200 3380.9000 64.8000 ;
      RECT 0.0000 63.7200 5.7000 64.8000 ;
      RECT 0.0000 62.0800 3390.2000 63.7200 ;
      RECT 3388.5000 61.0000 3390.2000 62.0800 ;
      RECT 5.3000 61.0000 3384.9000 62.0800 ;
      RECT 0.0000 61.0000 1.7000 62.0800 ;
      RECT 0.0000 59.3600 3390.2000 61.0000 ;
      RECT 3384.5000 58.2800 3390.2000 59.3600 ;
      RECT 9.3000 58.2800 3380.9000 59.3600 ;
      RECT 0.0000 58.2800 5.7000 59.3600 ;
      RECT 0.0000 56.6400 3390.2000 58.2800 ;
      RECT 3388.5000 55.5600 3390.2000 56.6400 ;
      RECT 5.3000 55.5600 3384.9000 56.6400 ;
      RECT 0.0000 55.5600 1.7000 56.6400 ;
      RECT 0.0000 53.9200 3390.2000 55.5600 ;
      RECT 3384.5000 52.8400 3390.2000 53.9200 ;
      RECT 9.3000 52.8400 3380.9000 53.9200 ;
      RECT 0.0000 52.8400 5.7000 53.9200 ;
      RECT 0.0000 51.2000 3390.2000 52.8400 ;
      RECT 3388.5000 50.1200 3390.2000 51.2000 ;
      RECT 5.3000 50.1200 3384.9000 51.2000 ;
      RECT 0.0000 50.1200 1.7000 51.2000 ;
      RECT 0.0000 48.4800 3390.2000 50.1200 ;
      RECT 3384.5000 47.4000 3390.2000 48.4800 ;
      RECT 9.3000 47.4000 3380.9000 48.4800 ;
      RECT 0.0000 47.4000 5.7000 48.4800 ;
      RECT 0.0000 45.7600 3390.2000 47.4000 ;
      RECT 3388.5000 44.6800 3390.2000 45.7600 ;
      RECT 5.3000 44.6800 3384.9000 45.7600 ;
      RECT 0.0000 44.6800 1.7000 45.7600 ;
      RECT 0.0000 43.0400 3390.2000 44.6800 ;
      RECT 3384.5000 41.9600 3390.2000 43.0400 ;
      RECT 9.3000 41.9600 3380.9000 43.0400 ;
      RECT 0.0000 41.9600 5.7000 43.0400 ;
      RECT 0.0000 40.3200 3390.2000 41.9600 ;
      RECT 3388.5000 39.2400 3390.2000 40.3200 ;
      RECT 5.3000 39.2400 3384.9000 40.3200 ;
      RECT 0.0000 39.2400 1.7000 40.3200 ;
      RECT 0.0000 37.6000 3390.2000 39.2400 ;
      RECT 3384.5000 36.5200 3390.2000 37.6000 ;
      RECT 9.3000 36.5200 3380.9000 37.6000 ;
      RECT 0.0000 36.5200 5.7000 37.6000 ;
      RECT 0.0000 34.8800 3390.2000 36.5200 ;
      RECT 3388.5000 33.8000 3390.2000 34.8800 ;
      RECT 5.3000 33.8000 3384.9000 34.8800 ;
      RECT 0.0000 33.8000 1.7000 34.8800 ;
      RECT 0.0000 32.1600 3390.2000 33.8000 ;
      RECT 3384.5000 31.0800 3390.2000 32.1600 ;
      RECT 9.3000 31.0800 3380.9000 32.1600 ;
      RECT 0.0000 31.0800 5.7000 32.1600 ;
      RECT 0.0000 29.4400 3390.2000 31.0800 ;
      RECT 3388.5000 28.3600 3390.2000 29.4400 ;
      RECT 5.3000 28.3600 3384.9000 29.4400 ;
      RECT 0.0000 28.3600 1.7000 29.4400 ;
      RECT 0.0000 26.7200 3390.2000 28.3600 ;
      RECT 3384.5000 25.6400 3390.2000 26.7200 ;
      RECT 9.3000 25.6400 3380.9000 26.7200 ;
      RECT 0.0000 25.6400 5.7000 26.7200 ;
      RECT 0.0000 24.0000 3390.2000 25.6400 ;
      RECT 3388.5000 22.9200 3390.2000 24.0000 ;
      RECT 5.3000 22.9200 3384.9000 24.0000 ;
      RECT 0.0000 22.9200 1.7000 24.0000 ;
      RECT 0.0000 21.2800 3390.2000 22.9200 ;
      RECT 3384.5000 20.2000 3390.2000 21.2800 ;
      RECT 9.3000 20.2000 3380.9000 21.2800 ;
      RECT 0.0000 20.2000 5.7000 21.2800 ;
      RECT 0.0000 18.5600 3390.2000 20.2000 ;
      RECT 3388.5000 17.4800 3390.2000 18.5600 ;
      RECT 5.3000 17.4800 3384.9000 18.5600 ;
      RECT 0.0000 17.4800 1.7000 18.5600 ;
      RECT 0.0000 15.8400 3390.2000 17.4800 ;
      RECT 3384.5000 14.7600 3390.2000 15.8400 ;
      RECT 9.3000 14.7600 3380.9000 15.8400 ;
      RECT 0.0000 14.7600 5.7000 15.8400 ;
      RECT 0.0000 13.1200 3390.2000 14.7600 ;
      RECT 3388.5000 12.0400 3390.2000 13.1200 ;
      RECT 5.3000 12.0400 3384.9000 13.1200 ;
      RECT 0.0000 12.0400 1.7000 13.1200 ;
      RECT 0.0000 10.4000 3390.2000 12.0400 ;
      RECT 3384.5000 9.3200 3390.2000 10.4000 ;
      RECT 9.3000 9.3200 3380.9000 10.4000 ;
      RECT 0.0000 9.3200 5.7000 10.4000 ;
      RECT 0.0000 9.3000 3390.2000 9.3200 ;
      RECT 3384.5000 5.7000 3390.2000 9.3000 ;
      RECT 0.0000 5.7000 5.7000 9.3000 ;
      RECT 0.0000 5.3000 3390.2000 5.7000 ;
      RECT 3388.5000 1.7000 3390.2000 5.3000 ;
      RECT 0.0000 1.7000 1.7000 5.3000 ;
      RECT 0.0000 0.0000 3390.2000 1.7000 ;
    LAYER met4 ;
      RECT 0.0000 2887.9600 3390.2000 2889.6600 ;
      RECT 5.3000 2883.9600 3384.9000 2887.9600 ;
      RECT 3384.5000 5.7000 3384.9000 2883.9600 ;
      RECT 9.3000 5.7000 3380.9000 2883.9600 ;
      RECT 5.3000 5.7000 5.7000 2883.9600 ;
      RECT 3388.5000 1.7000 3390.2000 2887.9600 ;
      RECT 5.3000 1.7000 3384.9000 5.7000 ;
      RECT 0.0000 1.7000 1.7000 2887.9600 ;
      RECT 0.0000 0.0000 3390.2000 1.7000 ;
  END
END eFPGA_top

END LIBRARY
